PK   ��OXϚ�  T�     cirkitFile.json�][sۺ�+��>�,.��1i;�4i<�N�`{4��1���RT�s2�� ��,R��+9m	�.��o���4�w=��FO��fQ�g��Qp�5�}���F�]=���ɷ&��	�~��a�������|�g�D�j��0)re�d�J�B�c�A�J���.�G�&�8r�#�8r�#W8�G��y�#�����- �H�{� �H���_�P9SQ�ÒU(�<	Ӭ�a�$Q�E���a<��q���H�r90�y\�I��*�$��`a�S�9�E%��k~��\&f�J���(�Da�RY˘�(*m���H����m{��C��8��8���Aj���6�A�@��z�\'�b�^��՞���/�C���"$7.�h��u�ڽ�Мy�눛6!E�Оr#②��\Z0��0Cs,��<��O�2�~c�_���p$\$	F�E�p�H��$\.)	�Q�� ��XИ� h 4�CqUa}'�9�'�A1�A1�A1�A1�P\U64(�4(�4�X��1�
ǆł( �A��A��A���ł�� �}V.pþ)(�,��T��s] �����7��/�o޶���`�쮳�E���M���m�)2��s$\$	F�E�p�H��$\.)	�Q�� ��XИ� h 4�9�9�'�A1�A1�A1�A1�A1�A1�A1�A��A��A� 
HhP,hP,hP,hP,hP,��;��s9>�l
�� ���)<����M��Ȳ�#�M��v�35����Qp_7z1��f�.'&ۚ7�n���ލ�4�\�Q�e�L �\�$d"�yUȸ��Z	�G�C{ъ��}GEj��x	9�/y��E�IYid��"LR^��Jf,2�L�804��+$�P����<=�
���t��`p`hO��e���E�1k��i��9.���BY���=G�������La��pլc�[�Q��й4�r&��q�����$�$�TC(�yСxQܳ�Ը{��e��|��>Nh�F�$��=&�ړ���g�u�x�w��$�ǈ�����Ն�T���M�7��������w]N�Y�Ws�4B�]��ڎ~	|]�^NS�p"Џ�W�ё-��(xlI�lef�')��|�e�`c����j�W�So�`k8x	���؊^la���2^ l�/��s���;D;����_���0@֢�����7J=vA,�@�	�roB|�2T9�\J������'IT����_fx�$	�0��H$� 0zkL�`��><s+\� >��=�		� 
<S*
	0Z �Fb`��3�>�:�R$�Y��K�Q/��<�Ia��bEf��>�+�Iv�Z� ��<`Up ��P%Hё���+^��4�xO��?������N����(�o��+X����Q�5岞uǩ���#�����.�'�'�5I/��Iϐ�
I!�c$}��O��U `XÀ1`QX���;�̶�a��8��Z���X`������paq��:?��
�[�u���)A>=�`a+��T`q*��T`�)� ���2��a�}|#���d�'���ü^�g�p���tއ�����)�U<��5�����῰���훀�>-Ĭlv��-�hl���l�ږ��v����l�`{�����s������R��[
Wve8n)�6��'p�d)���BX
W���J��`{�N��.�-���Z^[�+h{$����J!3�Z}LV��Q!�e���=g��P?�<˳ki��}@����J�W����:5�[�Qu��Y��5�,�Sk�f�C��&vq�.��K��ؽ$/��K��{_6�N�Fge>�{l��O���]��n&��̴�tM���N7m��K�o��/���إ�h� I�$�H��	�42�4:�DZei��2eH�0-u�\'Y��b��t|}��1>
�Z�f�b��kE�6\���A9��Y�uSL��]
��j$Ru=z�,��?�v�n�F��'�hO�튭�l�6����TCW��Ͷ���{�>�"��+�t�n���%�O/��K�O��>9��O+}�O�k�]����-yj[��}��������]��ߞ��(��|�[��-b^��t�׭G)}�����G��v��ﺽh�e=�l7�����Ǐ�w3�����m��7c����~�WG��l�����yIu�I������si9���
̧������ 8���B���|�u>�][����m|H�,�qc��lYeE�lt�O��nk�>����>t��@�mǪx<�13K�,3ѵ3M�!U�ĺ�1�P��C��8V��Ӵ�u��̙z�^�T�uP�F���熔��%�{L���<�ſ ��7�4�C����1Di��\�1�d�S޵���9�� -�B�,̅�Vab�0��вd`��(���9��w;x� ���-�['���'�l,�c)�uc�F*6��Z׳����y��2��P�+���[ZJ�E����x�`��T܅��`�%]K�� &��|��C�e#��rV:{j�wV�"˘�x�+O3�8ᩴ��}]�7�M��,��*�F��n\G%�����xF��o��gō.�w��y���������=�lC��W�{�Upv����`te,-k��z��t�^��:nzV��嗕:VMvA*�a�:�����=�������U`3�/չ�p���¶�]ڿ�A�� j��0��Si��5�v�~�
P~����L�/��Q����ז���3b?�V?K@	 ���Q6*� �Nm��m���^��H�FD�5���(�נP�ɹ{չ�[^�����uB�C�t�z&��e�P���)���}�d�i�~��Bc;-��Ş����o�xȯnL�揟�F����f�g���^��iQ=�~�>g�nj�z���`e����I������V�.�]?�PK   ��OX��8��9 z /   images/11b938df-2630-4b82-9eb5-abaaeee165cf.pngT\\��׎�j[�4[AY6D������b+��
"�@Dd�����(5D@YVT� �M�(�+#�a�,�! {}�!��_�S���3���������|���op8ܷ��ZF8��|������&��K�_Hg��__]��߿v=i��I=G��y�p����󄙧��%O�9w;�BQppv��p��N���>vDc;�G����O�P��Ĕu�|��vj�����m�w=�*24��o�R���惐w����)\�|�e�|���5�������/W��*���ϯ]��H;h�I��G���W�놮صr�(���?�ޒ�f����ok�5)h48!�~b��Gݘ�8?5L�>��ޡ�o��p,^����V��"T�-�X��;Ğ��QU�əc'�f^Mɍ"��-r���g�2��K����ٓ�9�S�ǔ:y�C���(b����Jb���zE�'"%ʤ�����	��/F��#��a��ҕ��1�x��3��=H�ކ�=�	�z�7�=���%4���<��g�[l@��[���;u���Z&#�g�g��wV���{�����$Cl�.���9�Of[�������j]�Xob�y��CF�b�f �~�)�'�"f"v��ҋ�,x7�=��Z�,��ԅOz�3[H#�´�B^�����#k\,-�C��x�7/�:j�:
��brc��H�,�1�c��T�l�G=+�(��BQ�y53���i���xӣްo�g�8�3��SF��T�h�͎a�x_����Q����[�c?��r��E���V�MO*�|4Z����#n|�Pd��ޫi�6�Q/YC<P��}���^�Ǟ�t�\�&���6���fɍ�Il�p�?^
�Jh[��klp�� �U\��>���3�o��zﱭc�S`hݤ$��A!M���������/���3p�.��F.�����qpSE��Byy����<zA�=��e3žk3�ß�e)	�$�wpՉI����9�M�C�ןM2&�軛�Y�g�J-;��n��6��0�4�)��a�ԱTȞ20p�T+R�7֐���0��r96�vsm��%�FR޳��9O��"kvn��_r0�vL������=Ց��m(��a�Pk�}uCCC$dt$`��\�t���JR�J͗������g���x���e�[�I,p������\:�BR(�FRb�r�"I	�{n�å�$n�Y ��/���/����c8���o���{��TD"�"%}��ɸ��Z� Kb��e��2.���,V�|���2��͈N߁�7°���GX�����e�9_�Q���c>�,F�J�D���ʼ�;�8�d�/�M��z�&���r��t�m�m�Y�����Sgi�����?>���u��Kw��6��|>|�G�CW�/��ٻ�C�[/n�E�`XѨ�h��s�k����.�~ž�.[P�m���Ȧ.�t�E���nnnO~�
>������;���=��#l�'�~����B��n���l����6�u'	�"��Q�z�63�u�lW��k֦6d�ni�|/ �è�c�'`���T�GR;�vMׂZTox\�ֱ�ǯ�Ʒ�#1�����E�&>��lbs�o���8�����[����=Gqf�;���(�<�Xra��6$\�{��4Vɻ��|�Bb�7�����_R�� ���_�VWWK�[YY]��h/Ύ�N��555�7�?}"�"֫N/LЯ�������J9sw��
̀��
�BA/��Y�h@�v`������Ԥ_I{.g���?��n��`%�����1�SO>��}$='''$�67	��~w�oA�ĿP8'��F}4:,u�˗n-���D+��$wG��kc��k�8�x�XE��c�uNcf;�S�Q�]Ҕ�l�L�v�Ǐ�;3z9�sKO��^9a�y��H�J��U�Rh�L���@J�q���_�j���O.�-��E.��+l�{���#"y4`����_�O6S�MJJJ�{g�����"���զp�mw{��}���w3��/�=:�
�8�޸w�^r����+�QF#�9��+���/��r�=�к.�;�~�~�?h�Â�Ni�Mz�Xdy��6[���^j#F0X�����Xp�2��JШw���.� �������wwLs�T��|L�'�,x&LFjd�9��%k.mG���L��?�����C(G�@qөŸ��ã��nf�{��ߌ�r<��9t�Cp�Ym?}a����rJn:X���;��X��2ކ���E��H+k���fRǍy�pdk���f��Ͳ��z.�;;;�9m�bϷ[�*����vj�fBӁop����=y��㹜�7n�7q�a��c3�p�����n�U|���]�gz�ˊ"��'Q�����ʖ�u�	��[�����ʕ�ά�u���\�{�)��]�Iyv�0��#-��,��wW��ܴ����K(KY��~~4_���:�\Nj$�pol~'�!#N��sy&����)��,=���
����)#q�"*��Ƌ��q9���N� ��G��f$o�Д��,�����Ɗ���dI��|���=���\�pw�s�^�.60�-����ptʃ#.g��i���6��&Ñ��BJv�����|nT���a��網�m�Z9����8Յ���Օ�A�4,�HG������!��g����8��u?&ikJl\(u�ߎ�<Ӹ�S]1gA���(�Ԧ�:�:�g�����?22��r���!�)��4�$y��G=;���q�b�1�ӣ����SX�2��~�����xP�)��u�����i��oa@HW�G��J��6*�i}p'?�:����Aq�"�P���Ak����U��Is��,֬�q�̻z���#tތ'��oQ�!���sQii(V��Xù����K�<F�"�~���&;��Cj�Ë���F@�ARFzn��|�8�mN�Y�d��|���Q��]�'M���k�����������7,�2�@���l3r<��_so-�/�]��0/�4�	r(�w��"�{iai��[��"r�cz�����?���a�';��ߍ�'�m�.�>5w�ǂw���x1��{H�iɽ�bgn���*��>���	���a�9�G.'�`N��@��]u��a���9���L�=	�c_�k������[�XyD�ٻ���*X&&&���c�ӹ�-����H{���{��h���=X|G��Dt�:�~�4Z�8�5dae`F¸���p��%��F����ö�/�"����˦�v t:A���>ڌ���N,gdkhح���FU��Ҹ��!�&�'�I�������g]mu�z}GF��k+},��M�ӊ����S���ƋŞ�S���"���f4-�������c��E��ҋ0�T_I����+�78�A�\�ƓƗ��F���b�:bsL;щ�M|ks?L��4YL�5��Yp���N�M ��ر�>$�yY��$��]�_~��@"t���L�������Y�k�j�=�q{Ҕ�������
�� ��|�n�:�d,]>07n�+����5Rpi�u����`y��{��S�0���v��տ�i�YN_oed��Z|  ������G��C�Q���`(�vVg�� f?.�/r/?��&�*�{Q�Q���N��5L�B���.���X,�XOq=][S3$�=O�H4�����&fN_�"��T�I��>0�'����C%�I�5�?ϗQ@��#�2���X�����VK, ���s:N�:em�[P��V��4���}���p�m�E�i,�"y�&9
X���Fdα(#TN�2��{_�vT�O�W0���D�?�!�)�� ���$�'�#�vd��4�:v�����qXN&M0���}n�*�_��B*+�P4�:u,9Z���-f�I�5�H.��(��$R�i�L��]�55+�e2���ʧǢL*���.cdkV.KlZ?����ـ����"I��r��!|Ov�㕦,FEw�XiZq���nޕ�i8^��uf�X揲���M�|Y��_kk�X�ce����I�zJ�wL���pA�}��3��%_|:6!h�O��#�&\<ރz�OZT��	��~��E�*�]0���0���=�J:<"���#�����M�*�'I�8,�i3�	/�����#�SW���$9����u@�h�b����}puk����hW�����i�������"��D���T���-��aG��}S��Q��d�i8�s/J1��F/�J����BN~�G��"D�E��R���7�5���y�1�;�r��u������23r�r�-�ɖ���O�0��ڏX{��Yp���#}��ǎ�Hr�&?��6�mF����J,��+�3����zD�.����8��`'z:V��K��
p��m�{4PLcEC��S��o �ѿ�0�
#��L� M�����k>��h��(��5bNq�`��?�P4��F^^}ػ���]c�྿��J�J�E���̣,����7o0L\ņ�ܴdH��0^jL�v�������Жg�aj5M�]v!�H��FR����}r����АƊf��u��ܿ���΂�a��yH+��'�r/66�	�B�=�~4t��8�(�ʕ���3� ���S�(7^���0J���@�%PomcD��{E�wj�t��GDV�E�=L���t"6c%ʾB�j'�<7ϩ1���\!�s{�;Tr�`�y;�n�u-4#���x �N%"�FS��d1F�v�GH����܎�s/n�q���e�����pҫ�&�L�M�E��")8�aSv��B��=�"���e�R��<��!L���
����|.'�`���c>d�򗋨��u=c3�����C�����Q�EiP���ɮz<1���r@0g|�TS��u���#��B����-��<�>D�a	�Jz��g2�.���{*-���8��*Pc$6�^�D��K\j���7�r9�V��hZ��B\����n�!%��)u�%�<��a~j8r˖-��ƺ{7u�#��?���f���閬�ŏ�_$�ӷ!�W��nU�dg��|�6�9\��4;;K��籮��]������S�å�8sN$�\����-���7H��=Oݢ��#�n�}˳�.��S[��KR��ʃ�H�}�F��-���E�����`���ݗ��}�Thh���^&�T�Rccjn�:����;�%�"�Nއ�zP`�I�J��ԓ�d<n��E���J�Low�n��?�V!�<�����p�SM1#�T�R�߇��QFM������<���/�c;�ѶA����%�7,x��v���k*0��m
R�4��#�aV�AYg����þ�<��qg7�����N�F�����ᰧZ����	�|�67[� Ȗ��J���\l�N\���I۝I^��@�;]��#*���(HY�1~�i��ao[��)�1�������mgtg]<<<��������9P�>zr����q�%$�wž�إV۩�j#H�-Ej�����h��᭑ɍ��h����0�ʶ����nwL�4����a��g���:~՝M��3�*�P){?��?�S�� �_%���+-u�]�oZ�z�:Y�2�D׏НG,xz��;���˺$����	s���[wy {Yl{�c�#G��]%���"�R����O�3� �)���*��Z,�WVGj0����9�r:�f�{!noo?����	(6l5��?�^UZ��L�-%T�v�bא�a���@͝��F�<��β���`�lg���:��3d��''+�#D��!G�����b���&�<��,��n���A�y�b+�SI�]�]�6���g�z��RW�w�� �D=���g�����E�	�Z�f�(�G�����ז�2>[�Q��-r���q�|�)��2� ˢ/>�B~`���S3��������H}>�P�:l��ۃ��s����M�r��{�8�N�_uU����ʿc����Ypb2��+��h`3��GGGw�.̌]�o��Cg���GO�Ӊ[�P&���[��TH(�zl�&�18�ǥ\H�,ҕ�w��&α��O��� b��2��C��1���$���M��3����;�O�ʂ��'�2B[�Jקq�'8��u�֎̎�Mr�/ہ8w���/�_'±Hl��Sp=�c{?1q9�X�����w��hJn��|(�F~�SCf.�ONVWW����"�xw�,���7�a0^B��_|���~|m@��H��_�(�l?lbw}���T�����!��`J\bb�)_R�ӱzU��~���.RL����;��'�[v��x���M+򖜎�"UCH�б����Wr8G�#��3�����X��e�Q��#�ӄ�P�����|��z���9R_[[��Yo���GU+��?Ć���-)�c|��1���e�@�*�c�\�֋}�_����gF~����]�s%}����� �䁿������
&6�����Aܲ��}�-r�/߻��#P��
�𰹣cz���u�/0��L
�א*�FW3��lUZW�
;�@�E�c��pY��e���6�**���|�I���ɶF��w��=#-��1�쀦�r,IC���-�v��Ӡ��q掓�YX��8p��˲�x�i�z�r�d�՝�";�AT_�	��*}ݕl���o�A�_YYi�U�>j0�D:ħ �Iw��W�`+33���?��oz��ca{�����D)Mߞ���>i�ل�v�W��X��"�3���� ��xEZz�8�P����Q��D�l�\7(НL���x�8C�5b���Q}#Kl�Il���d�]#P�ω�+��*�(�g�rn��{"�x���Gl�q������qq��y�%�ԍ���/���Tp.u�e0kF����k ��Z���E�.;�GX/x��0[3lD'�NJmȰ.R����+5��M��bܿ����}L,�)���cޤ�GS?�u?����������q1̨�1�(]RXC&��������/"�..�8�"g�G
�
Z��_�[~�[�1 ^�3j8^KR�w����Pi��[����3��:��=�$ �7?i�(z��J��!/��������X�����u�Q��tL�<0�Kb�M�`Y�8�e-�h�3��Y�`Ge�Hȋ�|k��ԗ�|�+�E�V���x1��B���]
Z)��'g'>��l�>�ý�f�+����@�g�a�f�T�r>8�w����Ϊ������b:M�8��ܲB�@.��?
]ZrsH0G�nf�����	��h�[����H��r��0��b��� �����Vb�qn(�@p0�;t���]]�ǋ�D�x�[��1l8^��u�%�8қU��ss9���v�غ�P
�0v�C�%;a''��N�Q��X����v9_Gz�&A�������N�@dz�y����m����g"E����
�O�>N}�.�{CTo�[�`Dgy�KǢ��^���3Rw�<y�
]0�e�䛪�-[��+So|�%�^�Z�҂a�~s�$�E�a��S�l�'[�����_��Em~��0s�{������xq6z�U~A������|��z*"���=�Y����\�;P��}0��9�\���O���˴�mv|�~t� �����>E�8IFU���*!ѥlq
��Ի���)�ФC�<���\�s�V*���1Jۄ��
:؎�9{�X�������0CV�/@H�K�4Mf�hY>g�����p$#]_�����),��w(�T��~~~��}���v�9�D.1�rrr����3�dIe�#���Ƞ꜋�U�\��Z��:���+��������S���x~��6�n�;��t���C�V�@�6��n�,��P�����59N�獀��<'����?u��~��� ����^9�5A�4.@ɔۆ�N;@\J����E�^��/���X�y-V,�˾����i[+��A��J���>a��3A�w�T5��ܽ����Ś�xe%ta�PT��**��1�؂]R���4�*�^��[������=E ��0�L��hXҘl�|Y��Vn0�:�:��,߉�����O<�>�s}�K���# v���.� _2�0������Y���b���\N��ٶ���[R�8�	,~3���w���ӧ	]y����+,�����\*���{�_[!���	V�A�D#�t�R0V��:V$��ô5K��\)�э�j�zW�n�u`�"�.�����F�9;���k�!��<5(�N#hA���a�]zN���.�����h��R&$(?!��%P�%蹲ER�����e��<ÝOW��$������OԝC��e�]��赐Wa�掋*Bm�;��^}]}�r ]�E.����a�dO����J�F��d�m�z�f �IL*<����Iw�V>$�|Ma�f�y��$x�����
�x�?��8.V������O�⥚{ʙ�J?+��rRAHxUG��T`.��8���@���2�]��'������G,l����8����2zFA��!6$vI2◴�˚��%�V�߅�#���ђ�����ސ͖�+6��/�'K�ڮ��]�=��6����_��~�֎�w~����^�:i�u�t�r�us3�d�οx	�kN����i�V���87$=��2���4?M;�#w��a晩8i���V��k{�B�$�V |G�B/&�Cݝ֊ۂ׼[ď���<���;5E��1��F�#X�V�p��x�n��� �U0"�G1�IUbi�f�;B�*j��G��4�'1l8y�G���'3��ݻw��<�K�/���Rݲ@_�ƪ�)1=��>ܕ�~�՝f��R�ؒa�|f/�T�n�����{�嘌�p�O�M��]:������ˍh�|t@��e��]^��V\�JX�Ekjj4�a�?@���VC$8�I����x�o\.����D�^F3��6~����T����g����*�Ż�����;[��?��b=�;H��$�R�:�}�9|BK��d:��]>������_��E�~��O}r6��k���<����IpIu������%f��\	��oPƜ=abbAӤ����O}2U4��yz UT�Pmbb"T���v�4�o�pg��N���躋S
�/�����ܼ�PZ��JU�|�r�Nm[��,�]��PWVi�OgL&_�|�Q
�����������H�}b�uf%`�\61��0ҍ�^a"WFig���[g�!��(�~(�d��&�š<'��������qa2J��g:�m9ض�^���`�-Z� nf'D�c{ �m�:4k���K���?�2[��{a���bǝm%�3�'�n<����w6v#H��SR���# ��7$��l�-,
�Di�e�+�(��O�U8qV�F��t�N�?߮������IB��Mw����n1�e���;O7 �7��c!:c�5@�1�j;,�WdU���������l�ա�O/X��<����_jQ�&ܼ���]�5o�ΡU-�p��Ga�t�_����Om8mk����?:l�Z�2��=]6�^@o�^@�>}�W�9	�����Xא7�'~?iVK++W���\eR3x�P��ZM��_��鎎��:�2�|q�Lr/���1߅�ڻp�)eca.V��Ю�i�r&lK����%�V��hn^���7hƣ}3"���槆Ym �����M��Y�9��i��#V�(~;XgL�ac��z��ȏ��9%�A�D�PQIccaf��6��0H`B�q� ����Ʀc'Ow����>p���I+��K2�ESOf$��.;,�iI�U�X���i�T�w��f�"�v��Hn��|�h�t��q��[(+�a�ڙ�b��W���}�&�T���@�������������C+ ���F���3� �B��g��\��l4�i�M��f���=��Xd��7��GpV���y��+�>�iy�9~�Ԟ��j�A����f�_))�o�u���!���Pjd�l��~U�Y��"jH�9Z��_ �8��<�v�!���\ΠV"	�İ�M4�]�M��BY�S:��0� $g�6�j�u�V+ss_'����y#���!p��܏�L321���rd�{�@ �=[AS�pp�A���ґ�MIqފ�F #�tJ��`ك��a�R*E����u�Te�G��Ə1��z�h4(�jy���g��g;qT�԰9�Qgce�0�[D�(bg#�G�T3��С=�Nܣ}��TC_a�`lC����u���@u�WP�b��3:��ED�_7��h��f �m�cP�R4�BZ�� �:^�8�1ɾ����~��9t-����S⇮Δ YK��VH'���wyGrZx{UNM�b�+�B8fL��;2?-�	J'�LT��Ha
C��Z�Z��d��� '@5w2�6�yTD%2�?70�\�f1JYY9�O��C1��4�wQ�lG�H2�n��4��zD2c�(��&�%E�XVie����h3%�����D��_�A��0�!T����C%���bK�AE�yA�f���MK޳w�0���	�D�s�4𾱮�H��
�6�%to419�5_l�u����6߿'tw"���3�[������0��$4y�U??{���|���p�@�[r��]��f�|��ڋ(��o]�u_����op��Ц����O5.x!�sP���wJ��N��L�cqfm2�=��=�6��Qs�1��03��_	��=�;��7�RH$�<��a�Z���ha��%����x~\��I����<`�;�����.Z�P�������oA���f�ji�A9�0�(��������S�>�a#�_l;�bp�����y̷ 5�ɩ/�d����P�����	;5�::߹�dnj���2��[���Vy��m�)A��Z=��/Al"�v�����MIy�����6�K��T
b,s�_w�ƙ��NV��B1C1�p��y����8q<K��8������y{߾�!H3�bC�c�Q�$��Oh��zz��Њ�|+^|(�h�M.i0?��
	��'�9�E�<���C�^D.vJ���Y��0nP$��D�g׻1#z�����f'��=���6��޽{�;_Rem��K�#�EE999�'�Kv =O�����#?]5�$�I�3���}�Z��-x�|�>��ٌ�f�Bu�f����˚��K6��&<L\�8���Ї>��nX�E����4-�>�~
������O��b��7~|�;UT�%0Cߟ$��x7wA%Ǹ���?���6��ט��H)�,-���]�o��w�PMA��4��\I�	G�y����t�R	� H2�)��� L &��.���u�q/�-YPu�0�@�t�K�����8?���-�PuQ@�J���mQ�n��`�b�Gq�*+Amy@&� T����c�X���ž\cݲ�q+��|AwPtn1��p_��&��,��Ү�
2���=��].46�g����Dϗ?�Z�)F��斖����>3�f#�+�dq���jR;gS�d���C�˺L��!&��M��Aϣ�-��P�˚ 1�&�-�G�+R��#��x�A
��@�	���/qJ$�4p��4��t���X/�@` �"�P>1ߟ�V�M��)D��g"̰z@򎘝o*§ �Ow�2�.����
bs����G���E]��Nl#p2���ҩw���i:}�|i�����Mz<5�D3�D�f�5����֞^�ꆗx�WT��P��N�������y�n�o�Gנd�[f�t��$T�Lw����ù6�A?l��R�*��*	�P�ܺ�?2k�K���m�JM]�RUi��}T	=l(Ů�p��EU�RyB��Jq���C��9^��8��l��&&���)����0r�hN�<������6}��P�7�����<�\w� �0�.B��`���cN��<i��Y�9z���_����n�g .��(#�8i��@��b`bSQV�hZ�����/���gB゙!��6J��'[�����%c��V_���� ��G^��PV� Y�L�a�0*�oo�8(
���K+����ʝY����\��G+��{-��[����>�_8�yY���Y�*b�:��N#;pT+,�ϲ�\+Г�D�w�s����aF<3b
J�aLUq�@7Z����r��T���L]��4*���@�7^֚,'�F�yGA�P�#�
{�bw�������4���O������1o88�&丮�&A[���������e9�E)����T�
����?�r�vg���X���c��82���>QCbs}�R�tf�F�����C6[�Cۋ!쬥yT�H��߅��z7�`cf6�E�=�����I�i�\�`=�9�>�0� �!�� e�O�ʺ-)N\wU	�3-�=��i�~G�����wԻ��Hw����|�X\�M믇��- �5{�x@�hF��"K2�A���|���\o�WA�!=m�G�u0&�v�>u�y�i�!k�60����m��,CH2N�]V�L�v�@�3�i��z��!��Zd��;���E���֡{�W��-�NܩZ�Sya�h��1=�V��EKu�glҼJ뱠hq2W2��Ӧ&����W<D�+�ɫ���/�_­��%B�'����I�'AQ�n?KI�����ܧ�ín��i��j�ÿ@�!��T��?dNY��r�
�g*GEE��B���PRe��ސ��؎�
3�OU��Bg�ʍQ�+�X�`�*c���VLM��}8Ӵ�� �z��mЇJ�03.?r�j�ҾL�8ٚ��Ǿ�ZQA���3�9&&в�� ����%O�|�_I���i"��v>w��a�έ��Z+��ǉr
4�k�,�ا�����|�����I�����N���בMA�ѮI))�'N(1=���0���l�x@T�\	���~2�1�Q���;{����jq��$��\�HJJ��V��pǅԈ��4���:n���$St� ��$�^��q��K���d��`R���i��{���,�� FP��V
b���k�fl��*AqU�G�:՗c���*�q��倿�"���e#�(3$y4���?N��U�6����%�P�������d7��O��)�����)$� ���Rj��q-A*qW���ʖ���&���2����?JQ;K����n\�n�|.~F��5H3��x�j�a�y�L 7?^�[(�;�T��lZ}���	��AO���st��J>EpJ��I���@�2�	�w}��w���[�C��/"��ʗ������t�ɕ�f���H�'=���d�N������/��kOw��%rRRFD�:��B�\��K��h��zʺbΘL�h>�Ŧ_�=QR���#������@�2�ß�N�}�Lw�H��%���hЛb��P�=ᙷ�u叐Aȋ#����;��))~�Z�GosW��ĺ̝���	r���y����Dy�?�+��⬜�� נ�%��̾_�✍̣�!p#O�^�� �I�h=�%vwӥ�X���G�� �� �EML�ʰ�\����IJ
̛��%�5s��t���uQ4�i'��Ȟ$ٙ�����0֙��	�k��FyP��L>���h�_(j1�l���=�9���祑�V�5�<�>}
,B}�^�Z���u�K8ͶFh\�OF����U/�?��%�0������z�T������_P#�P#b{�F���n�:�,�|̄�KҾE�GJ��ZU�yȭ۴y� xL�9��.v��X�Ƈ��wϞO��M��ԅpi����*+k8P���q���j43-��;����� g��c7�[�`��aE&��]�mztz>$6i�b��L#�����Z�~}d��G����Ld�?ۄ'&݆����2��7�`�����F�c.~��:�>����TVv�x�����L��E0���U�q�U�8��*A�p(ά�b��"�hf���BSS$H�����,	
&��7�r����^��Vf����!�}u@��w�4��nˁ��c��u�SRZt�{�<��]�M�tm���!HS��a�'����>!��=%x�~�p�^3�=�@�U4U��u�h�wz�68�dvD���
:r�-�}� ��M��\������*2�Ȅ����*ϩs������璸Wg̣�ՙ�l=(��l�+bne����A�KI����n[��qJ�d <��T []���5��!FC���NW�SG�Z`���VP���L��j߽��E-�=��F�ԩ������;	��,ͦ�_�j�wpp�E�������y�<�l��Q���n�D���Q|�á���G�2�����U���������L)ȋaDD��b砍��T!�		yS<�y9�h���~��H��~��]��Z�B���k���������PQ�L<��ј�tO@8Y�����*m-9Ş��lZ+���y�!2�gW���-��W�rjbe�[e��~V�7������v&w�z�����u�5={�c^3z�p������SȤ�i��Wc��@�0�E�ľt�����@�/@'�4�?rT�T�����M��ږ��w,�X�QAX�/*̰}�7��7���*�����4G[D�AЅScZJJ����W�(�E>Q�7X���X#[pټ�͎Re�k'�wz0�R�����GẄ́��xeaL�4ڌ����o��S�E��ߵ�f4l�Y�a���K$ɷ�܄)���W���t�ڶٻ
�y.�VljCdP���^:��z��������Y���-<rE�$����]�*!�G�/.��L�@ؓ�ϚH{�����[��ų�E��-E)��}(���혪���ﬥ�K��&����2΁�h�x�g��������叄���xJ`�V��~(�C�51�*�k�wZ����?��49Ȣ�v�0C�3o��F&S`����p����|_����P"YU�<M�y��)W��d+�!PTT4X�U&�8�`F��"lq��YN���t'���+ٗ0���4��r�k#�&ݿ���~��)�%F�����f�����2ݽ��_�!l��2zKZ5(>L\�t'A*Fy3iy�Ϣv�o�_W�&L%�Q�SS>��	�Ջ�;�<44T���ޡ?nbRJ��mN�G����"�/Й�0�;q'd
�3p�?X�5)�}ъ f�n���n0��?�8��`��i|ѭ2�U�i)�&CWQu�����p�
�IT q�������ZN(�q�u�P��~(ï�B�%
��L�	#� ��OC��|���J�',$���w��,�p!?�V9���v�-B��d�3&^g���<P:e�;m=F2&�~���3)+�Le��A�liav�{����	4ii���hZ�2Vx�S�c{��ܢ�E���Z���+D,���ՠ����dr�n��C��Sɱ���h�[9��h�M&+��~=���X*N�1i��)_�Z@[z����/q�Q�h���2�[%)r�c��'�X�����A�� �3x��`H=�U�
c��/�����DJ��߈�?w�}9�����.���M�w��H���8m��r1�T%8��)Ƈ52=�s�1@	pwa���K����#���+m9-�������F�Ӷ���E��Ϫ�a+��(�R8f011!�9d�F�V�re�0��+��3q���ae��yn���k�Ѯnr;���M��nǝ�*;�������U�K״X���lM��f�=i��m���Y�x�V�3�zO�驞[[��~��l���/��y��Ϗ�,��O,�\z?�·�X���Z�6߁��:p��������D՘�ªtč[il��ol���~�ܟ缼r�W��Z�D�V����2 H����a���(M��fd!�@Е7�����mZ���0{-���I���P��k!��/k�MfTB��wB"Í��8FUEق������sʉ�5��Bp�֋����7�d2�#�(��#o{�+oo�9�q;�+����(�0u�f�-��q��{��)���}�S�5Vs�3>>>/�������y�ɪ���m�/� u:O� �B�SRX'�s[�x���MK��ah3NU��٘���<�D�*�
{�h,������C\4v������ـ:�5֚c�F���Nb�����T��SZ�.!~��8�x�>���*��ft���E��+�}OV=��ý�J��b�.z�Æt�pP�|_�j�7�*�,��=��3��_o�N�ѝ=9�?��7{-&����S:|���T7)@���J:������N�i&c���7�pDW�������,���!A}Q�{�(j/��$�py{ ��k�E--�լ�j-y�������?�P��R�����E���xˣ7���3 �z�ߵ�}��ֶ�H��&����Z�����b~�f��3L�z���_���I��v`���ev@�?���Z��ޢ��F�~$�ή����s9@[�/����%A�Ci��Bt�|�bY���|b_շ��k�G�B�rQH���zS(����p��@�ǅF�*���`�x-d�"���ׇ�Ќڱp���`]ʁ�Z[y�U�0jJ7���59̌+Q��2�R�u=��u��_�+����֣��t�,d��D�|�_��b������Ǣ����%���K�����J�9�)$�q�>�_�oE�
f�����\�n�ղ1���ӓ�²�(���q�&&*Z��/����0y���B;�s� ��6B���A���c*���L���~�l�q�G\��f��q��������/���Oaw{.I�	��,�'g/LF�5=������8�q�a��+\�I��Zk�;�s��]���-���P\"��Qo�w���~4������틵�O�*��lh@(P�z��6��#ե��Ԕ�տ�I�D5�ӥ~�z5l�#�PY��j�O��wT~x(�G2�ɫ����}4��U��_^�bd5Qzٖ�U?�����A�-'��UlI�g�vO2�{����������0_q|��{���-�㣱��#'p����ɔk�~��`��jq��掎����#8���d|�B��w௛[EE;���V�i�d�e��-D �M_�B��G����_�����7'����GB�v�vrr�O���.Y�>�Q.���p��f~�ZVQ�{v������ċ!8�2��Nz���?'� �QU}ff�-�}{�' ZM�A���73/hfUw�Y찆Y�I�60R�&���(%���Z�XP7x��������o./\���,����a��B�u�Ӡ:�U�bly����0�����,�О�k��?%�` �o�6�P����g�0��r����a0⏡3C�I����I�t�z�������{o�M<���TT�>��+/���0�)Q(d����_�En}���8Ѷ�[e�?�����Sأ�%����0+K���|J�F'�Z YJ�P�9�))�������Cӓ���k��s��b�"�M��Ԓ�_��1�&�� U�H5{�
����#!o��U}�Kh+���R[M@��H���*n��X�q5�'���#Խ>4uB_P�G4Ss����9�u���N�N-Q�ج�Nu@��é�&Z�V�T5��P��+qCb� =S[�O{j����"���g�>D?J	�M��K->ר*�Э%�58���a@n9I��$K ����������\���]} ��L�g �p��,���&RQ��g%%�Ra�ҷhΫ�=���w���$t+�c_�d�5��ؔ�A����w$װ?)CIŁ��Z�K�+�m�PƗ<���_B{�07����#���7�?zN��f�i��Ȕ� %BF��1ȄE������_����a*��I�r
�|�Σ7�� [%(�aά`�T�*h��g�i�u�z@�R���JZ��W�e]�X~s�8N_���IDu����.���pJ?����ց�ǐ/�QpR��R���TU��<�Њ��G�%q�`yK����ϖ4�JAG�2��c�2���l�Ԕ�����ZW/�z���$�u ��2B`A]�G���?��wQ{fU8��mڵL-��?��ي�_@�"N��"�8;;{\���-�S�)��{-��5��y?� M)U����V����T��˨A��!d�i^��Pl�6��U��a���u���p���fe}̣�g����A��(w v$Ju�V��gV����A����>��ְE��>i<wU!�<5e�~�
����_M�):���AT��4>���Q4���8v�$W?F{9$�����s^K㪒X�":�x2a�S+�&����Ƥ9�y�Z
�0�{����*�Z��A�bW�0
��+y���[�t����7�:�!֘ś���O� "��e�1<�dT����J�s�KH�h�[EJ�V�����9 q�����b5ͬ^I*��t#(��Mmk�=m�ZUT����}C���� ��i��⎆�BW��.���ii�@n _D�:�)).4�՜Q��KJJ��η��(B� (�ܙ�_ ��e���M�H����/�ُ�#Y���|e�֧Ub��0�xb��dǎ{��V|�P*#�u��/�o.�TJ� �q^Cj�Jk�j��G5X-<�D`�7�`1kQ���.��z�ԺES_�Z���l���|I��(d��Vq�� t� ?	I �KVUk��[�5�j
#����w�#��������v��0�}u�s�W�EE@a� �s�2��ϲ��U/��@<CoU(=��İU�w�fb�	�(�-�q�Iˤ�v�/��IP�������^/�
%������ͺ��d��yn��Ⲣ���_@)?��[���X�]o�d�,W	�뻅�����H~O�� ��ټ�K�w�Q����:�:���Š�������&o��s�Ϲ�B'�I��Y�N�B.�TWU+��A��˹�7iޫM���1�bU��.�*��P�Ƞ��Q�+��`d���wD��u{X�6//�@�\�3_h��	���3k�Jͭ���BFW^񃧚a$��-�~Ammmŉr��w���D���W��&h��
���928U��wp�i��-���U ��w��5��QUN  ����|�aD�����V��{��?qf�Ui��ԯ?� A�����sI����g�:�{oV�����
q8�qR�Q"E�ѱ���th�T�4���&�aK4��ٕ� �L#'M��JE4����������{]����k_��:g=k=���_�}���+'�(b6�|���O�>2 ��܎��$���1��ʪ{�g�= &�CE�yB��'�a0hD1@1pܶ(6m�����L�� �0���h�/?�P�5�����K�,�f0�<���Ŵ��)����|�\P ��C�lon}K;�������1;�lY1�����>@K�#�M���#{����[+��#ߗXURQ�9��P�z�t�mU^����]$�'�YaPE̩�[jY�ux5�3��T��KP�5��׾󖑒G�KBɭ6��y��G��^����"�3�++�y ��0T1Ӧ�TB�u�wi��g����0��}�.%��`������� /=z�#�����=�v
�"�;�~9/�����(�D�Uw��)�T�ca���3B�I{+���e&��^��a�1����:qT�4��عs�2��D1�n�{h��(�Լ�����`�W&Cx&�CKQO�MU^"�zr�G����`4����˗�C|v���*���ދ~���}	=�����JH�ܺ�	�,<�m~#}���.��RrJ`ͬ<ɖ�4N���	�{���y��ȓ�3ؗ�:��?-�4���{�� ��cI<��fx�k+B��޻���O��F�]dXX�4�U݅#z��{ |��H'5� ��Qm�P)���c؜�t������W��_�tT�Ks(eon.��QN����}�W�.��><h�N�"� ��Ĭ��-��s��M[���@�* N=}���a^r����/�Mp-��k6�}?�:N��@��Ym��^ܴ������8����	bP�zx��1�wU}<wv��F;��CrT>g�n�҇�+���M��*f޻����Q�V3��)U�@CQ�`��ޠ��<�W7��x�.&��A���~�\�G�D����I-}� �zK�r�2%uV@_�QN
��������Yț�g9Y1�ƶ8
[�Y����ԋiD S��Vy���[t;v~�X��,��2Ej�{zv�p�,M50,kU��T���l�[\�3)@��_�H�v��q�������&��8{JQڰ{�_/�Z18���`�-h,�ߓ���9C��4e���G�(h�:5g�5��'4,��MI}���TgH��&A|V 7< 7th)6!��T�O]U5WIO��	8k������9����Si���,?{�st˛�I��
j��5F��������~TE}B�*�-��������F�O_@��RXcu���}�b(J��3�:�����=y��Uq��w�9�\�t,N%�]��N�f����T�f�1<U�&t��=>Ҹ��ջ�egM��:�u��T����5`�o�$dس����D�3fY��:�&0��a>X�L������ς�v8�'0	��W�Yn��wf�������],
�.�*/m��Y��h��s!��(8���F���#{�{��=�m3���O��7�bO_+�ڱ��&߀���/��W�F��51�o�����g�����%x�K�����/���bjyM������z菙��E�V�n��-�GZ�߬-݌~�p�]b�.D� ����n�ʻ��P3�t�����K�w�`�c, ��"� L��y�4N����~w���P���ϱ������b����߇`~��z��	�^6DSL�4׽�ҷ�����(���8�� ��X21\*�����`k)hF4�M4Lu����+��_��9jr� �Kw�n�J�I$
�xz?�H��]�t��I�(t^���Y�Ϙ�i�-�n���G�����79_oQ�o����e�В
�/ߺ�����?�+NA��&�#Tr,�O��Z�>�%��vȨ;�߽a9�x-�Z�e���V�C��F��H�V��-�'���ܖ����ؔR`Z%�����s�9�X��߬p��G΃\�g�߰h���`�=��E����G{D�##��u ��?�0�A���ܦѪ0X��\����%���	X�ϲ����zzz�k�~`�^�	��ca������Έ!���Qg��P�J���� (���08�{3��<f�^l�5��fØly�4Gm�JMG`.l�����*]�Cq�e�:�
Ϫ��"0{%W77.���!��gS���C����p�C��;t�>�$�o�j�TeH��Q����������~7�.��J�Ah��Z�>n^^�{gSb�B����uu�6�� �ԟ �@�wi�
�KN0���A@�B��1��L9���0ם k��cx��z�Xhh�q�ë�r
�H'E-�r��B�>���)��ǈD�&��eľIuG�V�ty��Xa�Sgbr�443�=�maO�Jc����6 q�G�4z�T�'-Z�z�2�=o\�u�leS�7�]%W���+����<ک��wPʲ%�ݓ�ij!o�)��X~#>TVA*g��c�P3ѼӶJ�K<T#kƌq���S)�����8�X�\���%T����Ӑ5�ʔf*U��X�� 6(�������4h�l�a���@�(p�ʻ��?��J���+��)�(����>[�uO�={�&)>�@�p<�>�Y�Nڄ�es��ra��k�y=b)�T����6N�C��I�y����#�~V�f@w�mZ��֖�x����яOT��{KL�ZEá>���@�1�3 qZ�Tʰ��W#�ӂ�A1�Z�Q�rr�;档7[^��D����j�
�F��)���222`�5�v~��'����=MBU74$ӛ>a��D<-�������t�2;iZ	�� Q_�n��&d��.�x���ߢ���L	�e W���V�pȷ9e�bp�.�Ź�n�Cb��z2�Umj8�P�&sI��%WgK�Te/R�_xڌ96퍂s��{�l�����\��J(�����s[��U��u�dA� �E��ʅLIoS��zu���1�okjjjk	;e@V�u�aG��#�������Z�1%�{�9�<��,:A��4U�@�{tX�~o��{�e��
��|j$�[/+�#w\O�i�\�C�k;�����+�t��~ݭ5��kw����@��vS�e~�V=��^�z�ǂDY�vJ��F��×F:~IZ-Z�gQZV��fJ�J���[E�N�z����b��kJ�����~[̾/�`5�q�7�z,HLjt"�'t6LO��m��$�]/;� .��
>g@��?m�*uX�|Z�D�������@N��[�QՕ�ȹ�/�pa\G��_��a�o�{����ׁ+�ˎ���H�.j R���їPVr�޶R�����	��	uGn���|��8�����<�%��k���>��S�	Ҽ��@�8�.���Q�э;���k�GB�T޽�А��u���gb',�������n4e��:ڛ��4��?�JZ+�}.44T;݇ؿ���bb�/O��Z�=��x|ݑ�,ORLU�G��tm�Uo�}��V�ז��^S�G���}�"��Si�ND���:�����a��S��:���F@�:�e뵙wL�077o������:�ݮ4mB��y_=�}�h)U��%	��4~���g�V��UY���W0l�T�����Dxk�����q���)
�w@azxA�5��C��~,g�G7��en�'�p�Όm?�������L��֫���r�����}�}��t��� �u��Ei�f��ɧn,�?��A�+���-H�q��sMwR��q�º^ i��d�B (��ը����ő��?�'Ц�2~�#����ӧO�J�Ę��C�����e'��� �[��a�� �]&��
xb�AP߫=�ȫR���!(����;wС���+� �U��В�h�E���S����d؛���<[��0��S)+5��2�������e��Wև#��2�#L�N�K�*y��D6Jz�y��
]�2��l����ë�����ɜ���y�����{6���4�"������ �C-�_߷����D�eM8���ޒO)�c�^o� ~ў5U�A������s2po4�<4_M]�k/6�kX�)��F�_?���������⢯��Ǳ�a]�{H+Un�BǃWT���5�|+���ePpN�J��'��v��!�Q�4*�lV2>pYs!lg|�b�Q�k1��:E��*�btz��q�����A��81��O�����3�E���YI� U��n���^��� ��VSN�p�>2�^�}�1�fs�����K��0M5g��H�.gM^S��|Tq������y��t�O>5��06�͸'��)T>�����W�F��V�'!�(�ׁ?q����$3�M�7޹³��j����|;��{ 6!�9��T�gJ��h�4i5_�1~8c��/�1/�]�,��!o=&��=�ϑ���z����jd)adT�;x�Rpi�۷{�jI����3�3f����o�?Ĕ�D������[�#WCZ��v���&/�}��Р)(�lƗ�V:�t)k���a�obX���'/�^�&��f��῝T��WF�i��-pf���o�=��bRF�Q�o+@ҽ���Ӕq�9��+�
��%�������_hC3(b�tᆇ�#��ݻI!�	u�z��D�@C�m=�@=�d�/�gq�P	6�\"����O�����&���l�-����Oŏ%�gp,KӨ�g=\>	�������������<9h��8.*�A�&�34���Dv��JJ�}\p�\H(�
�2�(_A�@�W$Ւ��UeQ���`/��T��8����ax1��MhR/�M���d��!Wd_�|�r-P�
�li#��ͦ� ����%���+�rG�z���R��eÔ4us�K��U��m�}x���jvs�i�"����
l�Q|��ZU X�(-P�*����&���$pX۝J9���������������;	ԭ��.��lXX�6��ʉu,E�h_찵�y��z}�	��d:4�����G���A��!4�̫6f|Hg%C4�^Y$�z-G!DN��c����t9?c���yc}|�L����/��lA� � �ڷ�U�~mˆgr�7���=�.��я#/�����\}l�� Ȇ�4�Ч��m����ZE:��k�7k����sȶ)uN،���8o��K�,��W�~3��z�"Aj�y��8�)��U��N�����W�����O�U�W^�U��;V�G'C�����G¿�����?�щz�sXj5���R/����1��:H�����X����tm�o���˷�a�#3�S�W�����r��qSir��+V��{�X=���{w��|�+2�\�����P��c�M�C
����:hq�`�碯b.:W!^���8�O� %f�"�p �.�����$&��{������D�W�ml�Zd����֓�cg��f�������~^}�|����_�2Y�<Z��ƮO�����WQ���ͱt��Q���� ;���M�g��y]�;۱� Q;�]=�/P�8x����Y�vƀ*�.�ˀI:Ua��̦b@;�fk?�����V���Y�$���Pg��At����.q]�-�-
�	v+y��(O�����
8���JRz�.�Q�qh-"����EEM�d�I�`gC�ӡof����1RZο��D�NUG�{���Q�9�c��Jo*���!Ƙz��!S=F����ULaTi�]̸�Hn�}�*�?���dy�u�?��G豏{W���t�ܭ��~��&M�ry��P�������b��l�
��|�N�D�>/P���%G���j����4��h��aGΦ��=ik��/��#����b���p�C����}5��'Z�PWGB6��Pd��	[/�U�<�[�Ro*b���N��`Y$�eS��$�������v�&�ź���E�8�(Jj?Rv�(̭��R)#R%��C w�z�Q�c:�G^ڴ��4���`A����h���T�)�ވ�w�K3e��Ts*A�N�E���'���p�K�8�����l��8w���w,pC�q>v �֜)Y��E�H-L\���+RO��؏�.'���#���cXVS�c��0��w�v�+�!����eg(P^� Z�I��,h^I6qD�<x��H��@���·���� ��n���;M�U��>9#�@�oZV�`���Aϟ���G��qF&ٱ���v�]JI����Õ,�򶟇���Q#z<<�k��RT��k�؉˾�e�F�L�Ìv��4QD��A�\C��g��1�te Lۄ��__��X�������\Q8K�{G�?��t0:M���k ���s1}V�Ӡ��0}*�-� ���XЬP$踤c֮��0A=�Z�$4��p�a9��j0Iq*s'�*�6�#�Sn�j {6���a�n�`����Rc!��������.c�h�F7c8���Qi�b������L)Wu�N�<�>�T�E�&�YA���06�@�	�H�U&M�OOs&�`��3*�ѕ^@��E�4��<\��D6�':�Klz�FL��P>OA�>	+�=�+F�$���p*��%��q l;&,v�	X��LrB�/�S����I�`��`c4�!M�x�C������}�tKL�2�ś�����"O�K 7�e�,��#*�=g�Q>�Ng/���IH"4c�߽�N�����TAZ���$Ӑ��!���UNW~{�
/j��t3`�q���6i�`j�D:Mx_Vtr�t�Bʌ/�~%%����E�qR!*���D�����XD>V&TO��=2���#����-�
��>�x�xL5PK2�W--�%�(�w3��}����~���,%��4@�Bh<ɑ��*�63jleAO����D�q3^Y�;�K��P������;_�W����AM�>���(,x��X4t]���	�]�GQ�ӝdWA1�F��xC�`ޜ�X�k ���_�,��jH��@@��b��w'��S�*��;#��;拓��,x��X��z����ͯ�yw0�:�����ɔ�ג�d��Q}7Z�۞���W�)X�ryĿ�k�5w��VN��-��>�� �.�B��7&�7'{�;e�>��ZA>�A�e��U�{��3� ��N<������D����=�B��L��.n���ʔt�Leq�W��Y��-s�X���K%0���B�~y[��}�=���={Ǹߧ*��;D���8��:�!3s!��a�~d�����μ���3���4a��V%gS��W}"�Xz��3Ċ��SicxY�7?���b���!�قXs��H:��}���}��<�>�7^�emN�A��Q=�Z�m��
��Q��=sӖ����@�Zx�q�	Q����.��<�������/-RD*�݋~��_#���7���b7�t�
����;|w�
Sr��٥k9�}�!��fB)�Z��p�u࢏�{�'25�p>��Lh��A�E1���s�\q���1�ӳWeP�d@n7�4iźE��h�U6bn<����� �C�_N�84'�E��;� �OL�t@����g�9��VnD�g����1����t�C^�^��?��OuO� ��ga*(	�8����v�i�Û�
��Uu��K�s�����MI�����^�M��+���R�,dNīWS�������P��8�58p�O���l����L"����K~�V�z%�VT�ρ�U���F�_E�Z�.쉈��|$��1٥k=���,��Pr6ot8�fR�\br�ө���c�C .�7^��Ÿ�cN>����J<��?��.�It��f4�'f� 7�8�$5�86��;n@��fmpQ��{=_�������n�(��*h�టő؊���?�w�J�1S���D%�4nޓL7�*��mY	Bg�S���$��=���{nj��?ò�"q
5	w@l�Q��-[�*T�DLcH�v������I���	�h�fg��`�>Y6����ۨ�x���c�81�?��u�(�T�����}Ζ��՚�Ȇ3�πJ���=K!
��?�b�l?x���ճ�*��I[�xӨ4��e�A��*'׳�)�x]h;I�Ɵ�g�vy���+O��N��VW$��i؄�y����=��> 0u�J���.��A�z�EXlq��Ԁ�bb̵�i�bl+����r�!�U����O�8U:�w��OÁ*d������� ��+F�G�?�D�s�
͊Z�z�dK��ȡ|"�����*4ɧ�V|P*`����3*���Ah �����Aj�F[��(� 0�zfAU��m�DU}s�S����B�����|G�{;7و���E��g)RUMH,m6�oH|2+� r�������A�[ݒ�4*�1���Y��'�zE�c�ޡ2���6u�QٚL7a�Gn�$<������~��ДMG�?�^���5|��<*�u��� s*��!��R�@�W���
��? �y(h��9��":N��4S�R�"�|�y�5�����v�6�y�]�� 	'�gT�-k�%�H�Z�M;���TBK��݆+����~��p�dC�L�x�yd����u���F5s�p y��N�v`[�R|u�^r*�����
�
5Z�#��:v���7�p����D��� �<�?�Ia���V�6�@��+&��`�pc�ƴM.]2S5!S���ֲ�Re��I<9~P��"��1�R�w�J�	L&�v�z�0�r�ߣ��3���9�m�8�I{CAl ��t5��v�����D�	�:D!�ճ�?��w��0�q�EG{U�6kO`N�Qw|X0�c8g	忭�Q�܆)���>����G����g��\�N�Oۃh���s|�@�]�y#¤�1��?⭌c5i��^%�y��w��ã�'�=�{��s�\��̈́�ß���A�\��B_���#Br�`��|�a"s�U^����`�9�ZB�B�S�H!���}j
t*��Js���S �.gEW��"�
��n��h�����5&0�r3 ��U�Od�v�n7Ű�O�^^�+[Nқ�Z�*zݓ�ڏĠ[�6�*��H0�΅��]͸Y1M4��2�5�(B�S�<&�Ok�p-���У��Li,:Vi�I@x�	�c�5(:��xtS�D�Ux7�(��@4 PȨagVk��?��1�~��%��d�����TӉm�?�0�J���~���wa-�8K]�-�
���x����ܣI��}�TY�eI�](��<{"#'�l.uwK��I�@|�\�.af�-4��C�8T��>�IG*K��fI��CxK�j�n�Aj]�?&�6�b�f��4���>|����N�7��d5c���T�wnVP�.���0�r��I]gt�c!	�q�N�~LtL�l�����H/f�XbR��]�Ȕ�`���t|	#	ӛ�^��7Kt�/׭�P >�k���-�]7D�?�M��i�L�:�5
�kEi�h�1 ���/�x~���#7��z/����<�H�kD���^����Ɗ��q�lo�!O��lap`�"��i^��MB��3:ɶLj���LA�ʟ7=��t���eN�;Н^1�	 ����{oy�
�gB�ʶ1��.\j3tk���~�3Ҷ��6HtbW��i�넅�ؖ�D�ZnE��.�ע��#����^|LxD=t<5	Nw�)D�#�H�}K��Ge�p�� �9����o��푉��Z����u^,�p����� ۼ�W���D��Ut[X�
d��FQ|]����)`x�Z�]���W��v��&E��et�����Ҟ���e�tY��]�u��9HTz z�ʫO����Q���M�o�f���s(��'��&�
 �u�ɛ����+G<,MV�e`���c��iaw%c>{X,}��%ů	ܝ�'w�-D����q�,o|q ��u�X�'�x��n�sJ��>_
}�n;"��O��K���m�z�n������,Q�5��OH��:{{{a�����fO!�PWAC͚�ر-�҇L�?a>�C3L��VVRF$6~�&����T��M���-4""BhB�\C<4�����x�C��D�5�GX���	0?��b�`1"�Y�;x�XB慢T�QR�
"�	30^*aD�x���	�(�
����,A�z�P2��R�Tey�����:�ў�t3n��H��L������b:����²a������#���#��c3�Vm+�.�ygUƩ%D��MI1�k#����� !�("��|�)S,4ޫ�AN�v!�{�t#k��װֳ�8����3�U�nD.��kz��0�朧�/�m�T$Rz�,�&Ye`��bx �:aÏ��?!Yn;|�R�0��y��-)4�,t�y���P2;�`�GM�(@�|���t8CQpW�x�\yV4$��D�#�Lÿ3��]������I6�{ў��r���Y�<���Swk���)�r��Y�AWHę���G�otP����&�����/Trfi<Y //�?�E3�txE�Q�v�¦��d������fF�u��U]�������&�ֹp�cݡ����I�/xpp���=}j�u�ⶤQӢS ���1�`�$�p�6�Y�s���;λ*ԅY���3��s�#���6���\:�����@�!g6��D<��+k�w1梌J|6� e��6�l����U#}�J���'C��9ɝ��Od�b�[���p�'r,J"�'P��1�;b�UPc�l���5c�d�&sn
�r�էu��ߐ�3�V!��%X_۟`H��"�*p���|���U�4�ү_�l��u��og�y�&�S��q���,	�d�-��lr��}�@pˊ��z��Z�B}����=O��n�|ɑ�##��oE�D_��x6{��A�q��]�r�W�_A,"��y����D�Z$U�����2c:2c�eM{��&��*��VF�r��� w�t6_}S��eM�y�'��	7�L䏬L{Q�̇�n²��w.i��_�e�L�a�,���$
��`�����E�&!���߶�?s�o��ٴ����3�D��ӚT�6���q�/�$��NPFEؼ pg)���
78���K�����c0���(�Jߡ����T]ڧx0�ݪ"�W�j]MCW�(�-C�;ɮ5=�`l"��;lpg�ֈB���O�P��
	o5�gA+N\�y&�TZ/��yiฮ�E��@�b��0��*FᏧ�sf�LCL��S�8��&x��
Kǉ������e@��96jo��JK	V<3��f|��`ϭ��=�=�mB�>�������>�1G�o�M�Sl�$��Vļ׌
8*pT��Q��G�
8*pT��Q��G�
��&�A���!�?2u2v�[#�.@�9��a0����
�r[V�gնN"vۥT�Ƨk�����숬�I<�k��V	»I�U}<4�%���Ph4����3���a���'�3��:�1��m�Ɖ�*)��ya�n벣��cA���F�_9R>o��O:a��fN3���#8*pT��Q��G�
��M�u7����u�ʨ�8�tj��gi��5�C�'��bS�j�B��t�]�'#4�2��kF�
8*pT��Q���/�;VI��'N��;�r\���6pa(���}���/���{_���ˆ_&ұk�r����I϶Wyy�*��V����'-]�b��fuE�~�qT��Q��G�
8*�������N������3}K���u�Wy������d�E�:\�
�^�Ou�<���,h���sg�>��8>B���c|0*pT��Q���g
H��v[�i���Mgf�\�o��E���f��ݷ��_�:����ە���n%����Q��G��7�RHV�CA���z��Ik|v���9	sD�=���Ï�.�-�۵�Y�� r����"Uu������8*pT��Q��G�
�?A���M�c[����=ݓ������U�08�++��LL�4�t��قW tT�$}�A?�իT�+��2_��;�6B}���
�?O�Β'5��R�e���. x��}L���;O�v�-��M�Ӳ%T��J��}�j��+����Qp��D/�}"���\.�6����C�G�����/��9�C�\W%�ֵ{k'�Z�醽�O/�Fm�b�u|�k��ư�Z�w�������O�b���oj��n��b�^�e�����V�_R�8z�b��%��u�g�WQV>x6q�ܜ�y�Ү�t�m{�:.[���sP��iꍡ�v"sf$q�L�K��_����_���XzD���I�x��f��px�:1�m*�o�������q�=��^�ރ��t���W=��H䄺#�u��e�p]���	ư������Q�]�Rʤ�cE^�I�"�8�WK�O�6Qʛ��L�	����zA}w�'�DK�
LU��*v�����KG�e�I���hH�� P�}�׃_v_�H5`�Yв6.Gۘ\=󖄅���'oo������}�_��.6���)�a�G�,��k�+/�/)�����bob����2�V�N��Hsy����o�n�Ϫ��Z�Rw����M%2�	�^I<�u7���X��{�9#�Sy�f
Hx�m�!�0V��fW/c
�*�E2�WjN|�k8q�%R��
{�f��|�{;�vb�iq.�����_E�M؋u��t���8�|mX��՗k�b�n���5��pq��R?=�� D����n��"[<�ŷK���Nb%H�]���؛��-��jY����;��W��%�y�(}�U�?ћ\�I�Xsof�ߟ�7��H�n�Ih��
 ѭzx ��@HҲ��>�}@bí���s��^5�/�3S�R!%������jwn��Nޫ/�"<��9����9ɞkH��7q�^Xy�p.n�*��R91��k�~���B�/���"������M�77S��� ���|�h�0 �̛��zl��:D&����)���Hvy���Sq(ZI��2�QG���&~1���N�Ԑ���.��)���g��%̅�I�;O�%��x W�������i�Q��M���2�ݫ��i����
�o����jF	���r�����]��>oc��k��	� ��IuIj˕!c�� �XWy�˒�3nΌ���}�A��#�<�r�<�$�{��72��IY�����ͅ�m.ZIFo�_����:�ec�ӷY���Ϸ�v�~e��B�g{��Kwwl'W?���J!Q�&��a������ꄕYMqy�����]�m�у�Je���/��al�uGM��r!*��L5�K�5~�v�7�D�3ҁ:���/{~CI_���j@�i�z��6%�@�:333�MɧQ=Ʒ�\�eP
~W�w̟+:Λ{��j�����2�iݯ�������>���P:�ɡ�y����!3����4�++�S���{��+�J3%d��}��6�#e5�B鉄�f*r���_˗�������]]�j���_a��O�a��ʜ8������˜0��,�&�"���¸)(����ax�� �\ѯ�4�8R�J\��e�L�&s���rb��G��ΒXv���;�{�{ ���Ǎ����'d���:���6��7����!Ҥ� p_�//л�=d��s{��W�&;F:�������w�[�t�iY�>��y��<|֎L�+�-�O�/�������[�Pz���(�LE���D���~����Hʐ���_Z��R�H�#c̫�RLFPD���@t@F�_\�m;�j��.��䰾��aV��;���lr�\Sn����qx`��\��h��Rԁ/`��O][[[-R��oΣgb9�դ�j^��q�|�?®T�Иq(�u O�mr��,v���b��u���8DQ�g�;f�$Y�����G�u܌�.��9��79_B_��I����gӠ�E�j����ُ��OA�j�#��]�!���G�ܖ�]�T�9���~gPLs�={�{Ŧ�5�rv`)D@�ʛ�@jUdf4vb�<��̙r���+'%Ȳ��$K>���d�9�8[�=WF�H�'&����v�s91pj���\1U̫��$��h��������:k��O����_ �B:����p��dd�+ץ����_x���ЎTA[�w�p9s*�ر�h&=O�n~�Kn��S@�8�J���7�YY+��nr����k�������2{����ك�'v*--�>	Ȍ{[|Q�ゥ�k��eΓ���ѫ��)��_�N2�IF�"`����ڬ×@�&�P�.M�I������ϯ3��g��
�<yr���K诬���5�O�,�<��tO�t���:<�²p"�����d��_���5�������P�ǽ�-۱+���@/k?����ef�N��aʒE��B?ހ���p�2.�}	��|������Y�Qf�IK[z�]���9c��RI2�3�LO��t�2�l�y{9.�:0�ۧ����\�hu��\�f��C0���B�͸{��4M�	?��'��:�pKH��`��}V�����qeP?,Q�:��82lpd2�j��PG���hwkzY��t���W*�_�gG� �~H�,�%��,؏:	_ъq;�Rm�ҹ૘y��/�@��ʷ|��)*��y �čf�`�����Pd������Hm�n��fa�q�`�6640�=l��B���(����َ1Ј���&נ��襮�+��d��G�r�O�i��j���c���g��"/�1�&���I`�$}��M@�$��W�ޞV�����Ahv�Ζ73V�WEV$���]a߾0°�C9�9�m���Xw(�πg#]S��qX�cNn,�#NC��*J*����DΟ��T�xȶ'��'͡��]Pˋ�@��W ~^�R�m�aמ�� =�3𳍽�?��LlL2��B(agw&r��!�������ne*��nW�s���$�����ʱn)��E6[&���Y�BV�\}ٓN�?��Eb�-��^eg_�0��?���5���x�X�u_��g�g��BJx���D�/�Z�;Id!k�m��(����CCC=�&,�����o�W�߁�O5���$��m��mD�N=�g|����U����	|!=�O��wa�ٸp��ݻ���^G��;���M��a�N��sA���k���Q1�R�3�U ��fz�)��ZC��σ+������uu��R�1�t_Y̤-��i#��{���z{�˽׬ĳ'������g�+3<�}|z�����U�m*�S	���ѝ��{=��s�Nn�sh��e��U^���j��ۥ�ms�퇜ن^K�'(h���݇i�x�-%8c�W�w'���g�񜠟�F��bg�RȐ����c\��D�������u�E��b�[���3yWD�ʶ*h1pTf���`_���Z*�X�QZ�A[�zu��~�F6����+������u�T�$�\�
�p9$?O��{:��D.�+a�7�y���hpiz��d��o�Z��q
=�0F/�mۣ5KW���j����0/�������]���R�W�sk�M�茤DN�#���-'��� {��/��#'\H�3�;����R"Fϧ͆1���ޮچ��3`�z��F�/ԋ��`�R�3�����$ڛuf�e~�65���P`� �tXaaa�2*۱Q����x����r�7\?i��~;Û�gm���?���|�l�,�\�S�*��.���.�+�����>���F�����+/D>�7 ��w���؀�ʾr*���Tv5�~������h�
0$���$�i 64~�O7���Г������ҋ���	e��o�]SlS2�51-b�B�G<Pͪ��=�n#��Ed}ĈN��ό���ǡz��>觙����w��5�Z��\t� �<Ul2�Q��ɡAJ�"Lȅ����T��a��?�=]ݐ������?�JC\&���TVU���`a�;�����n��ː-����x�a4�fk�O��"
�Ӫ�O���a��huI�Xw׳�ޔ��|ZOp�"q���ҐL�X`S��+���;�\�{����i��n�j���AH�{h���Q|	屘S�����	H����o�nc7�gk#8w�W/F�����lڗwo�>oi8a�7ȭ�ϖ����(���~�Q�- X�����O�o`1�Vf@p�Ç�C�}��J|!ugH��81p���˫+$�������K_�S=}ګ����{Ĥ�U^����!>*t����u��Pob`*� �Ȅf�5��U��7�6��$�ͧ�P-��簧o@���	�����E���Y��
Z��IH���T��;��ҫ	��X�A�g7b�ïs���G�������X��I�p�!H	Yw/x��}7�����<���_� ������������A�0Ǧ�O�,!e�&�������ۗ��i�ii_Cؽ.�)�.\�ƺ�@h�����n1�_�����z���*�[z��({�i?���8�>E�S�m���[���/�8�?�����^��F�&+}��](R߾�<��gū?o��@�zu��nn��i�����3�R�s[[~L���E��U�!�5�E����V��x���/��V̲���j�}k!����kR���tC��������{���<]`��&�}۽3*K�;|u�C c_i�A�
}�?Hq�v<l
�Zf�	z�$ZU���8��0$�;���r�]X��u4k�~���LE>�_T/'���}��=�~9��+�ݻ��<������w�:�j�e��?as�C��,#��^^aaa�6Ч2=�!���.���v�[�Y�:��Ȯ�0�`wuu]�7}���8��)�P:�,�V5�/~&��2^��=�^y�0����(����Y+耇G{�Z�\����ϸ<�/@0+`��ݻ���%��>>>V��L ٸ�Cs��ѓ�kG���=�/��'ӛ�SC�1���37�a�ܤ��(���qWfG<��e�A��r��Ѿ�`��55�� Jr��?ɯ����]a�C���O�<���U��+ab����y�1�=� ��K�
QB��ʾ7�9��0H�1Ʈ��{�t��}��Bev5��=���Ð��7@�����3��UJ����h�ɓ`=���T���!�@O�q��2Į�x+ʒ��vh���{�t�VٗE{Iu���a&?8���H³���vz�sL�[����v���@�9P���)'�����*��@Gl\�������g������Q6�(��jo;�<�ﳖ~�i�����-&�xC�����K"�ǒX�����0X&a4�fEa�8Ӻ�����P:�������fF�<*q%���e��kO�A����Bʯ'�b�+�V����wumq�����pv�V���`�)�[�_~J\h�rr����7��j�m���n/����{��c!S��T��XT�ٰ�'cL�������$���돻��+R5[jV.���P�͘�?��-����ߕ���^��K�F��=�IiK)�G��I�����ݸ������lv��laz�e<K�T'v�1�󵥆,��eJ���tE��v\�i�!3���5�&��z��%���hU��a�С�y���z�3Ϯ� ���̗�����[�|��DEM���H��N�<x�F�}��tn���|�aӀ�P�����g#P����L�]�9e��4=�z6��zUK�2��T��e߾��i`�:�����Mv�"j�*ﺻ���ċ5�����/�)6���]�(fR=G�װ��O���͡DR��K�wi'}����S6���319�����:�莃N�u!�@�)�%��I����Y��#�����eΔ%��z�d�^�!h� gFLa��ֺ�Mfߙ����'nq�P!����>��ׯ�W 2��n�ėپK)-����E~����w�3��g1��g:�� ����Ø��;�Z�5���li6=��V�CyF�NUK�{Y8����Wۭ��ԓN&1���/�0��|��(����̉ҩ���މ��U���;����r!�1:_�θ����c���Y*fe_��[��#����L -&���TNR�] "��,.��'�"��4��f�PΣ7퉎��p2%N�������
c;S�E�����k/	'��wQ;p����b�}�yˆ�yyy��b�s��wi�)�y6}O�j�(C��aw3��L�bB��ڥ�x28�S�O@ �w��+ؽ�5$[G@'���-_�F$��"�#��v�(E���C���l6���B����&߲�5�p�`���o#�@G��m"'�����;�G����t��~w�2�Ō��ԎE�Mi��ω.��L��J���A��,��-�1��ۻa�ӄ�|麟`�K�)�W��˝��UDYs=�KG��XS��ڹ���r��J+��zM��F>��3�u��$j5*���.� c�����tC,0�&�j�28_?|�jt�1���%f�`�^�>hZ�fI{�V�.���t��}���c��]n��v'm(���$m����3�ؾ
>�v��8��s;��ʾK=@'(z�
�r��)�^�3��M����`�Z��F����@*8���>шE��$rnfĔH��$����C��-�g~�t��1eK׾K������(t̗v_NZj�垓.IXx�PV�(9�J���zP>�1e���TU
P}=�����%N�@�Y˗/����	�Y�� U���T&��\� fҘ�,rp��s��l�8��StҚ��Z��΁ ��HPbc��,����I��3<�@~��m�9�7WDc��.���ҧl�u!�l-�K7ٽ��j������{����Z����t�g�K)��/�Й��r�AМ"@�{�����C��D:����l�y��~�;�U���{�̕�i�f<'�go��xt����f�*c���bu/���rr���7�*U������/�VA�Z��V;��ɮ��-g+B�#_���S�ҕ����K/��:�n�H~���g���a$��
�/;����	ĉT�B2�+�F�b��\YY	5 6�\hs�9 ��gڒR)1�i7�)&r�(.̞"��w���w�v}o��&���R��m�s�r3ʦ�������Ŧ����|K;��ɟb�.�w��]��K�b�]?��CZ6�p�_olo�CC�p��q%��W};ʨx�_�Ź?��c�b��7y��5;5��@ۉ�*��gg�B�S��x�oϞ=�PǿC����ǟb�`�z�T
4g��G��V�$��Ӟ܆?��+˵��c��*�:'�wOp�z�;/�hS�U�R�H�bi�����_�� 6GOA�&-66��r}J]�r�a&��� ��[��WŦC�wy150�%�e�oy��^���"0;��ǹ!-/o0��f����7ؽoIJc�m4����e�%��C�hϐ-#+��Qh���.�.���՚.78_Cm�b��Ągm����Mo�z��'��ӽZ�:�=vlp߲uZ%{��Y���˽�� ��2���3?�Xf���'�f���~�ZDO�?�X/�p�gc��L�W�C����G'�!��Y e2@�HKX�cJ�t�����?���Jpy���.!�$�2b�����s�t!�����+�Ɇ��O��l��Z���9�:�3�v�RF�d�u���B�8ؾ�7��y��$ۛ��-�|U0��j]����DNF���	������l6j��@��=���+x.��,��-��s�.ġH������#0�z���DN�)z(�G�-��4�^g�i�ۨ�ϵ*�4����ad�B�E�̧K�<�\C~���v�W�!�L��E���JA����FV������|l}��!�. �� �)@Ȉ�nu�y��[]�����(^:[W�U��, .��J�֭�2y�������mG$$���z��W;��\.5{�@Q|�)vRUU��#d�;�v�o���Z<]).�z�=�iE��dݫ#p4�e<ߋ`d������:`���l1𘩓��'Nt��5��>755�(��e �(�����#s$�$��m�Q~�V���葾�~�������y�xv��SF�����z��>��C�8#�P�p�p�o�}����P;�C%��Փ�i�����p[wh����𿘙��[!D��4�k�J瞷�$�]���X��#�^E���ep�[�G=б�!�I���e.$����ci������qM]������^̵*�ԆVM��2
�F��AAA N 2��`�%VD�j1�̊�(T0T�APA�L"��[������__�O�9���zֳ�����L�Y���SxO��ZN���G��N
��	^|�<pJ��3�۠�����ň��^��#�I,CP��LM�/��+�?����G��/�?0� .�XV�dh|2�����������Gث��|=yZɧ֫ҳL&��!0��2cu����*m�f����]�;�&s����:g *s���#g�m�S:�u��0�\�}�}x��4'���a�.��'lN���a�)�����V�Ovʔ��t�w�		�_��`z[Ҍ[�!��� #Kx0�\��0}EZ߅O� ��M��\��Cx�ds��g_G�Si�A*�����*�'�r��[wr�e�]�P<�^43p�,`�d����pM��%�kT�[ �?���.an�.XH\�A�{�+��qƧ����a|z�E06;!�Z��͵j��P^���������@�k}��u�?�Mc��5��|�i�Bړ�>|%<6[�I��	�5��M,0Qe�?��7�X�]Ӕ���1+ZA��6T�zt�ᙐ��Q�e)��N��m����`v���'!��	��ط)#���7 X�9g>��T��^O� F�wM�*kP:c�-�����݀������ܷ�&�T����\��I&���Q� -�Ak�+f|W�`�ҥ�8���I����9���3�;���^S~FY�f�1≚���d���9����`S'���գ�F�^4k�����N���egAޔn���1>J^q�l+K��b-]�l@S9 �bA�A��O$�]�<b�!|Cʚ�k�8%gL0Xq��7��
,>�=y�#&&fҜ�����eK��ZY寠? p����cת���]��X��i��#�v���6�50�p0p�f�P�l���~|euO#�9�H��Z���^[�	��o�+f���>9^uZ1V�������C��5檧8��z��ΝS�O�'߇C��%W����6�u͚�oͳFSp�!�����9���]�-zwx�MjZ�h9�tXW���o4n���U��w��T����������Xw4@I�%W�*j�r+�ȣ��°Z�^��L������G(b7�KB�2^W�{�tԷ�F�_�����GQ�[�����������v�j�{M�����u�=��uO��������{Q/���N�_�����u���_�����u��Y����C��#{����3rW���O���[����9�/��|as���6,?j���Yk�˲ϼ��t��DZ�W����#bΆϾ��U��ϯ��f�E�/By���	�w88dH'��9�p��`k�Le�}�k�@Q�ę���_����_�3��_SX�o�,���O�k�B�Ǧ��6��V��ٶ�m��L]����6�?�[�M����{�%�s@�V)���ӧ���F����&���@Ly~�j�@8׬'ۘ>.�5}#�����~GG���/�����gI��>#�L�m@8}�}OF�	+���z���bt�x(F���Ƨ׹̼�}=*�,tي�ɁL�ŏ�5�o���~�F��ܿ������
4���v9���ٷ�9�'�!��ۙn��^�~mpgDZd`d��?���eJ��ۗD�Oh{���̲�?V![2�S�Ϡep�N�8*�y�T�g�jGo��CP������?"!�K���1�C�a��9t��q��Do��ϣ��Gu��{�4Ķ0�\�ċM����yh��r\>v���hF�#@D�h����T��飀�tS$=��`��:8U�]��!����8�}�ԌN�8�?kkk��r�lf^��Ũ|�/�b�X�)��	1���z�s��?ߨ�1��ֹ���wCv#����_D+tF�������,O�����F�Ou^����*�az�9E\�%'�3�����������p��1@��󁱉j���%<$�+�Ģ�2���D+�$*�dg��V4�[�'�4������G����B��#�4g���֧8����7�j
+R�v�iM醴3�G�	�K�� ��KP����$T3��j�;��v�n����	)�4n":M�'��Fʺ�j.�A�^�}�1��{�{�/��ّ�D��+�^��$��>���l�x]��M&a⍏v�Lt��X8uK~&1����j�i�Lm.l�P���,���MnC+s>=�6>l�ԝY�R�kg���������Ւqg����(�
^s����l�d�����)f��Q�&�i��܏�8��B-J2J��-���)�d��~��=��u���������og������:6{�w��_��t�Z��i4	w\ł��3O������3Sګ���簟d?U�
N�̑���9:	"2�p�!�$O�.��?t�a�^lT��/d�w؄Y��r���ﮮ�Z�?���E/~�P�p^�����|7��޾5c����B	�՜`w�

F�9�3+��L��|��8u���Q��}��FLY���j�1�"b��T�&;%���fP�7g:"d5=C:|�O3?�j*��Mѿ�iuR���$gg��g-=VR��4j_��-�90���~n�!��˳��݄�3����gI��"�:[pz{�r����jbc�S|9��B�hyh�դ��7���8O"y�}���h.۬ƺ���PxA�
&�o؃��P�6�b�!F�h��#.e֎�
��c��a"n50c���Z�i���+�٫h'D�7Ϊ�o�q�����Iw�ol k6���>�-x�&��{H#���w��3c�W��&�$}ô�A[[�DY��n�g/Nu�}`}��Eiiig*��Q,T��p�#�L���P��V�w#Ć�j���-�No�J͍y������^q�_��c���4Id�,Y�P���6]ʲ���k�k�.�B�/GsV���Y��Y�C7� ��wk�b\C�A�|�f'纎]3}|�Z����>e���DEB�O;M�5����a��}z��2���g�w�Đ|�L���[Mn��c	�t���4OO@ZZu��0�:b�'�~���-ɹ�a�+�b��\#����n*�yH�ۦ��/f=�p�/`<�|5iAX�ʹ�G��p"x��a)|p=wy��]���bܣ`�`xnH��N2�� Y��y���[���ʇ3d�XK+������	���^�jFo�1�e�����$N�
8���Yk�U�S�Qa%�t��8�B
>��S:D���#���#d/��Z�^���P^O�za�(�{!���g.s�7+��9�����#?�b'��ь����_(�ܻ��Nኸ�S|yPik�8'���x���J%C���rkW���|I���3��s�U�_F�17k���1sV�8i��T'��!��|\�.)V��f�b�Q�����o�ˮ�9�ai6�z��	�BU����}���`��%9Df_��ڷCz��7���w2���8�6�Uw�[L;�b-�����G�v4U��)@�v�H�)�u�J�_��|��X7s��d�U�ܚ{��ߐ��"�Z�w�054ue��_��u��]�>$IE����� �'�u,��*�:3�QK �^b�[�\��VB"~���f���r[[��*�_�[�]"N��FB���gM��0��A�����3^���gn��Ө�Z��"<y=��KM.d+8Qx���������i�$S��<�h�����a���<��x",1A�3��R�I���*�i?���dTjn�^!j���}0'��?������<x�WC����2������bG�k�J���C��Ei�ָ�L[���;��Y0���� V*1�j�F;�-��Էu�t�K��N=&+�M�)�W�;�޾}��G9�C��kLdZKMp���*~�:�1Q� �f�4��n.��c��%!����B�_:g�ϗ�qvd���� ��Q��Ʃ<Zql�u��9�!�����Z����<��
@���W���(�v���@7�~Q[�"�6y�6+�WNu͚�M�h��jxC��3�J��Sd�����(��P;ԭ.���� g������h�&�f�B 6A���]�<]ݨ3���y=q��׉6U�th}K=����Y]Cc�d$��n��}|��I�a�o��!�h4�	���0i(kE;cx�.�,�1Hz�Co�x����F���K��P�e�XU��sTQ��c������ȼ��/Uh} P�wL��,Y}��9�\Ń��)<Ip����}��	�ǻ\��2Ku�=ň�U��N�
a���~��S|hnm,"v������M8�L�I�h�{J�Jg$/ԟ�"V�k���w2�b']0-�)W��Fʚ�;�#'5:���s�Q�?��E��a�l~� �4c�-��w;(�%e���%�����N�"˨�C���⫵ַ���$��bMM��4����i7�$���0���tĂ�!��p�,(����zP03d6��Kq�r-*gq����O�T"я"��'��G�3Y<�p�ѽM���G�������xʑ]>�M�S��s.�*�`�� f�8�����s��K���c�qIMv
˯-����-�`dT�`���i��qf��\��:�����Mv�oP!Ϭ}gblH򱍢���^������'N|�2&�l&Q�=���>�����@ď�ZC��#�6W��3�(�n-��i�&6%�*�<t�o_A�@���U�O9�s�]""�VN�T)��2vtu]��{oR�w��^]c=�F��5����D����	TD�i?�%��c�
�!	�s
��7��QN��Du���9�c5�	ze�DX�@��4�J�����/���ǂ�e��+�h��{�nH�]B�.�	�_�7F��{f]ч*�T����(x�~{���sY�,u�TU���Axa��֪?-�*��P.������p|�wASwa&�t�������b��:�@�d㔗=�!+v��O��}uGɔ��l���9�0!��P��Ԏ��g��V��Y�{��r�o^�EW�M�D3�`��$���j����.Ĳ?y8:B!�V"r#"�����["��O�c�yT�έ��C#����"�+h�-�|>�d�o����}���]3j�#`�8!��<�������0B�o�V��C3�Z_0�z~�bH�d�� ���t�"�@0��숏-S�G��
�����1���������E�� �����і��~��y෥-�Z�!V�&�3���~J��3c��h�S�D2��u�Ʃ�^����r5�"�~",|?�z���������F��+kk�Qf��
gx ��Z$BLk�f%��AE�7r����pK�����_A�|4�����i�|#�_����U��me�� ��œ5�!h~\+`��Y�޼t�&�*�Ar�Ko�<��ӷ�I>"�r��$�av$�@���zF[�a�ϲ���V���n��dR;����d����Ċ�;���둟?��"ze!�-ʭ��G�����]C�Td��Oj}��k���ca�Ȩ�ѵ��jA�P���P�ݗD#�
�E�f��j'�@&�Xx�j��dV�K̜C]��b�!]%I�I�25��k@�����i��z"Bn��+Л��Bn���y�������y�xǬ�F�$l,w"l��f�[x.�gcu`�[DKA}=����}��G������No;�)���P��n쨡΅Fhmw䊻�W���Z�Fn��h�e�DrG?���{1z���s��ju�3�=�s�A��Nar�j�l�x.8���ܺ�����b�B��#
�O^�׶���Y��Y�<p�`<U�vD� m=R��+pwV]�ۇ�T�@|�)��"����;}��i�8Y��? IMI��n���H*ѹE�G*��=C];z�Nސ೤>��N�u�uV%�W�0^�U�{�5�.8�t�j���UU�=�@w&�<γb~��w��od	��V�w��]�J�������ϝ�1 =9��\��7C��{��
��{3"�[<S*Hĩ����k��)j��c˱��щIEZ�M �Y��湘D2Plp9|��'���MU0��O�,p�W��'��u�A�!�Ԓ�7�����.�J2y$?��ƶxnm�L���\ L�~z�Ed��()��*�VY�K���z�����tp����<ȳ�`�q�ݖ<�!������O�U*�&<C��5J<�mV�Crh�vH=a�z��/p�x��|Eb�I��T��ص�Z3���8�����F>���=6.����f��:��z�ʩ���"׹�)��i!)&�q{"���mn�ھn*ֵ��O W,sx��6Br=������9t�C�)8&4e�k\2����(:\0��LAc���]�y� ��?��"�c��0r+�8\�F�A �v����
/����*�s�U
W���B��P�*���$B �d�������I����,��4���])@��vT�r��j�>�Ľ�$AEc'�Z�㼿����[�G��+<�]:68H�S�&����3����x�uEv=��0��1�F�'��k:}2Oq6`��=�n�D��Y٠LQҳ6���h:Uk��� u��x�D{�;���!��"�j�&\������ys�ۏ����'�e��Z�z�d��<�B�6q 5�������{�=�}�<y��zx�gQ�S|�9�[Šy�3+��}<;��J`!\��O���:��~�4�xH��\ױ��)�����F�#)�r��AF�}*�L�mOz���dZ�\o����w:gdQ�r|��ߞ\�x�%��+�@wCe�񸭭-���R�"���D�����v���V��D�s�����V�����C��V�������Ldޚz�!C���Z}�9�d!�{�����u�{ċ=�E� 8���jU��><�ם�~�$;����[B89u����R�%7����@��[*��2�������ތ\u��ӰЙG�Y� =��*
��_@o &X��oW��^k�k1��$�P��`z����d�L#��6�+�e��`��A��Xj��k	6���w7NQG|�\�����J��N@@����N�Z �a��G5d0�r�V��.l?t4���¦&�d����� &�b�	�`@�?���H��df��c;�(��9e��U�񣀂^Y]�- �JT��v4��խ�2�J�GE� <��{X/���/����f��Pu�ʅ�"k�2��MS�.�!(�ؽd�'d��'L3��vѥ[���+�	\OR�#�Y8�y��.�707Ћ��%��y�a�������U���B.�1�ălpd�
�v�e��5kB��IO5�؇w�r�h�~��)،9� N��9�1�8Y��.j#<��
��^�$jI�hy?����c�����b	� i������v����R���1�����T���f���rj�\�_��	̤;�D���Ŀ��7�A��1a�.��呉�"h���9w=��f���[��ڃ#{���]�KcM3Or���Z�#�]~4��ٮHR¯F0�b��L?‷��˝3,��	�%���i��*)UN͝ĥd����θﳳۃ�ɓ��U�;���ڿ�H��x]C��{B4<����%n�@��%jo�ZC-p��S�d�纊j���Yſ�G'�ן��T�*Ů�CWV����g��˷Я��~���7��&͙˔��'*G3�?��Ƹ�6gg�&�j#K�2Y�qF���%Ү�Y��cܰ
�1�b�H������j�$�n�eȟ,�� ����<��c��j��Wϭ+�Δ�m2�ـb�ɻ��ʓLNr�Ѻ�;�@q�|�rZV%�����ԏ��ķ|�����#�q�b�G�fL9zz��R�qC�J%���x�9�<-k��9�xj�	yz�59��������x&%����m�_���ᾮ�ݭ�X�f�uʻ�_�\��u�$�rv�Y��	�-��h%�h�(sӟ���i���2K�:�v�.j����S���*�}�\����]�`}n-)��i�Dm�uW��2pΘ:VyK����.���p}(o��>��~"��j+�]��V�-����
�/�:}6=�H�Cxƀ/��Y�GUH$Y�eN)	~����{�>]���x0�G�7+hy]ӑ�/s�Tf;�Q7(G �R��X��$�#N�-@?{��������"v`���@���1��V������  ����!���X�.j�8\%Q�?gJ�t;o|�r︬^Ї7������V�<��K��g�xj��k���~�X�����A����f�5k�4.�U�M�M�Gt��BH�޸�+�HĂ����z���he&��(���O;A^�m�99@z8�vБtʁ��"哜)��\�MYZ� ��&����Ӳۉ���0^1��N<����d�J�&վ�CT\��fB��;)���v���ƣ��4�P��.�F���^kk��eȈ5JoJ6��.`��;��ς��gΓw>��N9g�Ds�!%��Zgrgh�x��6��tz�;-��0Km�� �έ]�r_<K�2�����z��Tq4��"�=R�&�k�{&#=]w��G���q4㰚���ŭv��u]ح����D�d�P@(.���#��c�tkl/;�Í����OwU\-��
0�Δ��ǳ ٝ"�M4n���Û7x#�B�9��궓�
�ҡ1{�S���ܹ��i�=YH�]̭����t�lěR��>��A�X�b�8��S��z����窐���ɿ����ɝxg���_U�rJ�f��<W�|n2��ޑL	.�O���B�qq��x�]a�=��$��;i}�fL���r[�̾x4C)C�^;�6�CPQ����P�䆡�7�lw��(Gs%�+KR>�A���j���;�K�6݅AE��4 ��|v7�6�;�1^�4^��MA�f����C��!f��!N}�ZK�Z?g�Οs�'�R<Kxw4ws��e*��<wI$�Q����1���,����/���e"ea�ki7����9c.� ];T~U��.?I��S���p�52
�E���X���u��$��5�hdA��zn�n�5�� \��oBւ{O��cG2.����Z�F�P��[;�{)��n/�*p��3�5kV�Wz�q,�ꐦ#ꣿ0C��eg�3 Fʔ�z��.)v.]u	�H4m�����)\��L�e��kޤ0Vjl�.�tP��ϭdq�,�@��:��̬�o�،Z�B'/6��o�d��*j�ExqwT�(��v��S����oS��t�ώgJC�&���<w�������'�SsuW�d�v���{�NV��$�Ҵ�u�0�D�����n�~��7ߜ�|��W��׮s�V�}I������;L��şUM�S��_�L�^~�T3t�[�Hta"�,$!�5����*�ٹ�Ф�F�Mj|C��:����&"n�5��L��I�=8���|0N񶅄�x�/a�@:�x|��]�i�u����$(�R�H|����J�C�8�Fsd���Z`����T���d��`�;Y��999�H�l�,P�F|(nz�X�������D�B-�����V�)Y|�R7�?�y����G�h�Q R���,�K�#] 2]W)�����M���
���C'���+�DS_�b)D^��l����K�ńy�D��Ժ�7Jػ��Y@8�gu��<+��
�
r�;�-:I���S�{���lv
�*��������IN���"�h�irйy�I[��'�.�j��`��� �H24�M���i�G2�O�mm����zۭ����)�D��D����be�:��!��/�tr���e�q1hi֍Ρ1�Xr(�s4�9�0�N�8�O_���Q�d' � |%�THMgM�;��������$i�������g>��6Y��� ����1� ��}���aV���aU����� �'���^)���E�˅3�S͂�´T�\�y~��-�م��;��Z{�E���bKZ_%��d/��%���Ǹ2�ءx�<�u���o@oS"?�J}lހMW�ˣ�EZ�\0�����r�!G C�*�b�H����5/\���j��&��	*V��U��N6Z��!M%��s�����po#�������dtEq��%���]�5}�'U㊽��y���U��c��'9���Bh��>���L��M��;�����@�.�(����L�;{ɚu������jq�.��z�����o�tU��8@��ƍ�Y��T�GԵK|H޷�m^��#��f��ڙ��ښ_(��H�//C���Ul��s���!��Yu�Ν�)V;�$\�%R^�O䚺;8�7�q[ᷪ���N�:B��<;���_싻b��ڨ�k�OsTH�}x�숏�m��Z�Z~4��Xz[)�s���c��#���TT:?��+�b/��j��Xs�G&q���5�xީ҂�Z%�]f&��/k�@��I���-����nV�Q�MF��!��pwM�����t���xyc�P�+��<�l�~EQ�/D�c�9x�,ΰ�m�� [T�-����� ��l+�'���������*u��8�9�L����i8v��	/� ����<��LwK|;*J<�Y[ʭĦe;axF�w=���g�ٛ N<~C\�V�V����ż�D(�KX�t�J��cN�]����U���Z��`\��h��:�9��h�x�~������� U��Vnbbb�An~������g�7�����v��j��0�#� YWSH�M���c��FDmOҷ����6\@��AF�P�V�����/^�q��mUc��v�$}Y��v��� �a�U��Se��Ж��*9�	�!���x�椦Ǜ�%Gνȭ�d����jr�҇�T��p:�kc�U|���f���9�=y��"�*�U�35����-q��D����Q/X�1.A;��F�*O����x$�_���@�^��VT��.3��p�%����XyC���!����C.ZN�ws��a�O��8W�Ɋ���F�vQ��X��Z��B����{�/�����Bw�.#�_��W���#V7v�*�\qύ�ŏD��0�^L�����4���3^W�W�C�n�iE����"�\�;��"1���N0s����N��ր"�בU�PQ:�s�#�1W�>������ș̉"��u�PO@�0�6v��t�N��DsE�l-�w�F)�[�� �I��At��9q��ض�������py��dMN�^��^�u�P���Tr�1��ł�Ps�jHDrx�@Z�VؕR}G���:��!ƻ�/IO����16nN*mgH�ۈFoذA�!׹����;�?�7\&%��8�ܵ�5��rv���IM�n��l/�^�n��y����m�B-v�!'YE�E#�&�;��hM]��b��J ���J�"n֍�?n4o޼3�?۲gaX���Γ,����=��t7�ߙ��m����0Ƿ"fm��a�n���s�(�����n�� z<5�fEԬ�����$�a�ؑ0t�睇���(�ޮ|$�}�nU���V�/�懲?=��v��KD��Yuc���ywA-fB�aI<�x���xf�r�E�1�r`��7�\���1Ѐ���ܡ,��������+铹��F�����M0S� �\�~_[�5!����3_AzLK=J�?�r||\bP����(��c.v[[��������4^�*Wa���]{JC	�K�
��m�A�x��Q��t��t�q�DE# �� |
�O�D�,��q���go�<I�w�~Gw[>������%��)��c<�S��U����P>���J�i�%f�Z��j�h9��Wɟ�{!�Z��^��~���۷�3�RH�W%s�Ƥz)>_����ꋂ�6;:8�-���Ӷ���r_M����Էo��91��N3��9(m��s��~�Y?kE#[-�C��
zX�.���Kz$�H�Q�ACc������<m��7�?�$�1�qBU��]��)U��\c[Y8ىsIЫ5�����a���4���q��=6_D�Ưt^�O< :�3�I�~�o^-E�\0�3N���:��g����C��[^�^Iv�[NS����\�≰�����=CS��oI�	oܸ!��#`;�D�Wz�)h}�s���f�"H���ma�����nM����e�G�Պ�����N��.JN^�)��d.*Q�����FFE��nkq��)׸�~c[���פ]!��2��>3&��=C��(��C!�b��B�]Hc�o�8��LK�_�8[��.��c3��- --~x��Gu���}���0m�~}I�}��m9��#X� ��B�Ēl}Y�����r&��	��Aa�5HA�C-����R\剀�*ȃ�֛�T�ќ1|(��:�GmW17��^:�v���n��8��v�T߿_�W�{��.��,O���ػq]\BB�����,I��f3�-^�t�o�D���;xh&E��qT'Զ�������Ҩܮ�;�{z�.@_�s�l�X�ds�q��Jm�ۂf�ޖ{C�y���\S�=~%$��:�#>�Wo��8K�1בCK������=��`.�ؿ�!y��ɑ*\������}p_�i/������E
���$7_�9Lʄ�9N��X+�J��+���or�;��_�/X��R����;&@�Ǐ�l�	�\�!M�$��������kM��ڎf#V�-�t���& 
�X����*A����r�o��/�~5eO	��%��~N�^t����?�=ͨ�w�;̒�#_n�H�Ы�J	���$Y��\��P�ot�e�|)�e�A%�*N�&��u4��X�5�r��Ns�$ �8��l���F������e_xu�Cu��2���[d�-��{��"�d�=XQY9�t�"�ce2��	��=�~�+�t){1���z�6�4�2GDav��g��
�t�"��"Z�q�E�]����=�ooÀ������&�_]]2�F~�!��#��A&�願�t�z�h=ѫ�{3f꟠�Z��9(�"��jf�'py�#.����;B�������|F<h�jHC�:��%=�� ��=��*�~�@��5�:�V�d����T"�[��EP-�詝�{8��<(�i�('�Y,'���`�N�e�e>�?ϔ����߭H�*a)7��������{�lU`%�����/�o����gn�q���N8f"���'9yP�Y[=���y�\��A/�;l/���8Smg�k��3.쉷CcP��X�S��_�z#��E�/4�͊���TX���խu��Σ6W�� i~��+"@c9C�a��H������RS���t�'��IMN�G}y�״3kp�馬�.��k�LSn��}派>Ҁ��@(Z���J���'��;��S@�/���@��o�x:�y�9����qz/{�@��>���js5��:!ۘ���<���D�88:�R�p�@�uy1��Q�zL�C~�%aw!���-2��'kiЛ)����Ց����A���`��V��-�M�՝!P�w@-��/ߏ�	�&$�U�Vvu�4v����~4꾽l%2�B����J�w0����Z���}��+Q�M_+�]��N��XBs����䔔��4{���d/Q��x���T�Y���~�ǽ/������m70x��U��?��_��B��X��X9�� �yy����)
%����n��U�V��*v�����GF��݂���'&�E�L�jA�^0�nL�'�B0h� �5g.҈�O�AEy���޾}{=��k�z�k|{Z�P�E��7����VLN�eյk]��K�LJM}��~f#��o�6<���'���Y��Q����b��m�k2�����S�R�l�d��ոR�޲n�b0JB8�%[n��'�����ݬ���p[m�b�466�T9�+~��Λ�nlvB��\��"��b3��-�u��+����׵ҁ^��_�iu<i���ʉ(h���?��K v��V/+;�#gP d]���Mv~�;�]<hj@��2��'�F������^��+���)�o���ɉLNNN\F�����m���>.�>�@��\0�x��I��ms1y���)��	�͖T2�Ġ�$�ۓ>��w����F�m��p8�ug���`��㢘����?�DJV�dL��Z��V�%.5X͑}�%�����<�
�b�r`u������5461����TI�8���\㐢օtV5��oJ�t���~`+�ң�/k��5e�=K͎�N4��73$�)�xb�#�V�̤��ο�߿��x�|p�rՑN�St���������Q�8ȼ��)M��rcN�� ���.m
��v���;;�����UPwO��M;�%��\ӆ�O�)5�� ����(	�f��]�Ψ�����t���"�$�m�*��0'Ȩ��d��-��S��<Ez�{�9��;B�J$���k`zauDQ�S4򕙙��]H�ߒ� �\𢳅X����"e�3����A�Ԣ1��Њ��T������|x�l�QuH88�x5}��!�����-F�A���MTX=�!�+�U9��]��>l��=-8O���휍�~Ƞ�5�s�H�n?��<�D���}�)��n��#�pI����P��ӖF�/ ���Jt�])S�}�$�����V��Oq���Y��W���>>W�X�.B���[����jH�)&&Ft�#C6N���Sk^���U�+�ַ�n�}w����r����c�'�,s��L�Q�JM�^��;B�s$�g#
']�4�=ڹ$����۶�~	��Kw���$A���O�,m��C�C}(��Q�&��8�<���(�^�����f��5Kg��`�C!�Z�`ℍ�7į�!���"@1��5��c�菺C��L��NA�z9�3���e`ʪ���0�F��e[|*�7e�*6�g�M7�n�V�
��C��E)N��\���2kf��x��f:�3:�
ݍ�X/�O��>�-�ߏ�톊c	��$�m����J����2h���S��8û�+�w����^6�N����������r�V�aS16n���^R+X0�р��X������pR�_<�37��{��ؔ�Cv}����fnn�������~	1kf�MD�>��z�n����\yЀ�m�kÇc����s���R�$��Z�
�>���Fг�!}�h�h�d�\^� ٩����x��� 6,Y���W�LY�f�_i�;B���=44�CY��1�-LY�'�R��ݝ.���D��{��x�2uo����e�@�Gjq�ũ�!��9��sԬ�0��� �w��߀�2uqEG�b1�:�b������"M��)6���U�`Zp�X�f�o @Y���`ƒ�F��׼,�}��Q)�F����~/�e2���	�V��΍�:��*�`�%�9�$!��ipJ��q1��X���a^�񃤏�$��T�����a�ޛ��BD#�8q?��LJ�UՕzc����u��aFo�!���f(�� ��s�tv=��K��R���0ώ3b��
�ߐz@���G.���o��۰"T\倫�x�+����;��!�?x���W$H�Ɣ�	�h�ş�|��r�dT�p�������*��t�������]ςҤ�������HWl|�/1�h����省5���$@��F́%oQ嘰o��u������w|ZQ ��ݘ��L���n���+��p�S�w��0��	�~��-���ǕF��O�IB����'�L�^MN��s?nUD,� �����n�h�0^Oc� 4X]G�?tTi{̭ʋ%-���9G��K0m�G��D��2}��w>�u��c������q�{��	9Vq}�Ob���h�X��1P�=yv�C�w�<�]�o/)�q���	w�F#o7��Z�ͫ�!���a�ޥK� ���/]*�����4�#Ô�;���Vۿ♉K���ݚ<yf�h$��JM��6�������&o��9�l6P�2>v�Ҽ�[-`�(����R�̪��x��O����=����\������-r�e��Z%װ���Z=Rh.���O/��z$�^�:ĂP3�?���[m��`%�ǜ����ً1�nE��N�9Jk36����8�/I���ua����n����x��3��i�[�����w���Sg���eY��T�:\#��f��T��t�������epc��wx�����^�E�a�<���nk)=ʽ	�$�l���K$��20(�X��5���8 ���;J���y��,�^������x�,�K��q��Kc.L]-��%d��v�['k�E��c:����Gg�wے���T�s-o?-��"�+7�sT��U*p���Q6���-Ȭd1li��]�X�iZ)P�'���OU��\�ձԀ�W�Ph)y9o�<��Po�K~�k��3�#(u�4�(���$��	 ̖֗���?q�>ڱu�E|�/�^�W^����:�k
4�K���L��.��:>��a� �S�U�f6\7ۼ%$�v�k)R��o��R�Ӆ���P#(���T����k�<~�N���<@��n����oܪL�<�U�M���z/�6�i����[���Iv�c~8�?
K#�x��jP߰��gx{����ʵdc�ص6��:	���	Bh�+KG�0Gr�8�8_*T��z�^��Ơl:�{ֻ� ��8�$����ԁ��@$�ƿ�O`s[[�XZ�v�nL�ݩ.�6*,�r�����MI�k�t���ľ�>9b�p�����n�C3�̂�_�uCA*���>�L�YVJ��P�:�b�4G����1c�Ds�M�]�4���V�N�k�;�����b;�nvb�@�rlb��Ǘ	��%��ذ�n�yvħ2D����g�T�/�'=�a��U�~b��FL�1T`�&��L�{�J���4%w�M@�<8Lg!�fT����	dVpI�@�NL^�&�ZAXIx �M� �����OZ��2���J[��(R��nO��\��E7�E�l�c�̲T�����MS �?8uL'��׶Ҡ�O[������P�C�O'��*���'Z䡎Uo���� ��j��?t��_���`��S�^aSw�ǹ���=���K��d/�T�S|kD��t�H��)��dS-��xb9�4�����hn��d,�h돈ke����V�X����:\c,��73:��p�Ns4� dt�J]�P����EH�&�ŋM�w���`�灻�WZ��u|n��˨�׼�<�w�o�^�>���%W�� V��(���V�me�rx���+ў��"Z�]_�:�dmo1����ԥ��H��y�5P{��l���(V���$(�|,�*��k���;w�4d�ޚIJ%
� $�4H2���m�Z����>G"ض8���>=����ZD{�j�f̡��A\_�.���` ��p�~_�p��+�䒝#p��o���?Қ2d� �nٯ���g��� ���\~����[MYueǩ	ͅʮ��7Kȡ /��Μ�T��X��*T�u=�Ec� [d���t���O�6D�R�ee���GP�0f���1�.'g��CS�dk)P�j4J�*3HUӛ��'������r����>���CJ��D9�=�����L��s������A��vˁ��P���@}����I^���7�]�8��q�{"��	�����L:E�m���Ŝ|j���@1cI���50��^q���E�~aL�U�� ��ч�����L�ڲ_à� D��tdY}��w^�z[-�*�SI�4Jmv���ߜŃuޢ�yY�D�j;OY,��L5����'�����h�#}~���W7ꯂ�~��s�+�:��a�XH��U��m F���$�w�����Vi���[2�m���E��-n�V�sAW7uΆ8�b�eQpQsʴ�ӑ'9����d�Y��슫����R���k�9���{�Jp?��mn��J�<w�U;����r�v��!����=���=��ˣ��Sb��X�S�ّ�6���|�Q�z�WXr�;�I��l�	�0SZgn~Xeޢǧ��`B�+������p����E����i۽�"�)at��1_��|>��&�ż=�A�h���V��������~��W1���㏏���ԡK֓
׸����k�S�M�)(���Rv/m�,#۳����DRr�bt��ۡ���,��qݘhS� ���7�ꂨJ$��Ad��c��waԠ~I��&
*���fN��/�$p',ڻ@{Cܟ�r֗9�k��X���:iQ�t�߽+�і"��-��պ������)���t��"5�Q�Z���?�i���F�����{^�����}��`��"��
ܖ����J��W�qW���I��"z�N�s�AϡH��A`n\&Tq�h*�-�ɢ�P����A�}AS>�+�.xs8}1�"�m���R�̢x#�`Q��d�VG�J�,d�3b{���U�<O�yeT�,b�it���%K��|��}
F��f͚�.7}R2˩��k4V��h�W�50�|x|`~���d����Q1��F�)��9�C5�@iU�~W�ǯd*/�)��S�}���-yQد����{�r����g�mj]������w۷��Ѕ-[~��}�p��rqפc��������t7�<v����f��g׾����z��eI߰Κo�f󎸋���-{b�:��v��M�Z�T�6�w��0saa�b��]�y�tȘ��A-�L&rh��g!�p��Qn��	��A7F�U��K4BI~Q,�B]��J �_=�����C�]r��t�*�����g/�,�/r���Ц?����o��%C�*�]2*g���i�I��0��c��Z@�<�f��%�]�=���:mᑨ�o��[��\&���*�����v�W�Gs��G��"���Ȥ�T�|����"Lt����� ���%����%FI��l�o�v��������������������>��!��b�����agJ��5()p��V��z����r�����%��	��F@?1dund!Z�O@�?y���'rh��7O�h�0����=Β?ֺ6=��V-n�<�X��zkv�5�����f,U2��/��E~o�|��� /��A�`��:�ABf���?���bwu����򿷠R8���MSuz�6o��<�� #�ȝ�m)�(謁N �?���FP�p�&a��<-�AW��Ha8��!5�w��dqw��'S�j��cZ2�_�z�����Qm���AO� [����V�6d�qe�~fx�A!�u����=�^���䋹�u��0�"��KHm9�!6'�[9�{�kVOg�����^s�a}�X� o��<��	L��ߎ\��;��/�J��B�@e�9
�����T���9�Q���x���Om�Z�0���
4��Oos���I���F��G���懭�Ofa��o�>������l�)�T�Բ_H;OE���--�4���y�{cB��;��ޣC�[����w #j��{o����_KmE0���l-�b�*����FdqE���Z%nP5�b -*�"�5��!(� ��Ⱦ�gn�������>|�sg��Y~�3g�j�,U�G؈��2KJ\�I�����$
љ�|/d��6��p���A���_��=g�d�/	��{�S��e��K���P5���.��y���B�<G�!�LL���?0��hn�2l���zp�ҧ#X��XZ�͔�at���,s����оw7����%�l�@Ǜ����T�|8�\�����Iiim�d/���l�`�ue��D�YJ�<�eXQ�
�zs�����庽�]�U�y�"h��uIOQ_"`R4�	���@����.+Ds��~s1�M�C�l�I��V�r�&���'�a��z5(i�����W'^5a�^E�*hm�����z( <P�.�S��� �% SI���[+���3_ �}B����ǫ�7N*�w������|��M���~*U�BLXM0��
�o�A�y>�%R�v� �4��o�Bz�?�key����%�d�!J�\�,�PQF t�3�R�ͮqz�a$.�|���C�LA��W~��·�U�0�bsʎ�
���t�(�#�3�f�?�#wN�L���p��e���ެ�7S��A��?G��_X����t˛������Ouva����{�6�����49�����ZA�tǷ�ѹ��C�/��� �Ff�J���+9EQsxW�e5T��<��Z'Z�Y����O&��-�B�&h8���U�Z
��",�)`��U�
_�����`�(Q��5�xK����� ��������c*p�]B�ښ�|��)����|n�Û�s筟$����u6ࡗȜ*Κ�?��'f���%�*�����d+\4N;���k�y��@�9�"��\y�M�����!�Fk*�������>xJ�Oy��MA�'����6��#JO���D��dڶ{8�B�P��BC��iI)JK[����;~���Fi���$���5�?`�z��FZ�%Nq @����	
c�H�+����$������-kT�V_G�w�D@cJ�_�	� ���C\CŞ;f*�@����������%�a��G��źl�tj�OJZ杏�6y�,�`��Ot�h�ӿ@�z�ӭw��J���M�t\�<��V_4�/�HSY�3ԊTz��,~�h��iY�8�����5W�f�旹�-�v���]� �cG��N�e��1�Q���u�FDdJ��s)�i44� yd�4^�}�ě0b�
:IR�R��p<K�҂Ȍ�EDZ�i��:Y��ƺ'�
G�����]�L��p�kx����T3�����	���xV�ۙa5���#ګ[�a9����~��I���o��p[�ۙ��;��[s�j�DK�����i#d��`[�C��\I���
��Du����1��е�)�[91�]��cNE�����~�����%z��j�~N����� ���b%l9�%�(����:��L����7>fB��vF��<m�Z�)�~�q"�U�#��l�[����$�E�k�� �~���/��?��`4��4^J�H������C:Wݣ�aN����-܃#��	�Za~v�����=��,����Є�Rz��`
���_��E鹚sHa��Iῒx���.�J�K�{j?���PYFS��f-p��˖�X%��Zb��j��0�x�po����姥�	��q���"��Ԇl6�%��ɥ��Ma'��w���f1d�����at�}>�8���4��jn�Q���/ׁF\�?���P��zo��uy$�Hq��p����տ�1��T�����Ƌ��:��3�7�C�'��#t/t��0Q���.ӹm�FUoz�����,(k=J�*�d�;]�o[<YZk������y��$��O�xvZQ�xr��//�U=M�77 ��$3��/����C����7��Xto��\�i�#x�XJ����$RAN(5䅗���@W9֢o,8I����R�#�	���
AF��0<�0y�J�����`�e��й}6�B�~O��F�??����4Z� �ƭ'''��E���# !H\�c������L�fȁ%,�s���D�F������!k�ڣi�
7S�k�L�r�t}��Ѵ��N��@���d����:�̷��c���U/��9�wIݏ�@�[�����J�:�����-������N�����<W���{�����3�S��'� 0�w�����u5�a�szF��
aǊR�+-O J<�P^%L��5@d�|h.�F� �B�j�߽FJ��5��+�]D��,�i��\)N ��hY��]����&O�����؏�M��G1i�Jm�9sc��s*U���	���,�r�&�T_�P��uI�sV��>q���|l�:�]Q�� ,#gY���@��H{��>p`��	+B�3�:�_)}�@���?]�
�N��gx�OP�p�o��8���uOq�~Ϙ��'^��ƲB�����k{�� ��ܒ\������
��q�>\�b�Rֆ�)������8S�����ny>Iվ$'�c=sgS�t�*_�nGA��-�T,���a���y�ia6�H�j8pv�0\ ذm��5G?~{U�P�&O����*/H��P�eN�7g�����AM��UL@4�����T��~���e����gLr6�*����ڼ��7��##�^W~JJv����я�����:m��@;|n���e+�-���R�s���u'���	�V ���+�R횆&ԙG�7E���@����:UD�h.�.�U��u%��u��T1�nO	«�@ݶ�miɶp��AE K#m��Lۂ�_9$$&��Fvac��h����`K���HW���-���[a�#� ��:��O�1+��)p��ޥ�iН�B#a=�'�_և#kJ�����0T��1�GP��O��r��heKK��H���EKܽƩ�������"^���O��P"�Z+:�G.E��X.U��c��h_i*T�t�ۆ���	�w��d�>�ˡoy���Wz���a+AY� ���zm��B�����@�5�u>�;�K����~��>�����W¢
{�7���*�N���"�?���	�jHt!��3FlЯQ�bԜ��_�#8,��ڒ2��Q��T���S!oe�p�=}3K�/(	���������s�����84aq��c���W���KZZqN���R0�zT9�벗����o�
��Lx����N�es��0/�a��H��T��u�Ww�M)D�z2ۈp�t�R_����ut>]1��	�]���x���:@ٞ��Y+��v���֞E8���T�쩇��RZ�>t�xG�@I�!2��2�i��� �T��	��5�����*vŧ���lR�����_�ׇL����&��	��!F_����b�����j��x�3w���EO��V1F�j�S�Z���7n�(�Z!�D�ywQ)lAs�2�8�yd��W�㠵u�	��V� �K���ؠ�hz�>؁q����y��r����ͭ'�^�����g׌�_eݏ謻bȰ.p{�NrK>��>�Up�~����H�n��
���`��x	GN��A����=���MF�<�����*lIq.�
�E�¯β+�
�N�
�U\|hδ��n!���X��A�����MKGpS^����a��W�Ix������k1� =}��N+�A���1��ZvK9r�t�z�9Z�Z�5�}���)}:`�1�Ϲ�ynu$�k3�(_Mp�1�7���A���
�ow���HX���T��
I3��S����n�KI����?��I�u��S�j u�a�:�Go�_bX�Ù2#�c�L5]R3��6�+i�� �۸}��d6~%C�_���6�7���"���$E鵣Rlׂ�_T���e���VI�!�L.��-i�R�T�E�:��vzn>���*%���k�	�L��a���S�ߜ����]@��?�q���!2�Z����:�����k��p�2]py�4矌E�]�#����g���w����&�2�)��� �㑩����Hjծ�
l!i(	>��i�B*<ٜ/e����c�����L&7�� �������v��GE�PįD��ې��P���&S"SNV�T�5�C��+Ο?p��]x�K ��v\MA�\��7�n.A���0�zG�IC��t�N����i����>�o �4�G��f�RW]��̺њ�?ȱ:]�P�|��#��}c��"��`�U��"]zq���gU�$H݌�ᗷw��:�o �s�0����C@q:@q{a����$�$���O�:��G�cG�� O~���F���s_@waN���s����K�q)��b��N�K6hh̓)}���d�5��������9��+d�lt0���ѿh����__���X��%���c��yhUL�TL����!xᾬ��"���D��-���U�:�U�Y � /��|�ε��0���s�־xQ�Uu6�=��d� m��$�٢mfț��p��ij"W�����i��3Q3��5[���#ȼ��fleW�͔ ��G^�O	���#2]��+3�VI�|�<����;�����t:��(����,��6�L3"s�j�y\�vR�*KKZ�����g;�r�J����BU�Q��:+t�Xʮl��y��}�y���"UġC�L�d��E��#ҏz�6Z�g�����|��+��2q&.�Q� G�8č(poq6�%&�����!l��[�^�)D�!����ǀ�����s^sV�����P�?��:�w�?u��w3�G�v�g��g��>�ڬ��K���c)��<x��2�R{���>�}���]�����<ty,H$�^�K�5E��(�O��:��]G׹�sl&%F�2��dNh�3nXN'�����>|�K7��IDf�+���@s~*=��ت���(�F�5����m�k����ܐ�"��JK[gEq2b�	�W|;55�'s�[�0[mf|@�G^�1J_[�c`�aii�7En���J�XMH5b�
^� .�)2��z	���Y<Q��1Q�$�CS�Sm�p���/��@�(D��ʹ}j~f�Y��䃏��"�CX^�Ծ��y�'�z���$*>��O=tt���Z(U�C��s�aj�\���4a�v%���~l�M��#��9���ĨS��^r�U��o#3pQ�_P�t�R̈�u/Q؅��ܱ����X��<yc����:S���G:�ό��q@1��g���#�Z�Pw;n��7=�O�aA�ߨڒ��02D7�ā�-�5�:�X��vs�>��7N����5�"W�|/�A���"O�����2��	P� X���0���*�x��,~�(P�"��{Py]xF��#�9�,����j@�����j�G�o1��H���?f�W���C�8���wp!1����dv�䩇�t�w���F���y��4�G�����3�>����!k�����p��,m5`�v��ֽ��u%�vq�l��-���*o{qO���+��!zGM�d���9t;'��Eq���`�O�9�$fR�?�F�u�_�N�f�]0�;f��>� 
���x��)x���҉��:+h��d����m6�?��e�m_�&�����N��3�0��R���.]j��&����eSw9B6�������~cV_*,y�g���ǖ2fs�{Vd����n.����B����
�ܐF+�O�R ��������r}RQQQ@#�,Ȥm�����\jj�Y-_hQ����݌Z�h8�@k���0w��.���7��=�Z_dA�ŗ+������"�/MjYa��;��x�xkmo�~ b�pp/�5	�f㣴Ɉ��0���:tmqv�����1��0��h&(-&%�����|�
�����d�'i�c���r=)��F�ϛw}1��ʆ���w�9�ȧ�52�\D�۷,8�[s��r��N�t�*�[�����آ�^hq��g�:Ue���q�$�ׂ�̱�B�Nq�&�ԍ���m��K��R�����q�B��2Bn��(��~7E��Ǿ^;H�#9��5��� �!�����G,�o 2�C�Mք�t�� -�P�YX�'pst2!���HXf�H�2��BZ��:��J�y&z�	D�C��a�v��wԪ���("i���}_�3@y�!Z��U��}Y©�3ؼ;�ݹb��@��O�Hl�P35��;�uB{�.8��k�����%9�zn��)��;Kkǭx�}��d�ڤ���i��+ԯT����'Z՞�N�S�U�'хQ�q�wbƤ���^���w�2��u��ՂO��/����7� �>h�H��}Լ
����!�Iۆ�X�IŢte�	���Cǜͼ�;((�t���f,JeG�eg��z�ѳ�4'2�<t�t�)�b���y�^���9֯�1dM��k�����;Od�#��;�r�F�K�	Up8/�n"-'�kdzs��࠳���:A�����/�0�#h�O>' yn���_1B?UU(&��(��>v<�::�d�^4�1���#\J���Qɼh�?]SC��+��a6������2��6lHh��eY��Jc&��~�ĤLIQf�J���fO����U�ͥ�z��>�c�����]�ni��D��1�[�$CÊ<�g��N������	�}���nb�~j�RQl��j�Ym���g�D:'�W�_GP�5��*\��r�XDۖ��V ����ZnZ�S-Ǘ_�BQ&��D�n���ѣG�����hM��1Q�$ra�!ɘ�L�<m���Uy�S�8��L�Jc�`�R`qϡë_a?��q�#�e�-į��;V��J�8c�ApyL���}�s��=�����T���K�AF��T��o��,B�c���:��/�6A�v�	���y�A�=~|Bq�@B�Z���<4!+"��7sni�{F���|K.L��!2W�qFd��ʹ�t���V�B����<�ˎ[K�����a{�?ǁ�ި�Q!*j��]�<Td������-uw�`P�c���v�����gg�����})9������m�@.�����4��*B��%XEp@��� ���S�� 9X��a]����{XQ&���E.ǢߩcQ�#������Ӿ��^��n\��♰��P���%l޼Y��0��Y�F0���Y��qk�b�k�[�^9j�@G-ѽ�e��YA/Qŧ��}D,^�x��܏�dkFj���>��s���F�"�ᔂ?]5��0��Y;���1�$�1��VO��M�qrs�́XB`�C�PtS���"����,Q�J%�y���ϫ:z?ۗ|��\�~��I�WM��R���x�%0�C�)m����8�/Ļ�&_����A*����+UGC���YS\!b�xV�<'��c��Cɑ��16kn8�9�W	>�O��{��6�1_���4��%���;�W�d�KVڦh`��Aw���Ͷ���M��k������b��7JDG�w��nCOF��n��F^Tc> *8&�+�6�~Z305#�<���#�M|v�cG���#j������F�K�ڡDG��� �R,dq[�T��{M��kY�X��gi#��=�ZRd�C�
����8��K">�� uW�� PJ�}�s����5�R��B���R��l���D�:��W �c��/AK�ɓL	l�!��!T�x�s��ߞ����Ƭ'D�a�5n���5!�9�H��Z+Jj���]��{NKH��0���G:L�}����b�`�3���Yv�B�v�M�O�/I5a� Mi,�u2?7S@�>�^�Ss3�0|
�}�g�$�&f�b%C��t0['6���+���72���R�J�f�����+,�/�  ��d�Z--��J���oI����]��x��)w���l�0F�xE�_y�ou�h�N@��< X*o����k�9Ŗ�"��5��h� �8��ߡkT��S���G7���[M�+������E����#o7P��3I�������� Z����we����+�~f���z��^�Ύ�iALX!�z�Df���g��)�����x94�c�6U}t՗��8��G�*�ɔ���'c�.A�7]Ó�>�(�_)_!k[�ޚ�3�'�$�����`-n�Ӡr�B�-�`m�$?����}�60p5��7�OK��!`*$�g�w�gW|ς�P[�O|�������^����]��˧�r�!����w_�*��X����!��7�抝�Xw����1oZ��;��+�ě��;HX��w˯Y?���Ժ�xqz9OVC=��n��~ۆ�������acI�Ky�5��i�'ȓ_`;�r1���CuJ���O�����_�?#-����2A����XKپ�����N3���g�ۼn����� -�T�����h7�ZR4iK�D� &qqq�(�AǓ�)&Z|��ӆ���>�Q1�����xG�:�Re�~�e�3��8+��W�L�q`Mh++iv��p@ŦM���v���u?&?g͙��L��&_�e��ʛ�Hq^)�V�B��s�z_����l�`s������\�Eb�C���3&=���M5���~S�xn/wl��0r��>>';#o$9Hx��f�=��z��Ǉ�x�`��`Q
�U�2u�^ץ�i�?��0�`?ڡL(��K�� ]�=>_������b,Gp�N$�y5���d����J]��Xs�.���*�ȇ$��Ǻ�٨����z�!-)Vp�ӶN@��:B��fٖ���-/T�̲�q,h�D�"+���{�����?�&Ѱ3� ��ƶ�-���'5�(�H`�*���� dNE�w����C͕+Wdci��63�(	C{�ÿ�5G�pHT��4�:"�2�?C�IM|Ǫ����Gl6�+"� A����߿�n�i�U$}��M��lV�s�������`; ��|�H��i�w�
�,�re���#�q���y�lR�!U ���o_PZ�$Q?d�xٓ?�3I�1F.�q��N��=��kI�5q��l��d��uF�hץ�����\�����w�LE˪�oQ�^�
�"%� �,���݉�ͭ�99Y�I.~%~��LDʱB="�Ž���Q�5xj�3��l��Gy�/1As���_�L�e��WG4��;뵥T;��z�U~ ۞>������>~��k����E�N^s������L�7ջ�x��ѽy�'�On�4�]E�:��*���q��)"�҄}�B�  �+L5J�V����	��0�ӧ�=����+3�o��ֿ�0܍���2���?a�M��h��f���c�e�:f#�b#i|�׶�{A��O]Q� ��F�������fd��B>�Ȭ�"-��.���lMKZ�=9S»!�%�y���h�(&���T
��F24G�����������S���<��z��*%����v��'�	��ؽe�昣�7g���7�a�E�]����۷Oyaq��wϞ=+�T;�l*[!�b0�GF�~_�4u��IF���
�w�>�H�U<�1b%��՘Co�KL��n��S�k����ׯ_G#��&������א�OT�4�u6�̕�n��9�6�����kA�_8��>ĸ.�����}��]u2[���S���I@���߳�@_��##�}Nj��t�Z/��(���1�<@�UU�蜼�:pḮ�K����m��q#6^�df��! ]@'|C$���ŧ6l:�Fzt�7�>گ��j&1���RtQ�V�%E
U ��G�0��$ �_~�҇��9jC(�w�5�uG�����ESx<2Y�P����L�mfc��|���	F|�[���f�:��W�W�v�i�3��{DZY����_��!���b�nĩl�8[G8u�)9Hd���$|�X_Ld��5�w��e�z�g��':c_`�א�8h(m\k{\���B���� ���O/�t�����uՏ�)a� �re�tG�)ҏ��*L���/�䉕j��uDTk�P��A�U�F%	Z�,ɳk�w��7�*�g�٬�y�FVlS�;KZÏp��T3�`G�b�M�� 5�`�z���㧆��*�Dv�VR|J<�0oko�{��ix����\�pd�SK�Oy ���IJ�v���fh^�Ax�7G�l�E	���m�(~�D�9�1�O����q�&'�y~?y����]�o1�/�9\��{m���X/�����
o%��똾��ܐ@��b��%��)k;-pa;�d����MMF���x彏\�7,Ϟu��?Ocb���k;��C�߳���r�/&\�%��js���J���ǝ�<4Dz���Uv��`�[���C�� �C�w�� f�������3��[w��T������	?�E,K���}u�)�ba�6��kTˑ����6�̅�5y�K�	o�c��敿��g�,,+|��/����(�7}O���T�{AH��0:��jjj�J�|���[17���3��xVt��e�����&{Y�#��P��Ç;���5y��݌��<W.�h����Z<
ߝ�+���r��|��Go޼��xaZϑ�bhK�5�3�u�N������=|f`3���͙u��K���#~��y�6#+������,�H�^� ,j����l��������L��F��)��ź�������c=����*rm[*7�,(kA#(�QU�w/�8(���@s��5��Kz��f�'`���y�����%Q�HgNZ�G�t���\��1K�O�+E����~?t~�Z�E�󘻇T� D�A�a6���Q:��=��7�P��CKQ3�f�&5��Gv�{A�C��F���8W��dfb�"O�g��dh�Px�&�_p�fI��(�K������OΘ�K�L�>�S����b;p3Bw�'1�Z�(�)n�p�M�A�/;��(k.�{�3�=g:����V���5���Th�HS��IG��GoN�3R*��-u��݋�I�p�=:��l��{��w�o)9�˙zE�Bz�ҟ���q��{���<z*����2�`�'[�'�K����0�A,g��u�N��T���ۻ�0�B�c�\w?4�R�/�Lߚ�y67����]D�Oh3o]뽕С���3�^g[��_/��������?�a�� �{ʊ��w&O�*j >8���K��N�S��K��)F@����7v�0�߼�ڎ��^�ۗ�wB��y?P�=��/N��ƱMO+��9��A�~#�Q�<�ECA�e.�2ؕ3E��c��G��)+���I�7g<�15iI�� ѧ��Ҩy
�l����Ѓ���"��m�C%�F�������ܼ<×ݺ�n���aA�0����^v�U���r���o�2֋n��84~0�կ�J��wc��r�'ڶ\0���#��NT�����lF+�H�7T/���15a<&�Zߒ�f6V �1_��+R�˷�HA�����4$2�̝��VV]x�
�>G+D��G[@'��m!��ǂ沵���W�Mܹ����.�Y�<�7g3\yPy{Oz�<E䗱����>D�R�Nt�O��3�S���O��&1�A�ɳU��4 ߭$�ALv, ���`bĮ9mM'�NI���V����'�9�xsTn0��Q�^�_F�<(3-�j��ߛq��Z?&���)[�j'��4�	����رG>tγI��#��ު�����r`8*\�b�RB�al.IN�s3T�ο#x���M���vr�ɴ���ݰv��������No���	��_�/�{G�ME�,�����t-f�������5��k�k�ޞ�o!���)ATj����iu�f�ծU��Dr�ģ��Y��B���,��������cmj�K�f��.�z<q��yݒvK�����.��uVRd1���8��q#l�R�6�3u����v*{������D�;.9wUWk*�ם�w̰UlH�Jf��?�&~'�v
��+(�[U�CO���7 �e����7C\�zdlܨ�hN���N2p �Qi�юD�i&GFN&��[XV�KA����#m�@�[
�*�h�h�ͪ��%-��(:�� x���](/ΊX��ď�E��J�'_�z)k>;yb���A��q0���s��
J{��$�l/'AOs�*�Ѩ��2���͙� �E���K���6���8���$&@�U��=70�S&��ޘ��!]6��g����q{k�B����u=��\,�w%~���ܵ��^lS�/=�PuOm���v����=����{n��
&�ށ;�.����-�3�W	�zH��Ĳ������^ւ��"�IV�ָ�7k��$Mp�(�xlj}x!�m�*���Ϟ���YK��vZ�)�GWWWk~@�5����C�?���@��Fj��6o߹�PSC��PUY�B.y��T��0q��l��7�5U�,*������n�ag�&�!��������m�Ő���8����֪ܼ~=Ѝ\�6�<)N�^OWծ�-���cX���#U/�R�c�+�D�G��\����T�:sj'q�I x-��$��=�TWW�l��X��|S8,j'Dc#"�1L}l����I/$�<�Ƃw:H`����
O��9�sZ��<��r[���q��i�\���x��-ĳ}bi��?Ԃ�}?�Nv ,��CE_T�M@LJ��`�%��MH�޲+��ߢ�Q~�
T7L�9Z��xq>n@fLd�����֓���e<�,�Sq�U������K`�Vv܅ͼ��5�Qmy�����B!:@�v��i�� �%�W�x�Xj�v���*r�0b=�����ק��t6n��'��/�pB`Js�1z�mqU;�.+��rZZ���\ɭ��4���%�~�HC�=\���l��r����x��%�v�S��p�G��=��Jb� �S�e�'��~H�8�֎.i'��_q"�d�����F��=�S˹l��ޑ����Q�����4a'��r��cݫN���z"�B���.�o��+�c���7��<�ס�?,�8�Փ�C8��K�� �Q��c$9�&^K#���	,'�g;�[�(��V���EShim�������-�)46���sa��vf��)D�#I��u$���$�~	�t3�V�K^��b�LD��Wp�L��*���S*�\�~���dp�v0-��4��� �\~;0nҥ�P�F���
�[�n%�s�B�T	�.	,�7����fM�a"7d��W 1z!Ъ�W?t�)�&����玠�|�}���ld�!��3p� �#O��:��.9X__o�@����<Y�a�+��3�Y|�1�旧�!���[
p�R����Ƶy`�/�}~vA��D��6���z�33v�^wez��Y�5wLsQ'.[R�>�7W,�����$ܡKz���)�s4~%��-S�L&S��[מ�lm=R���ڶ�]�y�H-���S���K�@����\�.��@7���-В���m,U�e�������e-K�l�2�o{!�I�ٳg���z���z�	��T;޴X��wU��04��;�I~�����*M���*�Q:�ֵ� I�e��ھ1v9��a?ul�8kn�a�m��DZ�!�u�y#�WgC�¾(��,88�̛>��Gq���K�D��c�)q�ϢйN���7y�a/��o11��1� ��D%t;�m������p}7+�	%=������,�ʛ����<����t<����.�sr���T�fG�t�P&č3�����I,|����Y
6��І�5�ǔ��N'Q N���#Ʋ+U�Fy@1�f�}u�wѫ���]U)���X�MnIE�
Z[�c�/�k��闬����ݻw#cD���@�Z~婭�!;��Ű�r{j�t��Al����r,��16@7$�����7q�;�
\�/��Ѭ�H�.y{��E@g�G�M�X�겗����t@����0���p�1,�w�k/�b�vv�
9B6.�GbIލ�U��F����$�J�D��b��Ɂy�&ѧ�rN3�'Ķ|عUײ�D�������@q������)�ě�A�S}KZ͆^p�A ����7��1�o@�.l���,9�Rߗ1\�*�z9�ߡ+��q��(/,�d�&�(Kc�������g,�-��n�w�F��|���3���؊c��5�_��q��k틆�¤��C`&:�������5�����*�$��s�Z�x��BO�wɛ�,�*��]�>���[N�gk���UV߷ۘ�X��ly.~�H��Y,[�u~�:����ٮ�!-]?�Ə�|9��9�)���y�5�&�F�kO�|�2������酱�Xg������Nz��ʔ�Tl&t� ~�0��X&���xs�����nB��vY��O�0��U�����8�猫>�Ϡ�ȓ�Ad�w�~k<KE��Hd��%_������-���N��.j�kk�e��V�[qz�NB>�1�Mx���DIY��=He۟-�rj�2���7A#�D!\<J�v�p�'OD���C
$��{O८���2�%��7M"�.[�n�h��V�z��c���Yb�	x�?h��H���a�%�L���m��NjR0_��P�E!L'���\�,^��A�cOI�(>H�
�8��aMg�ys,�>����~;n�p�9��H�=Ԇ�^�A�!�9�G����� ��P�՞��@I^J���lgpx��C��8*��	Y��C�R,�a�?~�x �4�{d �����,��;k{��]�2t�Ba�n�h���Yj�J���4s�W�"�ը�guX���	+*cU"\u�r΂n%��J��/�0����_����F���_��w����u�I����i�v�A�܇+���b�m/��[�X��1[����YL�[5sQ��PMu~*��sR�mf�M1�Ď5����큘a���� ���@��zU���p����
s:�m��';�f�lN�����i-@;y;�B`����]�fo#+�J%C�Y��iac���+����K�bͬL�P�_��o)!2S���b���6�B���`ᄛ7g��'�s(�5�{4�_�H	����3�a@;8S[�ݴ/��+ �&�l���I��t�F������{D�/-��^ԛa�-[�� !�R�Ap�ͦ-�9n���2؅�Z2[���xT�_�x�hA���3o�l� kS}spPrb�>d��j�}]�x�?�KΠ�^�����G��%&������
��!�U��s!5�y~�j8�,=�qi���'0H*y{N��uܛ�P�߾v�AAqVvi�x�:[�&������مm�"r�g3gۑ|��k�[R��|}C�,�lb��9�qP��u3�Z<���t�%�"�����\��/ֈ=H�FP���-^�3)V�f�
	��צD;{8D9��V�@���E�ü�ʰ�պls��d�a�ϙAP�4D���7'��n�KǼUH�R�e0��k�gmQٴ��5-��Ӷy,߂i=*/��S�yj�"Yhz�r �>����:�0����Nb(�5y��OR���d��*�b7�P�6�Q�����C!��
���7ޒ��w�| �C�z8��ա	��������A��,�R3K����.�,;��;��-H�u��=�I�5k�4� d �ȱݢ���/��ЋJ-��\���j?Wqnx��˒Ƚ��(��=S��{ �މ>X3�)�dE5ʡ�v.��Y���Va�جP�;��Cf{ O���̲A�G��h�Bn��=mf -�>R��䰊����$��C��]��X����@��w;;���՗`-굫I<'�w�\�w��})�l��	l����S��,�J�ld�քJ�%���#����1��,��:�eb���f�	ÕH�{��ڂR���SCհE�%�eb���3�>���ϑ��FLHC��l���é���!&%,T����#RҬ����%�->���"��֪�oaֱ�>=��ehG�ai�2��v[C֒`=�̂D��K�ڃm=!g��ܛ[��a�q�W�K�1�<)�� ;��o4#ZA@�ӈ4�Nt�.�T 5���v7�Z~�n_��8��ff'U��޽{w�||�C�%=M�Os�=WY�Q �;��p��*ȐëH�U��}�&�e0���ŭ��Wܡz���R��X�[*�^�����m:�r��G��yM 
"MI<too��/|�Yb�^'+��&�ƛ]�gu�b�7����2P�}��r��p�T�ٗ!��VRZj������w�d���$[՘�us�~����X?0��^���/����7nd���ev{}W�D��*�"�'X�B�F�r��kf���z�D�b��k�Gw���gv9|�q81��`f��h��h
E;���K������N:�VUU5#S!�MwƤ�e	*	��[���t3 �C�iB�Sv��;��)帾�1Q`�){U�5�ւ��3�`�,�;tsO�7K1�~K�GI���D�8[�����tU���Y�c��%�*�<F��$	�!��l-�;'BA�����܈�F"����#|�c�h#��ݴ���l,��pћ������=����7�Yr�..��qէO�\�:Q1�c�7�}!�}�q�  ���}&�yP���Q�ekU��'�`��)�,1J�ꤢM���#9�F��y4�:��lKk��z`{�]Ix�XwYkmml���CQ�9�a�Ო2K"�l.����:1��Z��T��1��SCʅ*�<uUS�ec�����t�3���!?�{�n�G|f2����ě�_t^]��gW��fT��)����U�R�XJ���c��f��V�2`D[�w��P�� G(�v�l�K%���Y�1�6
�t�'-.v�?Y�v
�=�uߛP�S�?\By���C���~̦�d��G��e�5�G�W|ڂx�鴦�s_��K⥣��?	��Z�4h �a���|�}�>���<9$�zc6�=d������j%������%���P[kfZ?S���Q�?��Jh��,��[���|�I�rh�Ɓ�Ȅ����Y�tD-pf��\~�6��MnC޲��X����2/��:���rzO�?���D����;�/~8�c�޷���B.o)���(���������}�8�I)��底*�������q���R/,��������+�/fC��:��s؋�Ʒw-�O$�T�4��h.,��iyY�яkzū1rb�bxI���WzX�UG����@nl/�w�kM�X/��y�6tͲ�?0�p�W��n�_�^�⌸����E�FK"�v���\�6ydggW�닂�#AZ�)1�ֶ�kl������X_e'F̷-����M7�)D�!����ٗv�X�G^�ûV��Dol2Q7gf��;��`+ۘQ!�~D�o��6I�]��=��g����0[냙y���*k��g�m\�+�ޙC3N~5��6�r?�O�us���bۼ:Ͽ���o<��t�n֧T����a9����E���X]]}���z*Q������I7�������Q1��$v'�1n�Sq��l[☝�X��-v�w�[o(ě����I�L@n�����
U��Nu����Ʒj�')�/��z.�v��(���R6��gۖ�:����e�c�k���̓&C��S�gD��e:�R�yS�d���aas��b)�Ĵ]���مY���vT佰,��'O�4N�k���:U�����^�����y�<�rN���؇������{��1�M"2L"�ah���+��"g�)HK��-/�\@0ܧ ����-�UG?U�R ���ߦ���������S�~A��	÷���YlX�k�˨$�2�lT����~��s[hZ޸/ҟS�MΙs���?�)�J��F?_�m���14�O���$��/��J4�͵r�{����9�7==��2^O ��rm�°G�`�y�o��b�+7n�:a�9�Ӳ�z^��L�C̢�>,�<U���=�z���o�d�+���YVo�S�6��|}�6y���Z��ktnX>O�%�n3;��8m�׸rQ��r����(Se`/����~ �a�R�"�
���n[>?�����O�<�v�^�hu���Ѿz��`8�Sj ��mll�O}��IY|e"s7(��(ϋG m��?[��ڧO�Vg橋iy��V*YG����z�`/�`�:������կ��)~�a�g�kl3�#e��+&�5�?�{]���4��T����5i=��{4�����@p���2������%=�Ez��g�c�]4��ٍ�Ѡ��e��)co�R���-�~X��C��;�:7F'�E�׹�/#o���n�l�ZԞgG\]�VLz �z�pի�_�v�$�9cb�f�C�LF��p�2�����ބUS�866�K���"�2x�4�~�i�ymch�zrQ�Ϝ�W��k䐇�[hA��5<�&�����z�qi���pܢD����̤/��9��?k���%ej�n�
��h��bQ�gm\e�_h}S�2����&]FeD�?5�����?��i�����+h�o7�`�<��W��V�`\��.X �Oo�Mzۗ�
h���E@���;00�N!� R���gU�puum����T�����4��0z�OC��z���o)a˻��S��1zy:U�Nm��!�.Z�hmk@����3hJ�hJ�����
|H̑��^�f������-�Bw�g?+J���C��VxY+�;���#٨�WQ9��j�'B�ҽ5л���$�*�%Y���cJ�D*��$��u@�o�Yi�)�|�Qa���,��b����&�*�,�Sm���EC���?bE�x�����I����@� f�`c.q��9X䲰�ۍo)D���X�h���^������>��ؒ��/�-j�x��5�?X
{Yk�Tq?���k����@K� ������� �k&�tǎ/N��LȞ�| z��p�ݢ�]�L~�;`��k�9��U��?F�z�G��_�J���E=y���4�)�E%蹬�Ud�w09��D�ٴ�&FA//�$��f�%&xA��`�FR��ar�H@;�~�Z�8����l�%���������m��#��
߈�>�yg�e	F~Tﳵ1���mh�ݨ{Vl���WL�s�b�?��%�����o��Y�$��Z���_E�}�G"����o���~v|��.������_����]����u��M�ǿ�+ǰ�tP-��?f�����y��ù���̼f��7Z�m����,��1����_c����]33ή���GI)v��)���?��y~���+m3��Ϡ�:�f˵���^��CZ,�{���0;,{-���p��Mn}��g����f�}�[�zD��l=�/.�:�._��[\GL�ՠS�<jv���-���	�K���^�U�d�ګ���W��\�v$�{B�@y���ӱP�ս��nª6��\��	���%�~݃�D�}ՄA]�踸o��=�b���_�y��ZkZ�ð3'7w/�p�~������ޯ��v�^\��L���a�����
H�j��:-H��Btiv�k�X�TK��+Q�:����7��ޝT�Y����Q��|_̏z-�ݿY>j�@ݠ:���O=H���:���v��� =N����M[�0�;�-<�nݻWWu����ph���zOj�Z�]A^�{�J�!=�/׼ ���ֶ�����\����]�E�z�_��(�S����r�V.pvj�\[�v���O��KB�7��Q�a)��o��2�ʾ�Z���Ũݶ�`��� S�^{]�Z}љ�#�F�k�Fâ�t��RPG>�����Ӡc9����T�_�
JUo�^�)'����_`��Wr���Dff���`��f�����}�]w�Fłba�Z�x'���Ps�^�Ut=
�'=\a�MU,�;_�_.G��/���&�k������)�	 PK   ��OX��g  n  /   images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.png�xUP�u��{�;�)�AZ����C�I)�-����8��P��+�{���tw��Μ93�pfv�,B��*�  ԠJ��&��q��un���j�	 0�����z�Hj/�w^z��^�V6 ___>GOk+7>W��S) ��AMI^�/�$���Ġu����������1�6�b���w ����(:��9�A�B`hz/�抉���T�K����%U�0�2!54����+|������#�lI�)���ŶE��V�c����m+�h�@.�����9UF�*o�@��Qt&��t�t�DA:2�L��K�H�e0�j8"0��h�����A�a��/�b�V�D�o��휞�H���l	}� }L�~���>��t����|f?�Y�����0)�){��`��o5����1�䩩��-��&�{�6�P��54v�J*c�?Ν/�yޣ���;_�����WF��� �z����ܻ���1)�?�n��9[��j��U�Ҫ|[;9�K:�D"�m�R����7 쟟[�ެ�68��<Sic�"�lM��ljn6b:m�&L��}�pj�������\����ֶJ�U5�tޢL���n�l�)�ox;nx�TY �J��y�I�@��y?E�ʯ���zZ�Ҍ�w�;��T)�?'Q�63�������W��:�@��e���4�R�I`��V��ʿ׋[��^��FS��'kc��������k����$C��7HY�T���H�"n���v+k)6���2�& �gg���;�>=�y������SAJP��f,����ׯZ�:஀[�?�q���Ǚ�UGtY
~s��^�F)O�\��Ý.�`{��3��b�$�[��H�:/7(���D��Y4�zV����;�r�w�Jtw��t��iYuI��>~ɺ��%�^4%����o}�͊��!b���k����PP�N�˺���y^�i���	?	�<��횇
���<疗9ϺN�s���Y�S�nF��r4J[���松>���]!faU����3�:ːG�q_�
���?�君���g��fٮ��v*�	���P�������)��Wic1�&��
�*�QB�#}�,���Jt��Ut6�c�Y�RY����m7�dgF����w�9f`z~���������4�)�n2~��m������遡`W���g'�x���!���+�y��Dx���/ǚ솎q��0�ط��S�<�+�/@� J��,jnn6�FB�YW�1�z���0i��,[����zUiQ;�D���ϽL���HN[��|o�����\m���UU����@�Q�������g�3Y@�/���Xޏ�w;�s�n�%߷�WtMfI�0�c�IUr�{��K�����a�u:S�a�n|�IY��ARĈՈ�:� ����;4�JMP�64���g �6\]a~��u��E��5M�e)����N;�Y���@̬�{V��ɫd}<,�� rp��!wL]ה��V��`�|��L&�E��LJSKy� ��V�;/�w#����(�.��o�L*��P�,���L��f���n*��/f����k�M��C�I��V�{��f�9��e��x�Wڜ{A���S�z�}������:L��3�DR���5s���l��x9�o!�b��9�!��9�����ӖJ#v�2w48SݷwӤ�Y��VL�kR��NX�I��w�L��/�����}��ͧ���^��hx��x��|Ԗ�+�鳵�	��H|:Cu��*Z��j?|8c�{�|N�1)���.LCCSu����L���(���(]�:��@-�/!�7�?�X��M�-�p�.Jjߺ$�s/ls͂��Eg��L�8�:�?���{t	)�|��V�~ܟ�����n��Lu	�gAOB�����Դ��>
�g���xԂ屙�WȖ ��#�!��{�8ğ]�7�F�G}^���8�xڎV+/��f�}�X��}�,�<cj{h,j���~f��gi��Z�陟�`�c@�3��8���`̂܇�7�7+R)wQ6����"z���:�*��F��7�|l���nI�o;u	%�_�ۛ�?>܃�Ѩ&~�	 ��:#K��6
n�F���4epftg��(���Қe��M�o�#�a��%�:$�O(���SH\'dn��DN�O�)�Y��"<����?c�Ǫ���	Y��;���ª;�lH(�)x[t"�"G��<��㬖�r®�k0�&�`��C.�"0��<e���a��@�^�c��",N<�s�9q x���f�\WOL�F����j�&l�f� �����0����=�����	�@L�6Y�Ed��Cy]���N��5?'?_���Y�q|N!u�ʜ�s��u�N`}���$~��g��^�z�qr	J^b�e�T���ouVT6 R �zynZ�e���ۅ(�0���ȗ�<Y�/�hm�K6`ϓ'�L4a4��{�щO����������"�M��8�;>������m+2/�O������2xS_:x���S���P��A$�޳�l�ϞY�(���5��l���M�'ק*������w�}�����Zq(㪯��ϣ�,�݄1��-����E�w�>�k�O��$ܗC�@x�j�]��O��'N�TY���"\���Q��K�iJ�y��1��欎|��q��b�ӽ�#W��T�Q��ݪ�6�E�#g}v�\|)&�Π��!��S�y���k��i�$��f�*����˫"T]P2 Ȧ��$-t8�j�QG �7��XV��#�{��L�v�&g|�|�;I�Q+>T�f�b�+��s.�	�]t�ۃ�cm]N�û8��z���׈0=XX���8l����=�]��x9��^$9�m��r��/���Ɗ(Nwn��X���Ea��z/�ejǫy&�G�A�1��u^�U���e�Rv��	A���L$��t���k󴊧b`�x�`�`m�c�[m|�q����%�`���tl&i��{CwC�W���v��3zB��/�0
�}���j�FχY�e��QeUNh/�e�违:����y��',�[`�Є���l�#�w�-ܳ�ע�yRx�DE�����.B��l<զ�	�b(Ι�O���5i�K��Վ���R�'C�2��Ut��v���R-�U���H��Sh��W�\h�a3Kf"!N�PyMlOB��	��ɦ��T~��p����&��.��`�|S�����YP�H9B��7���'67���!�2RT��l�K>P�����F۞)/���� y�I���I� ݺ�
혷7������v���4��YH��V~8�(�y�E�l#� ߄ϲ�̲�'7@�eV�M �:P�����D���U9&��*(h���p��`�V������Z��ڎ@����Wu���T�xhT� � �ɣ����w|��n�X����7��`���PI�l�� ���}�wd��.�Dj�z�P�1�sB���E�!w���Q�(�����z�Y���H��-S+����D�Gb1N;h	���4A���	��73o��Z/	[)*�PV�"6ӱ1S�$RϠV�+��_��A�>��2;DU�l��
r'F����m��;d�7V�+�YW�H����4��5K�/���z:©��/ؐ�O��n�w���f�eD��<}�?�Ҽ��_)��dz����"��Y(v�+cZ%,�`�UH��(4���ٯ�P�e�+�靑A*&�4Xf�%�#��#�(�C Tq�j�YSu*r.������K�<>5W179>G��gf^~�Xݹ��������.+Ը�.��� �	Y&Ic0mu�]��;LlV���ֆ]2a.�|�K�FE[o=�a4�X85�=�%�P����V/AK�Ndb$���
���(2�R��t�b������ޜ��R�~�kbs�ۦ�]�{��&S��Rk\B\c��#��o��x��cK�\ۖ�1̥܊ou��p�rZȠ�xu	焝��9ȟާ�F��|nG|Wo�bhp�Y��`��sb+����IK�h�=�6{Ǚ:_���������ߍ����B�"@sMGK:�`P�Q��Ls��A,p|��{'�ڤW�/D?EWp�c��؊�o9M��
��M�'�c�{y�z��e�#�F�l<�B��]O��%۰O%��<r�e5C�f_��!>�ν���g��_��/gL��f�#�EgN()-#\$�\�Y���DB>'d�f��d?���@4�7h�
ǉ9���x�5�������:V19q���WxQ $���%��56��	�2��ea$�E����Ғ	�tlRh��`	d-f�Ԓu���:&�h�S�3��я.˨��v�ٜ���j$cT��	�$7~U4��Βy���&��=���Y��!1b({�o��rz3Pǌ�:֦�<G4�R<E�e�̼螪oJ�e�=��{�ތG���#��Mx}I�����G���1[g���X��p��ѥ,ߋu�e�&N��<.Y�WNH�k�|c?��M�
�t>�,�s|�2#b��-j)�������o?�ǘ�}�U�ˉ�V.f^��q�`x�9��K�!m'�������7�-�QMs�E�`λ�_Nz3
?�;�e�͊��~�]T$r�Ɗ/U��
}B^���c�k���~���7�jF�.l�g��^pr�3��+q#��)������{�{�H��C���c�L鈈�B��\�c���ġ��q���jh���@d^�Ѯii{���;p��e}w9��l�����YT�'_!ߚ;���¥HfH�+�2k�5�ASF�j�ʙ·P:{���s��	��d	��pT��!i����x~p󂭡�RS�R\o�"V�XLq/	@�U`,0�������""����*܍u�P�xC�|A7K�e#,�b�m��:��*�8�NB�������X��[���J汁w?���h��09qװ��~�g�(�5�׭�F�J���_�J���b��5Ƹr����z:P^��kϹI��\��7��������%��|�SB�/�[Q��"��ƚrK��T��(�R��T#����-K3uwUi�4_I®g����x��t�S$/�������v�"'V��c���)ʮl�R�Fp�I�xrQ'f$��[������X�%Z)	��t7^�RƄ��g��:_�ޘ�K��������.���*�|�!���K��s�?��Rl9g����fr��F���f��J�CrVZ��_�S���!�Q�̛��D'~�A����W�E�pP!.QC~:�/�y��$�c��3��4��֋��ULM��W0Q�v#�C/�B�9��q�=�݄	 S���E���}�AX��a��*� WMa��ə�qOu���EDO��k�ء��NF"|V1r�>�R�ʨ+1�T��@	'��x-x��ˏ�g�ea�{&z��6=O5���p1c���X+���cQ9bǆ�����dj���[���d-*b|Hvցޫ��i�zeG	{i�*.�P�a*`��!���]}߷NM:V�hR��~�
�v$|�RP����(����'�c{!��8�[z��!p`�����B��۟�֚�-T7!��0 ���A�Ԑ��@�$�9	��#��AV��ZO�TL�����N���V��@�2�x�M`�w����@T�'��B|�T��)��J��o��))��9)ӢD��s�a�!8t��le�%?'B��p���?�F씿��������_6_=UbkN��Mj��Y�d�_|�{1D99k6��Z8AM��ƪ�����rF�Aq�� MWZ��m'FM����;-��<|��t�mN��a��O߰�O����O�',���;_�h��u���sm��$W�S�HĊ��ԅsv�wث
�� ��2E��4���a��y��ܖ���䒺���x���X�>/�X������w;Q��kG��J�ի�q �6ǰ=��I�u��F$���س]8���3�F�j��)�/!ݲr��Ք��4��l��hgf����c�&�IK��6�!�Q0���x=��]=���,��d� ������0;����=��i�@w����sk).�sOvA�y��W��oh��6#��Mbۍ	Fm�����F�F�2��PK   ��OXhT���� ċ /   images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.png�|y\����Td�D�+!*ZD˴qk�J*E�B(�F��-��"d�V�j�s�!5hE�(��}�]gD��<�>�_�^��m���s��z_��u�3~�5�7od߈�`6��(��`60ƪ���/�싿��8����������7ت�s�`v�F��)�����vCQ�������/a��Z[:�_��$dcoE�a�`x0�
�u��}�R�8��w��`��&���`>�kq���x�i����-�S���q�A�rg1#u�]�u�\��ʖqѽ��D���A��뗬M�N�Wj��S�1N�0�����^a0-ⷥ�^2�;R���@�z����f����n��=S�u��x^����:v�5��+�5����;����w������;����w������< �M����R�̼��CwR_y��ح�|2��t���S���]o�[��}��C&-�Y�5�	Y|�F/	}<W�|i^u��b�ud�MK�e��W1�F�]����F�I�G������&Zꅽ��c������7����Ϳo�}����������lY���и�vKr������?���dfE-���aƪǛX�nd��z��"��&�99����]�ʎ>��4��u�8�O �d�%���	g�}��&U���x]a��{+�;;�٧xՏ������ZB�����A�ca投�B��䠏����d�������l�i
^�QHȤ�����[W����9�9�nj賍q����#I�_��Y�6l���xrR��Ӯݙ���\�/_�Ħ�:�|lB¾���FB�q%%r��~ۄ5�*����i;�)B���q`�~�*���;gF��:+�l<�'�%o�9�I�?�w$�+j)��˫�,ѺU;�_�vRU8������Z̕�~�!rMG bf(��ْen7�����^ &F��}��l���^
�ŚU����M����{���M�yWVRPPP2�9A-�s�[���4<��ʕ[����!ܚ�v�������lb��ˊ������x��e���fii�����C�{����ޘ�׷�u}xv�n��Z�iĔS���߄{ƣ��yL�Q�'L�9���\-q|���M�99G'�~�)��璛����Y6%-y�c0+� 6&C��uO��\v�zK�W��a���[k�L_���g����sRv��Ǒ<St�fF��d[h�J�l߯}Jv�OP^+5+KԺh�J�`{�����ʬh�}{��٤]&��oү[gnjʣ#�w�f(A�N��ŕe��>298##\Q�jtS}���$Q���7�|���	N�f���k�:9===���h<��uA"������o�aDј��\Y�v�
�U]�*�SSSsbb�≔C�An�U���vRڑ��k^�7ݺ�3���k:�H�WllB�ڔ�>8xnۏ?�{W���o߯Q1?\�=\<m�6���˽������^ϫݧf�^�L��@vp�4��p1���5�u%�m�B���뿼��/-�K۽����I1��$�]��WX�֐�J@���Z�;hTp+-�M\կ��r��Ü������~]�!I��0?��f���󱣃;��ACC,��������l��Us}ͳ	Q�J��`�mk�������\gF!�?77��au��[�I���%6��76oN�.?��֢e������b-��3��&'�sJ��{��p��;v�����R!ս����r�#̓㐣sRY!«
Φd����hur�����|r1�;�l���M�Qd:*��D"���rdY6g �&���^C6dQԪ�U0�h�i/�^
��]Anb�.��������?y�ĉ��Ϧ��Q��[��;^��\�Ӟ�,��_;:ǉ�w���>>"!Q�.B�+ڕ엘�H=қ�w6�t�,/X�	�}s����6Zǌw�ڔ/,--=OM�c���-����A���I�'z֐x�;�\&�KܜQ@R�.FL�Fʝ'�͇ۋ����b:R��Mi�;��)��L�� k���;'�MB��m������[@~�	FٽV�S1��Y��,�3���-	�'��j�Gf��ή��Q����RT`	l	�^�4�$i�]e@j/��~^��QQ�)�vLJFFF|I��.y~W�Ǹ��{�e��i�������335�M$J���6:]�,�4YZ�H���¿�n�E��SR���eV����T.f�}v�0�ݺ:C6��G!�Ĵn��p���Q%���uuuN��������/�Mca5�=}��o�G��~+!d7$��#��H��n��F(W��8l�d��G�V�8���.���˺֘�4����ݺZk:������Հ�q!r�,�"0����l����D����|�9MG�A_i���Q3Z�ɄP��������y=���7��[����㲑� ����Ӆ���c����m�/]�v��{�.��hW!H�g������O��:�8C�jr[a�XwM���=Z��;�vG�ef
���h�! F��-�a�� ���d5��0�!�sww�Y��ʺZ�x ��T�|-��KJJ[j/�.��h#��N8��JTfm�y�?��s�OԌ�%x6�Q�jn�'.[�TI�	�]o������ͩ'x/rߏA�-��6O�=�&�z�x��8_p����C;�ߣ��E�/���Us9V�ºH�o'��ЭoM}C��2�
m1Qd�c�b }��~�ª �	��'���-+>�����d#C[�j5)b�ޅ���e���G���V�E����mQ���7l狧v
��g�v?2b/�Ĺ�G&k�l�ׯݔ��dIOv(2!��jf����
�Ľ��h G_J��?��@ �h�Y�?�m��I�^[�{`|]�I1�ʻ��1�N^^Z���|���@E%%Y��j�^}��`q�����J �@��]8���fn�;N�'����������v��ф���1�@pnR"�6���O����z�Z	��<f��8���=�x#/���?~Fޑ�����8���f]�۠����SQ�v
s:��%E�%���tF�.\:���I��/�Ja���;[=r$ܥ��n[���n3ʱj�/�hhnN���Ɯ����oC!*~��A.��LG�[	h子2�����Q�uj1@F�!C�=���|�ܻ�.��5Y��\Z�c%�@o�:<\���	kD�<�/��ikk}'���o�!�v��% !��@)t@L`C���\��L�V~�X<�;�
V-�z�Ȇ[C.�?��4�Q��o4�p���-�Y�	6�cC3�V��M��� E��{ ��P���-¿��=�6�"�M4d-t�L,���jB��R����D�����Y�(	������$yp��+3=�<;�Oe����8�v�����Y��Gk7�!7�m�w��i6��D퀁/@�!��K�[�mpHyP��E�i��B����E�#�Kz'�nr��>���W7�?�]� >�������˓���F�f�LZڃRG��<W�~j���
2���]&�I\��^����E�x�g_L<�O����kF���k�a��?�4�z�y[��&�?��9ui��p�%'����uA;:Zͭ)K��Ϸ��C���X���NX>�P�D�:�bt�����#�~Jv�%�4�S �� �.r��^��B*��S?��!V&�|����(����2�b���kq��%�s����^q���T*?#jjj
t��O,�fVL3)�����F#��#�)�Q �Iѡ;��#a1{a�%b����J�|��q'���>���H	���Z�!R-[)_ʡG�e�����[�kܧ�X �թ-ɺ2�V��`������'e��i���=��c��f(��E(�W��sW=IZ��!x��g3�|��}^X(A϶�q����Uabj�*�(����4P��w������~Ϟ=kpeWt�?2ӭԮ��{��E��Ln�e��uD죭�(����KT�3����^:S)l�99)� �A�-�{��Π��?�í�կ��?~���Η=���CP��_�����"kFA|(��˿����dXN���m@��|j&��ʦt�8v�����r���&�?�OZ���lqn2�"��qf��r��n��v9��r�{F����wC��� F?*s'DN�z���H��_�����2L ��-RE�D ��m�	��8Pg�� �S�-�4�M�_�۾�
�7P�?V�p`rrr����"B�K��e� ��T�eg*#����l)�YR ƾ-h���U��c��xO�����uR	�8�|�KlT*�\�Fi�A,#U��@|"%&n�rυ�j�.�Ifs���qB�6��X��vC��#�X�n޼y��M�
���7W>���[%�l``@͘=fɣ�ň
Z��IW�l=A?v=0�V��?S�ɉ�
J��|TR'y��U4�jSG�JgV��ԹM�ʊ��/_��2����pE���p˳�ޮZ̈���{��1)գ��գR��FR[��r@F>I=�M�_�:ܧ���S���CC�ww��dX��WZ�Q�8�=C$\�� H9R�S�I�^i��U荌����39��s���`�d�Y]L..�����I���M9lkR�d�������(...`��)�CW��m�����{�߽��Χ�H�N�sǧ�N�0�);�:��^��V�WD�c��������!AduP����zR
Q����a���[y�z��sܫ�A�ժ�0(�I5?)�[��b�eA�X�#��G3-
>�����p&�rJ�o����%ub�$,��Uy9�=���c��׍ǚo�R���]�r�ލ��e��Ӎӭ�0^�/�+�,_7s��e���+X���NzN({2www'��5>e%X~4�d�ڵk���C���G�B�t�������r��囵tu#���x:5##��&2�nF�΃$�n�����R�	��;�ϯ�͢_([4�=�)uGT�D�5<��Y��2���=d�|��2�:�}�Qءgx۵�~�̽��h���ԟ��H�K�����⤻IZB�8y���PEP�c4 Y�N�g���i�j88�E]��9�r�I�]��e�Ϊ撩�Y������婎��ojj��ۘ�lIK�Dw�w���9�&T�,��))0��v�z�j�}͡?W!=\$���57�ܺ<�,��z����	���� �����Xj�F�F��_-����h#���'X�s�,�E֋�-��I?�#  (��Ǔ,�q�9^�֔��/$R��4� ��?6>�*=[�8��&hib�Gxx:��O���M�/�zӭU1��ꇧձ���7d����|�� �`0ã���|ڹl3�֌T����sM���#�&Ï�HK�����T�>���Jܺtqj�آ��G^Jj**��[o�z��y໧�؜r�E���x�!�������\*�XGF����u�A����6QS<�#�w�S}[H�/��YlBn̤�^2$S���B��C)��1I�d*�f-"��ɕ*�nn�<d�S;I�G�W��?��C���z׉�2٨Zl1UϏ�y�˖���HJdu��1�~�rJJ������e0}ю�j�s-�v憾��ٚ�0=���iC5�c��s�bލD��"R^Ϻ{�l�a�S�e��ZFFm�yTO~sdnU0�������0/�����}���v]ASs�y+
�<ON�O��n��0�l�}�Νb�Z9B��x�����H�#�g����S2��5�Ɋ��v?r��*��6�5��7�]m�率�(R
���I��^�"��L����##Y$ڝ�mLVOS0^4Wj-��n�M6*8���k$�7�<5Wz�D*[/�q�n�2�87Ox��S�i2�3�"DFFVs��	���N����d�#y�����kը4�H�f抗�j�f������v��z�M�T�aU8�i����2.:j�*�Q�q�}���r�s������Ʈ�m�����3�v���3�]qBT�,���u�������we�_,3��r��ܦ�ӭ�R�Q�sb\�9"���y���Hj0��jL�3�pv&�\��*aݚ`L�%^�M��Ή:�}p!�cl�K?�K��z���s��݊�á����J����P}��{0���ȸ�UR�ŷ�o���p5���T�?xP������s�[ �	2��u�̦zXdm�e]n����S{� x?�Qov!��2�|QؒD��"����A,
�I�cJvuR?@P^�o�娭0?�(.���������Q�˟�7�
O�QM�A�Ņ0���  rST�:�<̿�8����:��CWW�e��ݟ��+�;�N�ZGRx��E!I���f1�����8��Dq"!����[~�U�$lb'�@�G����d�E�����6R������pȆ�|n=]BWH%�T�3�i������c�+_~�B6z�T�Unn��p����!2B���7m"z<�����s����!������{8��B����qo�06����ʹ_3:������'r�Xt���39��������*���,����o8:�؟8~�833��ww+���1oxsO�03��(�K�����'����E�s�.�aY�DJ���0v���q���R�Xk:���E��
����Z�0���>��uuu!O�x���C�^~����CA�]��@0�c�Ν;�&���{<�<D�@�7g�̰�9b�ޠ��q����!��͂����Ό�����h���w�bcy�N=���4�y0h�|�8a/�&�]a�:g�N�g�Йhkk��r�좙�,������i�����A�a|��a�����5�[g~?�OmvCfLsYqA�;s���G>;q�����]߇g��DB"���%���k+t����(]�t�T���Ј��xUp�m�\�E�g�'6������.��/�X==�Wyyʎ�ӟ{ݿ���d;� )���l-f�>+�����7����&1��l����x䞟g'�$2��0*��߆ey./��zz��%:�EǸپ�������,-���{aK�"M<f?��Q>��+IL����\�_SIM��s��21I3&���	�5�k0�]�}��Μ��l�UU	�g����($QV�V���rc�D���e"� ���C~ʒ��9�����)�&9En㘟��>?U	����8�:Ɇ}��Ri��Rdew��.�ˈU��n��e`����R�0_	����x"ɴ?�|��W/�����D���?��������uH�x3�\�qDD�����d ��$��pH�Kٍ^����ۇK歁1I��ޯ�v],K�}��+W|��� ��4���R����"��=��T�/�c��JKw�,u�tR��x�= lX����:�S���qpp@���o���!������C������B��0>u���OK�`����g����CȻo[{l6646Vf��{H��<�����{xc�	gE�K`u�_z�B�i���� �:!�Q����W`�3�ی���K	�pهG��A�K����yB��dŞǸ�?׊CA8��:��y�����If�ux-==0��X?�Ą�}��c�g��j9���K����(���"��Pd �J�7ݺ�-_:ܧ� ����i��J�����1���QA�)��֛}yuUԼ*�yZ��u����I[D���=d<M`�Qu�c[�w�;85�q�d�{���YH:Y�c)���y�� �m��D�:�aT\��U�vr�%%�ggg�}�l�����L[_�˗��)$EԄn�gI3sUm#�]���,�H�H��,]�Ƣv�d�A���	�b<
5��.����a�v_�kQM���H�ud����,�Ůĥk���B�� cCCN4����CYכ��J�Q���eܨA��K����Z�UZ�|�tqq1�(qGN��c!�p��˾��E産C��* ������C��������<OM�X��rnG�M{��--QMM����

(�!���i����Ec���5z�4J~rʹ�͒:|$�{㓔���N�с#xo\z�!�6�
T��9�5���0��7nެ)�+�N�%o����EJ���XOm����]<��QP.��^9���խe��5ݱ%%r�܊�u�����:�RN��'��2p���+KaBa)�%�\�����p봸�=�B�� �����cW�C�Ҝ�e��l�P��"i�o?�������/I�����,��T�<".�X�p�һp���*U'�Դ�ۉ�B���כ�oF��	%]�H`>~���F��k�ޥK���^�I�̴���Q�%e�uأ�*J],��2�����~u��q�Z�_#��X�Yu�Ȣ@R�}��C�/@�qF�:Ec�k�׈|G=I����G�Xl�y�:2:wZ�Y�*�Cð9�PL�٨g���"��|��B�!�Y1��u2vB����lVgz^�?�'X�9HX,:nϏ�Rvo�tyz9��u:zqF]&w,���|"�uzz:��ӷ;,�3/ف�4
aꋥ��X7���"/��?�`��� �mY��I�F�ʻ�ө�%XHgz1��3C<�z=�������M�/n[#��%�$"n��j�kew^�������X�#��v��8��V��WM�=J:_s���ANV�;��y���>-/.��h�B'�)�� p�t�7գn�UsK����)6LLlv�*��̘M��&;��]��		␨�
�0��aW�.Q�Y�'�6Qc%�L1R�V�ER�6��������CB�d��|с�=C&gg��z�y�������I�A;H�(���r
O�y��	�0l�u�R��:��P+P��_-~�����"ؙ���|�׾mmmZ999Z�f rv��͞�/�a��uV���)@4���.]\@�9����q���]ee7He�3�l��
�uR��������0d�h�����_��}�Ơ~-c�����7n܈����>w�-U/3x��Y��8�h��:.�#~^�ok��ez�L	.��+�7�@��E�ĹI�h+2=���tq�!����+���#��0��]J�?�vHFN�d`ˈ(��T?�4�Ƅ�ֲc�5݈-�d�3�e�"j��J5dv:���$g�"�k���X�p5�,�Z��X�:��!;��͌ҥ9h!x{ZA�C��ސ�ɫ��=hX���%j�	斏Ʈ󉘛���s,َ҉�K㨬�J��F&` �o�s	��Zbe;Y_"d���@�b�Q��0��:Z����An6
2t=O�?JC��I1�Vw+�pJn�l�BMZ���v
�M����$ J7Wo���_���O�>m#�Nʀ��	�M]`M���|��nSDqy����%J5E�2���>��@��Ȣ�=�*�]����_� ��^ֶXq�W$���n��⼁�6���ظE-�Pԉԙ��:`���[YŕBvq����i�<�6:1q�yd��h5�/�Y�<.��Њk6B3n���Y�܌��4 #�:P�hԺ��Mi�L���<�q���[�W��ᦦ��K�e5b;����~�'ʦ
�5�<8���=�AR����P���T��ػ�xzQ�o�֬d��)oɳ1�׸�;�jD��

��أcccr]�0���);˼鸹��� K?E�Lx�9�=��Y�bH��4Bg@�Y}~�����B"��ZO����w�ޤ���j {"k4n]H �Ine�,;	�� B�{ooRm���uxHˍqYwV��`�%3_��гx��FXP?�ۛ�+�%�q����e�Da��z�~t/��L���5�3��>�wtǎLL�[Z7m�LZu�1�k�5,������wd�������)bB���Q�$�~��%����LiN@���^!v@��-��ء�84�;w ��>�F�������Ɣ
:�������/�Ə��r�V2#�H�5H��m������ˋZ��[��x+��g��>e�v$=�8Ib<!�-&&-�:���у^ޖ���G�/Z�63%��R̓�!Z�k��P"{�ñ�4�i�g�S����M5�jt+@�7蜭
9���D�.y���A��ao!�L��|�F.s�D���F�!ȓ�N0VfzL�J:�����B�l`�]w�p�}S�����4�KD�����3ޯ�9F>�A�鐺�ΟgG D������Hۖ��"�qi{����܍�!��jnOv�Yt�?�)w���|"�kvv69le���������q��v ����C ���}�D��0!�v�x"� L�����cb��Y�/�yu�㶈x!>Li�y��%RY�Wx��h�'
�;��Jĥ�
�}���:�Aڣ�`faIҠ�95�2�n�4��ЗH����B��WWø_z����iS4�ĉ�q�r���u�+D��s��c�A����h�KK5<�D�^�=��z�OK�}�UIVbGC�	��r0*3�b�QY�wɲsHX�����TV�Qؕ�Sͣ��U!�]����Ͷ��~?�v���� n����d�P�̑n�g#j����2�d`SI�(��f��o�*�ink�B�r2��܂۶����,&n�M�,��Oǰ���k=���'�gGa蟀�.�vUT��&��X&u��y
<y�%yR��T����VN�}����P�1�1k%�|��46�ST�:V/��ǔA�A$j����2�QZ�&ɁFl��¾f��#�)u��i��K�;�Az6��:�*3�7�<�;�`;3���Y�s���uA(�v	��4�=8�ʾ��>Dn�
j�E)`�|���!Sh8��X����hD���
p�����g6 g�����J�(�k,֑�{�&���e#�HQ���u�� ̻0 �E*1��1��Sh}�wt 5S���q��t��]�J���cSRP��WŸ����	f�:��G�4���_鲐�?j�꓏��L��Gb�uO�\���r�M�)ӄ;D~�	5N��A:�����M��yT��ma�sLj��&�zz���Q��6G� 	4����MN;`"~ZqJ	+<^�r��x�����/���9�pw�qP��{����сO~�AjMMMX�\YSSs���ԗ{����)w*@
Tz��ڰr�R&�K֔�ԑ��fj�DĶ��3J��p��'"��l�q�`�P�|��G�^�H�d�б����ZU{������~&�J��2#���6����S	{'d���?�mi-�#��K���'V�>H23�ۨ����a��l7��DDDh�=����b�Ce1�}��0���^)�G�<fPhݼI�h6rL�Ja��xuW��.��Y"j ��x��2�6J���>)�gQ�V����r�w~�T>צ#����#i�D~���¼���x���w�O�Q�d�Mu{�+���,W�r*H>�� 3��c����
�XY���� �{
X��=�����f`���E� �@�.��$�5�]�TUo����FY��o���Q~�va,��&��<+K5G�rf�vr�{E�� Z���=n-���RSfT��g��!��j�	ʚ~�l
W�a(^ڱ
u١z� ���' �6œgQ���y+`k` ;�F_���񩪪�<��"%kc����Q
�)dط��χ�n�`ع��.��Q�8�8ر�hW���@����
�e_v�
�?�L5�vG��kg��p<b�O�W��5OhSxx�o�F��V�\���<=]Ok�
�k6�S���yFF0%˰Ə��B�^\>dH�=>�j:�q���.�	�̽�>�*�PB��ѫ�L��x��k&�L��O������Φ8�����w�i��<`�8�pSF���/y���Ѩ�J����J:�]<���,���x��×�1n�ŭZ�������A6E<Q2�j��u�O��h��J6�z݋���ݫ(�zO�/�/44�R0�����~=pP�hkadHU�`�Al��Q�*�}  5�+?~\GWm��JFb��BC�Y�.���MX���H9P
����<�XEy7n�hV��Ի��ⅈ���PH����%�S_Q��TJO���u��c�GG���2?(�ߐ�bE��-v�{B/ 2�L��'�]F�`D Ea��2S��pT�Ӕ�����X�3�J�c�~�@�0>E� �P�?<\���������I[J[ZX;��:��DT���C��@@S�%��9�`۲��Rۦ[4V
�	`p�H�VN�<ʘ��{'��c���^�խ���GU_�{::6\��H�L|]4}:������G^�.�8+7��r#�1�݉���ʼ<�D��^^�޻uF�{K�X�	/�L�?�ޏH$�IqE@n�G��!���M��	����&�o�ܼO����u���_�%��q�������$��x�Ow�����W����W�&j�VN@��WX�踞����U�c�8�>0���@�w�ct������7��9�\D��r~o4+$��kAlv�/.D	�E2�hyxx��O-����Yv�T266FZ�1�V@�9�3����&��J��L����IO��5ݔbP����7�����=��8n��-��̓���Pj��l@�Z(��쪁�ch�V������\�h���իW�5Rvya|�8��s�6� �r�Yݒeny�By E��>���V$G�]6�S6]�˽˜ঈp��21}�j�@.�N��Ać����ς���AG�a|�'�ƨ| �>�J~S.)��%��6U��ڿ���OQ�r��Uកg�cD���GI�C8P��P�/Û�/E��s�{�h��c�!v��v�#�N�b�@�no�֜@��9v�9�퓀��� )G5�3�ފ �Da��_���9swf�t�R>�'�)�R*�6���sb����

����&@Q ��8���Vn�X��(K��]@5���mG�g�q���b�{{�o��d��.���uG�ЅW��U��ܞ�,�Lj�B���Z�ῐ�?G'�ھ�\������K�X�k�`���8\%Z;�C�䂚�>�4ee����>�9�X0&$$��=cg����߁�{������î�9��2�{���k� �)W��mu���z)))�0�e0�@�����.��b�e��H��b�d*'Sѣ�O�Ao���	���򳪨���AU�njlA�˛�e\B��_R$0G�k�˱I2�ߡ��+66���VA`y�⎺��.�ꜳ��4�ѥ$t��.n�ߣ�c���:�N�����A���E+� ��S�n�r�b4����K~�3=���/�aFU�ъ��r��-���Ы���n�1�}�|�5���"��Kl>�a#�YhnnyIm |����*t�1E�'�r�x��ȆXH�����B��:thT�sB�w���K�_����
��BB��@���kx�.��R��U�:�mܺ8Љ5d˹���FFF��Þ?��7�.F�����(�FA��ϔS�v��E���U���@G0ԯ� �> ы
��7���6̼��t�ċ��g[��:��k��:Ŷ�J�Y��}���c���'��A��{��7����X	���`0��l�T�%F�P�̼�+1��r��,�T	��-,,�����A�:�42 ��뼎?��9����D��FQnq>�f%���*U�"��|��^��Hq��Rί��ji1�:������L�H�Ofz��<QX��Zzzz�ʅ�y����M���?%��m� ���x46fO�H�\�~ݰ��W/ �(�4Y�4�F?Iыq_����1R���葘E8";c�04�>�+��b��s6ғmvvivew��b�0�ʓw��#���~y	�{86�����u<	>��m����7���}jh�7�l�A�e�V)�#�}�Qt�k�&v�=8�SD04�vw5�.�ܖ�;BJjJo���)'�`����!%�ݽ���=�-��9(���!yd��X�mص#�t&����A�������#�fdϛ�麻���3�S�x�Q���/�H�dmS��wWh+ڦW��]�G6EGI�帖���	啃dr���<2Y����x�	:GV> èV�N��O�H�.3 <ѹ���Tp�'ORΙ72��+sEEE3z��~9�{<��|�$�*UYY��-�t��v�Ζ;��={v�g+qT�L*{�P_��y�a����.�O��	����vS.T��]:�A,�F�NR��qv����xI����r��1���(�u��;�v,�Dw.�����R�b����u����F�G�tK�T�~ѣծ�(��EҖ�����T�/}@Q$��m��eSZ���[� ��3H��H"�4+��.Q��7��
���@����PzKQ���1~aa	ۻ�#���ZN�m5�!��"�G;�
��tZ��_�Գ���w'̍� X/�.N�#�~/a`�N����εs~,�pٍ����j��Cg�讽����\�h�M�A��x'�1\@���	�᪞����Ћ˒���9���&Ƃ~BGP+WFD� :����o� h!R�{�-�#@� F�Q��;�y�P�Z�����D�|�AO�O׊SB��(����h<@}��8nE`li�s~�&3`�_//N+�R��m@���*��U�X�6b%�t:�%5袞��(� �#����r�Z����Zq�P��?�\2}��f9���.��_	���� ըe+����aJ� �|萐xc������G`�T`���0
��T�^�F��������o/�ɀv.G�G�d��?{I�V����ۇ+~��5$�P�<�H^����;v��>`f=��y_y��=B�� `������/z�:���9�Ά]��Մ��Jщ2���gm�	L����pr$����+��%(F�,6����Fm��@�mQ��gՌ�5�/���rFyN$���#@����]j&sg(L��%�&����Ǧ���u�?QeeT��1X���X:�Z�o�������Wj�i�{�Y�~���F[�AZ/����A�:y���C�����Qy�H�cS��y�."��}}}*����$D�������s#<��EZ�����sM�.);��:�D���υ���7I/we��w����G�~�U�c6��~<��z����6��ƛ��C�~Dg���4v�Q[{_�?�o|4�{�y��硭���S=�Mt������M8�Ǎ��$�bZ����Bx]�#��~�ć����D�v;;,�@E�;�x���{"�o3���'c|��i6��&�z��<ʽ���1D|���v�m~}���x��4mL+/�-��k�>f)B�|�� p�E�W�kʼ.?K����$�U-w�����b{'DnNE��Ћ:,�Ѧ��e�Ś҅ {�t�3 *yDA�Mt,/v����Р�ݤ�A�:��������4��*�/��K��%�i�2��өO��a�F�|9���J�Erl:�ҍ��`���:v��A�K?}�">�%����*��!�O1Nk�#�z��{��$3���[�][ڑ�O�A�loLs8�v��L�D0�4$�h@�4��9jO> �]m�����R �#-��E�Ν;MR���ӂ��0�@1����f=�]y4#�X	t�ϳ����������N)(����wov��=qx9�/��z��z��Lt���Pey:�+A1`����s�Nx<Y C�;��[`f�1�z�oo�3���[�n.]�Z�_2O���vb�K
�c���=77��z��_�}�?�؎���������7)������dքH�kld�ϵ�l��!m���Dz
lW7(8�|�1��dV
��޾ͪ{�1*B�288X�UN��X�Ɣ��'�;��Y��_i�ndccs��l1ǽ�o��.O�}������b��6��dv5[f'��2�ij6�2N��=Ϟg_�s���\�	~=�����Uv�ų=QX�@8�䙇r���ɲ�ȹ�?����SH���`fjqqvm�ŋ�5��;�|���v-??�e����� s�˗�X&i"[�]%L�o�Wx�}�I��f�~�z¥/i��p�I���/*xΔs�1�Ӓ�h�lIe4׿�z�-o*�������#���XmC�O�.RU5N���cץ4�Ь��V�Y0�Ž���n�x|zZ��A������w��}���1K���$�o��6E�>��Yv�R=}ݑ&g���q�o���F���4"�Y���N���;�g�����t�u�>ncF�ǲ���Mh_�d���Zi�N�cRJ�6����r~����hwUa�89R3KR�^��5biɣ�9;G��] �@d�B���Ǘ𷈤+<��		��z��uz���Tp@Ȳ��^$�_p�M�q�����+7��k ��q�^DH���"�W�KZ\\<���U}qq��?�h"�b`qM��`zZ��E�_��20�@�ƺ-�/�l&&n,�T�����j�AG~u��器�y*�s���z;]̰�w���XŹ$Ϲ�ꏏ�Ů3�R_K�Ù����O&���rȮF�ib��bbڈd���ߒ�T��0� A����0�q�ܚS4� 4ū�M�:Q~l֭I
� �4ИFdgA��$rt�G�BGC<u.�ᇆ��v¸p����]�9�H�8����X�5��	���8d��[��~�M�W ۀ�����&6�RFaa��/��7��/H��T��񦦦^M�8�M�~Ih�J�d����g�ݡ�Hh���a��{id��~�̅ό=f/��c��u�v��,�2���O㴍αL�%n�E�a�m���H�� ��{�f'����L1��I�s.���|� ��F��}dL���kW�f�ad���Y��q���a�4��=F7�?�d�dD����)A7;vip��1�Gn�DwTB����x
���j��2զ!�tI΍�,��&2�i�,�D���v�Y�ﱕ� �O�m��`[��ۅ�Y��YJ�=�\Br�*0�<p�|������iڶw	��z �%pΗq�mhh�K�K��Y�	@Jj zL�]�t	�a���		��tth1s���!'MLb	�,g�TPp�(7���Q
.B�LG3�u�oJ;g[@��DY��=ʯ��o2��	]n���S}=�j�;��e+%i��Ra�w��v���F����J��C��!���l�!j���:�O,�2�������۷��-����I��)�v�~�)��1��w�d2�����V/���8$Z�̛�2��x��֕I>:|��ev6��M��D���9::�&�c��I[X�8�Q���){��T�cWY�ʮ^b����� �ޕ����I1M����o�U%���y{��� �y�<~�Kέ[~���ӷ����@2�yp����7LT.����_D*�D��g.���~�g����1S<���)[���0}�����e�m�[���P��8~�̀.I����#22VT���	���132�6Gv,M}����*�㘽~�}VZ:]�+CEL0�H�qƽ��T�S�y�i!��|Ȥ��*�v�â~�d�ê�<{�ۣ�v����{�fY�@�eѭ�[d�u�s�1�,�\���ڎR�[����|��K~��xmmm����ׯ�2*�	����L���{	�a��5i�1����i���*��m��~�E��o���?iz�m�}(Z�]���CZ*#]e/���I��G2� v�DS^I�2�{�n��ӧ�B@�R�����9u
�=�Y�1ʦ�^��IH��D������Z����x�@�]iLѥZ�ʅ(	��o�w����4���^�{�QUS�>~�G�e0�V��5U,���6�i@��[�ݧvĢ�s��UP@���.h���տ��p+��!��	w�ڵ��a�%�ג@�#�d�t����2��2}?~���ƀ���`~Y�i-�)�7@�&��Wo�VE�[��J��6t@�����yрf��e~7x��5<M<��=h�{��ly+���t��� =��mbB��6��(��~&�g��
�.�=>��m��}l�s�Ƥem׿��"��pJ>ML�dp������Qq�%�����@��l�/�۰xy�v*��ZXh@!�w:;�����8����1����f�{IK�hJ��˄����z���'A�׼���OHH~�ܪ�ȷ��e�G^�d0n�Fd��.��7��l��عs I~1���ð
��{Eh�@F UW�Ux��4NG��A(��[M�X�Ƀ̄����Y^��-�J%A�U�jy��t���x�c��`��,��bbaa Ȥ-����|�P>Y�r�wö-ws �r1��3��z3��у&%�����������k8)H��Ѯ�q]�K�0�ͳ�9@�x����`��V�@����QU]@P0��+ `!���}���?��4Uo?P5���b��Y`�ɘЯ��H⹊�\�^�*��x.!!a�J���&���
�A����EkUqpȖ[�1���/z�1�"�b��?����a� �����{6��*�����}��s�U�h(��0F�p�V�\u{u��o���ÿ]�_�����?M����2,M�ѵ_�_Q��jaٜ����(0�9>�q~��zLI��_1L`DoJV�G*�T5��%��F(�'Ҝ�&���Ǯ闸�g�&��'�I"���_��6t�c��q��*?Y��+�Y{ěVYhY��q�s�˰��ΝsY�퍸��6�[o%J�HJ>oLՃt�
�G$�l��3��/$B��%���dΓ315�ĸ�7<�t��Oi1X��Y>$���V4���2�)�UG��I��ЍQO^�� AW~��.+�e��a�n@���/.��B�`�QWW����؀fF�Rwlp�x���j���d�
Y���,�b���l�C��끙'�g�<���3O������qtI��6+���~�p�Sa���{�8l��r���u2gv�����������-Tɚ�*�7ک8� �}�Qf<vd=H�4���T�#7�#� �+]�a��v�ݻwG��d؛���$ &VP"���4��*M�R�����87	_��X'Z�}�į�l���1�O��t,@��x��n�s�Nѹ@��z�h���>��$R��jH�;}�=�Nd<dy&dŉN�l�]�	�hT�.:G��a�Kc���a�g���Z��M��g�StS��Q=�w��irLW@@��M�������D3Z!;�J�Yy�U+AV���I��s������g��	��m*�A�]�e�s���X������Ů�����֛�S�>���;�ž�J�TDYCZP�d	�-�ز�Ѧ��&Y����-�#�R�PG�Ph!��?���������u�y���y��k��~fZ���<�3�kr���T��l;��o��ߏ��Ղ�������0�枚˙F�O_�U� x�V��RV�	.6/9�	>�G�IJZ�@��xɋ��o�u��3��sѬf�?a�����^!�����	׃���ij���U�x�C���9oE?y��*�0l�t��/7���Q`ᓮ{>��d}Xe^DI�a3$���dZ~�:FY�#�W�/���나P�[����4��#_r��N��S[���%-��[��%�o=�{��?m��9���ϐ$Y�G���{���;�������7�+N慞)�����)����c���p����D���GC+׮�{�ҵk0��6E+�b.b��Cs5/~$��[,d�C/v������k��}W�k����ۖ�R�:��s�������*z�}�^B�IFY(�F]?�n�rt����O.���0[�ߦJ���mlh�˺<==<W���(�꡸@�U�菋7_b~"��6�RG������$\��+��~Z�IT���I�T|����<>O$w23�s�, H0l�Ѩn�A�Ӥ�sqr�}41�:X�+6��G̷��޵.�"u���6M�z�bbu�E�n���ih,���>!���ϗ\v�065�-������}�����5;"�Xk�jr�__LMҜ.R�r�|�s#�H�<s����n[�+8�� �yp%�p��Ƒ+�J��K�#�:r��������lB�˺�;s?8����	��<��҃׭(��~,ή05���D�.�s�� 8�X�_��Xtf+>���ߴ��G�
����_��;�z��Y��	�(�G��T���F-����)��]�&:r�����p��j����@�����2w�-#��ѭ���.���5###f�����k>�_!W��K-U;��3`�~��#�_��|Ω�':8,C�

6@���E��R>�[��f�9V��Q?��adj��7L�[[gc�r��f�_�2���O��5����P�����毚���/�6��u���=���Ϫ���FjEDD�����0���NP[��� ���r�y�,�����.����b4\�|�l�3���;fo������4��l�k�wo�<GG�)��l$<���?��9�
y��@IR�������߇r'�����gՍ�����\Z�J�Pk���0��nnYR	��$6AN���~�Q�
����u;���]01Ȕ�n��D�7�WR��&=R���m����|�Eꍐ��DB
�0A1���w%�
�*{���H'B<�=<��㋄��Y� �w�}�$����;�\
Cd�Y�[X�||.4�I��d;��m�����r��Z�	)�!�eʆ �x�G��Ā�Ʋ�FT?� I��ם���1�շdZd�<8���م��ѐ���	�˚;�y�����7A��f'������/p����>����ꁘ�����J���LW8/��EQ� ���o߾v���D��4Z(���V�`�R"I�~��_�1�����Ɯ}率K��v��+�ظq��o�}؆UH�M�ɑ�\���Sʁ���:�N��C��g�8�[b�ns�˚4�`�˗{ �H�ϒ� 'w�8�|sG�]>>�$%�֯$�g���i@�?�c���Q�Q�D�qX\�����m���@3�ED�	'l�ܖiII���� 'e#G��ڙ�����GMì�~�{]�,���+���L������\}�w;�����x8N�%�dU��]���Z��3<�			Y҉A��,c���J�>;�{�)|��A«�p��R���o�[�'n�raQ�8'��K����J���V�wy�'�َ�_�*4ݻ��fZ[W�w��(�~�r�����j�A8 �8��V�	~l/<�ui���f�����/����˖�kη��x���gq��#���TY<��b�������\ s`Z����Q��`do��9�/�A�Wo]i��S��*t���*�.����gϟ�|mN �8�����1��������c��LDm���U�.:�D+�����uu��6O�)a�#����a�X��� Rx"T�
y��	ϴ�XS���6���Rk�s�yc9hm=:*i�
!�@xq�������|;����g|�㟜����#7�����Aj!��D��l���9���{���4��:��,8�1�	���zg�;Qc�?67nm�ȫ,��_��U��c�`z�azix�+/�	�t��! Bۥ��J�*�~�T0n��u�~-�ɐ����J�b�iچ@�m�sihmy�|6o���u���E���ʩ%��+�n�1[J|�
�u��*\v���_fuD�8�^��K�46�cW��:�2w�#�����;@k���"��>���;w�Z��ܧ%�B2>��7��M�W�޹��wA�elf�}���\�!�u���#vg7� >ڛ�L˵�$'!ʹU�b�*�N��� ��e�#o]�����+�:�<��'�<��8�v�|�~�j
z�%��� }��/���]����U�Dc}���oQ3���>������.��z���U]g��Y|��E[�e*H��>�Ƈ�ԑ�]�l�Q�>8	:s�|�O��I����~�q�����n򠾎�a�+XT~��'kAjj�*S�л�[��7�u.��J�һ0Ѯ0���<2�⣼�$ �h�����4�Ʋ��<R���1`㕕�w��%OX���������?K������ �/���k��z}ĭ�l��qV���;�*�Sς�j��t"Z�ќӾ�m��� �������#���J.8�������\��odt9��c˖-w��[�����!77ܠ�c&�UC^Y���葿��^齺�DR �~��-����6���L�V�A}�ͭ��*�>|�xhr�ם�,rwVx8�IQGWy������]�bϧ��q*F����QL������CA�v*Y�9�;w�v~~�jy;XS�������	��1V!�;�F����V��^\*��@Bn,��o�"�uiH��\V6��ikk�U����1ɹ�=�P�U���ǻƳ�4f,�	(���3[ݓ:�s��i��	| Jc��ywn߮V�[�:��K��O��|�X�h�Ft?Y���Ĥ4N���y�֌�#�0�S��?
0quu}~��V���Դ�H�W��W�%j"���I���o���|>�tr$;���f;�4���B�DUU�+[�$nܿ�8�H�:��pb<��H	�qrUD2�����O/�[�f)mؐ���*A�;7on��/�����9��L�������M뙳�{+d}����ǊO���+��L�򙚘�R� d������/G��a�7����(������6_Ȇ%��ԜZ2>%��r��A�����2Ѫ<^����l��n<�<���������{V�6�|���Z��Q�%������j���e%m?�;'g�}]�}�ߚ��ys)(%=7��!8���s�'h�N������l�`6�:�q/�էDd?��?Tv���ݻ�G� �W���fw�3�t2�����d}���Kw��	�?̴���?�����k���oK|�!�^�v--.Nt@�VQ�e�Ye�%"����L.,4el��d�fC.���Чh�����L�nMN��Ȫy���߿L�ulP�o�����K����3��O^M��O}�o�2��K����̋�	�&D���kK�o�4���eN��
[p-���M���A�� `���ANsi�r�<l��4ѽ��*�{����k�e�'����ۮ��ד�w�����|}Uל\\�$�qpH��'����/�w�����hbgle������'q� j�AII�w/j�� ���e`�u���6����SQQq'=R�b����7SQ�����	�5��f��~�u�4p]�9)��ش헥��ʖ��~����YS��6�7�����ϱ��2��w�j���in�HJ������`H�����$<��(���|w�K�'��_`���kͥ�0C/�x����C-�d���b���q`sCÍK��ܼ��ug����������g�i �1�!���H�Qx<���9�!c�;������`]"%׳��/^��d�	����[=����/5��B�����o����;�����2g�rI����><�����g�r�����e�VJ-�o����@��Q��c7|8(U�E�>��K��8�X[gǫ������塀�����f��m�%�ȃ��Pu5*��o�}�L`,��o=LJZ��ڊF�|�����I�5�#�!We�RZ?�>M�tUwk��Ϡ-eH�1����+R� ȃ7�⮂z��h�"A_�pA{��pE�ɹP5Øne��[r�j�����'�օ��)g�E��p���[���K6�[�]Zj0h+��u�2D���K��\��耬R�?��N.A�\ED����bbc�8�L��Ib�ǿbժZU�54�?���=�,��$�q�W��	r@�m�)ɋQQ�ǎ1ÓkTY�;�&�����}��SU֢e����0��<�4�z�W��ADt��O�̿.���,����/g>u�.�q��dWГa��OODh+�=1�"�_2���ᑃW�q�瀢� ��[���`�#4b�!i��xzz�v==�ւE�?� ϓ4�9wm���f\�;%�&O1��E�D�܌��GYoW�9 +Y��Ջ� D�Ǝ��*�����ھ8u�FU�B��̭���Ϟ=362JvnJ5s,��$���de�G��R� /Z���m�D^m����-s�	<]�k$����5ı����i��F.M߰u�E�3fy驩�)))xBə�d��9h�!��������̢��b�u,�d*b����f�҅����Up��tnTlr� ,�ML�b���ۼT��#�<n
�x~]�e�N�5k���Ӌ ��7R��b��V�~�������"b�5�IL_g'']���vo�~u��z2�H$������TTT<�L����m�S2������7y��<6+D�]��@�3ٶ�$�q7O�)��<��u��q�j�+�s�?ʆ�Ĩ����w"����EڒP�P��ލ��X|o���9E��L�H��@��,�K|���K�w��?m!߱..B�R �Eݭׯ_��z�~�
�r��I�xR������p�ӈ<E_����08�k<u��K���F��r���t9IP�=Eu���7X 
�Cʻ�?�̑�������y�Gw�cy�g������[UK'N����Ͷ	�(`Ïϟ��i1-���ҷ(t313�ο��6�Fs�q�v�2�8L�V9�+Ʌ����_�ƁO=y�y��{ZW�^%ώ���9�	a�᲻{1y zVƖ�;�h���׫W�RS��V�r8��ڮ~����������ny�֙IK�X>��6����?";v�(�4� ��d)%ʭ�8X!��̥�B��?oߚc%K0-,�R�d�
��ۜh�]^�5`��x6��$��]w��E���RJ᧊t}�y��R���u)�ғφ���������D��b�Tb}h�C���`�-���xYڠ@��Mg�ˑTކw�&�3���vH���k�e �E��;|�i@��׀)"��$��ϫ���\�� �m��'d�xpZ!rsVi����]�G�W�̲e�/�Ф�����׭���a��q�	d�O�C2K�B�°BC�<w�&a34Vœ��"&�0�Z���\,� �=�g_��f>�,�p�Y�PɮY��n�FFgH*���X�\��o���E���G�JnV6���d��ITrK~6GFFa�}�r�����!���\Z9����,,,o�d���FC`VW�\!O�u�Z"�?�\<�$%�;������H;��l"������?u�aA��b�/^p�G�A�� M7�ڌƂ40�/�W�Us
�W���<�=u{���OXy&�3eٵ5���͂(���4Enɴi�2�	��Z�����==N�t���g��Z�ǅi�I���rk F
���;�
%�>-�]Y����`�J~a�E/AY��Qܘ'g��Bۜ��X�����5�,<-Ԥ��A�T����HE�����5Y딕oi+̀���� ��I5]���+B�iw��'�1�=�.Ϻ&���hXg���g�n���y,��7�I������2�U BCZ�����nU�#�R�mʘ�MA�kq��Q>�[�K��a�S!.��򗭯mij*�b��sf�ׯoWVj��� �|������F��qk�	PGk�EN�����\�
�@s HO��L���hl������M�]k��������P,�(e�2>��C�28]�@���b��2��7�<0���rN�<���Y���>>>�(��
�!G��C<�Seպ408���g���e$��gWF�~[��P��y��ё�+��Ő��{���(=9�B�/}�a�����Ԕ!���D؀�z�,�nޢ�����o�ۏ[y���@��٦t6�����
���Bƍ8�бS�[2\_��[_�!: I��c˳n��'Z�� �1��QrO ��6,��o[��,��]��ѣ6"�����W@`�4Uǣᐴ7��W���pOv?>��Ԋ���KT�,F��E1�j(x�U<Z�Қ�|�K��v]L�z���O1�*o�8}����]o�n�0V"�'��B��W$�x� ���
[DeC��k`K+�s6F���~h�;���0bH��CLv�l�ڟA~�@n���C���zc�N�B���ooAp����ת�� �C��J\�0;���W�1�n=�=��b/<� ,fd�|���}-f�h�,���QB*oE�������lr�^p��9��ɉ��!!�DY�Ǐtď�b�t+��j�X�=� < o��X\y3�������*Տ̧�s�6 	*d��m���ԃÎ�ơ��^��Z��E���ڀ�{���OD�V>��}�ˀW>�����9ŏ���;��-����?0�pݬ=�������ON���̿}�Ύ�ܝZXh21`]|�Ӧ��w��'�����zEE�c,Ny�`�ʌ�D�km>����͛7�F�������<�ܲ A�m���[�GL��:�!'\Pa��x��$9rY��Ǐ�̥�R�]�����H���x~8�8�����	&�&��ǿ�9m�nĕk�/+�q*^W���X���?�f�Q���#,$�G[����.����ߗ���x��� �l�:M�<���6$M=!"*�
|�?G2,�.L��	~�W\��#��Sz�L~]#Q12:z1&D�f�+c����m����ݖ��P�N����e��A�x��9r�ѣGQ����7�����!��� ��'!w����|�E�����),�OXke�eKy��z&�ޯ����)a����9��^c���>^j�03�~�����Y�Z�u�l�w.ã�<�ٌؙ>��X�lYuA\�'�r�.#��$�5���������̡Y\�����ލ�g ���� /�2utrbN���2��,�
��y��
�qtt�Cv�����'zS����p�O�h=]a�!��o]'����:_C�4�P�R�v@&݀VM���۠ڐ]ɛ���ޝC���e,�N��N.9��1>����x�(��9Q.�k�B?�m窔�#�dN�W����Ct̗޺m�ggƸ�I҃�W��cR]����Y����|�6�c*��M.8._W������%KT�75>	
�?�iR��l�uy��j_㇂��
Gww���V��_�Sg�'��&����0Ǆ���fkx��y�t�O�V���{��c��_�{�Gz'>�hzz��l��,m4}�@�S:�Is���~�]q�?/�A�E�)���J��}�O�##��Iˈ��ѹ�lm�b�~�C��{_��J|���9c+Z��%�i��2�{ڃ������X����`B��TI�DV�5�u��IB�E�����x�~~�J(2���6Ѥ9a�]ݱ47]��)\��Pk #` [�[��m��X�sj�g7���&����/�����/�Z+Y|���<e������S�X�Z���H�W�<��D,}�?]��BԘM���!�ZQ���|+�b���j?�d������H�Bk9-?'�9�������A�)�i;�V9�4�g��QOu��Dk`���?�S���a��^�|)(.~; EٛNkN�`�_���A�Xק��Goc�CL����u���sm�������Z\�e�ݿ����`���X�ï;;�s�lx
N�yf���_e���Oה֯���-�
d�������� �0L"2����ã�Ѷ�X�뻡`%l�����p���*,���ӏS>@�ߢ@� eQw���i%��,�2�a���Ԛ�~���q�w�K�v``�8�A�W��SwRۑ���<��to�av}J؛��2���S�/�!�v#􌤙,�o����1�TG�J���[s��4r$�N���_�C�b�)fMg���^)P��H�'��3gμ�Kh�8ƨ2B�a"�\��q�RҤEq9 N��Thm��e!�|����Z��^S/�lw�f�9ƃ"*�`��ttt�p�\bx!۠�*��g���?c�|MP/|��G$���g#ӵ
�w�Oj�k��⍱����L��ze<���\Ƭ�E�k�A�arH���;�0�i����Jh�qQU3�=˨\8�i�$}���Y&��^"����$o�����=�j%�qH1�`o5��|�k��^�>uU�̯*e��R��1�VvEU뤞cL"e�{%�&�~�)�C8>{�g`&l ���5I�i�Dԙ��?2�'{d�w�~�p��b�rFk�l�	Z��xç������a<U(n*�o$M�+>��1�Y��E��
�������+��d2��`sxC�Ŗ�xC䎔K�Ҹ����5�.�C�N�! ̍Т�B�c�A�l$,�,��$�kAK,�Ԉ:_h�y�I	�ʒ]s�@�rӜ����+�LYմ�v�D�W7�� -U^���K���"8���tV��"N���rD����_�`w0݄�V:�o������2��;	j�`+�ǵ�+8����c�/YZ���rB��Z�K�~���lD\kK?6jR��k����+=f-�6���JX
4p�?~�������6t}7�\&��� ��y��t���U�u�����? ���*���c�W��v�^R����*��=���c�ب{��;����b.ChNl-��ݔ�j��f�y&�YTJ<�
v��݁�{��3*� ��'s/���$_Vq����O�J(��X�OIS�8�����L�̌ցt��fc�IA�"m:^6�(�ƎrbA,̚�č�uww���`�噱;v<����bߵ�)uԌu�ηč��;�_he8�"δ|f�ɋ�f����R����O,��b��F�ϬQ���O�$ު�`����w+�SZi�&("�t�g����GP6j���q�ꆏ����U�!0J��Э�:� F2�Ak@XPPwz˷��al1�3�d����{U����*�|�yl�ڋ'�}��,��̽�V�iӇ���<����P�+!� *>!!aŵZ��죔C֫��"�g���se}�,y`2ҵ�����♈繬��ò߉|�z�I[�*e0��!�ρl�����#�x��9���Ǝ��Z���%�i0i| ڕ���gdx9I��Z	E~��Z43�n%k��M��+ ^��9i�)��0���/��7Nb��0gAmijk�~�05xh�J����ʊ u�O �H�1�	=`�~��4W�:� ��Ev%{�7��f�q]k*�m@` �<�:ᒃ<d�Y�$Bn������y��'�����-^�v��j����iXrk��e��=��
�k_kA�� �mDg���Ֆ���T���Q���szPU�P̫nn7�����j�� $:se�LO,|۫�p�4Y9J���e�5�ˮ�=�t��qF�LWc=Ǿ�Rt��k�[::��	�!���	�2�s�f���zHVn�Q ؙ�r��(�<�c��=���,��		��A�,Y��bG��=?<��b=g�;�"��I+��vދg&2Ņ��LZ�>��:h���R�T�5��ʎ����9�Zq�:{oFL���Q��kK����G|[U��3����'�V�E��^o��]�yA����%��ep���~���5�"w&�xn��BEM�*++��*���++�t���>���V
[�����hG}N� �Vj�����s��s��/�z��j�ÇeQ~z3�MßBBBH�Q�aXB�(D�|���O��fDb����[?O��f�w�t)0�mϋ�V�ӊ�kxѓ���H�jg���2_H�!,"��c�e�Z[ooE�v^_�g�Y�T3�2}�:|7v��3��@^�����=�v��L~Fp�nan;��CCC�߸���p�m�ņ�Xu�׊	5y�dZ\�Q�ˀz�>4r'Y� w�0���3)���G�	�/�w���[����@��C�5,��Y����&@��z *˴�/~��y׌�v�2�:�`%4=
!�n����*B1�g�e�/Tg��B������Z�`/mpk����[�2��G�P��B �~�h~x���S$W���p��niQrĕ�����x��`;v�	�����C�3 �;���.�"���'ѠNV1�&l˱����{��9�^gpd��n�
x�	v�gcg���};��w��ࣤr�\��<U [��qq��a,�����a5u�ŦB���8����f�6�L��s���
��7��2��71�N;ԝ�?bk�Hql���X����ʈ�6��z��1'D���;�V[ j�A���ͳ�|{��`t,����l��c��y�dD!�Hp�������f�n�� �/ 
����b�NZ�n3�l�Ś���euQ�e�h��(a�� E�Xy��5̀}���P���B��c{�����'�	`�T�8$�?�c#�S\a`��5vAA�@��Ǿm��a&��1�م�J0C��K�9ۻX�c��H�ӟF���&B1
���n�ʳ��c���J'��B����GRٺhZ��:~��)�
�]�v�3R�ՙ`u�m3V�x����H9,�k��5Z�FZ,�a5���dBA6g�.��
�#Y�[�}^�q��:���r��)'!��������������h,܊�Ϝp����#Ǿ6
����� �+��mutt�F��8���
��3N�f��Ԩe�>���J6Lr�s_���M�'�Q�2W�73��P.NNl�����V���?'��m�"T^^����P�XvycE�ɪ����Su�Ũt�D�`�&^��+�Z�m�\FPo�&qU��xFб�_=ܟ6�`T����us�l��6Fm����𺀾xx÷]ha��?ݓ�̫�n���׶��`����Y�8�aI����ྰ���4[q��W���mٙ!O	[��N�FZ�v�e81�����Y��1ܻ�^��r�����S��p)l�3+���dyE�+p����w%���U��e

��p��S��l�f>l��	+�Y��R�"��:!�F�)�k���:)Ǳ���������m�j�m�J��l&"�>M��}�7


�9$H�:�P�0Ya�S�	mq�E�v&� ���h­�z�X�j�n$�H�	 v2V�D"Jjj{��5�gī���Q[��K��	�w�bo�>Lb�����`���-+�$��ͪ��zS�-�?��FivNN+๊�؁�FӚ[�v�;+ 0<8�B��=aIm��_�JN;����:��h��Q�'#D��ɐ��&&O��hT����tEEE^P$JX 9\dL;M�Kd���K���1pF+r[�#���-w�x��M<S@��j���Ә!}U@7�:8)��4�b7�(����h-� >�	����qk�oΰ;xP҇Mq`d�K�]�^y��x�����HL8�Cv]	Ђ�i�s+�A�A��@�1�n�2�<�(�ܵ�e)j�ۇZ#G�r�D�r��-"���s��It��֩�
3X�g�uWyn$	��-t�f���>�$�\8c��~�������]Re>��~+))	{�!��߀Φ#*cl��=}���6WVc�� ��zʎ��DO
;�Y�oӶ����^�0�3����\�|�5�_	5P8������#�z.��g�C*~��Q�?�O���z�G6>�j�bK����B;ʽ��j@��A���:���wz�Z�0x�౮CT�vtt�ąr�؛\�) o�'l��
���[ɗ�}��ϨU�iǣ@�{	`�
Vl�	��AV-�qr3vnę3yY��O�3�-H����w�X vU=��j�	Uە�6	��D�$N�H�՗��9�a�i\� H. �,  �)��F3�s���&̟a��֬��7ia׆-��w� ���ᪧ-v�255��&���1:�G�V�����ؘn0�������(�t�]`H���y�&Ҭ�E_�~�Ƃ��틲��oJ� �[R�b�GY�����ts�����oǦ�e"s�>+�9Q�f����23�!�J;BJL	�i��s�:��O�GV3��2��`$�r���*�p+�T�еȥB�KԚ��d����x�!�`j������!�1�
�>0,/�1��896ޫ)~�X�ts��������lق��Ţ�$S�2��=fv�����h�M� ��p��1�M=�4Y	�WX����㕭h����#��:2:px�k����o< �E�&ȭ��dLz50��72*D�W�+�H'z7�O��E!�׮i),�b���|ћ��%Nd�(�X�N;	~�_����뜕����1p���se������ p��h�އ�v����|�+\zޖ�oW<�^-��D���M�H[?��f�j0�zS�~��j�� rlu)��%,B��='����ַA���3�B�Ug����?��9����g����I4'�+	�ɣG�<����y����K�������1֘xm�w��_p��ޓ�w��h� � M�¾�I k��l�VN��� ;����	���y�=���f��MMN�+H(�ps��ϟ�c��u���h�1�1$�"���Ò�3S�C��<�b���������ua�	�cJ���t���ߐ��ERHHֻ����̹}�������3G�?oq�qf��@�1H����q}�z·�)�f�8�^i/��`:6��U���-5�6��&�/���X8ۓ6���X�ct�f1�-ja��%%�w�=ִH*����uv6B4���L:d`F=}cA��	~���$����u;��,Ì��pw◥����5�m�g���`R��NΜ�����dQ��(al�c�]��y��ͫ��g8
���� mX3~=}�t��A/y9�HU���»Ӎ�b�Ep' rs-,�����Ƈ�Z[����%��vN��~����R�2������T⹨�	�����ۃ����z�!G٨��:|��,���0e�?�5E��΀�0��\�����y��11���1�g6bbD��-����d���0B�9h�o=�D�fv�Z���X�{��(��\kjs�����䛃PY��.����w�4���=���Z������([:�}<6��>������[�Ӵ��E���b�J��oP��$��Bü�R&�+^�޽{�>}��~��݃f���۞Ţ��1_��El�η3�%�}��+��"���tɕB"�{��tV�<g�s�;� �N��7��k�}�.읁�M1�ZI�<�������V�'��1�71�#� ay�Ϫ�132��`s���^/[Z JP� �D��s��@L��K��},�o���g39���j'���q!!�3�A`pաء��u�ò�,I�!�T^\���I�Ý!���o�r��X}�֍3Ww���(�D7s"��F�����[���#���ۀ��8�h�J�G��UL�HtF:�4"D�	�� ,�e�����\YlɊ��go�6���q�ĈpZ�s0TAHÆέr�56�	Wc�p�3�Ȼ<
�kc��ao)�O>l��,��g��e[��A�l����ӊg�}	�]P�<�Ӳ� �:��e���$�6�sr����IWά�9V��<0����z���åd�}`��އ'�f⪦-�����F��J�Uf-f;;�AV��|�u�aXƙ{�S�Y����z��f��"�X�Ǽ�`V�� ��:��^��b�!���b�i6�����cSv�#B�p�<8�mH��i�賰��5׌�-Lk�J���^����Q�9����ʊ�l�Ӂv�}�V�y���$'� �ʏ��(.l�bx&Y�����Ǻ°�i�5G ���ʿ��B����`_Zƽ��2��_�V��T��hF��ꂚG��t��ޕĮd`�ب�\:�>�xrrrү/��M�t��M��z�?o�!�f]U�Ob���0��߅A�������bj�w_�r���Ǚ�̫�@� �֊��K�ut�O
X�&�m�' q�&E��ܩ��P���^s�!+{�p�ģ8X�̜���6�3����2���@'d�>�#�9՚J���{�d[�]����gk8'�1@H�!<�Z,�#�Q �i�q�/z�����ζ�h��|�x��V)\w�a�2�y�=���X��b��ꆆ�$4ҍaTJ `s�?��<�
�{1�����G����x��C��{���y̆���/px��Uk����ث��z�77fgY9Դ{��E+�[a_��(��khL>��fu�V���_�o�0�������C?��G��4J���(M�⺂�Ʒ�Ko�{��gZ����"�:ܲ�Y]�Rg/��bUY��\�Y�?�T�_�����iuLN�Ǐ� W�ip��y�)i��gx������`؛<��}M�**BxԨ��F��o�85�5�N[[��O4��*�2�C���L%�ōWg����11>��ގG����/��~��^4&�RP�9~5"�Z��&��e�Eك'�^��m� �>P��_���9rD�>�м��7/djOˁʹ�NK��W��*}�n}
V߽��׎��S㣅�z�,��h�8fH��>bӠ?�S�O�&`��zj������\o����nę3g�G��׷�RjU���l?��.-��qr/���(� G
S�_X���\�Htl
X�Ǻ����"�=w����0�;{J�n
j���x�\���
�2@Ew��ġ�/.��X�.݋0�kL����e��7o�#��<؛[��M���N��?�ǫ��yvt\���3��|�"�8��L�|��t�@xż�)�޺'s�]]��<�
;����� �h�%��rMUa��+��+���=٭ ɦ��c�;::�F�M�]���?i���V>����B���t��	���vUҏS^X�������� z����Z��[����x<�Ss�t¿� ��>p�Õ�����q?d��S���u�+�؁��+l�'���j�s�ʖ���=��I7�
��z����{R��"���>�!2Pd���HYq�⏄c�N��Q�kş�RqD<��ӧ'�Tk�4���.EW�sZ���-�>�a�� �p@"�<�# ސ���޺���,Z[qG�*�/��O�/`��?x��5��i�c/Nn-�w�0b���~��@��!���q����3 �x�u׮]A=[]�.t$�=�3hb	fb���<,��v���|@1:*��+[�x�>�l�6�
��w���^��Gz�m}
�*��@�)�t;j��w���G�Ѩ�@w��$�$��ȥ#�������@E"~v�h��=�z|�+ׯQ�Sʒ����!��ޛ����Ii�b�yĞ���,���X�k����!W������N�gO��ѽ4B�6f��d�$SO�+T*���;֩=E��[vD���Z���L�Q"�!_�x�/�Y�w���Ɨ�w�i�Q���W�~�J��C19���Q^��ٱ&͉&e���@��o�!��ʔ��e��
"�YH;��H����@K�6�\�|Y~������	։��⢢�z��ކ=�������̟,�m_�]�7'E�;�R�>�*�/�Rw(k�x��߿�G�UVV�����
o�7-=[�0����py���c��F�>H��X���hZ���ʿC��'��MX_P�R����z25�g���J��"7,9@��G��AQ[[�����x�l�hS��]��J��o�@��!P�79Ih8u�'*8�CN�ih���)����p��C��4�v&Sl���=��8nȼZ���R��7&ዀ�!��=>�)�L��J�R�y~�O�T�o��t�џ�H�xI��y9���x/�`�V��3�!M���gv<��N��U�����
��m�U!�:����j�>W��9gqK��ʹ>��˅����q������\�m�ǰ������v�������C��)��+1�$�cw/�;9k��� ��~�냶�Gھ��{3P����)�oT7�U������Z���6h<�i��%���d��ǚ~�G8���+p
^�.��3�ߪ�b�������7�zh�=\�c��={�<P=Y~��Y��q�6��2R)���D��8��Zc��>^��#bu��}���fY�C^�����{q0BK���'�C���$��}xp]zW�.NN'oo�}�ҍw���P�����mjo�������6�����/�Ic3��;wd2��3=��L.���CP�W��;&�|��X�$Q�����w�Ը��k�b�v�̡�CN�3�Ni&��
�,D%އ�L��w%)�
e���S�^<�BQM-��I���ķ�뮿z�:ܽ|���e�d��Vel��FAN�5x3GS��@�����;$�zA:}���O֓��8�*�?E�ˍ�u����7�����!������� �޾�q�\#��d�����o�I�{^�x��rM���P/e�T�,jyb}Zc�!$��9���I�l��0ܼ{�[�������h9�ʁ��G!M��V�K#��ŉ�H:'G Y����6P�zB,�|%.Ж�\�?4�J�� Y���|p���1cu���ʢ�ᇅkך=��`@��g�AOOC�_5�rr6 ��({��m���)4o�l9m1�V,I8:j����E].��6�� ���C �A 8��P����e��W^�QS���L[|�~��=E��H	��φ1u�o�2W��C���x��x���X���D�� ��� `� �@�z�Kk��d�.2QQq
�Trko�w����_���(�V�D���~�F`��͇2�T�G�ȶ���}��.��̒��6M��O��=�Ѵ���e�%v�\���4����*��M�\6x��C���ܬ.�!��{f���oޘ%������XZ�G��L�G�b��q)<�+�NMM�US�k�{�Ň� T�-�<�GZMfϺ�p�OYA�~vͱ��o��Pm~}���{�+�z*,�/����{�/��9����\sBΝ���dne���Շ m��{-7wh���,*���܍����s���ۼ�4��Ws���o{|d����c�N=R�f˅#�\��jdd4���oP��[E����o�(�K�Y>�<��ĥWw�a�2��|��d=�իW�=���M �k߆��Vbk�E����/�o`9w'E���ΫL��[S!��n�0c�F�
M��@Ugx��v�k�?C�#�t4/��\�
$-�1��l�R��6�o��b)ؽ�V�#���ۚm������
b>�}��<
7��TZ��ԇ%r||�cbb���<y\-611��M}pjN�<���(w�s�$�P?�ɛ�*
�E��Z:�a�O_�r�l�:v<JK�1�`��
lnmM{�rϋ�ϫ���e�c�z�݋NQ��o�1�؛���e��w�#�;8:�hN}�<���9�8ٗ���<��o
2�	�|�W���D��Հ6���@ �c�����哓�.������D��gVev�(��{�\|V[���RS��-��e�үk;ӛb���&�/7g�`?0�� ��'��6aϽ��։�������Z˗/OŕS�򋻤|F�MFFF�mm7���3��3���Ibu�
�ۯ ��.f��͹��#Oߺ�����,]I[��`��5��n� ������].>y�~��T枟F⇂tJ|�6��P��.��+�k����k�^9r���{i]���~�"���\Ǔ���1�>����p��E[�43���Hi|�*����A�azS�LV�%W#�+ tJJ��_zS�'D�܊�E���r��bq�;w��ǽ߾}����R?P>>�1���a�.m���x"+3h�~�n!����ڵ���^�&��� ;��/�~�d�~x�(l"u�l���#���|�R�klhx|K����C?E��B�w��7e�����ޠc��M�4j:�i� ��� ��$5?   !���нշ��~�㛚0���P��~|>"��WH ����=����u�m_�`d������X�v�<W��-�~��/�&Bb;��Fl�g�w/�;�P����~�
���δ�����ڌ�/ޙ��?8���=�M޷�/)2KypS?��s�m	.��������U��oѪ-[��V���pD�}i�1PO½�U�S,���s��X�m�֏�@/�c���K1����F��y���Jv�x�[�-Փ��ӬT�7�����v��I�}l3��G#QV���}8Nh[�9D<���((h�(�L�-֪���oT�WO���_}�o�H� wT$Q���~~�j���"~u�qm�t�~�:�F�������;��6<�����lx�U��tYi_�@l��=�reAs j*��.ޟh^�{'��'��7���q��)[�bU	��(wۗ�5�4�nQ�8qJG��W�үg��A%&��+�������C�N|�+0�Q�_Ɓ�E���������mZ*����+=9[p�U��s�<��,8	k4�۷o�cr����zn������~�"0�݆=<��9Xm�c�TC�̓T;��ي`gh�l�v��IIe�o�ؾC�2�/kI�3sW��F�/RI꼴>���!���ǏV�0�&?z��p ����f7����b�
[��j&6������
�[5��1����?�5���QҔٵ��X�ʓl�l���{��K;����%0ln��r]�0lA�_�����g��aٌ�V�֋�t�������V��~�b���/Gb�0i1�xt�RUS[��~���ڬ�l��.Q�d ����2'�kP9+l6n܈�3דU��R�˿��u_�+&"ף�-�-[���5,@�N��(�޹>a�o��5;�൴�lc�L @�S�[N�:��8�EP�!,]�Y�*�@9�X}fh��~d^v�贝*�V�2DWY	fXX�_b�u �wC����]'�2�:qH�AL�(�3�ZP�xb�I�9��<�'�*��̅!�����dSC���]� t�=&&)CA�j�\]I�~6T�z�
X��(l? �x�9��8H�*y}W����}}{d��^M
	*"mx/$V������N5s��(���C?4y�oL�hvr��ց���Y:b�[�\��0$d��k���`�.�8w.���"�]���6�f#� ��򐈄���IH��g���+h[��r;%e�cmZ��%	!��X�@���9P���.����M�m��ނ����~4*<�-U��P�ņT�X�7��t�K���R�<��kc܌;����c�;��L�nX�U�	J4�dQ� eH��"9)93�"�JIr���$�Y@�9���'����ǳ�Qf����n�[]]Mـ��p�坽�0H�jۧ�=&��휁�#@
��Dn��Y[ZBq{�a�fg�w��δ&���}���a���H_��j xm���JJ��[+P���������/
�j��fh�b�U��+�*U��?v��6����+Xmym��?){�ȵ �4���F���9����U�!]R�m'T�Wl	_
&�+U��y���N|���=�9��>���f1�kN��`�����I��W/�g"�xh#c�w�H!��]��Nyyy��i{g�'x�i1 ���]oϡ^\?_%����U�N��`��j4��U���/'�:�������`Eݰ�ź!��w��gK~��y�
���b��U�����ͥh`��]��G�_�Y@��	�`�.e 5�����x�)�B�Af|�0T@�F�nA6����r�%��� :8}4a�0b �e 6|����2�I�9N��J��E_\�������|Ϯ$/J�z?�J�� ?�J�ؔ+ @ި
<�lL����뱿(a#m���[{��{���˲���v|Y�� V����Q���}o�e������ 0C�����ǏM
��d�z����g�GPكs��)����\���E�������|	�s�y{Պ]�[���Z{z�C�v>@D��eHp_mmmD�C�����w��6�MOW|/n�ng�#���y���t~��:���2������N�@R��Pel���k��iUxG�S<�q�R�2�nDd���>yBaT��:���}y��ki;�J��cכ믣��p$�S����F��Ҟ��iMM�Ʉ �9t�]iQ���:�/����uE"���*�F��0��9#��ϟ?aC@���8��g-U�'���g��:���n�I/b@� �3�:vI�[���|�UFc!lO&�����4B ��BqدJ'=���p<�1�齄�P��~�/R���{��6*q��!���
i&��%��LNN���%�7������k�G�P0�a�|��q��)P�9|������@W3���)A%j3�S�JP6��i�N��.��8�~��;^:�y^h��~��HB�C.X1�C�i�����2��� ��ځZXc�[bN�� ���).�������Tٽ� �F�JެP>���iH�����6g(������vnT�@6C��<*ג�3�E"��4�&��I�8��N���-J �rO[;rh��Zg����g�4���^}|#�q!�8\��^LB�����#�������˗�QB�'���z��Z++,�A��&�QS�_vP!+G�vg�7� B����Y�j���=z�Cv"M�VW�?"3���}6�<�/^�B	

B�70�)������(���1�����֚o���a!hX���@Y�77�T\z���M���P�1�40�	��KJbQQBX�� ������HZ���F.VQ=���.&	
</�êCR���`�=�&�}}|!�� ����|ow�9�n>��C�*4W ,���dj��&����� !�h߉������G�,L�z�v}�B�c������[)�䴰�_��a �C,,,J��-āW�+�S&�����g�߸���5�u��cx���;������
�K��q���
,�e�r�<(����.� �x=!/������~�CgExo�t�Tո. �a�0�	@�fg}�-�30R9S @�����d��)��Wƕ;�֝$um��i���W�~�������~���>�}�"d��e!�s´���yN�����e��C���$����d	`>��ɨ�Dc���}||�߁���)*I";�0�����L�"��zDRw�.G���@5@Zα������QUh���C��/�F����oW�TÎa��Xd$!�y%�H��7��6��\����G�3�s'`{Z�K	f��N�� ��}� �z��������\u_���@���<H�ˮ��㳧�����.��uN]���� D�L]خ�اpf{m���˰�"���a2hJ�ӯU숣�DY���*���,~��^XЁ`�mt���@гk����*(�OP�����yRԢ����A��'�؈���� 
��z��8���M� /��"��PƐ�l�wmmm
�hR����I)�Q:�6	DR���,m#�XwC�}Pﰋ��zK�T���sG4����5 +o:X��a{��u OJ�����G~�ػ�N�		u�·�'�В���	,G���|��
-��_ ��l�u�����P �@̀��@J�������\t2Q�@��KT\��I�b2�,�]e��wuYW��8I�!�I
��A1,,,%���7>�R��na�Y:�F�;X�E0�`T�t�
�oÛ(���;�Q��u++Y[[kf�ק�Q����y�+ѯ3Ka/bW�.gZ�S�Q�b���Y�����,L�'�n�;:����5�����_r���q����� (]J�7l���$Vo��>���y�����I1�޵vvj^؜t����Ot���#�� �!1����$$FH@X7����v��"���'`+� *-�G���F�p���Ā�-D�����6M1b�bG d���C<��M~"��b�:;;��v@�������O�āG755��O�
 t���г��wDxxZq��z-��x��ߪ}0���>,�t���Tom�Ѩ+q&M�$������9m g �O��i������;����`�C:����|
P���|"�,������ ��_�|�����ݎc=��;�מ��\ȫ��Qg)���r������+*C/���t7d[�f����>Ϥk�X��}� ���<����]:�΅Ċ
������ِ#�'��陙�1E��X��2�q\]u���=���a_��A4Z�L�F��sڀ�Nt�1���~���<z���Ψ��En�SC灷�X�~�n(
b)B༯7���:��&\:hY�br'��L��5�yp��7�8�d�m�YW`��ɴ�

bW�8�X�Zs���x������?�u*�ב�k��<��h�R3����[0٭�BAF��&lv���l��X��.�/����ܡ���˿�P�ttTo��;�@�Ng����qη��� ��� ]
<X޻��E	�_�B��+L�@��y�K��$����%�Z �28�3S]�_�*�m�;vjdh�))� .��׌<&�@���)�vD�=��_�5B�;B%�9���<�[������~yy��Q�0�.|�lO[]�\\K��\
�+��
P��a.ܵ�Z��{?�܆|�*|�
}d:溓T,�-�AA���<��OX��RIE��크`в��R���-�&��bو�l��"��V����C²xxdπ ̰l���%���f���o�����Jc�s��?c|X��������(��cA4�ar����J����M4�ml!i��mӐ§:�ٯu���H��f�='���cR���Z���.Ow��#��:�B;~�WS������f���z��nʒM2��4G7�����%n"E��yy�d�c�Q$��� �P��}��G���������y]\]��Ђ �:?�)*�8�r?a�X��<K��fWN������g����)�<�F��*ĻթBB"�pKO!��㙙��.���ʤ�e��l�i(خ�����A���ߨԹ��Լw�>i�g��C�=|�����@�{�uw�Q:'K<G��	�/� R^��F�Pc���<�y��Y+��p��3�;)��Ϥ ���3�a���H@D�	0u�:�%ȝ��,滉7ˡɍ���Ȱ���#�BK�Pp�Ѻ@� 8�<�<�Ȟ4�frE�L�{R��p�&�@ �^������n&���%�������yy��*�n�7w.8��\������6
�j����kddT�`�v��y���a@A�7�c�VVm�M�	���o��x���7�F���~� Sw��Y�%��ж7qm��y����o�r`r{�,\����%
�V����c��2�E6[O�[m�.����?p�YH��< X��pq���A:H��O��Z�es�TX?�r a��x���A-Aף�����l'�v�w.7x"""Rޛ�@����ʀ�p��n���M�_8�R���D[�4%���L?�@)�K�$bIm1�"=M�u{g^���J�&E(��L�&�l�c���*kȘ葟v���D��@��m��F�(�%xP�r?�㼿��x�/2�	#�^|��ׯ'�6��77�	Ύؼ�~�3�m�r������骓VO��)V֎��ʬ�����Ux�a�����߁�]�'�B6q��$[-()����S�������h��,�����^���<"��o�ʌ��vX�/%9��˱3@"���tD
�ɓ�F�n�TNB7t'��P��{ L��/%�Z��ߑ^�؂������] {#��^�{X��\�Fx΍��J��f;	c0��x ��?�w��ϟ�a2|��`����yҺ��84�9#C� �I��۷W���VQ��V;r�d0� �È��[c��޸��VUa�n3]���D��I������֖@/�\4�K؆�S(�6��*�x�RC^�����D1��Pɀ83b� sss�2/ ��HA�w"�L����$@
X�F�`%�K?Xa+�J�JX�C��q��DpssC�TVV�&NM�@{x�VPP|43�^2�E���\(߀j����x�a?P�0�7��W�8�q�}��Pn��Ʀp���lⱍ�? ?�`B�\o�	!�(LI���խs��%�}/;��Xܰ4���-������\�P��b�.�FTF&n�U�
�L/��^jr��6���<z(G�A<<�_�,z�%�.3J�I�P��N �:��Ba���m&҅�ZzzV$�%sP=%%��ɶ$���p�27��U��&��0Q��x��VW����B�J0�23�@TE�`{��zmw���#� ���HK�����^CJ�+&��@�wi�ۂ��iiJ�(��D^BX8�%��˙��@�7;�S��#]jZ65X Gz��w�%��2���cv�U��M���__�g��T���6�� L�?";P��` ,���G��*�i�Gڒ�����qqp?���aA�S�ɟ�
UI��XlV�Z
q��uH����g0˫o`@H/ANL��p��=�a��#(0R�ٰ�`��T@!y��L�r����|�e'�ԫof�%����,�92b<��8���1`_t��񪦦� ����^<��Z���g�����wO�k-tc�K6����LtW�q�~eK�H!x9�%w�����&Y��nOG��Ȉ��B�H��F�l�_H>�� /�+�P��Y�P2Y��E(�(:DA%��R ��Qd`߂1*� �A(��e�q��_R�!9��!}�~���0l�
�Ɇ��ۋX��.a߳I߽o ��ȭ��=��m��-S��W��[Q|(�N�Lr�����1�(K{��Z��u����4�AQ3yI�Q�j��w�H�"yS-0Z(P9ЅK�|[���A%�>����R�wkO~٣|y�l��g���Ծ���t�`Z/�cկ=��U���������W\a�<�qp��a�����Ty�ޱ��Ur����G�b^�2���ֹ��O���^	ȸR;�} �p�W�V򨯐G�
h9�wu���,�z�,p�#�+��lTu¹8��jj	&j~o��P02oi�^R�Z��չ7t)+�G���š��Ñf�:�QYu~���n�8�]3a.v�UGZ&���������k�@����*�x
}���@\��z^*_�����4*	QϠg�c�_R�X�L�85�϶,%�!P&���R8�'��u�ЫW�Ǚ�O�h�;s&?�3)�j��֫Wc����ǘ��n�_Y"٤�:�R���#�L�HY�����\T��cv`���
�:��<J�<���ϟ&���y�h����;@O�w�;���n*��JS�qF�P?ф��c5?��?J8:z�N�4b��u����N̨�JI5���G�X^e��˧񛚚�#a1�)�8VDv~h�'x���#r��<��H��NZH�pce�`�k��ꨓ�r� cɇ�L[������� 3d��y����������Ⱥ��6:!w�e?������\�+,�[��K/�~$j�pp�<�)��
@�2�cϨ�`"�Zb@��o�9jhl7�c��>�����e'� Q��������|����2ñd.@�h#�8����<~�D�Ƿ��V�5ӧ�����ob�=��{A�*��W��^�-��VTF��gs-�K@���ʩ����Hy�<�+ѝ ��e8�E6ڀ2�����N{h|zC�-��z��Pz� E-6���3b���gu�Nǰhuwz�٠)	Ơ��dm��������:j����Ð�I���U�|!�H�kR\QÔ���M'�I�d [h�P�.��"����vz��6�!:S�Xi_�N��2Ӗ��G�����[k�����ݲ���RR)�s��?W�OHX��[hτ8e����4�����r�dUWH�U�0\(l��������F�%ÖsM�x~Zz�.3�����5��"�$�5���f�\�8w�}�a'GXXY�['��ݬ.��ṈT:�[~�I����jc�qC��n�L��,���> `���[F*�TKIiEF�]��>^~��φOL�h���D���������*�2�[��7��W�5�X�K����_�N����5�f��<� l���]4�'�F�I�g�$:�4�����xԘI��]ӚuM�Q��/�a������L����������E�Dfٞ�A���堠`k` �~Nj
����^�ee�$��5�D�z4�(*!R� ws��Hw�o��C:�fGT R���������5�X4�Р��#����Q��i�j�q֥�++,��]��/�={6������rM�U�x��XD) �����LN���:�8�$[WW�"�㍬>�X*f�v�q�T�@��n�ϟ���Y�����Pє&B�nX�}kVm���XE+Go������X���V�p�邺��*-"�?Zi���y�J��d��+�x2�%��Y���X9��c ��ڣΆ��<�@��7h���\dV���7�(bN��lh_�g3����J���G�B)����J%�~�x��������sjD��+��&�c�B�ވ�$8X�^W�Cwi{xp$�֑g��`(���AQKS'#�O��^��yTuG#Ͱ�s�"���p-M�E/_�����5��ε'�YB�x>��C���|c^v��z����?)�f�!�!�o�jo@�y�0�8�bicx��e��\� U֬d�)Փ��<�P�֪�Jߒg֘kۤ�I˦�JϾ��Q��m��Y^̗�w�����/O�Dc�[��,�na��:,�C��GS����[��o��Y�;M�^��±�*�:����;c)u1_o.�1��������QQ���%Ml��/��-TU*�~.�K{n�p��ȑ�B��.��Å����,Z�u��5�.L�nIz~�h}����f�SD�u-pu���XO���ڗ�(_����pA���L�C�]l����LU+�"l��������ѓA�_���	"��#���%��2�2Ӟ�JA�t{آ��),aT/W�,�������;��
V�b��RB����Tq�F�s��{�޺.������?e�)��b�������t!�D�1P΍�*?�r�(J�,���g�Z�=�����ɺU��F�~.�p%>�J���`o��Ʈ?E�¤%�!6�@Yg�"�jx��խ�G�f���Xg���}����Q�������	�2��J���S5���~���U�%2���^�����ʛ�hS t��*�ۖ:��*��ٓ�1m{_=�\[:"��bar-��NH�����ď���"���D�d����s&ǌ�y�t���v�66H	����c��h`�m�y|�~y��ܬ�oV('A��>=���"{���ykc�fD�Lji�A�o4�c\���kn�Tт�4���M���4xs��rx�4r�Sc���Hz���!� ��]��L�C�O�^W����b��㛥O)#��Q���9ؑ��Q&�ӓ��s�bģ/��e���"ɬ�'c��m�%�a���l��wpbS��K@�&��N�gD�)�w�k���V�z�/z2l8��R��W�M.�ķ�����'	���@Ȟ��8�a3{�9��ۋ�M��S[��-�WKǵ��y�5�_���P�Zk���VYi�*��W?1f���!��*m��3�q1*_�\;�ؒEg���X�:7�q���/
sH���9ѷ�\��6V\�p��Vʪʓ}����ˏ5�i�NIW]m>�� |��� 'N����sԃ*�$N�<�=b�;nkg��x��1�<UuY�X�V����oDӏ�dwť�pڃ?Q���Z��*�4NB��=��Qǘ��4�Tš��@���4�}��H%S�l� �l��lO&���њ��	��'~s���Ri�|���C�w�37�$�C���Td\yu�_��L����$3YGL��C���� �&g>�.�����)��&��0>�(�⸓���V����XM�+�+��0���5�&����Vg>y��o��*�[k	`�=��_����W�N�,����j��O��CT\�����Mwl�=�(���%��>��I��s&&�v�I rJ��U�e�k��hT��?�(��;���n��\���6[G4���z� I��礖[��4,�[�;������<��F�&Bi�.Gww��[~����0\!�fUŃ�7v�T>2���Y}�i��G�:�}��=�P F_bT�1��+��}]�i���,:�C��]b�����c�^�^lޑ�/�.������G���l;���4xm�6��yF6�܂1�}�@��-ik)�%/ƍ�#���O��S!\��썔\�H�Z�D�wG��/ֺ�>P����Ko��"��v����z�R�ԸH��D����%R fx�x��6ְ[,����ۢGC�xA\<���[�at@A|�EEͨ���_S�@����e2���l�ӯ����;�;>��C8\��5s3� �R�!���ܜ������_���w��}�:����SL8������Ot�D ݗS�
�^��Tϰ�2�w
�9]����T;��,P�Lc����,�BV�2����I�q�իW�o+&����b�4ClR��$�"�?G҉)�{�r��{Y�o��r�������IӘ��:�Y����Ԋ����
��1��R�@,�G �tCW����Q���)��9'�e��U��F�IQ��Mܳi�wnX��P�����T7�O��؊4{��x����qn{K�J�^��y�Å45Ӯ��:]U��Eg�@'��W�e'�l��2X�i���-杙��ۂ������9���[;N�u��}�:mM�E�"�>Tz� �����PD"���S?Z]��IN�W9E7��{nn���'U�
=�i>�J�
�����2�J�&�9�'� �J��a\o��O���y5m0�&� ��7���7JJ�p|���8P=V��^z"'��п���g�`�`%�(w���%��W�/*�",�rqQ�?��z&�ag ��ͅ��k�q)'��h�µ�f�5һ��K23��u��%[������|+�5p�{Q����7d232��v�v�/���[��)/��l�잸*�βQ��31�;�@J��\�@�5���ϬՏ�5L\]v�Y��ز�9�B ���Y��7�61���D����ۭs#(���
9��S�.���.�;@�D� ^����w��=ȱ�:$w��V������R�=���hص�Z����IY� �h7-!&-�(M�(-�(M�-��&�v�/*Pb�Ґ��C�1��^/'m��Њ{Yn9�d�����LD�R��R���/���w�%���1l��2]��'Mt9��k��n;I73�2� ��/����S�\f�x��_�]�M�������ȕ�"�l�$LS����{i��ɋ"�s�;���Ҳ��m���`0����2c�(�,� `��9���-Շ���������|�+{�ό,���9���N9$㞸t-�n�,�P]�zvv���W�	f�I���蓵��)����Ӵut
�?['�yb��hh ��5ͬMcS?����͎���K>z�S4���˞z�X���p�<�w]� ��5N���/���)�8z(��1��V�b�7YY�Q�B%��ea
�uɯ�`h�	�]�CT_��~�� ��U��Ҧ^F㫘
��h�$}��V�o���Y&����=<ܒBl�h�s������jk�^X}��C��_cA0Q�gK��{���iOZ�@���}��aɖ9�^\�p�Wc�P���QVV��	->[��(�|�gB�#����	�Og�����b7�ucгL�+�9��}�)�T<��uO�bN�sB��Xl�ᯒ��/o����1%�m!��
��;��[ȸ⧶�7]51�on=ۘ����,�Jc䳛Ӭ2����z�vR'6�34�;٘ +߂?5�h�K>n)�I���U�"�ۡ������<Hy$��]�?�b�*�V��/�Ԇ�G���4���#��/�đM���$x��x� 2+e)Dqc� `�j�� e� i��o����럞dm�g��Txm5�Y8C;�/��
�fs�Ԧ���N3]v����+�|V�К��s�<1��[W)�rv|ثG�ir��<1��~?��q���z ������'&��K�H��iӎ	tN�<���C�NJ����B�#���qx�l�:���W����Qvz��}��lE�~x7��@��d����T9�R'v��5�x�ڼ��1b��sҳ{���0�SA;��ʺ�Y���o9���0�W���ӷ���w��7�-滖{e��%&�� X��"�;���<���p�g�H�v�H?�->����.�o�ɾ��xG��RrTǫ�R��`K��8��u�YI�)F�9�ff���v��������q��,�ʴ�N�D��R�qW�y���>���r;������__H3����:V��4�ބ�~���6I�dO�-2$M�����RN��.���B�U����w����'ؓ�6���Q����zZx�w!vn�*����s4�v����fD]`���ä�s��%$o��zqf�?�o�`t�n��f�̅�5�U�.H����!=5!G�"6]g�"������o������^h�{z{~T��d�����T���l��3"�/����,�#�Wz:�Cf���+ր��k�1���/�n�,,�3*�s�ڗsm�--!���U�<R�EM��Yg3��Ɲ�Vwu�\/�#��/��B�trr�'dǮ�m�/�.R1�F�b�n^,������4�v�<����8�#��x���c-�d��k�4?\ln�Fk�q���|?��{���|�������P[�2�d�s�����Ǹ�_vu��`|%��`�b|IK9�>��`̵�k�*��TM��?.��XЇ��"���±O_T\+�c=�H:�N8���o�zSN�����\e&#�����.��(oc.C�-FT!�[k�D�Q�Cu� S�>M.6�/�Nj	*)�c�y+�fљ%)+�MW�bW�f'�'Q�S5H~0�	'm�j����=��[S������l�K���mOr��ƬV�nJ�vdA$ZH���@G���T=.k�F�K\�ƻ�d%}gV�MԖ���S:Cm5�
��n=�[��9�t�SNM�gнYgf��ga:d;B�;��%���b�=,:f��T��x��1i���/�LFE��_��~������?�}`����0 ��3�v���Ng_���ם�y�ʜ�dZ��cF�r��bP�@�����@�0��~0�g�c/���h�r�̌�t;V|�o�U�uq������A�v�zc�u�4%�P�!G#��gg��d֫��"Ͱ��g
!؉�li������+���60�k�3���gy����y��`����9|�C� z,-W���W���H�I/��`;��?:n=�3�e�h�1B��z���`NY{��6�9 *��d �`�֖� �Ǜ�h�ء_]�`vL��g)��SVL������3P�.��}
�ea�A��\�j����n��`��k�J.<m�	�6������Ϩ�؃����������'{i`�����өy����;��O��k���8�s�f��8��B�$`/[� �澜C��h��+\ݮ�y�N�Rp|�����xjwt+p���W8y��O]�S_����Qv^ǣă@���<�1sU���ypg?��Nޚ��$�6{���v�9�����u�F���xI��hifZ�]dpP�n���i�1�R��G=�:N[,���β�q�����a+绛kg���Lk����<w���<cc8[��;f��g�v�8Y�.,��(&*���j�5�!�D5J�l�_�~���﹟
㓀?.���3Łu+>L��=qJ�
Ӳ�޻�?e�QL�+��a-��әҢ烵Y���v}�4�`��F'J��K�S��*����8?O��.�������2k��̺P�D̔�P~qqZ�EUb�"�I-)^YzN9�[4�Wb(Ki¼i��}����=TVt
��b�0Q��,�?��hc��\85��c�J��M�*uވ��"��h����^����� ��#ƿ�߭��0yasA?4�"��y��Lp�1�t��|�M7@.������g��#�fL��ڴV�5��
&�/6����� ����9�՞),D��#`K~nq<��N�����=�Q��r��3�cH� ��v����f�E��0����3�e��<�nK�r���|CߤO��_)7^wI�j�T޷wޑfπ	,�9���VPP�@���]W0:QIOwBE5�t�ǯg�,��?�d������Ga�����8���������j6ݸ' !l�M�'V��J'(6z#;O i���δ���q�̀��j�P���R-g��b6)nҐ�KC(�e{Պ�7��������i���L�6K��y������)�g��f�����#'̵Fa��q��@���-�P�����a���q��ȇ���u����8�T(�f4�d�h����R�vܒ	�Ɓ'}}�v���lAR�F8K�D,���ރ EuN&�4�� ��72YN�ӳ��֜�e�)+��ĝ���l��7���1�)(�7��V�}����,jy�1{����TT˂����W3�-��9TT9��D
A憘!^c�Q]����2�`RI�����F�8�s���L��x�.��";Y�;O��X�Q����t��v���'�J3�b��ơG$�ZE ���p��E����ƫ
�pٝŦ�&�z��kٚ���{3�ן{�:��n�j0<8r��}R��K�n�4�P/�Z ��yx8�D6#����3��+d��T=d�G�2���^c����8�P�u�E l+A���z�Ų5}�C]��ʋ������C=��oő]�����2���\��xЉ�f����Mb>N��P�������e�C^�|��qB�I��StH�9_��\A:.�kR��&s��0��؀���Fk+��9"ɺ =Ҽȗ�h[iy�����je_i��l�����F{�+FH�*�9��^�iŬɎA+��$�h:x'��f++��U?�v���Ii��������I���Ur"/�r��zfM'�IM4%���e��jYҷ�e�7��q%O�Ctן���%.pCr��u��>�B�� &	�T�G��P�b�iv�����\A,�l�Ȩe�n���1o��}6�$��t8[�e����{Ϣ����Izr�\/2�"�3ѷ`�'����Zv�;{����7����W+��%	>��?7Lr�X�!V��g�.k����&Cfe�v��ۮMuK\�����Uq�������?���x�B�� a�?1�T�OL!�Uo?���MTU�lA��Y0�`)ջ��ie�o�!SV���kb�H)��Qs�D����ª���kzm�_z$+I#և��W"{����� �e<3��8z�(\�:FM����Q5fvr�����QK�tA׮ )��$�c'a㙾������B��������Ѱ���M&���{|L��I N*��n��Te��@��ʄ|\��rj�y�	��;�<�]�Q�1���ǽ��JpWۻW�$NĻ�.�,��hx��Ӑhb��HGJU�*�Kkp����g\���]8�I�"��������t����y�i�ػ�J�<��y�&�!�p�*+��BF�[a�v�xz�6���/i*��Tz_�f�307�����P'�V��63�ʳy��S�Oߓ��"����#���2���kpv�3<���3�:T�x�v�JџM/����A?À`�q#�E ��T���kjY�z������jI�t�*�>\d��
I ���o�3x��_]��B]j�-��УZͽ��ٹ���,�R���]�f�=?^�`���<���ߨ̓?e)��R�''����,��u�|���
f��.;�}�_���J�VQ
��yrFT� T���͗�X_<ͶQ�oRà*���W*�w������x
�s�&��	g�M��t����;7�!�R�g1c��n����M�F�����׾&N }r���@��i
�Z�x��N{C�'1`���Ϧ�95��Hym��<p�ј��5�/>�l�R�0�3c�)ݨ�Ȍ�<�� �`�����4 nIea�?�1`VEX�ɴKL�b=�]���t{RԴ�=�r�7��V��/�#��a�?���c�`4�����ܽ8ͦ-̶U_iS��2�&�geLo�n�g��Ee�����9�0�J�&�'B{��=y���Zf
��2q@T[�Z���lR�j���;�k�ǻ�dߗ|#s)�f���ꆪ���O'�m~��Ɠ��.k�jO�)�:��������k
�P�'�G�<V�ÿ� g���y��S��SN-SK��-�@��uD�W���5Ͷ�?��FW�r�Z��� A��c�6��H�T��Mʯ�D��a������͸���)��IQv�EH�ՙ�TpZv�����[�!��7�)O��
O��ʯ��x��u־�T���`���o&����������]�b�ȵ,V��Afw�o�!�⾮W��.]�
�aQ}���(S�EQ��) 5 � �����B�մ���

��?F;�:)y�Z�֮I�Ƽ{����&�X��ĩ� 7>�Y"�k���9L |�c�	ƣ	&�)�Ƞn�������6���n�Ɇ� ��ȴy�X��V�@�Gk5�)�L�¦7ަM}�c^�b�K�4�m��)�[���B�z�TG�Z�о65-�01�����Hi&��h�a�iB��G������Ezp98r����/9t��VL�U��������*D�Дb�9��7��=��69D�g��_��)�̀-��:n�!I���B�Cj<�p���s0#��9�.
��/7�L�}��Q�M�*�G�c1�]&(�_'*����-��{NV�o�@i�QyPN��o$��ef15����ӫ�M�k�
����s�Kmg��L����!S�4����"%�ͧ$!,I�
�I����Db�ru��=���g�w@z^0]�� J����>�c�B�+�e>?ʯqFw���[�ϖ��fژ=�� >-�G��S�W��oɓ&����K�`�NX�N���zRP���9�c�J���\���>R���;-Ast����wx('��Y�;��v��}�0A�s�ӎ=�r�FJ�S1�QO�br(<�S1��ӤR3����X�[��F�[�H�X��7�r'���n��`��.iSL���r
3%���w����	u!C��m��ÿ(4������pz��0u���gJ�F����R*�M��M�x��yk�j
q�݊��h�Ĩ�qV�����^�?Z�>��5��":��,I�2�۫�w�ϾT��A'�)H <X@�%���l/۴a,�h"l�VUt�ٰ�c:�j���5�~攐�����8>��[���V���	9�W��_C�x}lz�Z�8� /��o�U5����"���j�*��	��9�����6�j3�u���UC�mZ�B�3�?�V�9�=FwH�sڋ	��`Z]����ȣ��ڱ<�lt����i_OO+��"uo!��.��Ƀm� �K8#k��f;�{s�|j}pl�sX�JOM@��v}�
7�2�������K��c�[5�)�򌧜�]�������S!~�Ie����#8�p�sUaLLL;XY�n�x�0dYC��
uo����;T�d�m��l���k3�CL�5�����Z)���.�o�k� �T/����m���2���o��]�UqUa��T(��{.KAUV�<h)�l��E9�R�{L�:O~x����A��Y���,z�Q��[As,���O�o�
1�Ƕr���W����v�>pq>���I^���uLP�}��ѵ��������[��_��|b<9�Ҹ~bSyB����t��VF�`������,��T`���r�.��igx�4I�}�SA"���$�rg�� ��yUL����7�v�M� �����S��ՅŮ��%�D��Vc7�nKS�l:�jLCD��p�t�
�hpX�J~��Ì��C����<oG���u��A��/j��'
*|��L�E�.F�JA6��f�*�.FG�~=KA����M-�L�{�h�}��/�y'��� w��|N~ /�+ϱ��	�vn�M��	��9W��mzӴR;�U�Pf�lLJf��n���H�IT�f��0c�bBb��>f)�kS�c���,�w.�U��	9�B�:�>Z��w#̀@���b�q�E�M�J]�c��l��gչ߻�[��t�xٌx�{�M<�UK(т��1���8�2��G�$�:�Zd��Iz��T�������,�#��U*+=���)�j(���]�LH�o9�0�̰��Վb���� ��A|��A��}l�*�V@ ~w-[,��tFִ?3���U�lz�����:��:������R����$����D>���zN6A]�
�^�QIЇ(Ed�Y�aRS�i���7u�ƙ�5\\Bb��?kve<�Ol#�X&�10հ���@!{�=A߬����}>�m!��H�y8}�<�G�a���	-���熛I�^�1M�-)h��-�3�-��g�5�5�O|I#)w;l�� ��?u<��,��~Ӛno��E��]���� n�g�#�WI��������Ku�
���\Ӂ��I��i�P$I��뤠��;@,���8-ױ��iJ�v�Y..n?�:��?6lo�4�e\�=�hͭӾk�'�&JU�����6����!/�q��p���,�NG)"�<��h��������#�����jfh��Jf�l*�[!|A��� �*�wS&��>����I�x���tg���f�k��w�[h !��:��O�^�9-�$7J6�O��v�E}�Bd��hB/ƇormR�F�&9�G�<c:�ri�3p}/f�4#�� i�*j]��YX}CC�Dٳ찲L�����Z ��ʽ��Z>o}�Z���orr�i�!i��\��ߘNмD������+-�: v/�m�H��!A� �X:�{�]{QF��BO���-�u����'�U����7�RVF�PC<�o��k� ��ş����Wk���D%V�2�{ Bd�I\s��R�F(�Ó[��� ����7�L�}�nq�y<|�i(�W�i��������g\�����b�+��>u�����苫r̓{�ȵp��&��� [^f��S����:��$2��F3�r攺�����}7�R��1�G�����y���������je���a��#�8(M[dv>��s���*���1���ǘ�vw�z�L��ti	�x4*�[XNc�u3�M�h�Q�f����	��;���%�o�g+Emi��H��|���J��H��p���M8���a�G�k�C�G!
�����������~���Ht{P#����V�|F���䯑�R�|��[&����%�Y�;	6��@+X	LI�� �_�c� ��j�q�qFKrP��_���g��Y�������/M�ca'K}�����u|��u63������ݯҋ����^o~v�"{p��w�ɞ`b�$���	��Y�lyt�L�Y�d=[z#]X0"�>�S(;n���a+Ol˪��=oAp?an���Wt�+���q=�b;�Э���TT8KI���Ǳ@���3v�qU�)4��o��n�c� ;��-�\�j�\��D�8}<��d_ܴEURP��\JW{�4���U��=�9_2�RK�@���������j�����ɦ���,=m#�����m��Q �3�w5�o����<q�R����Y�.�L����*v,�����h%R�a���6����Z�E7#X�mZ���.��p��Ն<�4�ns��N�!�0�M�`Z��0^�0���M�r� Q��n�������������ox��D��R�z�B��l�'�z�8�.��ND���z`{[�hoYd��
�1�=���/��:���M��R����(
��BM�D�$�%�d�5M�B�ވ�gYBeI�d�ٲ���;������3�y{�^�ܳ<��{_��)�y*B�f���K��������F�l���IIIFj�ed��߱��ח����Htkcr���X�^=�e��.|��� ϐ��e�ofX��Lz+��x�s�b݂gF�%��;<�ڵ��*׮��H���PMM�!��(J��Wod����0����o��&k�^9�?���Pc0��{<�\g�,��W��}�Ҫy�c��j�ո	�lƑZ]�u��n��Ƙҋ������>>uib�1���� |���h.ޯ���y�V�鄔#�I��r�u�᳻4D�t�T]k3;���������Θ1���v���ҥ|k������Y���u鴤۠4n���b���%����}�z�#՚����B���� [�/u�.&&&Fmd��}nӍ�T��d�l�k��4>Z�޲�%:�bb^$'>s�v~����������T�.��/�n���ԥkH�~�������d�	6�#_i-j�di�L�~���9�PR���࣫C-�&3�dŗ��Ō����Y��1���.���\�LS?�k��K٩<�N��h��z�7�Y�h��o��M\j|m"��%7��vJğ���y��Y�ً�n�)2�;��������"^7�:������g<�F�q�)~���p&�"��'�Z\��<g�6��1�l�����J9S�n�����W6�j�Ƣ�j4�_87X�LD+���tkLOO4ۅ0��y=�Z��s���t:`�m:��t||���=I�Ul���.�����_��s����ӓ�����o���ï��ދ���w0G@�.���{L��q���W�D(��=�s���/���=���];~6��N��/w��U,�n�j�d`⯕��.�Q���r�{zD�����9Y�-vx��z6 �%~aҚ��9��RJ�� _0��|+��c��]Z1#�w����5L�Xv=zd���B���k��,�v�P�Ն���v��5�w,;l7����*7#������q�y[���=����[��ol��X�����F!�4���*�OT�;����2��ܻـɩ*ߎ~�H}ˋ�]�@\J�<��·� Y��J��wzys�ߟ�ΎU�d�<rƦ�V|��]�j���dq��i�l���u#:�����M�ͫVX�V��Nc��_�����*/`��}Q~#X}��3Y��f�l n�����w]^4�o,;�`�_��6)8�:����@�L]uL�^���/Y0�J�~����y�o�bzƇ\/>��� ����=Lo��!.�=&�-�����+拄{��Wy���H�o^�`�ӿw�8~�g���6�:���/���Zt�*>�\����*�\���:rݰe�|����c�E2�j�.	H������ᙙ�/�}g�9�M�/�t��L��,�En�2���;�&!�c�3m��@�v�O��y�s\�t2�o�a�K�2no��-g~u>RNf^�������m��y~hP��������
5^�������%���/�S�%�r��mL28��-�_S�-}`5���l��\��sms���#w,��V�[V&B��Kt�Z'd�c��@QF�Pѡ���?d:�?R���Qxd>O,+��k�[L��x�8���,y�n,�h�i�!����~�����ꐐ�f�a9�n�yќ���,K6Ez���ױ[ ���
�\�xHm�Ȼ%�

���q���vC-�w�`�9�������(��)�k�~�L��|c�{g����?�׌��Ͳ�O�j/�tx�����=T�	����F-ZC�9ӆ�>���Ek��ۜ3���-�r��\߇aןM��\G��au�G�-�7��	d�ճ�ۏ#ڿ�i`zd��ЏG�wx��άʙ�'& 	��#�k=�dr<ȱܠL[�*=ykD�,�@҈۬�����~Y)W����.r�,�낶�t��8;���ZɆ�S��^[!7�'��?7ƒ��a�V�.�g����������ٺ�+mQ�v?�8�{�;��}�ï����*�X����W+3�W�i�l`z�L�S�%wy���������7:\F�rOrΙ�Y�cY]�A��%�IF3�2�i���<#/h���������Zﶁ<.�o�s�jD���SAY1;��s��f&�����"8 �&�*�8�rGw���Rg��m>=���]�-�-O]�9�x�i�SwG��ɱ��(h��p��Z��%�xf�~Y����_ڜ�·�bW|��?�<=)��]�Z[��M�,�"�BdɫrEO��aW�>�c�� ���Y�_�.��:J>��z�
g�9����tk|�my`|���\c����-��ba�M
W(ᱶr�cꔹ�7���S4��*� ��E�N1ky������O��>������0�^S��yӛ�Lҋ"_@�zmj��D����j���_[�V&���}}�.ݬ e�쥜����?��h$.��8��*���:A��;G�\�g���K1��*�U�w�o��f,~����Cf�92�-o��;�q��R���(��e{�E#�k��*�ҕN*]��t���9���,��x���&<=/O���f�]��,;�t�jHB��G��4�>m��O��"���HZ�,�]�Ƚ���v<�5##���Tt	�e�6;5^g��\��r���x���M,9�ԝ?1�w���B��H���RR܍��Xa��8�����������{m�m}`xFZ�G]�u��,�Vqu�20)�a��fYܛ��^��,���h��{F���6(���Q��rؙgZ���DH̓C�a�]�R�t˽��Ѿ߮�վ�O��E=�y�2��1���1*��:�#%�����6E=1(�$���~��ik��3�|�@� ZO��/�[�9����չ��rS)cm�J��M������i	�1j���"����of����
���14-�Ѽ����8v&?Sݚ�n�%<�\%X:@�r��X�%K ��m~Y���q�wtW����d�/p	K�i�c�4~JX]�>(d�ޝ�5�~W(L3���9�X�dĉ-��ϲ-��:9'u��p?X���Af�
I�'I�'ܷ}��(��`Luy� ��d��a���.���~4[���aE<|������I�vF�L6�:K�9��'�@�G����/8?�d��V�&S�Y��,	K��@#�4�0'��k���u�lw�	�[��}ť.s��GF�x!��S)t	;SL�V����)3�i���g���OoD�/hL'�F�p�xk~�A̯zg"����z��3*Jp
}z)��Ѣp4|�ڋK�w��S��1؜E�����`j0k��$scQ���@i�S� [y�s�1����5Y��|����(��H@����J����g�r���鐇`�bo�Q��5G���p^c�(����h� 7!�E�022�oL�����S�?5�S½�k|���i��`	��;._Xf�WVZ����+��GWY��6�B��ɓ�z������i�o����x�8�/ϼ9�}zbH����г��@�x�1Hr*2/���O��he�X�$�� �ffJ�'����h-�(���VE_���"��^É�1#S�*����>���6Z�:�.�,gn�o�g�u�(�Ýa<x���d'��lAJa:?���%���j���_ @�+�z���'�W���gn��N�(v��$��i�O��W��9���Uֱ��׵�LRz�L�SR�����u	T�-�5�w���I-�9SLФ&��l��`��_rI�4��+K�y:w����K�kρ`\i����P���p�f۹k��:��i3���"��[���W\��H$�3^Rv�Ȗ�"����&[���V��n5�
����P����m�	f,a݈!sƟ'�`���Igf<���$�"(���{m���7���[�(�4��_�c�Hd2rt��j���6����S;� ��D�H���G�=8!�+�!���)֜��Wn���J�cĥ�<���̕��x�^UUq�^� xD��cl�����r��>�����[�)�;Z�}�m5l��x��]�:\m����|���z���H8�OE��������O��n	�~m���	r7�E��5�>&Wc�L���JR�n��rc�W���u��6�/6��С��ڨ�3�;@���#��2Ĉ�A�J�I�ٶ�6���aT�UU#����r�>�sދ�	��vt�~UQ�v�A��?���Ul�qLi��6h��[�Hv('���%�_A%	��Vy�:!��[� qT��ы�E��8�%XE8 �E�;���Ȅ�Waҿδ��;��cvf&�_�H����K����;R���V�6y�NOѵ�Zl��{�Nl@��u"ٸ��U��샲;��o��hGx7NRU��V�P�HB�]��Q��Z/��Rp��Ԏ���{r�W��㾭���Ub�B&���H�!�����_��Fw���t��!��l�)�+�rg��R�����)ہ<</�p�ۅ���o��*�L_t<���"nU���#I���w��� �(� l�����@_�~Y�y����Zp���Lk�S��Q]>���=�8��~�צ�U��ik{@&:��x�h��'�����=Z.E!�~Հ��3�[	��x� �$��0��e{����P��ޏ��'�g�5R{΢��V����8�
�=0�E�:u��X{$Q�b�^���S�!a�t���n9�k��s8�NP��lB�p"�3� 8�̔�llB��B�h_'��IZ�+�dZ�a�NB���-��h��.nt����{�����"�:�Y%�8���0�]`�/���5������{�?��)W��g�h�b�ȕ���@�h���p�u� qm�W�Q�b���;�	&�?��J1�P�+5�YMU���5���OJ�m��Tay���������m��<M{oJ^?��$��t�%�@:ݛ.eG�|u�CT[8T-��9������<�.���T~tو�3Me��:�8��G���i��`����w�m��٠�>A_����R	W���&8��Q�eM�� ��γ�u����U@9��u�ƛ_�hf�*#�����h<�	@%�*!7��-�d=������T��?�Q�6����n��qzfB\��W��D�N��"�}ޱT$���s����bBP�UK �����.35�`�dީr��w��h2����EP�?�_ߘ�W!�,�5!B9l�ξ둹��E��9�9_z�l��@}���y�C*3��Ӆ�ڇ�/�L��#]����[�NAݺڢr�=�����7�;��`��Rs=;�H�4� k�z�E�U���x&a�G4�j{~�5�==���J��?	�����q�P��\ߦs~��v�C�&%&�'�~n�*�C��S*k��uN�[iЊ���AO4����H7`cERCُ��It����o���j�����q��\��G��FiA�
��p��({�0�l�ך��@�d9�j�
fH���]b�l˥48�;�]Q�u�ŏjG�ȷ�ŏ,;?�$|湚?�y)�A� �|P���"_�7�Wy��W�@{�[1=7=���+�B_�k�l/ ��Ϳ�*<uҪ�#}��Z����R�x)��E�yL,�Dx��g #(V��h�������T����6XHc�~�S��	@j�:,���/J����E?;Ĝ��;>}S�:ؔ��+�
F��rJ��S����k�i�����m�W�_��lGF1]����o	�.eR��">�������]���� y}H�
Ņt��wKx���{�Hl��Z^�K�I�S��i����*�L��@�5�ހcV.8�&>���E���;���ہ ���*T5�	�-z�`l���Q\N�7�n�Lz�����@����,L��Y]�:M_��2�y&�b�a�b�ؤ*7��${6��X!�^��\�H�����"\+:���m��f�n�sl�L]��F�� 1-?֋��xl7A���ȳi����J^5�� ����$��U$C?�r�w�oL" ��Vޑ�C�m�Q���t��_���`��YH�AM���H['ʥ��lX&��x���Rrc�|��@�Q�m�j_I��أY���B�= ��+�w����7����e��}}�~U���F���4���l�4�@z,̰�g����H�17�R�_��U�Y],�9k�Fi���JΎ(�^����#\뎊�B&U*@�M��O��[��̄#�*|����ͱ�1f)$�}8K�J��U~�5¡1�o��^���;��;�@����_r36��ƬAA��l�e�2,1�K	2���C�%LuY�7Z� �]J(��d%ˑ�PRV���}5>�"dJ��"<#H����WD����b�W�M�&vkm�g�+�L�2�T-;��5q&���N��D3��vg�T����aP����bc���0_oU�cD��j��D�qe�v�N�2���n��/���V3�HG�����f]�v虜�,2R�g�!�'@KE/�?Z�B ،�<�&�ylT�i�t9�=�it�cEe�(�ȭ�$ mF��졄P�[5�gF�a'�Z�q��Y�ϳ�5�o_��ӥ0}�Ɂ\�1��, Zb� �dL������*�4drCqZ��w�[?"�����.���j��'ٔ�h4�����Gp�ȳ��[t���'>�g�����魮A�L����x��=�҂�1z�ǳ��{7�� T�,D$md;/2?�]��w�ژ9D�����觗��l�gtt�x������-�>'((�$���n$�ð�"�(�]���{��0߻ʂ������[�g6e���ת��&T��Q��`�8�[e	�%,�+��񾺎�hu����Hv/qP�£�|�
�C�M%��[��.���^6������Ծ������QA�!8`���?P�ʑҲ��y�Unʙ6/-/�(w��$K��G3�٨���w�v��I̔MV$ e�0�H'%�L��s!�$���%ؓP"MsZ�^�ƨ�\�G��1�"���R��BUI�V����XO%��r!�4�lݿ	'L�����_���/���d%<ܞo=8�y�+���D���񮝩�+L������Q�ǳ7��`���v{�`S�x8K����I��@��4@�r�k*�D>��|KX�fV]p?���6(� V�T�w��M�CI&� �Yv�-�,����i�.�<XS+�Q�* j�D�8�G6[�����L�"~�pZ�`f��{RSf�+N|`Ү�W߀O�(�%)k��[ۃg�6�\gF�@/B��̞n�,!|�6�����%ȱ?���Q[k���i�T���������>����� Ly�X����"�^��R���k\{ .���� ɝ4�B��&>���}⸼�/4v�DF�����QZ�5`�r�� �#�;e,�� 
��'jD֗�O��Db���*X!{�hL��bv��X�RŹB~�B��2?񐔼-1O�'Yf�B{������0�;g0q���wl`r��D��;�l?�b���Ͷ�����,vV��9��\<��r��-��R��د�qߩP��j���O���>�/�1�,Ј�M�&� )�)�ǧ���ԏ��4���j���h,P�O;�X�wy	Pu$Yu��ʿ�Q����=;F��WWO\O��y?���v�$ڦ:226V7��F�Ȁ�l7�fLd"�r�H�ҽw���m���-�6���{ ,��jv$1\�FZ���
`��Ϳ�sIX	*�8��s�˖�N0��ig�D�ς����\MT ]�nÚ�x��v�anO�����ݿ�x�>�T�X1�@��'\_2��\tצ-���Hd���h����喽_^��Lu�����͚���0\J��~�9���7��&�:g��S���3fgj|�fNA�]/��q��{�'lv,t*V&X���߿�hI�w�_��la�U�����#��6��${�f4�&dZZ	�'`�N����1l�����"�J��!E�|�5��FFۑ��'�`ɀ��Z���4jPfo����]�g����������b�5��B��5b����[R'GM�x���R����&�0�x.���h¼U�?K��^�>�E��އHzh�#_�Ep}��p�6�}�S��I�N���߭�&�������8�L��uI�a�5M��~5��9.$W�w�-�Z�t�(���4P��·���' #mu~� ��s�]�$/.Kފ���W��qS������Y1�!�8��W�v�z׀j.y�y��W�g� �n�i��Ͳ���V�x��=3{�G�ǰEZ��0��l0�jȰ2�Նr��2R_=R��������@c���f���ysm3*;�w�災%�on��*\nPF�^��]��O�" S!#��8�h���:w�bx�
i�_��]N��	��/yksrb�%�	����q��
~{Q����Q���ݐAmX�a��?~v�`�L��wF Q�}��A£���;��g��6��A�Y%��e�p�Q����k;�$a0ʢ:01��`}���b�ױ��Ó��~��@���K�$Vs���>8X��M�X�&ڋ�LOx��ȝ�O%3c�}�-��I@�S�bWFt"(�e{o"������LKpYٟt�X��T��ǋ�~�[�ل|����+����3����U��"����>V��G�K6�)H��h�q#��8���l��ɩ���*�}:�l�dD[v~f�hm�au�{�vG7���dS�b�׷N���k�P�xı��r�tjD���>��G@���˷B�^��2�F�Ǔx����+����� 7�7V�٫f�y�@�h��/!�8�;Q�}��?/�X&�6���>߬��Q�#h{���>�wWߊ7a��ގ�rTL�@@}`����4Ǔ��I��:v�=�n^@*K��*!`̸���+xӪ����b\�M��	���x�>rc����F �#E�6:	vg��DLKV* ����+:W��vI!ԏ��kWi�o9�C0<���{��BB;o�:��O&C��9�홹|��k���զ7�3��b�V4g�	�v0�(�j��OQ�ݡt�+1t3��$D����h���� ��8��)�tVhcϥK�?ho���≶nUU�p"�F��k,	+q�n�z��:��{���mb���5�f����q�Ӡ��h���������Z�����,�h��%#���l���!_/p~_b��j}�Q9ܮ����s���)�� �u����י�rX���)�����ҟ�?J�Y��0)����<3理u�I�^ml���y��^��n���'ˎ�6�3��8=��P	_�f�XrR0��$�}"%k1��42ĕ�n�	w��dA]�Jc�_�P*��3�� x����'G�8�x
�}rrC����Vt%e�
a8�r�i7�`��+�-Y��(©49:�gK�ݐ�,Xn�8���R^&�lQ��.c�<�7l�28�6�C�O���| 4
��������;��
������4)��:DM6�n��z)�A>� �#bv:��ΚQA���eE�!ޗ�AK��$�����i��B����eSު��''>����e�Lj%�?�A���:���Ew��/���Q���]����� �<rɖ&�& x��ߚ���b�;����Xa��ܛ%
sB=�,:���ju|� ��Y7�:��-�9\��#�2Y�J�o�@��$kT�����������y���7�$~�jH���&��F4�_v%`����I��`JFת��T-�਄�9I҅����!��'�m���ī�)(y4@��pV��vk����/U.��;��7��-L�s������p���C�E�W��Ԑ|��F��QDF���"�����H"�w؛�M���Xh��Q�/�?���e�t��8�F,h�����"7c2��"Kִɡ@=;����� ���@��t�4�mw=�r��1�V���d\���c$��L���dg	p��_?Y1,s4w��7ٍ�\���g�Bo�-5c�nr��΃(��i�fɺ��WTdj;��L���*����ȳ�+�3	&d�SOȷb��4�}B�j!;�]ƨd���e�,�y�2Nd3S��.�9��_�:�ʖcg�-�W�{�#6�3!6���ur3Çѷ��y���FJ�`͗k+�i��z�x(9��qW72V�n.J�}�1�#�&������g����1�p��
�i��H��¡\~ҵ'^S9#/�Ӝܯ�8���Oӿ���ʳ0w�Tl���Ti���������w-�¼����MR*w��H���y��Po���V�&�^�kK!��j�h��-���&�^��N����k��[g�E���sPb)��,�!^���A�O%������g)������!%�󀾴�����VPk�?_���I֖˹m,))i�>��,�טq״I����;���+�-U�;�OC=�t���|�O�z,�Aޓ�3�$�_��kW���S�]f��?�Ĉ�(൏�����8�\��bdo4vC��H��f���7��gR��o���7$�O��T�S��9��!�!H�ɯ��~����v�7}��p�͙V�*3@�`���8CJW$���oN��m��r�{�*����ߓ���P��<�h�� ���N"o;΅h�{�9��477�
��O���H�N�A��oM��2�ID=���/L�������`@vٮ|g"z���ޚ�wDfw��;V^��8��< �q���@���X��ޞ�����󘗒c�~_D>0b ʕ��P�O"55��q�(=nj Ge�v1��t"�Y���TV~�y	����
��X����vv)0�H��.!�Y��[�J��ّ�o޸ͻ�m��W���226
��J
`L��H-?2�-��� �$�n�F���?6��{��ڜcֿ���ݫ"��k�Y��ח���c��">�o.a�74܆����G�*^���FI�: ���I� ���)�%*z����[�zb��yLv��q)�.��sr�ڣ����D�u]��\���� ��<J齜�U���V���hs[f}�S[[[�{f�J �"�,.Xs��tP\e��5R��^7���"bsy��%��.bN��"pd��hV�����;��d����\܀�v���d4A��\�J���߂�JC�#êƜ��j��o��CKpA��I�(�����a� �u�z�߮�R$���2�,���U��oP�%8��(�.�@n(?�_lS�B6r2d����J|@?X�g�y���!:E5I/�� c��U���^5fFĻY{e���'��?7Jۯ�r�
���+�PA$��B1G�t�Z��=/�S�m/���{����jO��%��M���9�v����7�V��N[�����f�I፲�ļ�dS�ɕ+��������G��bY�njnQa��i.�B78�����O���24���8 !VSB����Q&����?���^ݭ���������G�mNڼ9�<@q&$|A�J���mYK3.���TRo�A�{Kwi�4���˕��mETVH5pV7UE�v�ӥ�¤P���T��\�Uf��nl4E��'�,��B�e�wY��L^B�f�P��+�}�w����iR4��^^�輯��<�|�B��.X�a��`sI����D��Ŭ �$���5�q�N���0�)����ɒs�yO9lώ�S���h���Yy9Pk��~qq43�n�a9Dd��?L���.3C.���ޅ^E������/���b:�ҰD�&��������骷O{�(�w���r��9�N?�}��UܫI̲� �
$8�S���`�KēiNc#��gW�~l̲ѿ��H%����)����V�U3��?����7_��M�HT��7ֽ��h��W�:��~�|-���w+.:�N��O<5�%�<�j�'(p��`�/�����,�q2Z�8S�,$u������ �I��ԯ6 �#�#�EV7{����o(=ۀvI�u�O���q� Xs�~Ă����MDN3�Ej�Z7]	b����`�����$H:�.�m�?!qC�LU�[��H��MQ˿#�nZ����'ݎ��+���e������u��7�W
�"��W-,�L򐘄]SK��ۇ;��:Y`锛F노�k���v��n���	b���ݗ����S�6x�V����O$���ĸ���W/���7,_��yq����TF��TK���M5�����R!{�x������i�O&�𦬉��㛳��E����������?-���D�����q�m˺p	`�.I�ɑ����4���O�$��o~�y	��9r���N��`5^��Ϳ�#ֿBk������G<d�dj����$�;*�M������	o��^��sϼ��-č�m�ߌxn �� }�4��l����&E�ͥ塷k���E~)ѮTE��/��F�'�m���PT���l�m=��WC?T�Q�ڞ�C�h�m)p;|�`\t�T�����aH�# l�"�%cA�w��N��K��r�|[@����Y�C:��f�L����$y��6�^.o2��JUZx�S{�����C%TU'��&�+G!��VS&MPoZ��� 
�4�{���W�w���j�i%)�m�#�����ߜ��ͣ����>��i�K{B~ۆ G�� ���`'��*�&��'��z��ojྸ��K$=�d����V�5YY@��5 |�=4L6pPI��Iqߍ2^0̮�˨��F�],�k���	U2����WJ���`�ɂA9Ř��jr�P�y]'7��wHu��^R"5��8�ZJAW.�2#��ܣ��>]����RO�-r�|���פ^L��cCN,qj�A��7200 �ٵG岓i��Q�e���l�55�G��t8��&�T,D�?!�FF��6�;�&�#�� ���*�B� B= P0 �()R���H:ե�Y��oA�bV���Ѐ��/��h*�5y-"�qy���f�������*��w�+�=�a�v33�|�7�8�bU?��n� o	�~p�V�y�\d���/8����V��g��8�R2�
��W��*5�u"�e%yCs�!�-���F'\��{�W��=�Ž��o^�jr�.��`�uC<O�wc��:(���$��W���U��9�J�#��i�Zd\g$6�8f����R "�n}�p�.Pq�BR3�B"�Xl!d%�U�[�~O��_��Dk�Ϟ�*��s�X5�Z���8Gf����UBos)�Y}``���h�w�С'�b�E.a�L�d*ں�����_7��}��K����m�l/o�$�
��!���_��˯��R��>e�{��Y�nK9���P�n���n0��0�5!��7��撥�GX�h��t痜���ז@�rO� ��ᷚ"*'��[:2�!�u�y�))�!�(�=��Bj���s�.���k+q�k���� W��D�B9ڏ��O{�G��'����ɇ�6�?�����_d� �&���wE���,)�s9(X�PbU���dvR��˹�R7���w����0@7p[�ՕS1��:IW�e���L���_�P��迅��%O � �Y��P7I`0��7��C��'�.L��� ��Y�����ߠAю�u~�e�m��M$�]���V+�{L��1�o��M�/���������I��J ��з��wp��G�ӟN��i+�c)��C1�����?
��.���n)Sb36ұ EYL�^�7��u���?}:Ff���������ƌ�wEՙ�'�Bĵ�dv�Q����0���CAU���V:뭔-�L1}��su����7�����#��d�RX��a���^���u�A�~���n�Ŀ�`�6T�C`����#����`�r"23�M
?4!�=�O�p�dē"�e+�z��'kNZҕ������m�Ů�O�\� �i#�%��J��M�_����ad/�/������,*>�$���
�-n]@�klj����o���?�n���<���c�k^����}��������{�D�/��>���0�0�<��Ҵ��<�Y`z�+*�=9���nAA��p�7-+)<�>����ĸ"�L�K_5��Q.�@��vu���+5�g���o�e��i�#e���L ����V��|� �F��Q?.��4G/IH����J�%`&ޕ�����'�%��3)���t1/��4������ȇݿJ���T?��+܅�#��Z-A��3��q		H��G�,���!�\���ᦅGA��t|w��Ne6�E�#�S�z��lFvxz�rH!R,b�n�J�H�hf7]�i��d�zۡ�1")�֟��F��`R��X-��Q�W�^i�96��<�Y:1{B�p�`�_��@ 봵�?� 2����sӹ�R��F���y�/"Т'����s��HGQRNN0z�eZL��'�����P�����wzI%�Ԭ_C����)��g�|A�ս,�p�	�|>إ����>5��6�ih�i�ȍ�Nb���n��.痳�hnn�m٤�IMJMe�|����&�O������(ĸ���V�K��<}0�h_�sG�z��Y���;�|\\d�u��;@&,W<ȢY��m��#�����9O ����C�����(=��j!*7o*荎gڔ�e�1=D�����^��[�O��-]�M�s�&TKa�[�w�$����7cy��2�A�ڙ֯4����u���~'�`�����7D@=��Ө�t0� ����P���Sdg?�d�02�H:��

�r�����rvW� �ǜ��APxT ��N0�a�y���HQM�Yvdڷ�����.W��ICCܖ�fm*�RK5��4�H��漉0b\��P.�l�/�g�� _ so�~͵��2���h!(��X|��$f٧������һ�ZSSC �"�j��>k���E��Dz�5t�K�8���z�!9i��+W};��Y���L^�3.�K��X�*��z����dɞ�lK����2�s�W���ՠ� �ǅ�Ї��%��Y��B����aoQsy�P��c������E`����|X��S�fޅ�]SM:�n�QϾ�� Ϯ*a<��H-����������@����,�i��v1{��Z��&���������OB�%V
�:�������8�i�Y��e��`J_��|��[v���|�P;��ʧ�Y��O�.��jS��UVH��]�1<p$�g�QdA�7$n|xq����}T�o5�����"	�?57���'��k��Z�B��Zʵ��"UI��|)~�Cސ�2ˢ;�=��ב����*��r8�3�s�,Al��2��$xv��-�YK�6/)!| n;y;���`SF���!y�3蹞�����FQ�o�P�Z$%'?D��c���p�#�|�[�,�i8��,�Z��C��]x0{��؛���'����8��3�2�!*+�V�H�
�wu�.��!T��A���Ch:_�|������7�C�v�X4����)o�p�ᶃ���k�"#)M�HH�2���"�V	�1��!����q��:(x��z�|k�͟�S}	���&��"�z�1p���������B�
�q%�/&������}���t?�	�v9]�Q�|7���F6���@A5Nn�O�D�_^|���}�z����+��GG;|� r/ bYA}�t���d�������>�k���B��L�������/�k-_w{I�b���l=�nC
�i��h8�VVE_䗺��qj��U��'|�ȑD���ux��XB���) �]�%��Q'�h߃"�ׅ��F��H<y!�vI��j����M����A.y�g�ΛU�s�A�[j�"O��Q��b�Ή�2���i��°�u��KTBߗ����B�?����Oɸo�Ƚ�����*�]15&�I�za���p��@\U������#�WY)U9VC*�M�!=���W0UF�Dxu}]
���C�\ޭ7ZJ��[��xIÆ@l"A�*k�B�c��M|FRe=be�&��Jo��'��J^J1���9S>�* u��X�+$}����9���J&7;�}<�����Ѳ��//��#���V��m�=ڍ ���\�eQz�c [x��~kaCe)E���j�ܢR�jx1��9�Gn�o���n�!�p��?�B�W,���D�j��o4��8�]=�?_��p��,�̄�D�dxbL�}��� r�%r7rBFi���2�YP�4\��%++x�3�b�o�k�vus�H�#���B�x�1���	YY��eDR*܉���w���:�_hΰ�GL�K:72!������o��7�4E��]�/N~�8�� ��.�_�?��z�1E�)Ù�_��{dg����ri��[%LŽ$��P�a�afH@�����X�s��"7<-y"T�����J��a6⸡��۬u,�C�A������#���O�<!))k���a�4�-0�L��T^�F$���"I��t��n��C�C��1 ��>{���|+^�Hm���,�@��Һ�V��z��߆v8<��Saɢ ��̃3*g��Y��@"l�Fi����𸝧,nuSs��G�e�I���`�,�Q���A����!����[(A�ȕX��H��Wx�Ȋ'!Qkq����;Hf]�	2 D��n~n2K����+.Pg�XЉ����T !d;
\��7��[:耾���
�G���R�9b�Z��smz����|6/����Ka���R���Y �� XX8�J��� ��ꅈy�u���}���	%�6�
�x`�Ӱ���E-Û�Z�{����;(I|��yU�N��5���i.��h�r�|9p+�'v���ֵ]L%Ԟ��3�įh41c�h TIii�PO����h�$����7ϳI��WAꕺ0�&C���>R��F��R,�9U�:i�^߿�M���g?E絿���w��#��E4yoģD!\7]�T7�-�<�(�1�=0���ȍ-(.���'�4֣ffa����������>0G�'K<`�(G-P�(���E}"Y�������V\*������.e�r��T�y�H�Ql�Ic	��V��i�(WF޻���=��Z�����[�y��H���D<iY�$kѾl�c�j�ȯ@E��?����^s��W��_�R�>�Y�eW(�J���%���d�QO;���������Oi�s�Ο��ӱ���L}dS�a��WHGd)F���+��䑂R��ʫ�FD�� �*��K;��@�8��la���hl��KUB���O%P��V��͸)x!ǻ/��4�r�"�pƦ��V��g� ��sɹ��ȕiA�W���;����R���w�.��ޢ%��Vi�.� �b3<S��')�����=^w|?�Cb�(�x��qL���4��4YZ�A-vv� ���)d}K0"
��t��i+�ۃ'�gsgQ���=��4]��+m*De�AU�T�7��e�.��р\��ٹu�h���G�F27���]��g��O|k�v��a~�[`�۳7A'�����k̀���-o1��21hǔ��x2/�t:C	�iR�G� 4����hL��p�M%���Ӏ��� �2.fq��ݶf��E�Dq]V�Q���q���dhE��Wl�hW��u9T�"#f�/�$ͨC�I�˴�(�n\�ع�Np:�2��fͱ��k��b��6��D����gb�h4���L�{om����2���|~}�q�yn%��rJ���

�_q�U<�s�rh��ܙ�������]�����w�"2�2O�"�o$��(J���"w�8rQ�����^��<=� ��o��r�P�҉FF���\1T"�-/���Y\r$[�v�U��+�-��oi���͗��+�,n�}Ob����h��k�Rpe�8-=݀Z�q�"ДJpX��zKҖ�Lk�

	aK�
�]�����M��E���?�+!|��Q�������z:�>\C	a��|����F�1\�[� �ߌ��\q�F�f���`�����M�	B���ke�n���j�����QJ�ѩ������Q'��zd���C`��c_+M��k�O�]����9��l�'�h�����|�s�q�k,�RO}I5gW1�QP���ƥ��Ƥ�T,(�0K�"!ʗY���uu"{���dn�d.�/|@t,\��.���
��w�gv���"�:"am˯��Q�u얯��Ă��7-y�Ѯ��4�|:��k׊�^9T��M[��9�9�h��]���<����k�VE�.��V_k�w=���s��"m��C�i�i_�o��2S�IS����י���Ɵԡ�_��V�H��5��ٰ%��n�ꥯ�Z3Y��ьށ����\��(Ϸ����f*��[���n�3'hY�����QVsD�);�M��f�<����t�2i}�4�Gr��#+f*�gT�Qc&��*?

��Xrl�%Mg����ʽ�c�,�t.4����5���� k���M�]����ў-��+;�k���g����:�}���4$7�[)��P���:��{�T�`2T{a��O�1T�x�4N��fY̩��֦��ϼ��^%�E���������<k�cF0_��A2�C89�ɉ�y���-l�ظN��1.�olnv���k��U�&�Fh�Z��`R!g���Y���`��l뼷�Γ�Ƭ6<:u��b���sJ;��=6�p%�_L۴��=�Wzyv���0:���H#bܑ���&Vֹ��4d�>E�?c�/(��DB�x/��ʽ%7|1M��&O-�U8�ƲV�A��'���&��7���ivx�Ѕ�{ 3��[�Oen���1I��'K����HK+��QUn]�]�,$���?��7E�y`���7�,����J��~�t����������͍��ŗ2��1���y����u�FC1�:�{����'��c���~5�?l*�9��!�DpL�W/)�|�N����`��Gw-Q�f�T�o$�w��ѐ
�ӧ+-���Hs�!����0���E���󎮏#�feeᇉ�`����NN�-g�]�VW?����u	�������j��0s�Cn���V�	zY�,�ޒ������3t�#�_������,݄f}������~�s������c��/:Z���y�r(��������:{����T��|��k�!&f�Ċ������m��V�~�-���.��)�U�=>u�DՋ;w� �T�F�� ��
�sL��$�흛����������oު�;�󥵛��ieF)D�8ў�'B�`��T�8/����XzP	��8����6��h�2�58u��2�
=������ݼ�u��^N���i=��w���� !�#TN�k��:ȆD��,�����MT�"T�k݄p�Uf;�X��Py�YȐE�)���(���<M��R����'-�`2 0���`��J^2Z�N֒����鹭`��W���o���X-��
!%�!**b}j�f�J36O�ut���Y��T���7p���Z��\�7���;uu�<�ǘ�>�}�"��d4$�y����[H�Q���P��ezkh��h�1��u�\��M�e��2+�Q'`�rL%7��[l��'Y�=���wp� �n̞h^����G�u�Eut��F1*c�H1�(E�� �(J�"�� RX�^ņR54�Ra�.E�^E`i"�KY`)��ܻ��|���{����w�̝)�cd��W3=�f \����JR@��F��Vr{ �ˏޞȃ�F|�_m���qZ�V�SQ�:�`L6�37ڂ���w�%u��뭇���Y��.'�bHv�-at����U��nw�W|���nrQ6)!b����ݽ�y�J"�5��&;8}����Q��P��4��Z��1Gu��9< �9� �W�c���!�D�b,A�} �b����4���].-e��-LO��0�vZ#� �o#))��2�z>�]�\K
���r� /��Wc��m7�+q�"�wpvfL�y�U؏"x�zl3ei�ee���;F[�U�U�����|��i���R{�������NAy�#OMo�����5�R,N�xX��$�^�֫>kщ���Q�Ϋ4����@T>� �Vr	�{2匈j|I R��4�r@�EH�5p;�_��
($17�nw���9�-�Dj{�~c�_��ɖM0P�ج�f��)���nt�R��y:��]s@(dW�>ή��w�}i���.*��'�F\T�j/�z�Nl�,���ܐ�+� ��	I�{�\2
��&g���0u}lsn��T�e���js���>׶?�M��[�D��8p�;�����z͸o������&��� �* [�u��7�5���9-퍁�%�SQ�DH��'��)==�x&N���:18�ޓ���ڶ�ኇ�G(����ӊ�w���������U�M~<6�ڍcQo:' �n���a�0F�6�\�;^N)7i���a�M��!�:�5����/	L:4���~���X�<�_{�-h�;�h�z�`�l��ԥ�ը�����%,�W�?��Q�cSdH�}z ��=@A�[��ňX[����S�p&"Q7+�
p�����I��Q�Z�D���xZi_�z~��%��� w<(^^�i��Fx��J  8"�f $��,��'S�ǪD���j��d`���֯�	��b�Q���0�P��?� �J�H&�E�쎂��j�_&�Ey�F���"m�ѡ=/���2�y��\.�I�#60��̏c�G2���.yt����E,�� ��(d�j
8��#�p�D16���G����`����ޱ��GL�v�W���DTk�9����?Ⱥ����1P�S/����Ťo��2�5�Y?t��x��~�mX:/�U�=x�69Jb�\�$N%�
Ċ�(B�c�4S���C���G�����l���v*Tq��T	x�*V��{�J�	�0���L�f �=T��,__|� ����,���q#v��ΐ˟^¾�on�; =
��<^Ŷ��Ch�@M:<+��*䊠��[Qa�����%�*�'�;`܌�B�ؐ��6���]t��ki�;H�9�9���z,��a�@����^���z��~z�	_P^�t^d�F t!߸����3~t ��rS���['g�V>��hv*D��BPO})t�J�m��s�P%r�(�x� -�� ��N(ŏ��q��}2+�v��%B�BK�����@X��|��?��_�K��p�%(��=�
�D/3U�h(؀�Pmv�3 :��F.@��G�s�-t�ŵ��ʵ�/0�����y� .xTe'�},e"aw�	�������������6������.��vV���!�4�L[�L�a�!��&O�nG/6�<0:���g���f�}�<��z9yoZ�2nk��F�+a|w8~G6�c6)�G�u�<�"˲�0�QQP3W\�k\N��+l��9�r�؛JK�GOgI6�F$�!�E�(���w�ϖ�2��>�� ¾�R�7��!Z���xb���*��J���HN�C�m��=4�����E>���NA>�y�MXo������ �BP7^�>~����'pѝ�6�����]]	�:k�kH�P�J�zO`�=��q�zry�����6��!��S��Z��GN�����m���D�ku�L{S�$��S�v�`8g;�1��A�7�zR�Q퓟;�����O���Kn8!�d3��E��^���s*o��������`Q�`@��G���C������#W|
85��OZ��P|4�
�c���rP��S[ےl��h=M����z.�q[� RֺT��m�o;o��F�ah0_���A��oT�:w�X[F��3o��AD��7Xz%�7
��6$�=5�R�^d ׎E���9���+q~tC��$Du�E0��
��Զ�����Ц8ަ��oTP��|�M@�D�^��CN�����5��M�w]� 2�`�g��x��ax����(�)�$�����_� �م������{�aVݾ���&�9x�"P�	��S:��VOp8�̃����WIT��C�˲yqd�Q����\^7e�H�E��[ͬ@���ӥ���wN�3�;A�c6���mb*�۔TO�@ �������}^�fSU�LDe�cy����={G,�� ��c����I� �[r�1�n��9Iϰx����*�8�]��.�q]�	�|xR�c\��A�3��׬���2���V�N>�F?#���c�06��!��j�����c�ZA��{�G��!ѐ/Ҡc$���U��m,4
�����=�¿�h��34!�"��'��P�P���e���#������������q�$�W�2�.^�:��	ňXR������f���^�[*#�����	S�� &)2���/ρxF1��F�� ~�M7�Gg��n��x�mj���&"�sbGs�}����*���߶M�%,z7��5�)�W1�X�>]d�3�.���Q=%?�J�; ��p�"�[�\|Z�p��#�F�l'�+����xӥD�r�@��S!��A���]��czR��DJoQ���َGٸ=[����|ja�-�C��D��� ���W"�3�2:�5��c��3$ :=á�j�� �3��Մ�g��@���b(�LԶ�<=����ٸ�%�Bȓ��[�tZ��&�*���DoonN�}��b��!)���c�� �6���0|�����V,�O[G���X�}�Y�S�b��	���{7�6�Ю�8�cF����»�l,ԍ���t?`v�����G�'�A���Ui���e,��`*\E��<�@��/�;>j�PN,�4~H�SV����dC>}�]B �M��R�Wru�	x\�Z�Z�F�@��c%�E�UP~��F�a��:�����Uos� �P-? C��S~�C��l\�(�h�y�ײC |Oڱ���mA�n���x�>&����%�y@�Y��}	��A=݌����a��9n�����'�'�6�i�&2�����V����47�l���a5�̈́��D�;��#�����y�I]6Ρ��$�����F����x!��w���S���0�4������)�/�qd�N�FJ_� ހ���s�m���XL{� cZ�qy�+�/�"�VJ��}s����MT/���	��v�4
1�q5��t�8��vOJ��~��Y$*&5��A8��I����P�������)}��j|�[��ST�ȿ� ��D�@[hQ�� �c
(~Xh��&? �M�?�$C�!����&ئ-�혗(���V�r�j]��\๼��Z����Y�,�B�6�!T�Wb�~�8Gao�n2Aױ�ǧ$��ۭ����Ș�/���n�-cv8�s�h��J�����������Rj�l��C��/*���>�;ji�j�>����I��M (*n�+/��GV�����^���.��5v������^f_��A`x�G�%[��v��=�Ї�1|[bX10�.�ur�Z
rJ` �ʫX��K��������i�8�rA�: C'��D���*RT2�#��kk;�\��ޜ\-������U1�'8m�����ѨY3���}rH&�N@&Ƹd����`NW*>P�'��$
e�urU��mRz�t��:u��C*F��a<���s��m�:��#z	�^b :#���dol��h	����:8����~�J����a0��V9]�+��2y�4#�Ţ,��Y�$��[A���	�Z�����4a���kA�������B���33ڮ��/��"�h+Ȭ4��w��W��x�mwP�v�|�'��a��f����BxU��p+��NN	�d����Fp{X��)�����q4�bbx��~(�����P~,74�Ȓ�"�q-�r(�z�r�OS9��h]J����g�iOY}�O��Xբ��U'��ɳ����2�0����F�<%��1�����Y۬y	�#&s-�ຓ0Ћ��}6��t��9�1�������C�W�6n�"y냱Z�qۤg#H�  Ɯ����Yn���`�2+��� S��3�bj.��d�B���f�z��7al��>=���b��(��Pu��"M�o�	�μa��RTq��*o�vOG��妍���"��NM,�?��ۯ�EׯJ�6@����
`3a�`{#���ް�l�| ��ڳޛ�u!*�ʣ'�h�p��1ٲ��A8��]X9v�4.놧�j@�Y�΅�Fο���Wu����]	�6���X���VS�T(��ܧ�����Y�N���m�C�~L�߂�%�%Zo��H����H��L�dX�ķ8K���}7�n�C���\�k^�]�y�mр�>|�X��(&+�H�� �P~���|k6�׋����
�>�ᬄ�م.����>[�:]0�4n.d��k���F=���%�����	�X0�!N��8|-*��nY"�Lfe�/T��٦�!թ	�'�&g~!���}�J��8ݎg!�o� =���`J6涖�.�1�C��eC/�(gi�|�Ri����z�ꉻ��o����d�+|���o�	"6�L��(�̻����J[���^\��"��wo"�
O�R���˧x���``�i�bY�Џ��r�^x{��
H��[ȃH����	xC�k�e��v-�r@2��t�|�M�~�����i���q��on��t�oY�,��~�睅�8���H���L ��?Ru�@Ner����6��2V��#�&t�� ��j�B�O�С��"�)2�˧�5�e�B�ʳ(l��ͯdc���,�����;v���o�,��k/��6y��B��0}���~`9%��In?h"fU�@f&:�2���L�4�z�������h��&�%<�����\����*�!`T�Ȩ��	YD��#xL�B��yc��gv焴"��+h��zr�V���`����
�[u.���l��+�
?w�̷�̫Vb�
Jq
��MK����ծI������F�O�iH (�MH`���r3L�:wS:S~f �jC7^����A� {��q��PJ�f�����|ł���;�a��w�c��a�� ��J��R��[	��W�(�F���6��.{.��F����n>Xh�M˥�)�C�1�f�� rVrr �[B�AM[\XN���R� 1	��i�oy}7���Y��Nt;Gx�I�õ��m�����g�>�lh���� 6TI���ۍ�Ehu�7D0�����;��"v*����B"��)�5������	&��+,���{9q/I3�����އ�/��V`��6a��@r5_O˭��I}�{�n�^�@�_�<�Zxj�R��N�������(���}�]�<6Qu}�~�����c�D=�Ѐ�8{]�l،�/"���X��z�P2����h	Ovv0	�q;L�ݥ;W�F)9s������]?�{���&��^+�2.'+����¢ʁ��-oz�})Q�WJ����׬��/�F��2e�4&V�FO�f��'M7%\0�d��ؔ�ed�6�誂�cOS�a<���]9�XJ�T�x^*/ ��d/�
����t�b��ls���6�g6i�;��"�y'��Յ�=^�$�fp����v����ۧ�`�L)��hbd@���ꮔ�E�5�e�j/q.�V��Pd@���a��8�mr%UTWl��$�D��������F�]X�x
�R&$��z�X�����$Dૼ@ �~6x(߹���c�(���f5ɻQVm��!�(T���"zc]o,��������&R��b�zϲ�U��D��Y��Z��К~�ng�FS�S�����+���(���&��F��8�%:��q�K�.ho�V�������\	�O:�����6�x��Z"�+((�KӀ�J��h��Ou��>�<r�"j��=khcʣK��S.(�FG��������+��n�۰�8��zԵ	�]�y�����Znn��j��-�[.�jw�F�eN}(������WυwD;,��g͉�+s��5�H[�#���WB����!1�{��/#:�L�9��c���i���fz���n%s��o$�������m��=��.%腣n�S���-�ߕ���>���@/l��]�j�<l����;x?%V���$m�z��]m�)խ6yPtD�S{���{��&�9�1M����t�G`�,Y�1%��؋/S�Y(jJx��[|.I��_c*��w#C�� ��b\jʶm�[��`I�N�������N3�����h��Ѱ>�);9}�2xכ�[�n��L���T��������m�pJ�Q��4>t�����iW�u���Zp����e�O�>o	��;����>�*�I�'c��tf�{�>��H�����n�|��w��������/^����^Y�.�	[+q���41uV���(c6ЯVJ>�u�\��8\6m�Y}#���۲�F��%�֭�����"��5�[5� 81.~0��t*]}��낞K�J�dk���$*�8�;<{8H��KDҗ&�i�N�n�q��Q;n����q���gQ�aF>����i��$�<��ކ��l�./��N�;]��~e�:��Ʊy�����𳌇	^�y�_��4�I5V���u����8�=�T�mQ�U=gN=CY�\F��&H+&Z�%[��YSq�zd���/t�����ꗹ�0�O�����k�~�.�;oE�٣,`�p�C����}ʞ�!��4/Mt�4!�[j�&j����CC�?G�
~���Qd�e�z�))�<",.���C�1�-@=���#�����Y��*�"�H�c ��ܶm(ى��0@��"�T؅6�0¬����:$�y��q��>��,ا-q��ˮH��f����z8qdC;]ch����!i�Q��@�qg�YCBB���f�̧�A��#�s��u{��@8m��z�#�&(p7�|�t�]����� K���=��H+hÌ�!M��2,�x����g����I���2ܶw�OP??���>��U'�c��f��Ð ~b^��Ky6
?�P�y���)�{�,�UkƤ� e� ��5��.�|��+zj�MY�hw��|������,�z��Q�!����s4������W��.(�]���KS�˟�7�v_�f��o2�f�T����%ϻ�Axo-�$��.Ι�n�-s�"�/M�e;L��ͦ���+A��L�ժBDAT{U���`
RK�:�����P{^E���7ڥ��(}Y>`դ��^�'W����Z�e�`��r�������ǵ��A��6�&��`������H��!J檞S�z�&vL��^9�&w��J��؛���)�FOO�,����ƥ%+�eJ�����g��Oc�q��;|C���|�2N��o,e-��3<�܆�����#���:�����r��J����B����T0���O�u|�
a�\�|vM]����x��˶�]1�'V�%(��Y*A��ʕ���n�%b���v�^}�9�ZY�Z�����?�#;�W2�G�@#5`�`�4'�/[a�O�Թs�w�Ǐq��W�h��#���$7��7�j��	�} 5���VO6��N9�`�m���N���32����vl���˗|Td.;w�����^��<읱�r��:���OXT-V���--߾]u�}�8�}?E���
�y痧��~��-�?,�D��C�`�=x35R-� ɇ�ŚJ�Bl1/%녇��x��ִ�����U�/����o�y���"'��^8���?�����f4��<7�~8v�3L8��r��.S�~[QJi�{��K�ю~θ���s��0��~�0h��B*J�*2�p������.Qڇ�o�a��z�:!**2�o�����Ń�ū�2/���.�߂?�=�2U�2qc����n����DU��-��ƤܥpR��*�n^1A����Oo�j9���W�^{m�n`iްM������s
K����G7��*�4ͽ9���K" Tg�|	ʑ�6YY�˱�[�;���h���Q�9�k<@����d�u��҄5n%���ƻ(��mch���h�p`�9�����Q9�LA[q�e(���O�epO2A��0!n�f��8~p����[��P� � �A��)(�>��o������=N2��"�/���Ԥ�ƅu��M�́O%Gy�ρ�5__��<Vd�溷��>\ER׷)�J3ٝ�Ln�m� /+�/N��#��A�qV�R�%$߇]$GJ�7Cl���<���h��<��B��
��{��u½|�g�j������u�w��X�1��_�F!x}��[�z�����K̞�: �y�" �A��ƚ��@v�JV�w��+',� Y �yfD�!@@����-/���l�
v�F��<���VnJ�r�({��B���C3���Q��o#A���J���������X��엡ܦ̓�䚹9�Pu��i��˗A�tt�ݗ��C��1�:J=[���ш��Q"���:���N��E�$��6�j�xe�����2��Q��>J��	��/���7͇�q����@i����O"+����oHQA�#�����7��/��U.1(YJp(V�l��]��G��!b���3Z��W�a�:��	�C��.
����_��������guu5$�P�֥����qL0f7��8ߵZ)(���O�̳���P+���vx��ƕm�x�L%M����fR��&��D�xȡ\y>���KzO). �Y�z���N�z��ϟ@Q+3�A�B��\t4�V��n�r��'f#���]~B�~DP�A�8����!�K;E. �h�u��&�Ck�����[%7�j�ع?c�Ƙ���zf�3�x>A�g�V-Ŕ s �o���\/�)�p����?��Ck�z���=��̒���ȓ=��OIC���f\�7?ko׋-�U̏e�|o��U�tm欤, dv��;�D��c:hL����	L�;�B֓�C��1�L���%m~�ing'ũv�!�˿���@v|�e���Ok�u!��9z��xez��h�JxD0�Mz�.�u�wƱ�ޡ¼۴V�,���p{N3�􃠒ݻ\{{8{�r�Նz��eo��8�;��e�Z����[�2o_���Lq�\m���"��U-4�I�ݞ`j�S�8����m�����is�֜��g=n����S���7y����m�G�2��&���ՙ"�K��)���?�n@�W���ya�7��B+ֻ�KWG'{��� .���DA_���[����O4�< $���2O��#���-Ŵ���J�k#zR\S�r������O�78�Q�)��	� i6�(�2�`J<���Vn\���=2�8��7Q�#cc�a��"1����{Z��,�Î%�H-��T�j�#������|VN�s�����=�w��ۅ��֌�LԽB_8��NvL��<��+��;�!�;'��]Lj��}�,� ���a��R�R0Hy�}��maX+7�r�[h+�,rw���Q��{��nY�.0ԁ��|LNQ+�N�c�׬�.��i{{;�EPq�A���W��CqO��������{t�8��˱��kv!��P�hZ{�g0�kB�*�&oNu�y��� _�.�Ր7���SX�����Լd���_��r�HuR+돷d��	>�2�ڡ����57Q��$�<F�@&7o!4C&SM�Ug�����f�.�Ⳍ�P�ڊF����7��CFq���9���e���9qD}Kx{i���[�{�\�C��"����~W$�Kʷ򅷓!���\���*6['#��}���;lZ�ӨSJP��N����X�y^�&+�QɈ�f��@�^\�"*�7�q<����wl�B^����Ug\�: {�ŀ�{(8�L-bv�:�"*'�����LE=����2'Yށ<U*�:8سs&�	���/��S�0u��鑎�N�4��;��+˯�q<8���R�T�mڀ����R��e�J�C�>5�D/��;���:e����hy��0{�:գ��Pٻ���]� ���p��5wsC���]cR`'��`_�l�����;����;�ĝ������L:Ȇ��G{e��j�_���9�d�^TP4�<��r�I��aC.:���u�6�l�g�W�K*t�RT���v#M��1c�h)�<�p�d��k����0��R����'�,&�!Vc��F��a�\��&�Sa4Lk�]6⎅]��|�47I��:��i��UPל�y�w����];d���4��L�8���Cc����D�Au�ڧv��/R�&�X�J붞�l�L�t�P����%XB�l���(������+)�uJ��D5�bf���SB��K7�ߺ�n�7������ݿ;�Y裭�JroW�Ā�Aŉ�&������KWg�ȆU7��'�*n!��:<ِ��yG�㬴��N����7���S8r"g��*��M-LtB����WPJb���OZ[�����Fљ �ߵ ���|���w�R�}<�~t�
�8C���4�=q�h�pP-5u6 ���[��ؼ�E�[�PPV'�bH0�Q��R�=mȱ���3P��D1-p��� �ݟ�r�WW�����%K�v+�X�z�:10�6<� ����$J�*��8�ʆc&�ݔ�#��1hX
���"�Tr0�y�a�6��f��r&a��� f|��`c��VE�X!�۴n9�95eo��_����$� HCb�?�sB��Q�.N<��;%�dw���d9���o�1�nNY-�i�w轢�o�A�OE��=����F��k]�r��<����� ��N��q�.=�u��l��YB�ؗuho;�~eks�*�F�J��2q4 U�5'G�&���N���b%�3{Z�~�r������4~DE�-yX��������- {dd��hz{�D!0�w�l��L�q���~'_�_YA�Ǿy����'�U��Ӛ�/:&6�vȏX礆�'�.�'KWMPL�g� ��'�J�F���e}����㊡�څ~������3 ���x�n��Zr��Lo��OY�@��Xz̷6��4�$�] �&��
@��+��&��Ç��e�l����7��gfϞp+��Rl�dl.��R�I�wZ|��������31(�ʋ�;���5�"_�D.i��w���#
� ����f�����]�I��_P��:��xnC�o��?�Ր��rAy�"�W���ݧw���W��|��!" ��%"֕*�m��L���W�7b� �)��ĺ����.���- a�蜑j��n�zDn&_,E�3_��l�v�tu�Z�,*|��s���@�5k�C5�]/A��(�U:~QT5��9�)����㰌|Z�60Z�%JȠqWN|��T@�? Z�;�8{��K�577����UjQK��U���/J����t@I�UN��V�%qz���)�� ��(8Y���F��..y���<� �ğWe�׃<.�(�M�%' Dv+$�p&j�����r�5�MZ|"�(:dȝ~�e�/rl#��H	�����0�+�f���&���.��CՊ�5�Vko�Cc�+3�Hy)�{��P}]��h�R�b�j��.���/\#��I�>��j�bd������#��@^',K������㦓qg�l���_�Fڃ�O�F� �����luT��O4X(�es���b�Rz�K꺛;lӨ�E�"���|ʸ��(�#V|����[=v���Z�-��۴Jx����E~K���e8�\�{;�g]��c���Xeݠ:i��_�	7Y���D��:�H"�d5${v����[=��xų�m�kЛ��s�m�1_dL�*����f9 ���\�(ˍ<J~f��띜W�ٿ�*�oF���oP����4ǧbګ�����鍊WL�ԸB%��p3�_x8�����q����x�fF��{�8���ݘL�=�Zy6�VRd\��!2�i߫�\7V�ekM�|ƣ!�2�b�^��T��[�tUu�� �TF3��<��{۽�r�]W�?)=Ǿ�wdⳡC��W�k�p��ʃY��e:$�6���[]1��?P�������i��.��X:�} �
�^}tN�O�7��O>fg�'���؂52���4+�b�!S�x��z�/� m�=Կ�d�)�;�' ������$��^�q=�^?�!A֞ȒL�l�ך�ܷv�%ߜ�;�x�/UM��e���̃x(��(w�)�' �6��� M��&��Qm��Ǘ�[��U��Y��Lʞ����'**���v��k`n Z$����T�ou�G������>��g���#ܭ:)r�V)�vS�G���Hާ��)���+�,S3ԫ9�m���^�쾱� �<��wCnl�͏�K:�����BO��y�#r���@ x�G4cҿ��KoU�M�(���@�x����`rt}�ۭٹ��L���c�0��N��R��k�P2�\@$>�hv�4w]�B$�������!��ׄ���&��m &�6Qsj�0N8���<�89M�'L�i�g��1/<x8L��B�/�� �QP�:T��@֫!�q����W�Ѧ��n���5nP��շ�T�e�K���� P��-��3|d�/n�1C�<b���p5B�ox�?��.#�:�7'�O[P�{�K�!�F�s����d�0X�4�4n�F�����S�Es��d�Yy� m A�����m #��x2죈:��YkE�l��Y򶟣r�c4�N�j�ơ�0܍(U�b�@�:be=�8 km7~��a����z?ȧp���	L�qBF����k�(� G�fK-��Afhj_�'Yq�LoP �=c� 2����&KS��2�*�{��������M�	0��T��0��Ғ�� �\�46�פ�a�8���|R�a��mb��2Rjr6S
��o�)�_��Ю�TtH�������-�mp=�ybH�\ ��7�+UAa�`@���n���	�i�w�F�Ͱ�O8�����[��h葻���E�^_$�����ט��^: �rJ�Y�SG����rN|��R�C����w� �j3[4i�IU��ܞB�GDh��E["��V�|�_Je�A�Xt�%�͚u���9
�|_��`�Q��&j���-�NfI����'����^��$��@��w=�K֍��S��_�,��3�6���u|��a{�'�}�u��ѻ�e�̉<b�1C(b��s�m6>2[�Vil�_M��9��	<\*Cy��gUP�d��@�Z��^|yni:��j7'�i`��|R̷ɋ�\�@	$��Ʀ���X�o�K
�Lej����OS��1��y�X�E#,>��y���Zh��O[[[�|t�ʖ�zĩ�o�;��7���ʔ��zES�?j���#���z��}��\F�]��L��FY*/�G����� ڂj�$==���SP:G�G�������ny��7R�K����M��W��V� ����N����C:yS�<wG$_�Z)Tn������"������Mn5Q̗F���wl�"5�����(�^kd�����70B��qZ�ܲ�a�T4�)���2:��rj$�KB��>��/
ܡ��4u��F՛����/o���go�O�9 �T>��A����i��U�8Sp��0��iW�;��_��y��~8|�A5�l��8	��'�)���s��Nj�ڍ���|�SF�s�Mޥ��'���<n0[��N­����!�uZ����1���(�e��c��+�(|R����J[�������yൈ�J/�8;��ZZ���m��p�68hG��3u��@��0�	�E2$[�I&�׉�g�q�4(3j;���Y@ПVW��=�
�h`&�B��
����D��l?�]X���G��{��
��T�*Z�=�d����WN����e�t������rQ�|~r"1�Loy4��Dz�4�Ɵ�{��_I~T9�/:�疝0+Ss��`g�Ǐ�q�݂�a�@�U�@��?�JCí�x���1��r\Z�za�Z(��E�����L����%�̠�Fض-9Cv��փ�_)�oLZY6t�2\yd��1T��F���XH$�.��k}�c����[ԮK}<���ԤYuS�;��-�9�
�#��m��j�;p�۴�R�&q!m�Q���<
S[��*N�ӊAx�Li~�-�*�{��O^��~�\�Fa��O�&��� �a� ;t�CU7��5w��91{t�fB\B�K۔5/��1)p�����w{�6�����Jg`��^iud���Fݶ��R��3}hJ�%AOl@�介�S�ܜ�����Ef��7�L����J�B�P.e��Õ^ �;P���B�CIm���se��Z72��!������"�'Y�6�[`��rs}m��V�n`/���"v���]�U��Y��xm��(�h\4}::S�>j����9�Id��(���i(Ń`:00 ��
�W�/�_����'��{S���y�Ά��{̔�����qބ�����`�r��>D�q���e%29h��^�a�:�q3j����ԯ�V�xv����+�����P��e~(���:�b��˦ nɆn���������b��뺷�ˤ�$�j}}s��DS�
�+�f�}��q��p���c#��\r^��viD����S�����&��A��T4;�Cm���A}�x�����߰딨�F6Lb1_���y�}DͶ-�GK�¶I K���v�"0�@�G�PBSE���T.�	n��.mRt-$G �j䩟U�ޑs��������7�9ܭx�<Z��m��A�^Sw�_,s��'�-��F�i��@e�m[�Fx䱟�L�g�s��s�<���r� ���B�q?���w���M�6��#��/h����� �`G�N��=54y��������M��Aզ���g|�z�c����%Wd�I��3�h` P=ؔ!n����_��)TZ���P@���v���,Lt\�<.��w�����f�
+׹aq�|���z����[:b�3��R����F�9��)���Q��őZ�A�;� �(,8g�~Ě�CKV�I�yN�p�����^Ya�Ǩ}Fjx{{��f%j�����H��z���A2��&pK��D�+í̋��]���¦&r�k�P9hR" �j�T"W�����֞%鑐�?Ev�.e��s�5�ޅ�ل��-7
c5U0�6�m�ݺvݚU���{u���������9SC�g�	��r�(X������Xxb�t�;A��+�b%�f.���N��q�g��T��<�*��&**)e�<��+P<'��x4�f�N)�������3���@�I=}���m�f�۟_�ȟ��CG�����7�d�uW���-����",�S��G���9��/i l<�GTDD��62���y}�wѶl�!�.kKC��7����
��_���N�Ww[��+z��q��#���'�J���� �Qj)���C�޲RW,B�׎G������^\~�*>Y�*�zo>��u
��-������K�0dＯ��+��W��M7��.�_D?+��z#^FG@�r��r�����9z��nSS�v�S�bRW����g!Pb��L+�).u�6��K�=x�D�7��4n��P�k��=E�����jF�#�ժ��$�=��ސ��#�d��oViT%�]`�xC�RzkU�Ű�l�M�tN)QF"��٢�?�b��e��놮����?�rA�/0���hd�?}d�A ����s�U�$h߆$s�im���sB�c�⩆�S��J<����AHs��kR�㭳���֖'��Go�u�ͻ�C7�|7�<��u��FQQ1AG���	���KU�(8fl������B��*U�![���)[D�����~�f���E�MU�����l/��L�^�G��y��%t�]<����)_���,��0�޵�F�;�Qq�En��::YP\�mc�<y033�lRg�I��Of�`�pO��³_�X��@�����M)�8PI��U��NB��9��Ř8%C��v�yaX�6�f`@���Sn�/��NjpO8�X���X����}a]�=/ܐ����m�����ݫF�ۼR".y|�����o�2(
�Ğ������@�ߛ�1;��^#�D)���%[�EV�漩�K@?�G�vk�dK����{�5�;?��j#�a}�Ő������C1�t)#rssӥd~HI����.��y�:�>�_g���%f���.�v������~#��A�~�-#��pC���x�\�2��� ��yK,�<��*0�W��B�D�w��K*�;�ϻG�>�r-���<	�AQ˙[֯:o��;Ք��W�1��5wAc�5 ���k��kwq��rny&)�4�#�xS�0�)��k"�;�nu�$�
���e�����ζ����g�l�4
\ťL{�M��9������E�/�*���b�cR����[1v�Z����*�|�w�ؘ���>K�����u}_&�*��w�jxxx�ٮ;�/?ž?(ix�n�`w~H��_�����Jd��C7>h|�Q�jr�4G�Aː������Ðf< �|��x�����q�#$�<���b-�@��U{���&�g��'�Q����X������D��;'���4��K
F���R[M��hgx�s��u1�F��,��7�X/z�]�
d˧jP4
Xg�.��𐮨�D��"oι��V/={�Iq lޏ��:���&���/�0}�_ж��� �e�+��-��6\����X$:�s�-z��#����&��L���hV��fo���>R�h�%��Ee[�0�����D��*L�۹�q��:gay\Ո��n&3��S1d��b|彾6~�J`,x�ȅ}]6_v����ʴ������5u_�
.6@ GWI�A*Z���9@Y`�Df���s��1��ͯ���v*l�#�໘H��]jU�;B�V�Ɓ��UMyo�,r��Ï����@6nb��㮱k�Nj
�S�S!>&nY�����{_Pt)�mS�3��o-.��7-�E��k��q�Prr2������u@��$�Ҍ+_��M/���@6��\鳐̇���z�އ�W>�`�Z��7�?�4���YΦ�Z÷�.]�"]3�5�����]�6�6x ��PUx U�W֝�O�<�X��2��f���2.oXS��Q)O~ ���FKk�gec�D���v��9����C�1�c�`�{�ۦ/�D|��+��*kf�B�(� ؒx�<��̘�:��*�W�#?R2	�tx��zɯ�˄�=oo��Ĩ�����4tIv���1ј�C,��X��~{�\�s����1�@���v�����ݟ`^t4Ee��G~�n���ZU��۪f����rt�3)�q�e3@w0@ � �ן����FE]�T6��͜��� �]aQY�Rr��I��7RŻ]x�k�eA�q�<F�zP���!A҇��t�;�t��r�����:�i���l�u?�!��b����ɋ��� r��ҏ�=�0ԗ�O�WuR�^&zE/87��>,�&+��c>~W>"�5@X����=,��~�ر��W�~	620!�.@�M7�O�X�胸ۊ���E�^�WOpe��<	>'>u�<T5�5me�'%�K:<��2�����H�&dÕ�<�/Ͻwp:ɧ���~�B� t�BQ�U)��~�RO������1!##�����x�m���&�$�yP�ytE��W�#�}$��~�Э}O` b�B��h�5�ҩ�`����*����G����O���o�T�AH�DM��¯�� GӅ�;��i�����_��4�L�@��?����{���0�����H陪LJ������m^$m����(�(�������Ϡ�_	
v��ߏ�||4�2�i7�#�*�T���#eZ�ݗBg[4+��~E�u���?�;M��`��m5v�Qɟc�6`u��m�ԉNt���:į��t��]e+z�)t�i� *�1�3 �s1s�j��09�&�B����0XP@Q)��=��N��%u���w�g� 	j���w�n'�;�X%�ߎU#��������K���f��mn��t��ټs��v��J%�I� �y�$\���[�uc�b,��5[��4�2���t�/���~�Qq�f�y��ɖsF20BFa�'j�
J���iMew�%��6�w�զ�\K�1=��/[�Z�K9d=$�Sq�k� �bc��. �D��.�l�މ콹���˻ޭ	R�5�������{�3�:LR8yO%R�Vz��r����g	�	�#Wa�rk�^�ZH�W;Rs�`�~b�`n��	�[۵�
2��uF;�X��V��;���E�Ʊ�nǑ��|7����Kn4�0qx�2�
3�һl*H��8p"��#T�L��\[G�Є2��^�3Sz�hhz4}�s��8�!��!��=ExNЪi�dG�K�r=����1 7Nv����H@��uu��� ڍT�!&���ݏ/�za�T�q����u�&���9���x��CR���r ��ҥn��][С�|0��b�&�n�Owv��Kъ<i�
��C�lV4�_��nY��u�p~�10��v�L�P�Щ���q��n!�?D�@8��1�R�N���Ӱ�����P�@޷�����M9��]T2t���]Q�o��'z��,e��$x�6"���ͼ����K�{R���^��c 5�6��W����A�������M]�j�[�-7�W7N��F�j�Dj�{^�J��s��f�䬭KV��6��\v�ҥ.2D�	�Ni;>m#�L?I�9��nyOCHtPKu7)_��J_��9qFS�fF� DPċo[���v�)��9�N*�ZTWQQ����c��t�%�,��?�K*��v�%>�]-�E��{�s�L�l���w�0{۞���k��u�w)�˜�Ka�/37�8n�����_Ż  �{������^ߊG��եP��Y��Y�}nV�	��˽{�{���5��3��/�S\y1�����b�N�0E�2%���ۏ` y#��PT곑���HIA�4ȗu_�${�yy/� t�m�ked��I������jr�o:�JYY�'N�9Ȇ`�/B�>#��ư��p%|�x��Q��qYf[��p�����R*�*H�c�"!! ���� ݠ�`Q�H����t)!"% �t>R�����~���}��Z׺�����w{��ğb�/!3(�4L�J�rq@��Ò�,��YN�/��8��~P��+*��R�S���>������#���C;��ɂ+Fp��YN�b�@�U����.�]��0���f�$d��C��i||y��Z��`+ *�W �og`\u���}=_F������y3u����^����f�v��ϼ�V��Q�ٹ_=d#r��|d�BO/	��Z����$�' ��}�\���mJ\�A���&5U���9A��D���)*)]?�3ښ����tt�Ed	g �	�<
�B�ɦ釩�zƿ��6e`�Zp�á4���.�i|o���r�#]tf���uDx�F��8�\d���,L�P�Y�eA�ys�~��Ă�!^<�����է��n2n%���g��y��(��q�������k#���F!�i���a
����I~���*�U�.R>^��D?)� d��o�GK��aѹ�?+��dd���}���١i־Z�il�X��q�Nq\��'�"�j�����d�Za����I!�N���!���|����cB4VWm����Y;ͅh#�Ј+!��y��`~�Ҝ;u��C�օ�n2v��`�c �I	G��*[���c�?>]������~w�r쏍�8?�9P|��l_7�caL���.e��o1��hEj'0�$%���?N�/Q�W�A���2�
�
�:ζ��^�&(s�MʾfǬ�Q��]k�lԳ$vxK��9=SZ���Ņvj�q�#A �����db?����l�%��^U���&f%��+��x�a)��+n�cw����jq��f�9���ȱ8aINi� �:���=�������Ǐ�4�2vX��>���m�(���R����F�T��|pآ�c��<�\�3�5�<�M<��yR�M��|n���~_�����ʺ��%y@�ǫt�`e�T��k-���( GL
JB�&�ivL~�	:�k�vK�k.�^^�13�t�-e����Vd�^�.B�����4`"<�]��)���!(x��) ,5y*NB�9R���!��e͉�[L]��|��y�ӑ���滪$Wڠ�x�%��{��Hy��?-��V����u�Gz���_L����WڟO,NV�ʘ�౐J�sC�>x�ZPJ�hct9��fmm��f�� =�Ԡi�]�o-"�r��R����ț�'=�����VS��(i�H�E��[:L�����_��@�;L�c"�t2@��Б�����_�_`U�wv����ؔ��J�����<W%(h�U��]�����H̛_Y���$ux�ή�������/mY�ب��p�f������>=>HpJ�q(6��H�(�Xk7�V5f��l�P�Ԋ9`!�CBC�(i���̆��+O��f�h-��v1���]�9`ЛfW��L�#�\S�Y��]r��!��fO��d�;��|b�u�l�UEGGwg��WTq�A���hg9福���6��=_r��5<
�&>�9l����S.��g��D$�T�E.t�t����p\!���hcŢ,xO�R�b����܉@���Ts3��7Р
��V�M�#���Ę٘f��&K��^�4�k��۷��3Z�;"��즳�gk����m���ϕ��8�ɢ�4�b�����0��?��qX���uKk�9��!�Q1C\&J�`� �ņ9�ք����ރ���{� @��p�Q>�F��GHw�Y+
,������/4QSX�k?arD҈[��qa�='��G/��5����HT�O���y�\�\��p�` RJSEq"��Ȥ<j$5�|��"�{��o���wwR4�N�P(/���prFdoYr��$g�y����α��a1�`�G����j-D�)r�[���sK�T�����LWs����z��4@+��mK/���Z��k[���F��@S���H[��dd��������s�/��ݝ����,>ZX|=���̯�2O%H�CNW��*(�AHb���0�����F�Q:��2B
0%e%O��q����I�݊aFFF���+�ǣh� ��ўc�封E�����i+ݨ�ݱx¶��yp0���篸�j#�Q�Q{s�rᜆ	M/�'�.:^}�l���ʶ,�cslsBn�(�:�-�2U�L��K�ؒ2?��������8�m p�������.�꩝�����M����\�4�;6	kn99�!y�M"��S�\W��*�@@�9�o�///���{��D�`��DV��� �
��~�r,j�Z>>��m#ZePvD���,)��/����3t���0�E]$��;A)f;��K���fJRCva*�I�����|@̑����w9@l�v�{�,�^�=�88�K�en�ΰ|F���'�@�"ɲ��%�Q��7?�����Nေ�ѻ`��og|�N^bۯ~5���He��>lt��oNnk��V�m�=�\����R��@�'W�����UHт�r�|����}��]��옃K?�޿	���H���L��?�;EH5ygD�j���f`^��r�����I� ��uʯ��؏瑴r��,*e��I�l�a�6�nл�+v��46+&]��1@>q��Jڍ��v ;H.����Oԓ�6��I���~u�F��h���4o��+��il5M�f�u�"K
@4�xWS�a?&G!�X����m5�ZZ�������U���)���[x��m?׀ڍr��Ò���7У��|eh��TD��u�۩�g���L ���)�ݛ��o�iʥ,Q/'Qk�ٽ�E�CfN�N��-!YV�J��9F �t��/�$��ʲ��eJ�~xz�S5,��y��C��yh��ڰ$�dG�������0���j�\�IB�ל��tD{�k��H��UR2�Wh���-B���ùB�9��"6�;�d-s�,Yrs>�"-О��!}?��3�+�/�!H8�f>r.���w�̷��p|� ��v�X�������L�"_���B��;�v$������{�<�2ov�O[�"�����f&��{?�Dه����q��2�ha�4�ITc��N�k�]EoL�/P�A�bd�n�r�q�F��	��#�����l���/\����Of��l�)�� d��ȯ��A%�-y55��u��u�u�;��S�1V:�yO�9)��EeFd>\��Fz�,�b�x%_��<���wfH����|�h��3��0&ܑ7��H��l��`_?/ʷy�Y��Jx���2/cs����,I��9�E*�J�I�E_����� 
ncc���KI���������y`L��^��IW�L���}/by*F��4�l��g��S%����<�g���CJ3O�[Z��5��$h��:LV�Ի�W���|�tX2Һe�늡Cs����c��-yw%��,26E�:�0Ҝ�
��7��;*�	�wOyG=�!� k��OxY�-N�^ݦfP:?|���c[�QՔ�w�i������1B߂`ZmWD�C
#-=���ѯ�֓f�#�4j�Ә�~��&0�2$jd���"<�ԑ�d��I�^t�Z?�\G����q'3�e�*�uk��u��*E;=�N�6��t�����d�JnC
^��Lz�+7ė�����I��<=-e[��CǸ� �R���^ W!�V	feOpc����v̚ۂh\,��%�ڄPOz[��d�yaF�X�����	�zVSy&���ҝ#��gee6o+�-i����`_��ƽ�b���wwfC��������������o$m���X�Հ��ҥ,�Tn��')��I���Tr���&���ÝƲ��cR����hhtk�{���(����~ץ����C�ny{R=[=^=�\8�T	�����n�L]Ĳ0V��ba�Q���2�_ř˟���Ӛ�F�c$�Z�mLm??���DL����of=]E�a�U��09]��0F�Exz��n��ݘ��]�Fܳ�X��[9]�Wְ�����4��pC �YDh>�]_�XN��q3']7�`�옷�d�U���za�����con��Gޡ,p+�b%)���{�|����(5��ח�4S��G���c:?�p3��=���@��I1�y��f�j�?�8�$w7l���}+��}��G"�`M{]�E�cܛ4�
:�L3��L�P�A�q`b)�>.޷�a��Vk:S��\B�(Uܡ�E�DT���م�A����xn���Y�iۮY!���T~�>������	X�x��\͞�*��b{�!�z��!D��u�<} P����Z�;�-�*o#��#\���/k����ܘ�Z�!�X�*�GqY/aʑ'X-�x�.)'���?����Zy��,Xj-�f�L&u�ؑ	,J�F���	ׅ��c���
@4="u����p��x�ߎh���Ǉe��r7�s���ܫ��&��$a���1f����.Ї�UZ����{�ßo!��q[�u�Ѯ<���s���u��=s��
���NW-Q�݃F6�A��r�FF�6<ɪ.���߷۳�����i��VZޝ�p���M�Mm �/��Z%���?AA��}#�Wԛ���H�Y)`d�v�+��ӽ�N`/�p6h���ٔY.����u�b�r����KY�A���Ʋ�P�����.�m!�+}�$�h7��ܨ���9XៀqX}��kcN +�'���z�d��1X!��k���m�<��:PWoc��4�g���N�y����̡��9�k�$]�7���#Uv����m�j\W�^��,�JE`��Q�T�oW��A,���'�|=��'��ChRK�denњ���8� �]`a=�1��:������̗����������k߃�ۏe��a*�'���U�^��9�g?��Q�>aR�b�XYYy�[e;]f�M�w�ߑ~B��r�@��h�����Dc�������0��ɫG�_^&��Pv��ݻ"B��R|�B�F:�o�+q��e��O�\j:g�^��<[^�����/����'C�O���l�/v��Xs���%/�'%v�©� �啾�n��@y⑕ҷ;Nod$�ؒ[��{��Z"�
�X���3M��2>YG1�����#,+aR�ķ��]�P]�˅�����b�]E<Kwv��`�U}�폖�����]�ew�2s��̕i��+}�����A��E$=�P����������M)�Γ���xu�y�D�N�#8��͹�0�@�O;�ߣ_��V���$�A��+����*3혧�쵦�}8�'�W���_��9l���U]N����a�)*(�`����@+�����׍�} �@��M}�ͱ%
��S�����W��.N��4�1YB/��vP�N��[������ޠ+TqG��
f���谰fP�ll�n=^���4n�,/��	X`V
�e�{du�+��NsZ#F�>"gr0 %�&T��T`Ӥ5�|� �/���ϡ��/Q�r��Ή ��7=�Z)�}��.�C$�	��z ����-A����\mz|/z��{�9SZh*����Lڞ�q�iA��S���YH�H�b�!�a�IH#������Tp�09=�	�h@r0�=L]%nNbZL�#w���l�)�S����H޿ؒ��d���m@r�"hw�i�)�̋�2Yo��jk@�{`�������1<�L��l��$H�nT�vM\���y�My�Ie�@H0��Vҭ\�k'H�yOTF�#A�W22�խO���w�e��(9�Rn�@ꌧi���!=$��f"�7�@�!�5�4�8\��ԭ�a��f�f��ee1W�߭��>�܄Fo�q����|�TY�+�*"}d>��Fms��f�Oa��B�����%M�t~�ޭ���8Hkl:EM+
�+JÝq_M���d�-0"�M/�ؔj�[���VCb�h꥿�z)���l.�}��<�G�H޲}?�f;}�+�⥥s�W�y�h--�����ZF�(�~���?�n������Џ,"o?�Jk��,UZ�x��v��茍�U�N�k����s� -�Wօ��.;��Ӓ�J(TO�����n׈j7+Ò��o�;�`��h�5ګ|F��@ui�f"��lي��*����]��>��-��y�Wfq�㛆/�#*E���xN$f��d�����ׅ��
Jj���_gV�5ԕ���
��֕�땪�x��������b��i�)dyG����u���v>�Z��<!�)��_���Kߴ�����^��n;$%*^c�2B/���,=�����8Xq:][1����/��H=���:�|_M�����	r�b�4��"�����	(T�&N8p6&&�gE)\>��6���L�D����]���blC�y����g�A5�4�d���%0�2Z�Ӿ�ʪ(ڀ܁Iե���=�A$�u�5��	�M�}Q�d����NY������B�-���׻����X�j��a���)P��뿇�&)Eˑ�i��an���+�Mx9��tN�M�H'�0���WJ�9���vBt��!����u���6#,��G
�j�\�vm��@LU����r�sq��ߵ�;*�cb~K2�������9mgg7�������ű«�yLxKFW���ƞ�K~G\�dl�g���]\Ssa�3ɿ�ߨ��+p�LX��|�~���(���j�k��-�Y:i/Nz\O2��Х��}�7��V�.�����zX�3�LF-�^9�ir_������2�4�,�f�U�4�ǩ����ScI�i��y@����Q��NHvNN$�Ʀ�Q;��F
��6�b2/�,]}��O)|6�C��>���$"o;[.*�I���Q��4�t�b�q:d�&�PE
�Ν��(�<���2�nrfܾzu_�������	�J&�+G(7B���I l^>�{xG�r���"v�]��&?���v��U��S�J�+�X�^��d�Y��X���ȌQ��7�������[��Yvw�`}}:��,�v|�8R��ق�%[�h��:ٝF�_]�~6;y�١l���i{�N���A��޽
-َQ1�%7�8V80`r�R �nC�ve)_\��K>>��F�:��S�M��
y2���koW}J7$�<m����A^�ʥ��.����=�w��.+�bUC��}�I��f��� �`�8X,��hF&��h�#�������2U9G��YlK)���^�#RR��K�E���	/������1��/����r�7�>�EP��&�R7x@�p���ano/�s�xj�#CYF�t�f�zc�жc�*"�[�B�x	��1E�¶dIH2��Jn;_1]O�<�5W�C�=��G_�
d,{���Sڬ���-��mX�K޴iSI��0�n��{����
�TE�b|���"?��0�����|�	w�g�.�F#V��&�>��l'{�7[�]9m�Y ��%����[�6��Qr����,��2�DZ���\�����_<F=����y��۴�=(b��Vbx�F��[u�����H��\�c�=1�@{>�@_��aJ�'��!U��q8�al�ȑqz��W
s�v) J��9�=��~@Ѩ�~��N�p�v�)6�}T��f|'����`�*:��R25c��>2�&C��*za�`'$�̟�v�Ŭ�����A���.��,,�䣞�3�M|ؠ����	w[�W�}����
�B���a�"���`#�S��Ĭ�ج�;��£���0X�^�HiYq�ۄ�g�e�c�TI��
�4�M�+s�M���8IZϨ�PDr��ў�����K�w��d���Ҽ P�)%�\)���!��/**�^��}$�>/���G��;�l�v�˶SW�6�������D�w?�Ea�r"��u�K���v,e�HD�:E�tݤ���]Y�M��.�R�,�t��'�����n�|����^$e)N�E,�{��8���-_����;?-�4��߮�q�f��%��ڳa�%$Z�Flww���5H.1m��{�r��I�!l��;w���7�;���0L���O��k����9Ӟ��053#���<�)xLBb����:�) �)^��7���{��г���Ff��8&d�%�3݋Ǹ�n���$��I,���k�a�E��(��-X0��=�g�s@��8u.�����n-����z�Ny����� ��޹��G�AR�)e���r`�ᙃ��r�>J$������CO��B���~��Y�|3B�7'��t��1U�����54�pqq��� ���OOPaxA�t�ڳd^ }}�x�6�5�L��� �'&n�F�hfE
�� ����<��H���>5>&��hE���4���Uss����j�'�c̋�.0�ќ����L��B��;��<q�̈́q�d}0&B)��<h�ƍ���@�Ѫ���e��6�! #�w+&|�1J�9ި��/���Y!xF�X&(qp+P�,l������"bV�
I|h�)��ՍQ&A�e�V5�T�X�c-��f�g.�O�����F|�!!��@�xf��4�����Q��7�2��s,{��f�>�pbeeg�:������a������
��NzT���Z���x���@���-��2��}^���]�h󪲅��\�֡�1o�V@�7qq���uј$B1���d~��
~�F��y��#;[��x_|��j�hw��v�+Gl�Ϟ��k'@�� L_�a���.�I��)�l�w#Âa�c�O���8��-7X-�g.�BCp���nX8#{�9� ���HE�ջ�28!zޖF�{::\��+c�������h��ڪgnn�]E=ѹ<��S{�S!~�VLW�7��$�,��s�wtt�����\�c��{h4MVz�\�=s����6p�݇��===_à�����Փ��)���M4'��i%d�t�D�tyQ��d ���Ъ�<7�!�H��*�1D�6!M�d�ک����=@Y�e"|�#{����۱?�5��-���T�R���|��cf~aA�g�祀��y�> K�I��¾>&���#���jl�UE�h17O���vWtt�	3y���C����;x� V�H�G�Gr�����[G��J�op�m;�a�g��ҬR��=;����8��B#�@�c��1�o�n+�+҈u��7�b��8�SH�*k�WN�G�����d�q�����14Wֱ��lM�Vɢ��˄�S�a?�]����>�촶�����*)I�F�6��fؼ�4�hn��N���}�\+QT5��?�:�6��t�Tm�D�F>�v�3$d�m�V�fb��<1-M�gv����]��������JryW�:hh��x�UtG�?A�"���3����p�6��\h >ؒ��y7�j� %�)ioz���6�i��K���+�c��Qe|B!�bء����*����Փ��B�Wh�N����K�������'0ݍ�6��L��?N7m$P@�1&��%�'�FT�(��	:M�?��2���U���}�����k��� ?%����U�ꂉ�����������*TcҰ�R�/J�\��#pB�1U"*v'��T��H;~������-����0����=@}	��
ВA���>����=�F`rF���1�E�|(�SE��m�@����6�C�rtrR3vV
��|��sW�;lX�|�	_Aֈ]�3��i��?b���q!t/��[�����m�xs<�B@o������zu剷�� ��u?�Z�L��[����?E�����"f9f	�����A�8W5���>�jH�޼���y��h��OW����P{^��$�"�:����X�p�`Oqo\����`dQ�Ճ����C��6I-'�bd�-?T�e$���##����Kg�b�iy��چ���|.�!�m �ސ�wF���{DpP��q�%)��V^�́ժo��XҚ���:��.���w,�#A�<� ��9 G҈U
�G���8�0F�{d�i�6��J�0@^<�>�O�LA�# 6�����=�U��r�?��Z�?�`c*\�fFR��v�A%����� ���zК�;6��?.���ۢMS�(3c��%� �*��-F[�)���g�hy�f3��Խ�6}`x��/��:lO����Q/���n�w��bn2|��2�W�1��*�V&�Tَ4�Z&�SB�!x�{��E���b.\�t��r�;�%�N���m�����A�'T,��$hhG�=�y�hܔ�]��������rG�ٌh�_J���^����.���ܙ3�Z|�Fb՟ _>-`<�٘YY+:y�鍓�'_^0�j<h�H�[0{���~?m��7�g��I,ި���������I���n<5��1�����2�.ށ]��_�����
b�,^D�>tE��X�,�8����3�����Zئ�_jeq��4]ᤠ/��C0����2釉�;���V҆�R)�]� ���0)�d`�i?dsO2_������)E)�NI0w�%Q#]'�|�`�	��Yc�j���eה;�3I#���e$��r<���x�&KW)��Y�Wa�+��B	�;<+vF&B9�n��'ɽ���&���{ϕD/�����L()�hG�3;SE�RXx�WY�P��k�g �M���\(/	N�W@�`k�2xz�{�&���=	z{>{�Ī���x3]�DnS�5��4�VQ��R�m@ං،T�����4�`L�&���{���i{��S_��a�W/1�O�]�`o�w��Gц�ڒnj�+�D8HX��'f|�v�'jj��>p�5X�M��� ��|U]�B��K�6rG��b���F�0�#""\Y@�HU�����9�W2�\[��)���1�W�����梩f�ٙ��D��¨����m�)�����
�Qs��+n�זC2���������.?�aw�B�:����L��6,��w������x�VS�O�C���YԺ�=f���[00(�~Orr�2K����L��X��{�K�
���cOR�-����� * �֭�4�t\&�]�� ⛅O�
�ذx�4��f�(�߹uk-D��)���� 8x���͛K�*C$]�ª�u��}qNN�L*ku�\6�fJ�#��=(5����Z~���WBq�����/_qv���d�y4i�RD�Wp�c^�R[�T��U�q���ۏ�F��	Fb��ѣ�\gÊ ~������7.'�~~��3�1Ug� BQ�n�/�i�_`�9�O�I�[q�yR�~���H2tv��/��	�e(.��E�6�!���Pr�L���,���v��s�;]�b��z��0[�G՚��U��z�?=d��-#����\�2)2?�N���ÍIxM��s��son�[��a`�c�ð֧�2/�L�����7zA�Z?l�+H[�vv1U��۳m��W`�'o9v�ϝi1%0�k��F�b��zϟd�qzg�N҅�{aU���LR�`�`���7@��T���M����.��'D<yUR��o>�=�Em��?rL(�L4x~bo���(w�����6r�N���I�NEr�B��8m���<%��[��'��p�Iw�/Y'7P�%�������x�e����f��Sw�и������;��Mu����X����Ζ^�l���t�ȕ�����3ݎ����,��R��^GȪ��n݊�/`104�_��k2�Kx���8�n$%)|�Þ*���m-�"�zX�R����.�	�Ô�2��u]����v=!�`0������ß�c�l��,K��i����"�+��vc�I��\�4P�:3SϨ�ÞH�L,������"r:J�8_�Wd"tfEF>�L����� ����p�����$Yq����$V
�C���2 XՄ�)�t?)1���B�B�b��l?qq�7��V�>w1���n3O7�W��@x� 嶤-Ex�*��\������[&��7� xE�8D��G,�h~ZNP��M�SB����Y������� jO�QbN�e-���H������ `%��`��8��d�3$!����}*A��;@�G�l%\�.؄k�􉲜�<^?W(~�
�m.��<[�	��i|a�.S6nKӤ^�T!KכvڢQ��YM��a�y��/���$���������6r�b6�7f�Bv�'��í|����v��A�h�e��š��4֍nÌQ���K��G��,�Pc� ���ާ�Aߪ�����`>��q��"�Y�� $�ԩSy��||"�rHp��vb�@`�1-�����|����ĭݟ �xR;��c����^����;X]�����%��D��
�MF$mdl��~B�L>��&����&��0H�a�)<
���O�W��׫�5��*t�=? @��yk�E_���욨�+�q�uu~i/!��&�}K�`��m��ok���iʴ0*�΅����{�f��07��J��w7[�t�C?����,lYdAp�s��I�ֹM�F	�
,|����=������6���.�2���5y]�֮X��Tj&�d���*��:,�ȏ�9<����%u�.j�]�v�e����a�g��5m�N������jٖb��_�� ���:�2�=��@\"���g���KՔ��%��|}�fh�?FÂH��'\#'P��4IF��?Q��ٵK���<��)t��SXTTt��<��6[������2��a������ק�] SB����a��A.)z�9�p���Czk��X5���R�:����Ae�]���7p���
g��a^���C�����7�?�J���_��K]�W��G$��t�6ƪ��C���槭xpU�4�ʻ_g��ϱ./u�Hs�w�{M�����ux Q+��Ex
�2)�u	H8� S�
�t�/�7(_�����SkQ&8�Ç�Y�\+K�Sj��d9~u��\�q��VG�8ѕ��sr��ج����֔��\kJ B��
%�ӌħ��u��[�-MF>%v�y��^�ڗ�<?�4Bb�c�����aEz�Ios�t<:4-7�_lҮ����!��Mf�?��_;<Jp��R����x�w5��/��{� h0 �AJܙ�C�H�%����"�y��$� "�òt��FO�q����� �:��(�����<����]�W��>��.�LSK�,�|�o�����9�M� ��<��*g�N6Z��.���	����ծ�|�f�/�{�t�X��?��6»���Z�.�w���tϮ�.��Uu�����66�%� �Dn5�3��tU{�g�T�{2�D�E�2y��؅m��MN?u�����Q�U��<���c1{-�]]�!��t�zuz�U�<�5V�������R3NLL$M�"i˙!�ś��2K�� 9 v̆�u�r/�zI=H��u1��͕�0�т,���i�������b,�$*W��=�@� �O ���q�ͷ_�
�I�8o�z�VK�!�/М�S33���0�od&ӜMZ�AfھZ�G�lW�5��ķɥ;��V_"�v�͆��z�~ٹf�,�}#����ov�WZ�nd����a�������Ӊ/����������arP���,Tc l�tf����`�r�4ʋ��QO�ż��b���>H�6>->���C@j���,��e�}))�������o�myt��~�$dvq��^KP�L�'�ج�m�W��b�p�O���Y6��NҪ�-5���G��NM'����j�J��J{z���%6��r|�r[����f�����Aڡ�,���f�C|�y�w���/o����޼sl+�L�� *^�n���2��%K��)R#�4���2X6��֏�}9ߤ����+x�2.�abZ�,`@��4T/V���%]c(a��7<a�f�邚ȶ�S�XRK�QG��a(�3�MX�)S�č�:qi�
�����R�v�ik��rt5�*��'��v��aǘ�.�]�/ΑNL�C���:����[ Ɂ�sa������>а�5��0׈�/�*֫��M^|(\?QH�P�`����Ç���R&OA�cͰe�5G܁}�eD�C)�#6�o��`T����l�����y����@�!����x�ei�5��v�lW.����
���	WApG!�i֦v��������L�"���6��Q��ӳ?�-�Gn,22RE P͸�PӲ�eݲdH�K*"���c�����C�E�v ݸ; ��]�[��?�~�R���nA��OҴ� �q?"�thy�s�dn���E	iF�hrrz�2KM0:�@KeW�3���3LȚƋ����?.V�Bp�x�315WE���3r�\��c�/z�~>`F��ggٽ0��[��N`���S��P��ʂh��>��?ءw�(Z��h0���)Y�399�{^hrE�������%��"�������ץ����٬gGy����j���]Җ%&�	K��MCq�ef?F�c��_�빟<�4�����o�0!k��վ�2�7��2�s��`��?^�J5Vx��J�c��Y��lI ����	=�@��e��!���o>*C�<r��?�h�-Ja>r7ֱr��������S��vE�m�h��9w�)�{��]��_ʿ��߶la.׬��#�UbXG<_���d7�h[��y��7����$�rcQ�3���J�q�d��:8k��n�Fe�� o>Q1�HTR����z��ʪTzeeէ�Ƙ�߀_����b3H"�yg<	�N�%i�Ƶ����A
��lŚ�z�"ۑn��{����~��Ƃ�*1L�򆽎�h��YDx`��Y�^ܴy��#X����w�B����ğ��mt�R~�r�����+��y\����j-�#��oE�q�yze<�q�&��DJu�Ԙ��� &y�R�,f1x�4"��s���29vb-2u�ϗ�kע�'9�v�vt�]���G#v����4����	�;+�Ԟ"�_x��={��H�c�^��Xﾚ�D�ۀsC����>BySS�=5|7��Q7�R�����i@�'+ӳ.�g�-�BWE�ZѲ~�,�9�ng���=:\�2�;!3$k'ç��ꂠ9�Ֆ�硝�툛~~H��kݧr3f�u�8���^���jO�{-��o��v���@V���C�&d7���m�]����ɑ��Wó/����qi����W��d�nza>B+�e9��lm�bz@�;��o/*\����RO{� �*���"�y;�HY��t�I�mq��T"�K��t�,�:Zl�dd\�ZZ�@�:���콵��$t$X�_Cҫv[�$͝��@@��"���U��`������odM^(n�V|hx�j3�@E
���Z�IiF��U?l�{m�j<����+�~0s>&���q�R�yk����P'D����Wc��7~��⪅`I��ɧ�6��'NDG`��>���%NNe�8$`�x�$˗��� �Ng�ö���px�4GG�վh󪘪{�a�xyy9:���t�����^��O��_B] ��7��#|��B��˿�W���2-�����i�31�0s����T��(��u/p�`	3�G�[�Ҙ]����`/��o	:���	��Ǉ����rz=�N��N`n�P����j��x��\��ҵ{u�W\��މ/����v��� ITh���C��� �1[Y��)|xϞ����p?�J��d�G�n��&��mYV���7�8�B��l��4���T;0�����~�ؚ�Tx3lV(u�?4!����f����V����
?�=@���;u��e��ؑR���yٌ�kƶʍ9m8_a1�A�ѳ����s�� �Y���9ݤ��6�f�T�d������a1����Ax_�����^�i/ͻ��s��3���@`
f]�Y^���q3������s�~f�����8���ǹ^:��_k֮7is��sj�)�|�mq���Mw������ռ�}Z�@<1.��fz����i���^D�����R���rN�Ä<�[�M8��f@��_���d�� ��t��ޮ(�����_���_#R�O[?mgcS200�_p4�ʺ���m-)`���D����0̰3���i�F$�uUXn4pk�$3'}�	w�}���bڬ��rcmO�'{ܖ\��Fg� 5�X�P��?�l9�FUj�Ȟ1;=M*�Q��$:j�QUA����x,�mH�~�+ى���сr{'@%	*���	�zp X-@�8����C�nq���#Z�����C�R~�L:
��:W�ֱ5�����c�3�?��^A�1�v�x:��x�E�r���	F5��X�.�����8��'ؓ#F�qc+�'�" *� ��T��~�V�<f-'�:�7(]Y6qsv�Gs�N.ߠFq�`ǆ�y�6_	��c��9]�D�ښ��{�Z4��Ar\1����M��ã�6~��l]���uia��l4т����9�]v��=�ѕ�7�k�A��JQtJ���|ie�����l��ů�ܾP���D=^�D���,]o�dQ����)+��řV�?��[p�hZ���o���Kc�Q�@�}��Y��P�����FU
��h�2���xg.ʄ�p�R�� ���gNoA���+�����g[J��4rB?���X�Nf����Q��7vyɱ���,-����-�q���e��:������xX%q�;:XCfaayT��+x[zYĲ_��J���,c�t���1��]�(W��} ꖜ�Y60`�V�ø�:"�T��Q_H�o�N@�����iǡP�hX���X�Uk�AG�<���V\iC��+�kp���)+�z@ب���e�X�^yNN�!����[�WZ� �)s�ssW�e<W��&���,l �ucc�t��-ȭt�����U �.�g]w��e�Z%�G�l�IN"W{w���jQ�xL6*���P�|w��y,�~�L��Az���zÇ�lj'\��;v��m0&�%&&1
.�t0v�ZRE�]�䴶��6Ņ]llؒ��׀W��p�[a�=�l�y�Ȯ��X�|8}��@^�*�z��ږ��
sW�9a��̉I�����1!��%i���� �ϰ��1�4ܯ�V�h�����8��ݕ��Z�\$i�����a���缼pزߠ�<p�N��g��<pK��{��s���x����E[g3o�Azz�pS�
ox��\��[��Z���}5�w)�&���=���9������ޫ	x_�^�>Ӹ\��$��߻A؝�j�����k�I�Z�mڷp������]㛛{�������ݗ����;�R��~^���/����&�e��z��Go����(�Cڕ���4�d���+�m"�����B�Q��c^|���J��׻���BB�`�����ɰ񁮢�\��A�/�;v�<�å�������sp'{��%i�����tZt4������?8�Pe���>lQ��l�樯�M����&�?��'L�g��Nxz$��fUد��z�Å�A�q��ә]
 _i;��ׂb��r�&/O����g���K����9U[�j,8���Y?6�ћ���H�E�]s��=x��eJ�ȧjr�-AF��i��˯�s3Z��߹�ٿU��9��)w	a�-Z��ˉS֔�i��y��x���V�wG��G���b&=n���j*o�tPTT�Z���J�w<G�w�aL��s=�A����}�Z�2d����ǞkE�d�W}���_�ҡX�	E����t~�K����#���*akN^ay ��i��O՟����q���w�|�n�ڷ�3&?�p��3L�M?O_pD��ʥ�nJ&H�b�9J�ܥ;��'$�Zw<�}������c�~��s����Lѝ~o�����=���c;85X��Ln��d�o�a5�G̛�q`��`\�������ԥ84sڿ]>���汗Ns�]ͻL�U�/)Ӑ��1&_Y���}�(���#nǦ�=;�+�X�_�pџ�?��K����O��8���w�w>xI�v����I 5Xܟ�.N덜�b:{U/�o��9ⰵ?���>�{�A���9N=���B
L)�Ռ^3���wa��gnf�5(N��v���-O�s�x�=hI7�rf纏����W?j�0>������/e��-za:�b����{�k��������5ΘG��5ȍ��l�vy�V�7��1&�_���j\'P�����
;S?�m�k�gbb��4pu�{�����8u�FF\#bMk�Ӵ����7H�H���J��@���٤������`���|Ϟr?��̣�����-u���g8�K�D�]A��#v��_Ue���+��y8y�,�k��f��l������o9[2��%EWռ�7d�j���d�CSk��w�9̤�OoR�]���\dpD�C�tD�p	����_�s��I��kM�7lؐ�8�6��z��܇I)�G�v[F�O�2;�����*a����g��fh�!����p�'�r�˧W}�UH��>�rwE��cU���6?����0��qk݃+�Zo5�ut6HV��L�n�������Mo9�x���1��^��?dF��ҽ$ey�I�i~������G�!p����zS��)KO?��*��/c6��� {�y2F)LU$�Ar<7���� ������٤;����8��<=�����w��eFe���[�Ԩ���M߶�%K��(o����7}�?Wi����Y�����3�b��W�W�d��9mC_�UT+1�}*9�奤l���'1���Й���aw��g��x�x+h�5��uKD�nc��$��W+�z���K;N����r��
�g��A���D��-��k�v&q�m�-Uˈ-=�Ƨ泵�,cy����>x�-���~:���yzp:%{����gk	韖N�j+
��=��b#O��*��𒳡N\��w�4j+9"vҸ�=����uG��;"��/�V[['���	�&I����s��ǫ��6���`lM���zIQY�g�3�iv(�?��u��˻�i��.�R@���oUcM\\��9�������C�*:�����a�+��z�Z��G]���(�LO�tsVAd�id��L������)σΪ>���O�ˣ/��>����
�L�����=��e����ۼ�,3;�j� �?{Eo3S�p�F����7v����o�Iφ�-=����/������4ڜj��0�.�6�����R���p��}	z�jit��_��$ ����!Y�������`~P�m<�2c���8�$�k����x�n	Q��޼3YKA�Z� �����\�յ�~����t���<mӮ�<�9���7�x�ݹ�7^j�F����|Pz�9��{�ii�+��T���:��>���r����t�qю��M���A��בg|�s/p��!I�Y�G=~>>��'���&��g���Zh#��\�`LؽyE�VU	��SJ/�r�@k۬7���v���&''S�L�cZ¢������;�ͫ<�*˃�lb/�b"�1
�4�����=�I��= 䊨����,��ߨn�D_������p,����T�$IFG�
��le�gvvFh����l/�+�!!��MIVFF����}_�����s=׹N�����s>�w<F8DM�b���~<s�%��������Č쨳�S_S����"֓ٓD/����<7	��<����Q
m����hC�=�K�~\K� Q��7=e��{:����*-#�iA~���}F���hD~6Z����>��IG�:�������/�����b�2�ѽmQPD$�������@g�@�ӹI� [+Oi��L�� <��L�zg��S)ޫ�G��=��o�����ks��T����Mon�0{s���-���Or��h�X����:������r��N�_�
F�sTA�9^%���f�	�슌���zeBu����������{�K���oԉ�B��=��H�.O1F��`��Vj��~G��T_OQ����/�[(�NVp�b���+�MO�w�/<�Yj��C��Z�����b��ϓ��n�.r�"��"�_�$�IJb[����߅�����Ӑ(\��9�vs��P=����oԅ��F�B�kK�n��L�P]Q����>�}��R7�
JK �x��?=%/��V9p�'�q7z�ɉ D��Wo�{���B�}�6!1�B����)��|���)������mm7��4�Oy���5�T7��`?��8z�<T.^�(�}`>�m�sm�.^�"���_�!��gzĚo`b��־_��Z�������c����Vy�-)kG0�x��,��fa�#��	�iߕwB5~���^�Q��-�8����s��P���S�"��c���5���Nc˗��6���q�}�����pl����9�i�����n�����h�b�2~��'u�Lt���@�h��q��06��Y�H��R�zg&�*����)��1��)���	��o�OIVqfLN�%���v͛�{�g�����i>~���"�{��彩A�נB3��5���k?��sO����f �L�����I�����kP��U���������U� �Ag F��C�k�]���M��������s?�kfr@�:3_L��W�'�q�B���`T�@gg�6ɕ�J���G�D��3I�-^I}}�?�����
��jL�Ŀ|��#ÒjR�i��؜a����z����/7�gU�6��s�,�s*Y��Y�<��:E��W��P���{�����賓�����߬�!p�C$Q�nN�W�j��Y����aGʫ�ˣw����{��FMvq����Xx�E;!G�^A9�p�<�_�mp0�������''�B��|��!R�eN���}u��_	2�Z�p7Qx:1^t������f�&A���,q�ש4ҹta�%����p:����߮��<�
qz����bu퍊�D������Qξ���݇�޼��*��K����#��:$�O~{�ܽ�@��!�ԏ8hC�������{F��L���Ui��k6�rZ�7BЉOc˶|=e]��Cc�6/�D�H��{��s��S�vΏ��~*ė�*�����.����aA ��C|\��Q1|��9K�e
ܙ[�2<-[O������=�BK�����^*,g�;��;�`�����T��cK�<�Q���D1��t'vxH�߯��j6Zhw�`�6�-��P(���K��\?�.�����{�K��4<�Ć�,36�}6�����2'���y����������|q�}�&�ϼ�ӦW��Ry��lB���)�	��p�4I��/�c��g�M.���&k�(�?(N����isy���Ə"Zn!��{���:��Ӹ�����yj�P]`]r��O����$^B��+�A�C�,�iѨ�o�y9�$5L��#�	���zc���_��`�����_�ec��W/��1�`�>����$�`������:�
O^�SG���������f��L_�����f�4��H%v����/����D�|�F��k�89S��N�1��]5��:m��!w~6�_ ���q���2�MW]M9LxAQK���l�0G�J7Y�I�~]=��CJ���p�������Rm�D'YG��q�YT������6'7�!��f�Kh_T��]M��|{�o8����EMI
=�����_����_�4~?�@y�%lowp�c޸��S�F;���=�g���z����m�����w_k�jre �rӆ�̷KX�.�Mod�s�r'�� %ѻNb^���0\Z�.p������en�=AnR�lC<	߶���x��LJKο*!� 1#�U��M�cHW�9q~��qΔ����Զ͡��L�󝕄7U�'2N������Iݺ�"B��(�Hcؐ�cI�}�R\�C���f�{��t���
\�?��ü��;��P_��QL��X�{�ɵ��j�i D��,�[�/d��hO��9(���؟}(Â�?���uʸh����N�r��a�����'�����sE�ox�:�[��5��Kr���i;��;��;�)��w��G��	�~U{��9?�Sx��v-Ƿ*�p�+ �0!�1��묐?������]��ݿ�xl���G�|��bhl���Im��� :,�q���$���_�o�
��4ϝ;�,�9�O�0�JjN</|�^ۄ�\.��:�ȥY�B��h�L{�����1xE\.ؠ��k,c^�������V�7�^o�/���$�{��}�sR?�h��*�����Y�<��\��d�5֗����7S�>�ct������m#��W'P�p�����z���TI�"~$�C��~�3>|t"�6Y=U�nʈ�c�`�h����@j_��,���`\���X� ����c��qζ���'Z���6�A����d�6�o�=˶����&Pz�,Y�⟠�����P���Sh%*ɥ�Kr��[�xب,�J*̚�����������9h������v#�<�%B@�{��鹶	%�?yT4!%E���T�h�V� M�J8�>һs;3��I	י��鱵�t�]���ӿ�%��cup}}��Νݩ��_|�!w�����"sߌ�{����'t�8=�;�a����h@�)bzi��u5���J/yT��C��A��8�!G�Z&�*��<���7�Hdй���i������O�l�����'�ۯ���}�;y�Vi�M�b��fT@Eo�Mz�+�d]�v��d'��<��|�&�����W�v��W�Q�TU�{=W��<��ɦ͚9A"�X >����neg}_�{Z�]�'��e�0�#�^�r�#:>TS�co<(Uy�QP5�c;eX��,�B����=Ē��0	��P���9��Sd��_Zڨ(\�W~HR������K=�CRW'9g�(;ز�5���^*�[X�*h��Ə���lm$܍��ƅ����w��8��q*?I�bf#��
R6����ŕVT�XW>Oq5^I~=FA�v���CGnj�,��[���-���8
W�a^�F}/��z�MT�d��㕸�Z����OD�3����K�LF,N�9�
(t�o�'���Maˇ��-n�D�	�k�.�G�Ug_m`/>��v�)I:�$E�Qfއ;͆3�10ɝv���NZ&ݬb�QQ�i��i�d�S�{�	��&
'���ړX���@�J��U6��u:!�VYy1�����
���֥�q��|���o7�.�R���㶍�����p�T�St��Cn.����ȇ6���Ʉ����\��WJ� ��^�*)��e�����jGЕ�@��G�3N��{"��ݸ��ݟko>��|%�jw\��a26���l�7�s�J�6�]U(6Yi�:zݐ��/[ƺ�V��m��$�_P�NR�+���1$����~��8K}@��(���L�=�:Ÿ�FE��o��:��u��WD�B\�I�/1p�P��ipSnu��u#����Z�d�Fvj���ŵY�:�N�y�uG��|�j��=B>����$�mk��D��V�� ��[���4�;��'�h����#�� x����.̼��K�]U@#����vR*��.""R�RT�H]69%�5���$y`ʯ�����G%���^�/�7��rȰ��q҇�;99�:�^�e
�<{�ӱ5=��|T�%�p�`F*�ϩ��5�_�ܴu���!K�x��N�����L�Az�f	�n������_��o<d�&��[�y-�455˥qцN��>=��J&?�=���*>���+/+����-�3c��&�֪����s��E�v��l?3�k�PH׸o������(��c������z�C�$1ϩ�|�����2һ׼��{�4X�cu�A�ʜ�[v�:黎�mVn(��u40������H�uu�)㹄�� ��}.s�j�L���J-v{���ч����:y��os��-R��>ny�v͟>�*�U�ua�6G'7lYg���N��hP�]H�uU�v3�_	?���~L�k-zeU�A��ӽD�;3��"���	�*�	P\���x�pQ��f=��I=�mY����$qo��Ռ�̀��Y�n<���z�sdt"��dUԦbo��N�v�	^���&^o*6�ލ1�^�-����m_�����q�%-vzj?���j��ێ��IM13�_�u���s�-|uyhS������������F{8���Ƥ<�������=�?cވ>��yû�;m`m�u�qi�/���#Aq��kV����j��g\��7�ϱ��'2,GQ[gm����u�֓��2��x3�x2�ʆ���-�7n��AJ�%n�Qr&�ۑ������}/��Ctr<���K���/=E�V���?o�<�u���V���O�I����w�����E��ͼ���̕��=�� rvlل���蜦{6
�*_���]��ݳ�ؠ����I̸�����m$\8�~���&��e�Q�r�N�DҞp�-.u(�M�n��I�	��ڢ��`�ݜ�y�l$m��-�3�!�7ؿM�B�|vݎ��faeL����w/6���pr2.e7�۵������h쉼&sV5YH�b���X���K��#A������+b���;�(��!����n��Ι��:�7��&(�վ����%��îD����t��b�0)�t!�&mllB�k�g-����	�h;ym"=Τc}���{���bC��کjj�F:Ž�A�/��]b��Z�_պ족��D!'�s�U�L6�D��Pu���C��T
��d�K�/���:��������DH� ���5i't�f�4�
j�_�8_�L�9��Dr����L�b�~�'�z�)
���X�ʪ|���^�K����ָ52*��)	���0RڄN�ٻ
b�϶-��y����:���+N09m׌29�Pc����D���H�Wzhg�Wz�_�3�d%w���Ҫ!5��W���o����T�.�g�jRn[�PE�.t����iY���K^j�Ƅ7����s��� |岃��MTM��N�r\RU,�Bq
��IZ\����1ڪZ9.7J�R�J=�O>����這�C�4 �1���	�	�������:�Ie� �#�%�s�b�??�D(��h݌u�5(p��}���OYaQ��)
\5�'�0=�kd�1a:ame%.7��1�V(��Ԅ��P��j/���0eL��s$�Q�'x�@�|&-N������E�?ST� K�BKo��_��Q��ڐ����P����٭&A����{|(����5�m|�j6�'`X#�����>%V�CR��'�;��fAg@�p��t��ri�
�ͮ�^~���������IҒ���ȕzK�L@g�u��&;}���).|�ϑ�	%eeΨ�O��:;n���?%�2���,��&�m�)�7��R���D��"�}�4�QH/�"�p��+�x��6���}.��
&ٳ�������7L��Պq��i���˜@��$�g_�����L�M[GOq�	m�{����,4s���*Kb�o��/�(%�/-o����C/6�����ͪl��*�@7��dt���(���V��S�a�G^�Hlm.�Snm_������O 8f���[�����:ۿ��S��|��궷�b?D5��:�[�+�(���-��P�C���U��i��恱��E�~���Kl�)h���Ռ	��q��s�%?��R�2F�("�X�$����+�m�	 �+���L<:��uks}�xK���8�3���e/��ۅ|@WkS�i��Xp2$5[O+�����g�U{e�2��?���&3��)�I�h�du��]E^��'yau#��ln��he\S�#��<Ċf���7����'gʇuꆩ�;�57X�c��zM�,����:���V�S/ֆ��u�+Æ:���`�s̑=w�f¹�b 
���{�k�AH���	�4Y	
	�f_����<�vUa��'�����`
ϟ�O"�����Q0�v�6�� �8 �����u��*�!��ԝGQ�D�������.��Vsf���x�+,c����L�m�`��]Xm�]~���<��ْlP�S���T����EM(�j%r��9]Brr����/�#~9�{D8��U��0�*��l ���������I�JA�A.�YNql-�ې�������??\��i%pRr�W����"��PS�10�,9U�2�3�Z8���F���#,\�||ƼǾD.��N�ۃ��
>�ɹJ�J�pZ<\���(:�x�ȍ4�6�W���u4#^N�+2��.0�����\�-��+�l<E���$���c�ȇO|M��;�[RTD��\�ͽ��)�$
���t���O�K�c�Vs(���!���7π��7x���{��onڔ��46<��T]w¹��eEd�x���9Ӆ ��� ��yⓟ�����X����K^�ڼ�_���`q~x�r H���0�[���2�n*�|Մ�e�8c� Gm�Q��|ǃ&��Vd��w싱r��3>Q���}����͉<��9J��d?J�̛�A�,�ϔ/�����1�Ӛ.$#3s�'Y!�)�ZFb��2g���u�pa��ӛ������EW9��.�����.��v�e��K`�y2��}}}5�����T��7�W�HQ��j��@�3‧����i��� ����
~�����:��8���x�����9.VS<�~&|j����f��.�ȭ�L#޳�����$�ʮ�K�H� R��p ��we����Z����Rkgj6��O��~;��s$��,J�h����8J&���5滨��Y�§����]��Y�1�1�3����p鯿�Zq���KIu��^q��S��&�%�nLHH��>�?�ArQ�!R57�Q2���M��Pu��w='��x겇 ��a�������`��6� ��7d�ڄ���!��aZ�)u��jA�=��$$�'&�����@�&2mK��h�0��P��Hm��[�H9쵃��N�;e�ϡ����7k��`��!�r�w�D`�S�S��Ԟ�������a�d]����eLXYp��D��P����4L_�
 <÷:MJ��\v�nqE��1�Ǎ�ޒ�hfWb�	K䧝���t9�ʏnen�)��L�R' ��;����;�]Cè9���H��SKk9B�k��ݺ��|c쉰O�b,�ߝ��8�z�2����+�I�U{��M��\���)/S�ou6mU��:���¼�a��n-pR?�Sy�
GJ�Ebd��ZA��&R,�������Q��ĵ�/�
R�s����+ks)��/���:�?�Ҭ:^x3�S�<o�A�C��2��������{V�{�M-��4[����u_L9�qq7Ƒ3|�'m�`�2�}]賓%~�Xru	��>�9%�y* )A���������ǐ�1���]#)tk���>CU}���~�Q�x����b�5����2����3��o��5���J���g���ůt1Rt�,�l�1gᙳp��:u��?�)�[w e7�W����hjjB:(/�Q\���� 57�KjP�?�yb$��ai\q�r���̝(�<���� ������#Z�e���Mf�Oc�@���<��� ��ϕف�ԏ�l�R�(;?��k�۶�Q��!�b,'N��^�|m�?��S6���T�������b���0U'#�� �#�no����_�G��iUM�Zm��ˋ�9���VC��4u���i����lQב�����L^�Sg�k�V����լ,��m����E<p�E��e_ӺT:?=P��~m_B�L��W9�<is�+U�Z�<v�L��dʰӞ�q�c"���Zw��5P�w=�z����:�����w7	hF���~<D`�dChh�yc�S�4�N�(�u����,&��{�v��Ё��'�n�esi�8���� ��Q�|ß3q��$���a��B4�	 HG��O���ku��:^j��K�,��i���m�����AZ�����W�1�4�/e���6��S�|��}A*�6��ތMq�B�K�ē����z:>�l�d�"�zV幚T
�e1R��������l��S.���\ް(Q��k��X^^~=J����`�M���e�L�9���7�4�<�#G^[�Tm���y�w�K�0Ĭ!�Mԏ�C��t�:��~&����F���kN�W��,�{j�X�Bvz�=nO�^l�2O/���.��t9
�۲D>�9>�]�����hsH���%v��V�݌��-c�?h�}��h�
�B[��<�������c�AcA÷-jek��"�p=�A������64����V��|2s�A�s.�旑E��js붖nK��f��?�=Vȉ�C���)ᴸb:��J(�W�9��|Hh���4�!%�p��ʰ�B#-B*5����=�_�{qq��.{�H�����X�������/���5��%�������K�5֗��~H�խ�yl�-�3��>�a�H抃�C_O�~��ˠ��arP2A
3�V���@���&���:�K�x�����E_�_L�a�zU`�_F��+���8����k��5^�:���($�N]&����SI��� U�j�±�k��h��J!�66�Ї��M�	�8�} �O��ϟ���kg�i  0�_��n���l�˰�����k)۫̄�m��?���.�ޅ>s�a�E�M�co���**^3}B;�\�G
|~uZZZ���˛ߨ��͞�=�[��h�K*�N�qb~�����@Tᦣ���
�W�e#i�ND=��\c��GK��7�<ǚcΙzx3��'�hqY�A������Z\铓v'C\��3���9՝��%E�3��i��Z3[�#��-�;��D�&�|___,a1b�DB��\��u�~��T��d23E����9	Kn��c��%�N�n/��VU��k�Y�k��(Ґ`�%U,��)�鵅c���=��R�P �G4�;�۽�+�Y��[��~u���Ի�\;]��]��v��U%14����Ǩ�y��	b�뭭�ϖ2V�vd(�>2���.¸ۿ�J��UZ�ײ�@����C��)~��{.��g׽���sT�����UU0o�?��8�_�Z����UnQ�LNN�MǧO;&K&��/h�YWV6������E��Y��G�e�B$���zn���K���l�<o�CF�P;1�U����yK"���<�,�<Fd-E4�i� ��Y�j�� \ԏ>���ٱ��x��u{{��~��B&�{hԙJ��ȕ�ohU}� D��?t9o�Q6�rii>��r���/�qg��v�Ѝ5�������U$�b�Kf�|�(�x%���w�>66
�?��/�"�v�yϯ��de��2�е%��@���qr���$F5�1	z1[����e�]]���ʪ�����֜ԏ8�(��~� ���sysK����&SJ[�SYvv���]�x���s(�U�����?����n�Q��by�>5'�+��?aaa��9P���Z[[�R�8���V�6��CR$�_��tEKQ�S���`��e��A���s� 3���c��|@�/�QD7{�ױ�7�eL�ϯ�����E�{���`����ٙ�4��,�m�k+�}ܧƤ������dFƟ�����uy�min�SYd���4�͝��;�\�#�@9��W{�:`�zx�Wo1��վ{��Nx�M`K��0��z�uȚb��~;U�:��G����y�>�y�A�8P���ۋ�l��6Ŝ��G�� EEEe(̡��Qu��畼?ޕFu5�.Cm$f@KEb]��I��nC��/I�]���ᜉ�	��^��111`��ri �H7~�d���KY�:%������7IY��ĵ�$���9�Ž]Q
�Lz@��y��R���
��w�WDcZ�K�~kk��sR���T��(��2��WVZ�U�p�ޗ�0O�R����YJ�h@���oj���WR���YY�����)0���ͥw���S��a�sW��(�=Ĝĺ�+��:;9b���MV���瀨�)��������u�I8�I�s�֠4�ځ]����xJ��skj����0���Z�^@�o��;�"pl02x�-�gve-88gZ�f�~����/2�ɉ�\NLLLPH�Z���.6��i�M zK<-�:����s������Z����=�7R<F��A,���IO��a"CjL"��E�R)p�����#p�YB�j�}��{�h���!�G /X؈KU��vB���Av�9W�g��uujri4�����^GaH}x�&�����Ǐ�}�� ��G�C�A�xΪ���ru[U�l��'[3.�>]7\�Ǔ����u�>��������`��T������|�9	�{z��M'�N��\N�|E����%�1�'�)��f��/�Qx�tϔ`R���MĊ��w�~Lm�f�+5��CĊ�l��*�mi�S�e�I*X���r�8k}Y����p�p5��sݦ�O���M�%���|��+�}}�<���X��g�uPH�6�'�أ����g�w���y���o�Wh� �����|^�6�¡�������k�4'�$"�b�X���<������9�g�����]Z�=0�lR�^+A(%�,�]��_j�_�{�Ճ�j��~>>�h������*����AyF�ܺ�Z��u&���SQq�|�r���3$5���Y���3��n��� �������6b# ��1�G|w���� U��= دP�;��s�.�L��.��M���ʻo�(�Cg�� �T��L�yS��@�|�'�~7��`��Aon`��wȐ	@wM���ߒ0(s<Iذc$���.*ػ��Ƥ ������%�2�F��`�-	�A�~��j��3�������%u��[	H'��s�a�ڵ�f�9�,G��i����i����>�ַwpЄ2����X�a

B�댸Ujik�Ր�7p!� ���m�:?]�]
<\[k�ض[�����O���v�f�jVu�a��G��� �p[@Ʀ��aH�'�#�}H	*l��?�*�+RZ��9���-������ʱ��?o����YS�u @��z��j������A�h	:��*�[3�o7�(c\L�59��>|XV�A;���2p��2a���U�M���A�o&o<�.�pd?\��n��ek52��1B0��)��p������q�B�;�Vj�ف,��fe(P'Ooog��#��?W��ϟW�8�v�ߴ4⍃���(�|E��[���ְ N2���(>�?&a�f��Dt����Ç��zMJ��	#��oIpqsG��W���&cX�~��գĞ%�E�{
�A"zx|&��������cccP�_���]@k�1som���Vr��x㦋���kk�Nõƀ��H�f���#�`᪕!?P���%p�����8+�:�ekvv�h�Le��^�g�k��P.2�ձM���90�wΰ�"�Y"t\�Fy�w�����@�w��̴�p���h�^	�(�� :���f�&&�&������naq�X��N��/n:
.:
�5Ӟ-EZ��و���4_"�8Z��#�)����+��g��@�C�l]Z*<( �2F��e�/�{�N���q�*����7p��<m�t�D!�o54���k�wq!��YU=謭��Z $±c� �3�n���~p �M�:?�z�bY*�Mcf����rn�h	{���%j���89wv��5xh��W����y���������q��Ou�5g��!ii(��S���3��/�9�5�J#�/⣍��!�31u���>r�C��ݣ?yR�=�<��P�R���\�w) ��^(p�����2���9~���t�.Dc	^�щ!�=zgz0�8\3�v�Y��u*�����9A�}39�8�ר�Em�j�nnnNMOR��Y���mh�[U%���M[����kG��n�9hkU��`q^YI�#�%>�S�ҫ��Zr���
����g�D	�|���g�޷o�ǟ_��KKY����_�4�sRG��ۻ�����ghz9'?_�['����ܝ==Y�-��[8d���Y�?�X��Ç=㗑?����S�;~0���7��,�>����أ�:�L�2B=I*����ZO��������U��oy�2�Uɮ.�)�$��Ii��CKa��� �Ǿ����
rgsw)�"{:Y^]�s*ZL\\�9Ǐ+�І��6� ��0���G�}a�c+��˶���SSS�SCP��"`
v���ay<��!K$����fp��&JVb:ğ�B�B���Ag>)L�w���� �������'/�xH�4��Y(��便Bl�TK`�h��:��*��X�i�|FF3p�������q�|����*-��b�J��|} 'Q��號bd<�o��ȷ����]����;Q������i�!&h/:��Ǭ�J��ݞ&���:�Os��f�?!!��DDr�I0X7�$B<c���n鹼��%E��Q�AL�2��*�S��zϗ#�����:B�7��>Wɤ?u�s�U�e�7�����F��o�^^^^��yS�=}��ȋ��xZ������� ق��*I��yH`.=B���'�,�r���D{����ث��Ej|KK6}����Ȏ"몠X����0U�$ǌ��޶7��+�"&ְ<'#����K�������Ի�C����)�*t�D �h���9PM�ܪ3�va(���f*݃��7E���t�Vx6<��������;���j'�;�p8�m����ϐ�JSGL�򅱒t��U��NN1���4Kl�q����$I?HUnG$�Jؚ�x@�e��^�`��u��=`,�7�\��6?[��!�E������{���t��4`X ���!�<�NS�~uV��+��W��d��Q�̭�P��/����� kD�%?��ohٶ%k��F�$��kf������ཽ�s�TWn�E�A!!��o7��yf	��Ş�k���v��҄��3~>�Ga�,�DaD�U2q�j�b>���Ô�\��<�Natx�J�k�"�]]]�..��o�����":���~t��ڒHJ\!?91��*9tgUV�ࡀ�FE9��(����(���5��������H4`G�`�����C�[�h���X���a:EV��ϭ�-0��{����'��v�:�H��hiI�pcHJ��Ȗ�N.��Y�����Mԏ�O�q�n)*�_u���9��� ��0:�IM̌�#��F�����L�jռ�G�s��aSH����4�ݍi���@���o�.L=�����^ r4�����έ8,Ouӎj h�g��߿�]�a���rre)G{;;u&y�g�7�=��|
�n�ۛ�h��''�����V+I����?[�����$����Yp���Х&}q��;F�y* I0ߏ���d���Ǵw�.��c=�A����E��[�q=]CM�1K�A�߰����ʃ���Н׾�<]�:*�����a���J �	��'����y������9<(��FJ�6wK�����F?��]�S�-� �7X� 3F!�i��L�ݹt	#��w�''=PU����B��EK++�puH6PC�xL�km{\z�c��]/�#�]DY<3\g��gF���#���u����3?>�sEuZ����s��[[�E���Ԋ��0z�m�P��P��}��J������eX�������bԷY����,c���"Q}a	z�҈�1kB� r��M������A��� �6D Z��\�H�Uշ�04��?�ԦV�81�ʖ1of*�7S�M
t�fw.��_��)�el�mM������,�($j�	��Qƞ��ݭ��a��K��1A����kʘ�Z#�v�cd�WQ��O�"D���,
ʰ�BK(��&^m�f(�����v�c�/0v�����ۺ���g�ߑ̺�����|�7�09��]!��LPkOd�#j��D��	��A�*�/�9L�ǙX���A��/�3��)':�"g53�KKˏ-��F*�d����Ff��ؚkT�&��ֻh�D>��7����>��8���ȣ5[k�hyճ���6E� ��>�6(��ԑ犿�e��=5�3�9�����f���X�]IA���C0����_�@�A\����e-z	����/Q��� �|$����:��+W�i\ �uMok��k&E�=�7Q��ϋ5���`��i����~.��&��f�w����>�\E�Oz�z;�.�e&��V�j����oq��G5ѰWkz�cx��|v.�>��H��[�2O�ݽXk`-�*�� �֝�Nr1��!�'��?7(s�Gqk\��Is��CL{�1�x�a�Z���ZP�a�w�/���h�q��m��}qt���e�������j�`�p���+J�fDVm����p�n�	(�0�����ç��.b,ht.����7UPb��[�{Ṣ��䄺@�N}�-EJ������`�h�6�K�v�DV~~7��[�	@�ܤ !�+x���]�w���u�&K��@����ۅ��ۻ��8�r�@_��b�ȇ�	�i��nG(_mV�p@�߃��8���C��]Bc֔��%p��E�H��t%�_�e�AO��o�{N��P1�E/6iq�ߒȇ"�*��g��7&slQ}��R�#�� �E<�GHJ*�-�G�W�R��^G(?�C5~]CC_��1������+o.��u��6��ǀ�K{�����41�����:K$�X��M�� ����t������5&��d D�)��CA�P�����Ѧ1��8W����i�hU���ap�-�������|��]�or삂���W���v@��ywJ2�|�W�, �6����l������C�@h����c�n�����}���@��j�,����N'�)���{����Ԗ�Vj��
��<t$�Y��_��x������B���H@h���MQ����~���!�;��O�m���%��<_X�9�"�!F�zD?6��u4��S`�$F��F���(�fc����4�d�����h+�P�'EQ >���#�� ��A�P?�I��eU c�{.�.����#������B�^kq鴙��V�JKK[[.�B����S�l_3w{�1�ԉ�J!�P�t{�v_���0`ǨW=x{ep�1z�y�T������n?�����&h[�pXt] �h�I�$S�pKKK)<(['�{kO���/�)굹�-���";���d���2�~��~(#�3 �zP'�	h7�\\ 9�����ugT� >��Y̨�3��`҆lz��*2{
F�dU�ߛ��	�.���l�u��r��b��
@#��
����D�)����\k�H
��MF����u}hEjf�&�v�[�A�� ����E���0�=/'G�y��|��P�秈F���+M��s����ǏOe>��g�F{�� �e�F��(1��B-�|�\��!������!MU9��{{����������l�\7�|�+gaD�2ꐉT
�¥li'�<�2�6*�e	�-1��F�7N�ҁ ��qvg.B��J�aI�a%ǼX�1x;�m�7MF	�X$&ϝ;0-��6}p���!��X�q�-c�]/�؛���53��w�Y�T�h��s�\����U]@�:+���j�T�<�QM���9�����
��)m�j� ?�z�w	qR/�&��^���,��_�T��S�4�
�F!( ��6�9� �ޠ�@?��|2���P}��J$, �;/,�uV5��\�0�?qҭr�7�l�Rs�Jhf���n.U,���)����Iw������*M��������+uۛUc��
�����#�����_��Ä��Q����~���7*��p��%��7M��b���^�rJ..����H�������(�"�����ꘑ,-� p�U�f+�i2(WUs�����1f_��yxyM��&��Nr`:A$-��4j��a�Kp#�Z� n|e%p� x��8�{�s9jm*�s�!���7���y�H�q��HzUj��`�az�+�C���ZÄT6f�Ez�,��|�ׯfb1��.
C##/���@<�x�`Y�#µ$�$�_adc����ը�ӧ����j��lS�t�V��#�}46��ꦁ���3����(��E4���glчQ��%��IU!4mE�cS�[b�B;������%)�$wb���m.dT練IU�F��4�C�;Qxٞ��lm�(d���+��W,٣8�3�V-c�d@NqVT�^I��=��+F�x�|XlH�|�T�m���Kx���1��?�.xr��]@�*�$ IV{�r�3:�k�ϸ�~7�\5`!�_ -�z`����������S�&���O�F���+���c?wa\�m3!R�/����
jH6�ps�oxbD̀|��UUU��fz(F"#n��r/�N��!Cfac��>+����L�aG���/��U�a���Ч17r���(� �s�ږ?6h%���1)�?�1�U�WG)	+��+�����G�2��2q�[����m��
�1�q췿KQ�Ԍ#�s��~�� :� I�=�7���Y��2�7�.�9����d��p�7R��М�F��y��@�o\"�r7&�쓤��e9
���}������P�Wi��%����4�f�b;Hߵ	y�3� �Fh��GtF,����W�(v0��޹|:�z�}������188853��C�	!3��I��9@�y��;��IG�ST���[�����`%y�/Z,hZ��NM� ��~ q�s�u=�+�l��5 ?�9iiW���#hB���?tvuM���VQ��,<,<|jidBW�^�+�k���x%�*���Eg�3yB��9�]V��:+���䐆P�(L�ʻ�����ZTPD�i�fl����O��h\�pL ����{��ҁ�{�o�����e�Y;�3��L!�G���&_2�燆T�ˬ�`oN^jΡ�T��x��"�E��Ў�D@;��^���^�RK�TMD��àD��1o\		�b��ξ���h;���r^�Z	�D�A���I�L|}�
!nA���\��!ڛ�����[4��W� �K����A�L�n����m��<,]]]�#w�;;:,�1�@k�x��F��~�nD�Х�߷$�T�B��<ף��0@��k�g�*��+���M83��XF� �e#޸�w����JlZ靆�Zs�h<۹�Ś�R��HIؚ�(�5aɼ���%cE���!�U�%Y��h�{�p)[��B@ݰ�7�����jHH�S�B�c�%�4Hj��LN��Tf�7Œ���(=>�]b�c���zF�ӈ�E�3�Ä{*ʈ2t�-������H�4�z���Z�.W���ʰ�-Jo����&3�U�}�����%(�ă-�"��i�*́�\0�T����=EO_����8mF+&&��Ƽy-�|��.דQ�>tB�s"p����@4� �� ��c}�|zk}.��7~�r��VRQ��X]�����<h��Rmcn	���KK�K�*�1-c?7{0�*D�x�ҥ����]K�H��@7�@H$�/\G�	�ߛ������堼�?[@
?;$�Kz'�I�bCĪ���_�ҹ		����?@�9��q�D�B��Zً^bI��C��Z�����D�:NNX����y���0/fg���Q�����<��$2K6�y�Ə���N�����<~�?ʼ]���:A��mCx�|C(�S�/˙2�V	E��:�ќ�Z�L'@P:�u���)(�k���x� ��cn��!��&�UU����׫�S�R�/�{����'�k�Y� I�֙)ņ(0a8A�JH���a**#�ZY����$J���IEa�"Zx��XE[;���k� � �*���}3GV]����<�1��04[1J)�Oef��,*���EzffD�~jCb
�kN��/����u��� 4A&=|M"�!reW��59�a�:��hE[�3q�f�Yp��Q����������^SU�i���
m��b�DY	�2��8裷1h�֮�������H}���gO0�*�ٳ�PSR�;:���̱}��}��� ��`�;�\ �����wq��/ ,��^WW6PA-�,��O׉�R	;%�iv�
�4ik2a�<��k_x�I���EX�z���:z���+�ߒ��Ё��F�C�m�3jM7>uz�|������������|*�!�=0Ѩ�b�NOF�Fx�)�ٖs��[?T�U� x��Mc�/g\�'!�WOq鶕Z<�ScBL��
��vu4i��u��1�:Z��#�n]�e.��QҠs\��Sªe�0����G9`�3^đ�:���e;����%�To��c%�2�QR(�Ch�"�<��)�H�2��IHu��d�L�#!eH�B2d.Q���C��߿ǽO�:gkx׻�^{o��n~>��d ʮ��u�� �&�����`0����u6__�=B1�>��2\k����v�����p�@D:Gj�oŮ�گ��|(2�2��7߾=����'�"�e�A�I�K��@�Y�����`�qf�YY�Cʱ��i\~��&�_1o��Q�t������\��_����{䨪�<�QDx���ȿNnT ±L����6��?ξ��k�(:��^�j�Z�Z��H�~�9	�����9�~O $���}���š|7X��Fz����>'�yc�b>�)[�����]w����pt~�/��?�E��|��n]�n~QӏO&
�(w�C0<,Xq������\�"tk^9Gc��e]��{��B�/1�va���x�oh;�7L���ϯ�a�{qm=�3�Pm��`g�|� �2�8:�y��O��1��E�8�2���_s.����1�\ �~{�{������WRi-��;�O�� �*=,C/Ni;��j�y'��߽Gߜ�T�4X�� ����\��~����?ο�~~T�oq�o Xஞ?Z������l�-�]��Mk���6\�Yl���-�/`��¡��v"��z/�+���1^�u�!�r��	��3��(Zs��,�0�rL�=��-�j{��u6��y6Pd���f����$�g�C��J��>�+~�C~zE�i�w?�~��º�#G9o
(m	:�2=��ȥ��3����Ą��rS8��Eb�R�6��M/�_�_��і�Q���x�Q@�qq*+W��vÎ�1n�;#w�Uε���������r�^j��a�!�5��=З�dR�ҥQ��ĝ`��A
(���� ��I֊�.n�ԋt+r����[�XPH��+w� @��#~oU9�	���4���r=<,,�I�p����M��׿[_w��n�=�z��b��#u��#�m�_��f+/�	{.���ayG`mO�����&�e���U�M]����GTT0(m2���jd�H�,m=�R8��0�� ��|�9/�r�i��v��{��&#���a�^����c��=Ƶ�cƖ�%Me�l ��!�3e��5��SЊ���T�Q�\ �����Q��!��bCu��̻��¹�/l�����:���he2�2�x�7+�GQ,�����\��|ZȔ���_`���7���9�+�:r����ߖ�"�]����Q�yY����q##�OȽI+u�v~�6����G [�^x���X��p��-��m��{���z{<8�p��sO� ����������p����B1d, ��0�*@��ó_��f�@��4?�V�qz%IU͍���j�`oi94 &���D����RG��|1�X��.*�@/a1�m�D���eהk�$覴)����b^)[/�:���n��(�������#���
�Pz�Gutt4��6t��?���yS��&��2F���� ���ϟ?ҹI2��U���C*1�&?�/?��B_-n}t�-y9�,N+m���:Y��Zt�`��&x_Z�������P�U><\)���*������9B6<i���^XT��It�M�����`��G�_��{������s�]ʡ`��X�ƃ�ې��~6�6U���������v�����|b�tXm���h�6Mk뎴7i�e�1�_'s���������
�>^v!ݼ�av�!D�
H&�:?S��Ӄ4�OB�K��z�'H��]{����fF��+�Ph�z_�C�d]n2A�__��W�j{�h��8�"��r�o�����}A��3��Q��m�6l��7 �p�/��'�]�g�a�em���n���Y��{l��yI�0o�}��̸��&���o�kd�U�`����E�wYVF��b�g���싘��j�*߾�1�KdR�D0���e�_����:t��r*_��Ҽt���ކ,��o743���Դ�W����P��@���W��� L<��G�.�&'���	"�p(�?J0���@t�	d,�?��+Cr"|�a$�BƤ�8��ɚ�ˆ���p�ݗw��Y4jjk?{�����i�v��ޟ�x7y<�,�E�m�Y�O�6,�/y#˕=�Z���n�|�BB����.����ĉ�0Pp�-`6�:KB��7:�~<��ڟjQ������"}!�ئ�7T�5Y"���
	�M9�M扺 ^լaa�T��o8��M/،T��w���놆2�y'䖵��c&�,N&^��-W��M��*�q�+m|l`�u�ǏG�u��J066�����%d<��2;����nA�ϐ��ٔ�LF��#�ƪ�� ;��@,ܻ3�
��5x��K�`*�m�����4���32R�&|� W�t���܄D�6�g		���Y��#�4#�:]����lxvGv�����*��Pů�eN]j��/�~B�u(�����9�D�l6�khkG��jI[��x�L��f`]7�I.�����p~o�������6-��X>k�Һz/�8�YE�ӧ��c��4�͔2�<��]���ǚ�����~L4J��
�r�Hw�H���X[��q���T<�ܐ�Pfr|���(���{#cno�s��;&�n�wr�������*�z����N�AѵL;_�8�������Fr&o��Vsf�ǥ��_��ʲ��Ns���*�Bׅ�~]�/�tL�������d։���B�v�7AWrr�w�z�GeUՓ���@�jsv��p������l�H.�9j�j��t�=`����A�w �p�T�u��H6����p|����^z?���O�t�k_�Z*�:9��ɉ��5ww��9�ZL1�J;�
2�����艺o��z(��'_^� �p�4x�*������s~w��F�P��!�d:��G�M�����¯�]w�J��B01�����"1��&$�z�����6(�Ι~�S˛x4�(�������79�̴o��Pr�
��g�{�%�M��rĐ k/E�{�#\ggh�j�g�iQ7.��5��kn缩'@�|llL��`����"�@G�ɜW�Ź2���E&�MK�M��?��:�����A}�'~�;�I`��R������h;��{R���888t�?����^���ɱ�ɾ`�9jjiu���E,�������x|����rSM��Ǜ��k���e'K�P�L��y.�0^�U,P���j�U�����ɜ�Ef�N�v8+���n�[L��)+���p}�js�l�R�����C7zHQUՏS��)�����+B2�i��T$�� �=��UP���*��+
j-�Jz�v)�wl�������b��>�X��׮��ݵt�>�w}�a�9�5�)�1�eÆ}��K+ǆn�q���2��[2�&�#VC|۳�=t�Л���A����2j�j���6ۏ���]#�c�0)V�2|���Fp֔����,?'��ԏ����1ժ�~E5��Ɇ	��?�	4�2����}�`��T�|}}G��'�����(�'{!y���F��Z�j�,X O�O _��Eb���	Vk�D��8َ����1R���bd��e��w�T�ģ`XR������g�T�P�}$fQ��nk�@���j������h�		5�j��#���/�p���M<����Yk�yv��%R�n%�g���U���ޑ�����)��(���2|��]�T���T��ѭ��Ј��\B6䓊t�#1����[9!�c�&Mf���ڴ�IN��-<���t��󜤶J�l�xSW��u��k:t���V��F�K�n#1��߾}���s��#p��t��X�_��ű�~��:K��&.�S[�G�jq	���� p��T�v<������G]��k�l1�63��U�d��6^J�)&��b�הzQ?x�#���ֵ	Z {������3�f���D	II�H.J�K�5�?��*a^L=��!oN#7k	���M �p��,xeޒ�/N_�$�G3���iڴ����WQcc.n����������}�f���@��ޗ�'���{�]@��A��=���˛uɚ8�N�������K��`��|�B?�X,a�׸qe�-}��*��j�����)�	snY ����=�s���W�+�5c�P>4��[ׯ�r�W[]�{�#ŚF�����V,�8�[D*X��9H���ɡ�U�l�:�>���������������g��}ddd������
P���-x'�=	�`�CG���cV#������ݧA�:^ �e��`��K��5d�		)ӯ3<p�S�����g��;LZ��� Y]m6g�w�y��%���nZ�p�YCPx��� �����"��=�@&TƦ��G�eFD�{�y���Zy#���1��n4���=��Ku��F~�OƝ�9W�w��~qJ3-Z�î����/پ|�Y��	�Dq�����[�frVX��5��C�y��O���]����n_��v��]]]5<
&J��B^:���u��Z��$�L���|���{2N	�rh��ƲiP�R|a�"�����@ ��V�]��ȹ��R7:�?�a���ۛd}g|tT	�5��ԏՃ��ѵ�U����V$�g��`���4�
* V�y��3o������q�_B��whA�'<n��Ө��v��K&��#�*H,\M^��F���;{�g�$k��>\
�s㤢5�ߊ�5�{m����>��>�N�Ie9'��&��U)��E���#����3T��o��]Z��o�G��nDMH$.�9�?��i��2��\�p�H� ��y�y�*ס��5<�0�������1.��ц�@D�]�+�����6�����h��x>�F����O@Nl�Ui�4-X��3�^^�]�^GXL:�u���X)�4ɕ4��/|O)�O*H!���k�b��[#=��[H�}����emR~s���N�R���#���='w�.�'��4�w��D�����]"�����"y4>r(�k�����$��E\�		g�j���Y
������B����_��𥿽ie�WXX��yi=jB���Q�@����V	��9�� �l���0������'%���x��#��> ٳ�b�aӏ������u����8�<S-+��j������ey,�y|�k�f�!���\BB���`m���u��c�]- �C�ŧ(/]�x�cﬅ������-JR����a�=֗��j �;���Ѫ��n8�.u��ߥ�8TF�K]]B[��'���V��.���W��z+�}b�����B[���K��ן���KKK#.iij��^Y���P�5��OS�ֳ70��c	����ۮ`ۊ���Aaa��˱����{�V�M�5<s�A�z���_����t�O�������p)��;!<� V�P�<�'^?���%k��ȑ��uN��l	��V3����g�"�H��2Ӧ�6�U��C�?�v)�;�):R{6������X`\�4#���U&���&�8��s7Y��ϒ����Սq Nv�r	UF(�"6���h��>.[|�#��R7�b 0�K�ܼ���|1Xb��$99�y'/9��/xxP�~v���7��ߗ��_�!ر��� �^GȦ�/	�8'F@�7iD��h7����c����F�%V16��D?Ö:�ɇv��}��gz h!YYY�8�xr	��'Q��A0�81
���3�q��ڼ5ܷ^@��%��[�"�(^h �8W߹zI'=��d̩�$H�0����_p�ׯ_0l�7���m"��R��X�7xpX[Z"+��l��p���q����l��H��ƾ�Cy�쀛������27��wCI6��[��b$G;t�uyrŴ���&D��`��CDt��2���DF�_���`t� ��������IwVZ�QQ��u�^��AgXH�蛬�G�D�!w�n��������	��3����}��$���M��}����%��?K�0����w�Un��ԑ�.w�0�~<��̏�4��]	ET��cX���X`cҰ��(qXY9�v��#���g�%?#��� �a �n�÷����XƷ��� ��IE�MHa7����n<$-l�dݯ���/�:���DA���=����g;���Z�u��E&[���V'�8Sm�D˭�؁�`�NuC�������)���y;i��KǛmR(�6.�Z0Ȑ!���Ԕ�\Ν1�inum1b�Н� +w@S���~�`���С�����*f�o�_ ������ݳ�Ȃ9���<u�N�"�X�����'j�l�v� � D�3+��	��+H�(���kK�k'�Q<,�OS�&67FI3FJ��9�b	�|#~�Q���AT��e�B`�׀w��g���!�PH|������L]��뎬>˳v0w���.	���C��� |��0pi�b4\5߹���(hC;�RL�$'��9i���L���L�p�DP� 2�s'HK�gnB��Í㞆,���s�G����YDs�D�v<%Vq��+@;e��G�M鄼��""�\��g�X��=WX���i/^�H	ω�Cx��c�u=�:ܲ��q���h~O��m��XOJ_) r
[8�	ȰZ���_*lNe�jR`u����v���`���k���2Q.Cd01][[��U4S�p���X�h���i�w�$��t��UR�2�yP�#�l�F�r�yv g0��Y�mZ~b��j�����>��lf����F���j�C��2`N�[BU���G��.~�������5�D�E�ߗ�{�Ҭ�GJ���?���2�P��2	��{عO�29��J��K�.���r�+>y�R�&pA��Õ�h���o޼�O��
���ڪ�7m�'�����b5<��Q�}Q##��
��M��
�� E�X	�Nr���̑���&�y $S�����3�}<��˗�%GBw���ɂ!�K�����@���������'���7
�c[ed�pKi�ȏ}�;j���aR~���HC����i�Q4b~b�G�}+q�O��_]�S)�~�Y������֡7ϴb�jj�g���Ǔ��	�V������0� +�.H��s��0��l�J��<�;6Q����%n}L���~Uy��]�Њ�֛b�)>���.�7����V��j��$�22�$&��n��H��8@Ӵ�L]�hUjr��
6ρ/?�t������&�n�5!����m�c��_�׳��v=��߿���"�)���J�5iZlx%=}W�^J!)�
2M$}�M���E�+�����&dd� �0N��|��B��ӳ��,��/��iffV�C�Mț�:��:_�ĉG�E�%͢�C�g��ӗ%fER���p�3��G��Y��%���,�?Sx�"��`�f�փ?����ſM�CDV���`���0'Q�E�cz���㫿��T�hhh��i�.�K*���}M[������o;%����m��pVٸ���Q:70�¼Yl1����� ���g��c V�x��<o̴���i[��2B��C���Ϗz�V�$��OF��e�3�9w<	YS�=�2U����|�lJ=�y*�71�1~��72:��sr������ѩ�1t;��#s>���]�87���oV  w�!�+���(�f���Z�RF9xuﺶ�l^ o<p�ӑ�I`EK�qi��.7�,>E
��I�F!VB��{[��֋vE��d����5��x؁7:�.�x�0P7�Q��˗x�8�Ltٴ]���F�Oj�)E^�/�9׬Y�I���	�_���G���2���`R>~��~���y9��MC�3g���l6/�_�b��mp�	-#��}����OX�RQq�zb���?@��C�-P��4��:������iȬ ����M�r�[��b�-�F>4�%�@��&�v1�犾����Z>*������~�� X��=���)7�v���������n��o+�ș�^�Z_oM=qW���ǉ5�H�Uyt�-�IA�>�>B__�G}LK:5�̹M�! tOO_��ˌ=��eۻ����Eݥ
@��<��5�u��ub-�T	�B����x�=55<&
#�Rd1���
�i��JBN��0`[�͢^J.$]������(xCn��9�:̇�+D>i�ֵ�T)��y�Y{i:�y����ԅA/�V���I�K���d3�]}xs���C)�ׯ�|�soI�o }���� sC�+;�N�B�OO�� #������[@�h4��:����dރ�: }w�|�se �e��zhL���!���X�t�ҥm�� ��Ӭ���jj�D�����\^��Y~���L���Ԁ�H�8��ׄ�6 o�$i��Ջ��q�s����$9N6O���Ҷ�������������<����wG��ځ�� X޽6Z���Gÿ�|!�f�q���]Gbb�y��GU�4���Ŧȏ��wT|���~��� d��D�5A\�g��V�gu�����6��>%%%�E;33�Eܐ��?c��H{j�,�"c��ͧ��{鿅?�,>^KO/��4 ���S�!��].$��}&�KAwvԙF)ρ�K���Z<i��;�k��"4�����Aj9��X���k��sg��[�f�e=�O�EI�x��9#�x��F��۹��S���OLO�nkk��g�/���<�o`�D����Yk`�*⫴pה��~�Xё���ӬC�/�,;u/�� �gΗ������ƅ���%�&��a܄��@��w΁ �޽;\]S3&��x��A������MP+�o���:}�	 ��74�Lc��Ç�{a�sO�����i�����=��-W��t�}�(��!�ce%�37���\�WcX)�/��;26%-�4 >>P �T�rz�������x�!l�����Ss�˚��M_� �Ά0���Ξ?}� ��,6��i���U���NH���(�Wd�n��� �&iZh[��*�V�Ķ��ŋL��hoN�)	&#�2�k'Տ�7-���3K=>&���Ke��v��%�	�K:�[�bKEm�R���M���n�o�=����?>9�J��$�my�������iI�A������}e��
S��R�E�w�� �u����G}F9i�����"F6T��rhh(���wIH�� ����R��b�r�.�>S|��`�%�R(����݃37 �m[P	�ھ}W�'�z����P|{���F�OD�G ِ��HL�E�����p��8�$����Iv�)�3��H�,OǤ2����pIl����"a����C��N`\Dث�}}*`�M����;��׀�������������Íۍ����(I�!.G��hL	�`�QDI�m{G�Z$ԗ����9�ӴӦ>�����a�_k��R�@h`鎌��T�@�"0�������+^�)�潸Q�ބ!<OK_��d�]�O�N/y�h��O�t�O���ˊ}�K���q�΂��,"���=5#��k��U-���N���*GV~/���?s'sM�`ֱ��^���\�깐�׹�x50.�0Q~�3#�&���v�`:h7D@��Ǐ�.Z�$ X�0?�Y6���54.�i���V�^=gI�� �?}��|�x��*�w$&)y����=���###�E���v��<�v��6_E[����P�?AF�ٲ�a ���S��=HMo��E����]�B`A��f��u��=z��s�mii۟�F��T	<��1|���8;�XT�����HC���f�wgg�z�H��7,S�O?�^&�4�ge{�����/y�s��u��i�sg��^�L�#0�C#}�K �c�R~��e�"#�*����[��k�瀯!�R�A��Α�D`¨`C�7/�SE�|��W��(�����{&��<r���R9'}�����2-6�u�2�>\l�K���b#sY�� f�VF#^=o'�'H'�*�9��n�Ց���a�Ϸ?c�O�q��*�#S�������^F}���#h׺����K�g�P&CO�0�:r>�ii1qq%�Zb�����kJ3;uʲЇ|y% pPv<j:��
�f��m�ٗW�#X�a������ů��1m�SX��9̲9�Ep��*�]�:��<�Q'W��=7�pd$���;�DcHKK�	 VU|��sC�,�4T��Ĕy���P�X���f�Lu!���)y!��S��l���O��� �F� �� 	�Ωz8�����Ga��(
H��)��ɉ��4����E��T�Y�p���M�=�஌S�@k�v�'��̮�*�z����\�I�V��{a^��*�j�@qկ�<��U��<7��R��:	��%ȹf�Y����O�JH;p,���[G��r/t�?�Ek�|I	��S��ZSw4��'�{ׁg=��?��J����C��ҀSXO+�k��w��ie������0�u�%����OwW��$�2n�U与�Y�cl��KVU�­�}�����ѪT|�������E�����P�*X�dA�^�禔377ϖ�fX�>�~�L< T	*�!s��VP>.���jJ(��D�h*$ `ٍIj_���3�]��^YWW7w|'��v�B�)͗OF;������t kb�wn 1(-о��j|�����7�ֺ<��F�<�*�dFe2�GC蔊n���o\�(|z���0��L����I��wt�Da(���K���zD�~gC<�e���t�eй��C)%ϔkr;�e��`ֆ�'��O�fFm&E}��/�hg�p���[�<��,�����/$��0�xb����}9g𔨇�b��&�X�kC�r���n}S�ԿDLtai������kj����������RƘ��3�����9���P�}~���uS9Ӝ����h-c�(ط������
d>~���`�u^�6m:}�L�*�Ģ�;��3�����x�᠟��T�=>D_&�����jp�,0b�����ɏW��H$�&�<�/�j�6H?Hes|
qP�eͬsQ<4��9�R��K��;�j�#�����',��ڦO���(�ǎ��6]�k}
����]YYM�U���?6A��р�I��<
�]Fb�,���y�hO�q'����'/n���75����.�b��J�HB�a��8�}ۄFA����w�ϟ���N���9� v�]�1\�X��q�d���o{���|OO�±��S6? XM{��(U�3Ȁzěn÷�|Z� \Tf_��Aa��~��Ã`��Cŧ~���ߓv�2/��K��)�L�{��,!s��Y$�S�	j�1Ϟ�c��5��ꘄ�Ւ�Uߊ% �D�b�H�"}��#��A������� _�w���`ݾ�+�WlV9
#g[�0����O����ir��������s��s�!��0���yE����-C�8 Rn:,:S�
:���ӧO��|�x�1�}Hc�1�.վ �A!!�SChӁ�1��l�`o`0���RWD�ْ�>_,|a�q�=6�,&������D}N�(-qѵtk�|wA�����b��H\���Ш�u�m6��pnb��}�Ԥife�ڽ��G�z��-��t��b���ׯ��Ret$�#0�\�8�1I��z��PaZ�=̡Fό����x�YP@�	*�Z�{���P��|���|�w�ڋ����;�^rs�1/{*fq��u5V�
/b&#�c�=D�>&��2 4��(]p~�+Ȋ���K*k!X�,���A_a#B���޽{��ٽi�o,�Z!�y P�.lV�����d��ƅ����ץK/!��kP�4��-������E{v��$ǭ���t���h��\|��5~v�E�Ԟwj�K��K�����Y�VKHa�
kc�����C��P�/�����s��B�I��M��ÿt�ط*	��s�(���2NY���|r.wg��&Ar���s�IJ:�{���l�z���F�/4��<�y7s���ظ�S�>���TFc���? կ�B+Q
PzCZ$XN+p���_MuZ��`^FNN��Q��b�'��Y�yY��C��\��N�)���>�ym������;�T"ы�K�s��5�5��tp�D�/�X���N�\U���� ��a��@�ކ��[�</�\Tpr�Ԣ٫�F�%)�r" @�&ا@��s��=MMՄ�A�=v�׊���������}�����k�)�i�O�7|rjgq�k��@��R��&oo�̆:�˄�T�7����ƀ��c����]6w��-y���D��=x1|um��P��ġ��xf���	y���3u!���߂�0�z��ΰ��|J�w��4�'�ݕ� ��	��Ί��~2s��lć��
`��ҀI���<�|�_����&���\�|�1�K���)_�hx[��Y�V�*J���>��@��z�Cw[=�F����L��xtߑQ�����߿K s+��c߾��T�(���	n�~d�6��qL̡��x� �p��'�)���+_ZZ�UP��`_�(�$�Ű4��;\��2fyio�}�I	�������c��s�%�>�i޳kh�df�dfEu.8f���57�]G΁���U�1w����y�y�l<S76N,+S�a7ܜ�|h+�9=��x�O�8 FX �
�L��V�b<r�'q��)���>��^�"���� ��8���C'���O�뾸L+���QMh�����'��Sċ9�c1�l /�~����LPLLO@�W�]f�I���t��˗+���r�M3��=Q1l��:l;���` �X�2�A���3�#6��a��T�Wޫए�K�����;��-�o��� Г���p	<s(	UG�=�Ԣ�lܴ|A��u`����Kxf�ˬn)m��'�}��O/ߺm����k\�(�8��14�0`oh^����'��i
�>���z��B���w�p�pN�v�� �m<�>}���ns���#)�X�︊���=W�E�B�qW�Cc���L���N��;��|����lD�ٖ7X{g�	�IO�!1V56&�?��O�1�}������N�$]��r����:2~�������3�z%D?�B^'7:Y�k���� ��'b<��l��S�U#��q����@������EC��!#��C��'ΑU�*��ij�k�4�i=�8���bA��tڿJ�KZ��� ���MSȾ��9�H�RL�b	|����/���ȿf�^zo��]j[_�H�j����½]�q���N�'�2}�i6��c �rǁo�+)IU�׺Qp��3M_�k�y���̰�:v,���M-]ݧ�M�:�[�7:Q��!1�ͽ3� �½vVç�I����G%�����p���_�P>22R&��?��P|�)B82!���df�g�ͧ�Ok�%�~S�����)�|�����f�����>&�|Y[r�������C^������43sjǘm#���ϙƾ��OS��%9
 �⫪c4�����dUWV�_9�'���H�#�e���0':����y=��@IԦ+w���#�Ꜹ�FΛ;�����.~����� �VS]I���W�;S���591zo��7��J,���qjl��*E��9Q3ā�z�P�W��c��pU�L�x�=	嬬��!.$���X`V�����O�� u��)�z�\�#��E�@�1�GkZ�[tlG�, �<Р�M������]��ծ��Ճ�^���4��u�j%��
�z*sC�'����)=|c�!�]�~��%B��|�Y�zW��ĝq��p��[b}���EZ��˵����Wd���*c=cUF��w]�Lg��>~���<���MWel:	�`��S�l���`Π;w,���=q�)a� ������@X(7��#`�a��z����{��5�������t�]߯���+�q�c9�oii���,!1��7�
ֆϝ � ��RO Bifn�=l��x�ڢ�Qh'����6l��̭Ӛ=��G?�
�C
�s�����	Z�l|�������l�j�'0��K�cuM����;�Ұ��_iS4�cJ[��ǋhZ  j�U��d������M�0[q��TEO/75����XS�4��.R�gJ(DOo��������5��I��TjF4 l�ܹ�[��}�����k&-~��$�����I �)0�[�Np�Fn~^��G��_�~[X��\Fo�'y���{ϥ�T���թ���=�\֝��X�u���L��c��/k8Ԙo�$�tܽƉ��7k���ڞѬ�o�! ^�u������V�Q=��*�$����<<^999o��9��HAf);�����ʰ�&�3;pz���6ױ�"��x�.[f�ݯ��?0|l#�y��Ή1
!	��5]qn�iI�5�	��wc:��܆r�������D
��4,hd�5��%s�����l�5k�=z���Pw�	�ԛ�<Pq�5PM��Qs~8��H���&G��k=�V~��%k���Z�*jk�"""pN[8�b*��	��,/��t�p��Ȟ����p�5�uRΑ�$��� �1+L���(��}���W��i���;w.�40&%�R������V���/�x��T-��z4��}��W�h�`l�SO�Q�[j��}r���(GE�%K����⒒ѪBBk݆N�ʹH���AdR� �M�T�x2lm"�C�3�}b�yb�#�ի݊b��10"ҏl>y7ٜ��E��H,O�����~u�Z�5�<��,i)����5x�'�%������/��F«tAL�I��
.y`���-xuC�9����c���'��I�^�Y������z����w��?�c��,`�.�'�3t2{����Qk���p]� <5*㷆�?sVC$�w�^�����8��|����97{vvw{WTT覝�*�'!�XWKT4�L��eR7,=��/�X�f�*�	g��o�Y�8��r���-^-_'~|��tU�����h``��qWM���Fe*!�[*���}$�}j������|���S�gL���;�:B�DqH�_������Bϟ;�������Ñ�ݩ�X�/��_;q4%
S��̛���*���e�r�6���S*��Wnذ;|�������mt�Q%�$�f������[K�^������jM�8؍eY����	���sr�'��=�ÿ$;@%�!���]�}���t��v�n�H	�ft�-��ڧre�{d�Ђ7d(O�(V��Ek��c��ݴ·0�����7���@��������,��P���ɹ= �P�m��[���ÿڎih��.�;;6�!��8oi��tDޕ���]�%G��@؍��<�����*��o�!F�kǚ�����8l�OD���7tfzWӓ��&1w⢸�D��G}||�<�v���&��?9�CNN.�x^���������ud/x��r��&���N��:��t��.j;/��!s��IU8+feY)�-1�a�xkME}�j��Qѥ�{O�˭�wk���+g�\��O�t['�]����F���J���h�0���?_�U�] _
a�lr������v���G]Z���/�ǃt����m��&ɐ�����͠Q�
rs��<�P<]L���U��}h�|F��P
�+Dn�/�j�-�"?��(�����vq"w�;Rޱ�"����'Ё�}�~�Fy�OmY(��j��lrc����������I�u;��
�	G�
��FIػ�߾��V+Ry�!�j@=5=�]���]�V��<�!��D��HEc-K�m,s�0��fů�i��8�
&��߉��:���������ٺ�Ŵ��-�E���ƙ������W��d�+���8�_4m���<Ϙ�N�M�s����':��V�7��xr����C?�����y/8�o������Ԣ����@�bd'0�M���w�ΰ/^\���[�F�1tL{`�<	�C�-�`�R�'s~�#�������g��Ƿ�>79�[�;�>�Ym�R��%rw�[�~�N2R_�T�E���g�5���|IFfr L����^J�p�tG<����|�3�9:�}���u��Z���u�GF�ۀ�D/��| ��z�*��8�������|��h�&�D#�I��6���f�)��I���</�.�lE(-Zsi�v�!���iEc���{���@���� ���_o��^�y���+�d����r�W'ˆ�Z�[�b4b�� e�ޏWz9���HL���9�}Yפ{Wk�ހ"�Ы_oI�#����d�N��)��#$_[�Z�U?��i��1��,������ϯR��?���C-̟.m���%����x��s�T#fy4����kݸ���ϡ��bA����ɿ��&���֎T�C�n`�x�LQ�|= iM�?����/}n� �* �,������osfR�qп�5��Sq�I�GFG[�B�U�,K��q��	��L���L�Rt�<��0��.���J�po�QX�R}m��,D��L97��Q���|v�?6d2J� ��X=�r���d��5�t4��3�V�!h��X�SP�a!6���6�"Lf\B�.���n� ]|cq���o5���0
�iu����?�����A��<ΒK�½��	���\��+3!u�7����^0�-����s��A���߸��K��<�MYD=��@9�ļ>dz�3J�G�풓#1l.X~�p�p�~+�O�nW7�V���iI�2�	����$1+�WO���:3���-ɉ��ʐ�Ŭ (;[f$ɰ�gӯ¯�gct��5�t�̙�`Bc%�S��%��IXkc�>R��wf ��i�Mˣ���	��3-������6�d#��m�xӔ8�e���;,8�fz�.
�м2��9Mgr�^��n{�Gm�����?#k>�O�:X�ŻThsٌ�44-&TN5���?��孃@~pG��.���NL�����1�Y�qM~�m!��٘�ɷ�'��j���8�r:�X��N��-�m�8�6$te��*8�c��FAo�m����� ��0�6�XAw �?�?��؉���&�R�=�>h�cin�8	���>TU������9��C�2JvLq�t�m�BB��?���.���.�E�S������G�SI�0�L��o�1�?ZH엚^~P
�<���@�UZj*�@h�~��S�J.f"�^��Mw��N��5�����޸v�Z�?��@�o�8�5�8]�
@�N��2m.�Q�G��ZM�*�9%A��\ܐ�}d�1k���3�Xڡ�>(�R8[���%�	�u����V���:{�0�>�i~��a�;͙���������刍߶MM��@>�5H݂ �.t�"�����GsY �p�C.Ғ��t�^�M<�-�^�5.)����JD�"���|��
�[��L�3�m۫�*#�N6�	{'2==��^��2ߓIwILe7������y���`Fƴ�H��2*8:p�cF���Q�u�uLBB�Lt{o��8��F�X,�<s�L���bH�+*������~�.,X���}���OH��RQ ��U�s��)%��|�4E\�oC#Qm�k�;%�!օ����7�2�K�Ȉ.��6oR�M��8���Be J��dN}�FH<U������v[<}���^VB+��K��n��=߿�`�M�
�<��8�룋�ݳ�KXe���������*�Q��8u���kl����_/!V�yoA80*z�5�ʖKz��Y�g� q�hR=�����=�{cc��NvO�.�P��D�mZ�~�z��23�a�_�P�}�_2;����|�j7�#{&?d�>aaa�1�n���i�ijr-�8���!��;χ�ڐ��`�z��0Z�2A4���wV"Ȯ&N/����jz�$�
�L��&�M���眜������{bFL+�w�}���I��ro1(x���>�`��Q}��tEC���]�`dF�$(I�7�fJ�*Fjjj0�mF�R��*���zW�&4w%N7Tlkj
Q��Y�^���u}Dq�[���g9tDMk�-udd���ɽ��Aڂ'@+�b�t�F����ψ�l������қ\"�Tl�tT,�6�|�hu6Ǐ���; �@e�_��L���0X��zw�h��<�����+���M���c���] "�q�_H�de]ݪ���(�uK�O���.H9x�!��+�ٶz�� �F�������߿�  *FFn������ G��r����͞�?���l0+k٠B��X:-S�T��"|����D�=|�s�/v.;m.4���i8Ԉ�ݦhllL�hV�0���U����*�]ӟ*Z�Hջw�>�p9�������'����ʜ���b���9=0� @xA�ϟ� 5앥��sgZ�O����Q��d�{�R�VΛa$V��W���[b%�hق��B�W��9���iS�t�t�fP0õ'�"�;��A��z("��P�THj����7-`�T�ȝ�����-�M����߮�6w����/�K��8)1?&�˯US�<���\L��.�8�笀�r��g���}o�Vx�����!u�~�����L&�s!������h[�\�rl�Գ)0T	1{| ��>�aqέ��K����D���c���V}����!�!e���`�LN�.����w�]eZM��[j_�|���� ��@��ݻ�-]j�ċ��%o􊔼�n෯W==-{n{�L������*������/o����h C�TZ	tٴHX��J!��Ȣ�(d	�BNjZ�'''�6�웓�cim����677�ئ|�ĵ��7�OFc�>�Y�����8�t�>��D��<�Yjz�N���ģ�`�[!�E�K���>x��V����������@20��@�f��6��py^n��	���^��0�ǃ+0:\��o,\��ld�������t��.2�,-J"�#1�_��Ѳ���B�Y�ظ!zC�Y�B&���i��u�G%�\bH ?I.ÿp�̫%m��O}rA�qn�q��dkkH���00�6K:��_XЊ\~��[����n�;@Б`������o@+��s��n�A���&e�/����V��#���zմ���@}l'��K2ՀM��T�]h���O�N���d�v�a�" 
>�� <�M��]]^���0��ջl>5q.�r��-��-"B�q7����P#`����]�adOOߗ�S�&4�X�D?�����|M����>}�E�_FP��B�l8<�s���u ;��e�>q[�&����x�A=��"��í��o��ˡ�r�\Ļ|�s�mK���F0P�B��������bw�������mWˮ��7f?D�gF`X��*`��l�Rg���:x�D!�� nr��6�7�[�~���g����-y<�a3[0��n��>���Ba'k��e 	�.��\	����I c8���L��<g�i�b���zj2��́���2A�b�o��6NhR�޵?FDX̝��4-��)�MgO�?o�Ic���7���_��Jy����jժ�66��R�2N���v9�PyT"a.��k����\�����&�
�B�T2;�S���I�<ώS�Dʔ��$���n��3�e��3�w���������/g��s�^�Z�u?���¸�vsV��0]�jK�=�qp�p!�9�����\��$r����� ( a�{Q^��"�9J`Zg�WM1�UeeM
v��ia�Imu�A�� `�/
�X̢-�*�C9R2�>�2ӚW�-��r`3sss8��o�'���]B4Cv�^^�d
8~��OY�cT�)���y/� ����h��oݷ�>y�d/Á����J��-��X���MB�~�ԃ!����u�Rʏ�J[�d��OP����)���6�*�i:���|^�Ao�|�c�Y���ӎW�<�ry�-e�Hi	�ŔNH*6t��;���A I��>\�'��Lu�&�@^���-�����wu�u�I�a#W@-��34�wY�ms-.�6�nhbT�jaT!w�3�1�,IZJǡG��:�Z�v�a�Q��k;�I*�O#S�Xhw% ���4�CSwc�Xx�i��x(\���Ҳ�j��ȹ^1���
�5,,����w@�9���1�8�%!!KΥ��j�Fr
-q�%�����!�:�_�F�W��)Sdɢo�9�������e�e�s	|��W��k����,�� ��̀	d�$t}��5��]Gk�����D�x���|Ȉ#w+�'�!++�OmP��ò�%����16�\�Wu����R���S9����0��Z;(����y|ͪfa�Yp#���\˹~�$ƗqdM:zzy�ڄ��WS����7cjkϓ��Xr��� 3u����G}�Ʈ�Q��x��ִ�tͅ��=����l���~�@�Lk1U|����GC� <��.-=�e˂���?e``��(ר���]�lvB6ݼߕ�M����rճD�q��jvߑ��!�7��(��T������ݳ8+I����	qꍖ={�����ft���*�qqq�x1$���8��r��EY��+��`{��:�:�q��&^Im������7���-.,���@+z��������t�+[�J�$��a���'wRT�BU�x�:.·w�&�S>�Ҥ�˷��kt�Y��N1㗅�/*�����K���9�g�����\c��Q�eEL�����M�g/0L�#I @�B��!j�OIr�Ww�������M���N��^
�#����h������I7�/��|r��w�L�<A�*~~
�YB^�͐��/G]�6�^�b�l7��ހ��&k/��Vn���b�uh\m0��4D)eO����[��&o�hyww���Rn4e�UW��xU���x�w��ˑ�%!E�G�� 0�`h��Z��XA�A�".�N�Yʓ��k8�tB���餴�a�s/眡9 ^0~��w�_�6��3F7+S���zr?�)���⓾�l�<A\��ek��g��Ţ�����Fm�]��0V���+����ԥ�5������gl3����HW��;7��9�). ���/�E|�);�f��#WUU�_Us�^���H�E�i=�n޺�T�IyM�r�����[�eg3::�����I�㫸!��%ෟ�(���"\���P�,���bZcT'�Ny� 0�8����7����O����Ʌ�,5�(���!`��ٳȶ����&*	R���ױu66�=��q���%�]�aE��a ��7�Nn�~��l��^p�]滇�b\��R��Fݥa���m��\w'���$/�} /�H�1ta���ج�f��O^l�5�|�^l�YS�\ t����@�cR;�Aoˠ��T�:ʚ�1O����--O,�����q�C����ݔ�S����SP����"q����a����~�F����TUV�ƒ��o� [��i�[@Bnpὥ�]��2�����X&Ld)S����,��/�5jи�+���Sa��--���\��qǉh!?���C�D��C�Qv�r��7��{M�[����7����.��s�n�̱jԨh��?���Aު�7t��3&���w�#� P蔶G"��@� �a�v\����_�(��"ۦ��>7g��аPW`�U-�`�]ܖ�R��"OKؽ�yX�.���L�w��z�|���o)F������5��-5�EFզ?qq�f���<1������ |b&����GiC���W q���
q������Y:�~?nk���hB�235���4�EȺ����0.��o���`@�}��$��quu��y� u�d�P0lѩ���'�1;�*r{�ې��w{z»x6��J8�����B����(TmC�	+$���I�ס����� 5�a^o@4z������5333����yy�p�3�zAƅ����d͏?��&���O��3�Z�G�[�Y��k\�-��Zs�Z�N���,)'k�b�Rz�毄�dPu��ٓ�
�8�"bA��$��	�>�%��i'CC��C��ۉ��� �DA�^�elll�+4΢}���' xV]A��j$���b��)u��-4#
�%���^s���U���*�5�E�j�7��fh;#�Τ۵ ю�)��m�=K^���-�h،����(�j�}����-�B���k�T�\�y���^�~�ݘ�m�O��!���2V��G�#�����W�I�M�B�d�+��E�p�M�.���^W�3~��n��D��dj���?:
M�Țȼ��Pʰ4j���_^.C�ۈpxP5�(� ��f�f;��.�d��SVV-=�	>� �H�@��W�7��D��:�4;9�6�󤘘�<"֢�Z�#�"{�����	���f�\�HY!I����������y� �,dl��
�@7i/-�,W���?&��pp�Ɓ([ �-;�w���d烇X�`�e}����P.�6�$�����.BJ�CI��@࿦"�-$GV���5*K���͚l��ic��_8;5��D�~��D!�=kћr���O�Nۑ"\�����7�����GmB�w�G���P�^��*�(��,۷C��GE[$	,��i���Ve� 	0j;�r������5���``N�0� ႁ�<�Z����D�N�iB�p�%�R�^;;�Hy�[��'7�SfV�҇�yڨ�*!UNQ�y�Ĭ�3hܳ�ewvv�@�nyz�y��/�y, Yʏ�t��n��
�����@\^C�Ӌu?pB���ID!;����܍������b�h�3;�l},�����F��Ƃ�'����(����BhZD��A���D��ᖁ����^��A�w7��mも8GCk�Z�g�q�^PXD����Ӣ��,v�����G�!Qÿ�t+�zv �sݸ^BRtS��.B�H\��+�L8s��a%W)��I!O�0����$ ����=Z�E�u>���9ȢI�aq_lEhl,�e���l02)�}.쯿�"�\yBE���3�H��ʲ>n�0�a^(�ښ�h�̶�R<�1�v*�.�#E`�
�9'׋1Q�p� Ty+����Y���Ť?�Mc|��ڊs�Д�ɔ�ag!�S Ehs��� �	�����ؼ9"*�S������CD����m&�g��Ͱnjg�^����6���yӄ���ڹ�&]%}��O�HJP��W�������:��[��]�*��p�^��a��B��U��'=�k�^^KVڹz�L��>N�s�R�:$3-qf�a����ؚ����
l8��t��$�~�4n&x�̸����������;�HJn�d�����_�˫��O���653�DK��B�	y��͛n�PfoμW�1�d]�L�{������U�zzhi�b���|cpA��7�O-1 ���/υ�7~eQ�KJ�L��A.x/p*ـ��o�k:fAL�'�����d>az���_��
p�4&�L����׍�࠱��.��S]�A��J^6��P�]��4����~���YBY���˗!{B������A0�|k�<��Md��틻�!�i��	a2�[�����K��K��j�s�!�F�3yS�@�[:��y��9{ԯ��Bl��7멐�l3�B��_�>ыI��W[�j҅�F������,6���4i֕�oa�e�s��Z�����օ����ߵ^|RS��E��8�o=�ɵ�&�lVW_�%�SJ�����%�CVRJ�3�.a�j ����)�������	�� eO	����.[L�S,B�Z�9��>݃,�5����ӳ�F�lS�9�/����ޛ
�k`p����t��i�	~|�ۓ���(�J
/[Ԛ����P �<� �ŁB�DO9�U��׃«�Yy�{v�G�r?�K�ý!>��� [t�|���( �-"##�{�F�a�h/*a��Gi77�pj�o�/����Cv���>����������;����S�����k��D�����`��e�4x�y!��3�����Pг�v�_��D|$rr����4�ir�HS������;uOI$��'��č{N��g��v-ҷ�
���fgvJ�l��f;�t�G{�ns[y�:l��+�&�~Z���~�:�����ނ:��إ��D��"�wڜ\AcM�VT���o�� {tK�?ioH5$�p�����{K#�&�X�������fo 6�Á!�9�����t7���W=��+"�^�����p�1�����	e�[`�~!�5�߸'�vm�a��;Ӈ��Nn��#e͐�\ٺt�֨����_B�ۏ�>ccc���{���W���b�#AP9|����4�?����٥Pg��)�d s�g�"���v�>��M�o|�����/>>�v�"�8B|�Kym��*K
�j�)~�;L$�<:0e�󬰰���x{U1.,`^)&�����1�>Pboo�-y$������Ե� ��<���(���s~� tZ]�ABF�C_����O}d��,{!�\6�����!�]�^f5j�,:�������H0��"�wKE�,��wo=G0�����F�[��+/>F~9?B�PPP`�i��0�֭�?at6&&��޽{��D�� ���؃��F����|��w�D�����S�4���4s;��g�����_dU�:�1Vp����D�3r�/E>U6�<6ߪ>�!��a'�+�U���T�&� ����Y@@Ey9��0�|����� ?Sè�)�b�}2�6�"�o�q�b�~� ^Qm\q^0\������n�=��p����T�5MM����A����<<&�l�^[[�Lh	�o{wP9�`WIH	�`n��f��x?ga�`l7��c�!��+(��R�A<���Fq�Q�`pk���OL�n��r�x���uȫxf�جg�O֪�qH���l"IP!�ߐ��,�~�T'vAgvrH)^Kz��ا��HY\��Kb~
R�����O5��^B`����=�|)b��è�T������&�4?
���%,H����/E�����)y2+����x����D,u�3@^M�L^�0�=R�
�;
L���'���oH��Q�o�q�@�sI0�����n��r��&�	��@�0Q���4Y������xw��9�/R>b���3��_<�=��HoTl'�N[x9u�<#p������>Aj�N��_�S@��W���v���<�����D�^��
�1�_b�?���$텪�Rg��b�� ����!��=>�UңL�LO�Q���_6XEk3�J�V�����&&&�����oU��cV-N��cU�?�a0\�Gyno&�!o���czv˝�A4Z`s�Y��旇�ώE}ݯ�F'N?��K,�%I����Z�C?�qx��R6npݕO�F�W����?jѼ�
��8��e` ʄ�;�~$�dAU`���l��>�,P%м������׽W�S#�$���H[����羢@���|N`���`CJ��y������U��V��U�t[��y�c�pT�Ƥ��D,��غ�С$��Eqd �Ԗ�D\��޺�)��v�lllf��D��6��a�����VC�嫄K���v��X���3�Px�Y,H� �U��⩥3�@�i��"Yd i@D1���G��w =s��
ѣ{�]�jR?�J@r�]�Kl�U}��m(b�s|��XlG_p���駿Y��5�l��]�3���oZ��'�4:�@y�Pk�<��i=֓��xwŧq�����%�JĎ�Y��X��G���3�r��J��.��/ y��B2>Q���v���p
���:��S�_lH�οU�&��N��fVo`���n�ϫW�p},$|�tSiIUMM�Z�ɿ�����.]4
�.�;���+P�!L�A���B�C>"���R��h��q�P'�}[�	MR����Y�� ���>x)�Č��At��Kn!�q������5�G@����p|ρ\C�1����,���;�531�0C����p�0��fL)�8'%%e>Ф
=Z��#�^� �	�g-��T.�{�����d-�D�"�2 �lOY��"�0v�������d��h�]�iRn�9��k��\�&L�y�?���f
�\����ʪ���Uʹm�v����vN�<yY1oJ�v����-T�h�VJ��%h��ޞ�޴A�c"2��%7�+���ӊ����ۯ�=	�6)d��c��&��"�B�����#�T��ROT40�222����/{;˒��gjKn4�A���|�͠�M�Z�jk�qE�G���� 0��=y��jbLMM��^/���1�|6����!~RA��xG��Dnh
��(�@x�TZVSS2���[}rW����aFډ� �%�l^{�6EPI�F�'�H~؉�PJL���o�h���|�8	����sD�,� i�6gcc�)���P$�P��I�yMڹj�̧����|�f^J?9�sE9A���`�@O����o�>��yyx�b��b�7���m۶�o���f&��&p�U����O�O�4�)�@�����d3!�@@����4�t!��jT}���p6�
�Q���$
��OdC�F�`�e� �>?9"��)���
�7�yTP+ ��V����n} �G��Bŭ�1=Y֙`]����.,l�Y#h��s�QMooo�Tcmԥ�Lđ�6�al�Yq)�� �`^�P�?FR����^?�PZQ�Ѷ���}�.�rU�!S�o�,��|
dW}�em�����q��H����ʤ��V���
��y�" c�p������3\[b<d�2�A�ݾ�8M)����>���K25���-�+��,�;��؅����T�8cc�;?����~q8��\�x���Sȴ[�LZr=JB��.tv��ܔ�}���E|�S��H����f�ׅTVW����Z��[�6i!���ë��p�B��.���鯯/���j=z�����R6�w��Hun���\�=��X�
V�폌�.p�6�b��R���c��7LSi��	�dJ�Y�|�/>]��p���SD$ip�W��I=ڑ7Ԗ�vao9��q��dd8�1<<<�QRb��c�Dtt43y�Sٜ�;/d��9�@E"6f <���s��m�st��O�w�����	2��V.���� K�mO�7�56k��<����W��!Q\�E������L�w��	�����#�.�h�b��8�!>�'ۉ�Ɨ��n�����3 Ԏ� �@� g1s��\�>�>?�=/�n��-�z��'s�w��&]����R�I� Q{w:��@@b�X����i�jbe�tK𚇡֜�o��><��K�C�-89q>�x�c)v�������<�O��o(�H2�*B�:��hW�JG"z
�rqad˯���
��8��g����$�FGl8�h��R�$�F����y��ā<r�!�0 ?x�j�z a�o����@��c��F�<��OVS�#�%Z#�EPK�\L�t/V�����#���ő}�3�qf����C"O �	����5 �WJ�u�J���D@I���t�D��a��y�S�Ne{Ǿ��!нʴ���)�K�I��G9zo��W�-<�]�/yK7��{֋�)	>~vWȤ����Uk/q{77u�JjL�r w�L�06<i�@�Q.��K�Uf�_�t���+'��Sa8�e�\⃮z�]D��g5^�3�y�l��8�S]DǑN�6�t�@����^�k0c�3�i��#^������O��N4�X�R�f7��@��Px���VEA\#"�{lԧ -hP�UsM��l��mhr,p}���,��=�>�N���'9��(��$dV�ӫn�aV?��_װ��v�7�.4/$�����	�~R3~mV��UĎ��ԨUG���d�2ż��>,=]D���en���92�4�GP�����mO�۷?�E?ĂlSN�/zvLo�O}^S�zH-��8G�����Y4����q��.+6�0�_�h���
@���c���H�A�Y��!6���"��HM��&�~"�s
�� -j3�LԬ{�q˻����Ǯ�@�0\�Ϡ�����!ߛ'h�QAA���*�d� �F�#8+�y)���NN�o���� �I7h���Xz��V�Aќ���fͅ'}\�zյX��& �Z^�/vٺ
R�e��\����`�NT��zl;|�o�	��t����K'�7�S7
��ޜq��0�/���i2@لX�*� `c~S�M0(�K���x9`i��
`,��X�\]�>��Ԯ�����m@"}��F�JJ@
8�gq�1h%��?�(�ع"��i'�ֳ]�!�?�W;��%h���^t`� ��1�],�����qJ	r�����H�>_� ��<t���_��͋( '���y��=W�����!�m)�y!�y!Z@K���9���g�l�
�C�I�5j#F�9��q!pK����f�t�sF,PK<����]f��yr2s�Jf�U~����m�S�L��o�+j�=���d��ma�	��ܞB��B����z��^�%]PP��usyMӎ�%����vf��APǖ��s�|߂�C��x��=��t@O��:�kY��)L�0�x	���o�fpQ�����}.k�U���D(pg�THB�'4�T��-����� �q��6�w����)-V^�W"��|�1������x/C��	r4`�����^�\�wI̺���von�<���6"�	��ː^@f�N��`p�bQQ�UbM�f�#<W��,oNw����s�AF(~��p	��ϑ����;u�N��^�u% U#�|:]�A��m��!0'=~�U\\�5g�^�10��� O�k����P�^���1ș~�H���X4���Z��5۹n�*Uh��Y�e�c^�QJ���{��RǪ�M��F���WG+WTW_1e��I�������q+R5%�I�s�Y%V#ͅ��K���Grc���ZGr(@'2/�Б:�X\�[�����M���8�%DN� ������9��O�AD�W�*�j��vs�XWI���=ni2�,���������|��a�@䍍�����L\���<��J8�= �:r��@��?������3����1����z�������,[^GF�M��.��5�G��������v�k1�C/]���ZgkApiiF�����W�g$�<�K��8�E��X��\�t�~�Q��):0�8��'��H�~��#�]vX�S6�����\����/���逵��b�&^�sL���2��!4�cѢ'�h;0�^]����x�I2�cйZ�o��O�S�Ĭv��!V���m	�}0�g�����^�*�@f�A)"�~����X�6]]]��w��M:ρ6Y3)bi~��.�[�wcmt����E4@���qڝ[x��:!�NaA���_�*���3j�g]���r�*�a{���I%1s� �\~GL��c2�)� @��-5ʻH`P�qd�� 낂���E�L��}��W		𿙳�c9�UA/B����3຀`������A�+Wn��DFF�^VUm�?��	��U%%�����i���^ 
1Ԧ[܍�ٞ��@� �Ԭ������g���:ǂw�Y1����6y� ��5����]#x�~��A	��K-���P��t]}��t_�Ns��ρ�|�JV�0�D�����@�O������6��M�J�DP7��'�B�k�Q����Q��H �_�Q1�@GVU�;�ׁD���:	'�\�G�(�^�O9�~��D<	j^�|đ[�����j#0���U����ٌ�P�!0������eho�eHp���y�j����~C�Z�q�� @s /�7�.s�'k�kHOK����~{5��X�g?	�`�4~�� ,�']�l��q!(m��~꺪��g���<�����ׯϜ?_t7Z���
z7�Cڸ���d4멯/s���d��4k��	�֣˷;8������<�Ĳ��g>vg�;�:��a���2�.�=����#�˗3;��E�/\�|���
'� ��w&�QVq۔�j����Z����S�tQ�N���׎��y�3h�@\���d���v4�˃�n�]�߆�?s��Z��g�(��*��?��ϐ���7�oKA� ��Ѿ���#8�0~|Sf7[���,�~o���w,m�QCY��(E��g�����FG`J[c��4v�1m�5+U)tN(��|��֋�ڛ��P�����ձ���*'��h�<�Y�G��/�ߔ)�(�G��Wb�{����3�j�Ӵ�YRt$�aЗ���T5�h�$[�^�}���7�f�TY�eo#8�h��%.�K�t�9ٴR�1��x����z���9�a/��GM��3�9�؊���+�8�V/?#)Q�9"�S���D"��X~�t}���q<�C%*������(�f:������MOOo����6��/�T��JKKn";�m�Z�����3�t���~�J4n\�X>�	�!7���p�r��$.�L��u�k ]�VwP=p�'
!�������H�:9>�w=U���G�l|�I;�oY�&�^;�����ˍ���� ^��i�v���7��`0�l�XT��!@XD�f�8�m�0�Mu�x�ML�@uZ���Z��C8�Șiܯ���3jB��TM���b�V��I;�,�ö����L��c��uc3Z��%@�C�TL�
�P�Ĥ��<ΐU6��ĹҰ�H��{͗�!���\��љ���S8��r怣�Y�P=$
��7{V;�9B������ t����C��s=��~��&z*�l�p	�#��'Xv����^���'6cS�9@�Lk3���9V����<$&�n7Z&>�}��.B�0��W":r.�1���F��"՘;�FˤLȳS���h'�NՖ����>ק~��:#7��8�Y�|�#��؏'��S�C��n�3u�AYV�C�&��v/�N L���뛙ͺ��PjÅ���W�&�@"�O~��j<�~��s�)#����!/<7�6�@}��-����� �M� ��Y]W�,d���nc�:C��@s #s5�����M�M0�	ҳg�Q�PW����ꍌXs�[�v��L����e�3�������"�`����ٿ�ĥ���|�^KSU�7N�Z���5((�)����?�0��moWF��'?b������%��$n�q+�z����C<P���e�õ�����}��F�~)��
$<5�ŋ�O�91�+�jA ��~�Ձ��"�l���\���:d���Zl`/�����/������޳����@�+����\��`1�_�̄�pc}5�AC��爙�m���6���i��/cx��is�j}��ky���)	!�a-x�$ԋ��k>�z��%j��ުS:4�pB%k�� "!!aiuei:~�&LEeOG�ZX0��� ���_��@�<yb���G����!��&b��awf���X���܊S��S�b��KR��)� T�x"���dTF� �>b{�M����֡ͽ$R�E�H�k�q];<
$�	��e�/i��X�=�kq�^Zs�����_�3�-f3���m^뺝l ;@�/���~���w��xrvD�sy�ZG�;�&&& ![�{]ʇ�К1�	+�~�fD̘���藪�$����\�)��?��Q��5(j�K�!�n�i�p-���ˁ��ƥ�S#]n�S�<~��͎�v��
��¸����s�b����9}r����_#o��YV��/�=� @��b�K1��4Ϩ����aI2�.�ʄL���~�.p��9nj`~.���_`Y�`���^�a.v��YX޺0td�)�1\7N�	�~�5����0eO+Ld7{i�z�+�;�4.��"�e\T�ub�o��������)�=�ů��E���`�����9����p�}��@�sy�'�=���;]$f���f�(��|��)��T�
�_��m�#�v<�ي���aX���O�P&T�,?M�g��.8�n`�?{D���cf?��.��y��Pw���_�S�-���U�C�<��M3��؁��o&�S��l�\�������|��� 
P&�R�@���`xv��9�L�^�j��4��kl���X��'��tEFs��]W�dv#�ƒ�E����C�q
�>$��������y��.�[���s/�zJ����w?|	i�ܶ�G=T�/�~/hQG@��ʂG�ϞH�l����?
� uCX�C@>�����H8����mm�w~X���Q�	��o���f,G�փ�����8ÁgS��뮀�Re��!wʤ*U���U�d�'�~����q���(�<���7����g�j�[�N����NX��
�}�����t���z�M�6nz�f�|��2�x<�!�EKϨ���]\�ݵ����j�5\d`/@���Æ���A7Qkk3fPq6�f�C}�ϡ��B�/C�G��:����H�����yj>�\�������
�f��C�,qf���P=N�^)?��@1SPy,k����i��CJ)��:]�	�}��%I�aLS�nZyU2�^c��k�/���}��������J�P���t�_�{���\mv�]���K�rgY����(��R��H{X|g��2�N�K@jXW���XI�	n,�n��������zf_>u^�}bN3�G����J�����20���O��l!����ƃt7ˊntww���xƐ3���{..2���V������^��W~i��1*�����?~\.c�ӌ����}<�8H�Edd����w:�1�}��ܾ��#�bﱟ��EB� n��%�bTC|��Ѣ�}nf"��]��+��8'������fև�K���U�pch$d^�UD�>q%i"���P�����}��pHto��C��\�/�鯫n�w�Z11��JTN�|�uc�#u��/.E>��ˢ�����a�!p4��#�4p8�e��l3�Ɍ',LOO{�S��ٗ�\�y�\f���]��x�Uz��+t�z����)1j��Цd2�\���i��v cπ�w�Y��"�J����
7�М.hλ����|���DϖP�����������#��� 0`�'+I�?����1?���nsQ�l�[�W3��y� ��߸q�l��#}�$(ˎqMʶm���R�������Y�mR�vp�ioN���}9����ǫW�~����p�8��ˡ�=\#�3����Ƈ����Kԓ����2ǉ��:ũ�N��}�xN�ߜ�V�l�q6��5��Ά�U���]$>8�����s��mLa6e������ 
�����)�۳g����c�aX�9٬pvv�3�)�mk㵩����{�Q&-���LK�g�ka�3 δ��R#��BT��T�o�b���4���@��-�_�1E�g����w-��;��9jZ�N�F��e>l�b�?�Vw���f}�9 ��=�Q��3ý���Y��+&^��F'7���|K��\	���Z>ˠ�*άn{�����CY�ǻk�|�o��2���R�_B����E`t���w������]�O� ���]�d��+�W�pZ�3�I���#d�������W�0� �^��ō
�z£3���b�������K��0�[��w���}�����W��:��7���8�5#�3�n���GO8e�X�ۍiǶ�P���#'N�H�ԖPn� =����0$����o���Ϝ��>�#���\%�"�<���T��׊	%�7�������T�UWo-**
_��� �1333�a����Qn2��GC����X)�;w�|��EԶ�<�^����ge�����b��<����<��ێ�'QWF�5뭌�̓�߄GEFU���V7t���1����a�UR�Qז��͎'���b?,$�d�8�hǈ' =~���[��5�J1�)?R��,@�+�"�UMS�ה:�Gj�O�x��|�n��x�i"�O��b����n2?�=,*�b�f�}�]0�3���f�r*�Ң�30��LO.�����������:�t��OF�=����8���s[�v�/8?_] ��ҙ�hl�<#Z]YɄŵ�
iii�x��� ����?�)f}Wz�D�^a�*2uNtn�b蛦�w�20E�DU�N����-x�Nî�����N�lV�b����啨S��qP$�r�gZ�������� ��/��il��n2:1��׊�>��[{"BA8���l<l�aVVV����[���Ш�����y����	�A�@1��Q�M�RF� ��J�6<_�zv5����	��E���~� ��@��P[�,(8	�U��	���Err��N��i��R0w������ˊmQ���|�ÿ��u���se��©ٍUY��MȔ\�j�,2q��z������O�C=��m'g;��K����]Ij��S<9]��Σs�*:�h��/��H]��N��v�P���ÍKH����R'����9�Jo�8a֫Py+����J�(^R?��g��Km���=D]��i�wK�����=��BMx�iݺuq��'�}�w,$��2>*{|�o�n*+��y!𾿿?��^3�>�t�F��N����t�q���K��oH��ܸ\�0@�Qg�?��E�盪[=҅{VX\�'��)[�I�[c����r����]�^?4T�l���-����>��L�Х��c��:��J�ˤ[Uo�z���w&�rܘ۾�i��ֲB��"JlL�������t��GT�z�.`!���x��I�m�9�wRn�ō��QWN�����L�޽y��A*����q�n��VT��C�\h��f�!b��'��!r�"mGݨ��7;��3�:ϯF��
��d�a,�$PĂ�{�F�7�O�RMt���渭�[F��y��VP~xf�	 ��{St�u.�ݼy���z��v<)p��QZnE�7� ����A;�����eJ�=z0%���8�����������cc=���9�Y~��]��@�����{w��IWq�ؖ���y����H>�	��	���ު(̊W����Xu�u��?oK�@�Jʚ�9 �w0���W��ek(�}㼼�Zx�3�s�n���_ܷ��w����ϟ�X�K�������U�`a�S{H&�''|�_I<|H=K��իxH�E	���Snge�%��g�]���R�;���K�Q˴N=z&*l��w����׵��B����f;5�O�x^0��]ӫ����oRX~lY
���p��Q��'Oᰜ�@~c���G�wv ��9k�D��@�>	�K#<4�A�C@���-<��q(R֎�#NM����2J�����fx�4�-�Hr�����S.��T3Ѯ�y���K�>�zeB�&�g"��0�	lO�=z��)MM̓J��$������^�O��o����2aݺ�1��?[��Uu����C�%P���p�����G�3�B1e�?0�a^^� 0����o=�J�Zu��ƻ��H=Dp[խ1�6���\\����}i��J�g~܃?�p���s�#�2g=Z���� ,�q��@����BɒkVPٽ�!�J%z�K����ȴ�
{/wR飝���?����w����]��*W����U���w����]��V�8_�V�����A����׎$�OLW����ΩǤ��4�+�61P��������$�_j��K_��@�ܕ��-ZMG������w��+�]���
y���!\����+�]��
W�������w��?Vh���@zL_����=a��pqպ�߈"��M�-��IwB~�����G�p�o]߉�)}���1i��� PK   ��OX�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   ��OXǐ]zd� K� /   images/972a987d-5ae9-491b-9c1c-35ff468aee03.png<zUT\���n����6xp'�C� �� 	'��4hpw�����ǽ���sN��N����]�j�WW���I�	  p�e4  �������u��Bp��$���< h
2��^&'�h�����*kE�g3"��n2'�5�k���}��z��k��Qr*��zQ�E���P�AU.%}�����	�;ޓ�k�EA�������5��Y����� w�+H�UhQ`�����	�dC��_'$�Hn���o�)B�х���Զ!b�`�[�������߰5��:�r�v��khL �t/�����v��K_-)��i7�8yol&�ө�������;�FF;����d�^#��D�a��|�����i�2���O,i�B�K)����SJ���	�d�`�-ǺU.��I���_�a+^��G�+�X�Ǹ��K/R>2��W8G��R�%�.��*ou�G��/�H�9u��{<i��'�G���'�*KR���k��n3V �6\�;l̊�n��K��x9���r���9�/�J�h�~В,y�t��J����L��H"ˊ��r�k\�}ff�ƟgVH�a�
�q�,T�l_V]z��)���<�#=�B�6f�z!�]&�5��.;ޤ��V�������r�{�n���������)Y�km��~��$�� �gz�����̸YN�#�f��x��~z:ٞs�t4hӨC|rS�ǅ�9?�UFr��?M�?����|�>\�5En�$GF]��O�=�_-;���>|֧=�!�����X�38x߹�s����SǮlћ���ۂW"K��� �r)��pﺐ�9��_��vw���ֶ�NW�Η��G�ZVe��?����Qۅu��|E�켙Qz����̮�+N{�%��U�ݪ͚D��L���Z"k��Ǆ�J��%�k���< �z1�*���Jy��DͶ|Z��1��3��
�ٴ�d7��[�7�s��y�j�sL�kH�\�o���H8��t:�5<�+#��6?̮>`�H��&)ο�P111�WwN��ڧ���*$0&}h���:%��d��d��۱�5���a쳨*����'�A!�+��G3�)�t��]E�0G�4|�@�����]�=�'n
3ާ�����0c�oi�-3g_����Y��8;q�t������Bt1pVc9#⣙�tӷu��p&��������(w6>�T��i�
��i�|4��@k�lHش?m�J���敒9DX�\N�(�
<B��T0�+k�.e���3��	��!���*���l������Fυ���w�o�Yz�]O���)3��P� �������Y�E��a�k���VUq��in(��L1q=�5��s��,'{1��L~ ��d���<m�t��n#���y5��ξȸe�N<�B�x�h���0M�}��]�C����4�|�ʯ�;~�\���<"1F��0���(����cCgK���;cqC�d�����5IZ�ln���_�Q�����Wnr����Y"�ٞ=�%���������g�)~-�����O���%ȈA�����cRdR�}t � bn�����8U����d��>��i�����IN�_?!�}Â)�ӃfN�j��z��{	�E/�vj�-��gBrh���F��FX��AꜾ��h���G��I[�l�Dds��if+�Ṳ�q��>�l^kE/ݧe��>��߀e����·\\�������<�!���GPeG']4��k����F����?TE-ݐ<8'k+s�0��Ш�����x]j��U`C����]�D������/��M�'��⚊�y��26\U���~@
ش�+K�S��CZ[w��`n\���p�A�u��h�x��fcƷ��_�c��N��!/���*~G���Le�Aċ��
2����!"�0m�Oq�ّ��o�v��'���=�r�1Fحt�i��BC���يO��]sB����n��@����1��VМ��K(�}������	�}�(��V���%t�p��UI'�^�P�7-��K}�:>bk������Z�S�W��T��sW9}���}#�>�~�����Q�bР���bBt�rF��Z%~2�c�����������B�!
ؙ��μ��pu�S��Ɏ�PF��Yۅ=�5�[�e�J�$����sC�(�"�tc��2'v����%�A$d�9�z�����w�TmE��꽍#�)LP-��>#��W�.vw6=D���
	~ �l��"�n=w����p���Q��Q,��j��LK�7�vU�6ϔKX����{�����3fݥ�VH�����W�+�s�ȵ_G���fz�+L7�e�8�n.�Ґ5�2���#Λ�N&-�Y�P8�CC�g��|-:_,��{���4�zb�Ð���Qң��P���I xP��� �@��pR�=�� �Pm�3��|��l�Qd��5чV���A0�}�v�{wS�� ��jX �)�s�e��"E�"�����kF��/Oi{ �n�*$�<氿>�O��4Hg_!1�fc�U�8�c��ke�R�9)y�(�6N��T0�tUi�ܜv��]�e5씪�ٓ�f��%��,�b���Ǝ��/CJ����zd�(���!=����*$�G�kq߄;����s�r� �QZ�V��]��zE-s9��8���ɛi��侮��չ'~�A�s3�TU�����#�(�G)�-�K�=�m	�S��S5u����U�ܮ��T�}[n{���H-�Yc���~�ը��{�����=����\�����3B-����RNB��_i�J���8v;*k��g�ܶ[����AU;F�$]���2��.dA`�� s�w��8h���~��x�~?Z@�뚸��\.�pD��O�����h`���@��X�~J��K����|O�_�᩻&i�1d��>[�7�:�1�6]�bW�RC�E|6"4|���l�tn�#]��u��J���o������a5��/����o�{���-i�{nu]W�; �z<	���_��(�֫���F��nM��d0��۵�@ ����ˁ�2�v�t�Oܦ|k)>��+4� ��=��o�/�%��~���[�92��/]/{N�ק��}���ވ�&���jwP
��dm(�AN���z8����%�Q�Aܕ�����@�/�U�s��D���gK��N�����WL�G��un���!���O�U��f6�2�*�?`�
ui����^�q�*_���ٷ� n1M�	O�����Y�|^[��~�R���_1�~��~��|�;��bP���"�g��訬��b3,{tt��� �O^)1aw���rнvZ�q� Jʗ�)�5�+0�n��y�4$�5���Ga`�Y���H
e�5F����~<��Z����s[�a?����̴�P�^{���>�r4�]��f�+�l��1�tߖ��o�W�{q�����0�Eد�?�$E����.��;w5�R,8'T	�?qepF��zf�!�UX.�i]Ͷ��S�/N��{i�����Ǎ�����sEc�7Za	����B�	O͐�Ւ����=<J����fE���s*�U���2�
�'�N0���ߝ���m���A��՝~���~���ߢ~M��ņi��j��LŊ�k��x���f��{�s|s��Κ&�K�-z�$/�g~���T�5~*�+�gr	����>a�܉b�*��M�J=�Ӊ~��^�7)z�f_��$�����5������o)�Fp�MQ��N�B���u/<��ڬ:z���='��?���J&�:��8����U%���� Oc1c]�O�z�h�/��LŶ7�h�\!�~�7)�II����"�����S����y�J�M�`���]�m�MN{�xh���Z�s��ƚ�u�������/�D�r��s�2�`S�s�7c�>�	ճ�'�}S����Ӥ$�����J���WLV�����5��t�����K���x����q�kd8U��4�?��?�O��¦�T��_�L�:�,W�^��l��H`T�3��P7d���3�����(��"����N(^��S�Q���+�K��������⼋�Ѓ%��	�y�9����݉���~�}oܴ�&k�;\$rw�J�`S�����A�ۯ'�u��n�|^ú巏�㧳n�k`�'��S6fV�x�M��� �����v0�ړ���*"�9��
ٸ_��`n���9x~ �e������\o��:���7�%&^���k�?�,܉V/�B~���Ia�3�q�=N ��t���=������-�dU�w�$c%���>~���O����c�)�#�O��4���w^�H�R��I�Jq7�@a�E*o��u"�E�F�L����̬m���M~���;��J���S0HiJ�2���lB���b�����OW�Lfz�g��T�m��ԏ��	������-����;��Ґ�(H�I`�.[�%���(�<Pr��8F�"01��>�/T�PCS�:�b���(x��[?��I�������_��5O�)����� �=�m7��H�y���c!#�Xm�p�P7<`��EPD�����Cm�?!���[1�.��^���l����p�6� px:v�ⱡ'8T�,���r	��X?b�@��@��&:�̛�L�*�׹��4�J�e$=�{�
:~|g����|�!������:N��$a+�9������*Z����j[
Kg�����}Eze�j�lM������B�Ϝ*�I�@=��6�/�N���D�W5m�}0�� {a���W�q=?eHP`9�!�����VQ�?����*rJ9�q`O,��L�H�����������K�ݱER�a��@r�ȴy��P^H��`P_��u�������I�U��bD@?.��^�Mv�wN��n�p���[��a,� ���B]X5���?�qzP����I���m�wcK�lE��5���OYh�,e:+���靏b�HA�^eo���ybW5X�9��YBޑ��T�Sb��{ni��z�p_
R�o�4pc����i�Z,����`v�d
ėbv�W�!�4�wj�N�*���y���3�A���[�/��&���fX�d�oC4�
���+2Z�B��$R���
 YSu��P��G��L�m�*�+���mVp�]V�ix��%`�/�]E�-"�w��M��< V�7�ȣYL��k0�P�g#��ڌ������`~o4�c�0q#Y.�4z�������e��� $4����㪙��f��zǕF�S6E�)�+T"?�Sq�P�ߚ�(��l�j�����{��w_W  ����K�ru���-!fjm��18��="K����ڿ���Q������k�uFDgD���?j�KmTk$J��	α �X�����$5�1,7��~�����d��]k�����)p�\�n��.������F�{�jƎF�d̴���mX�dvg8�����3WHC__!�ԫ�[��[�	B+>E�2��@��3h��5���'��f�}J���zF���6>/M�9�ϝ��^M��b����[�j9��9-��*����Uʥ�+M�J�m�l�U���&��7�䢺����P�b&�.��_�1�N�y�>\�z�9.[	���ǫ�K�<�����Im��:�m��?�+#'?Q���ǟ� �J��OXgv�>���{9��=/q%l��C�f�:n9�*)&]��'�j�LNz!Xkd�&me�<Ԉa�J���O'��O@��4h�wL���ZYխ��xQ�C3�.#QT��R���ٚ\3	\Ԥ���ے(�����_�h�
��}c���U��]�_���Zj~�jr2eec+��d�B�:B���I��^�$I�#� �N��0�fe�q��gOT�U6���� �f��]ۑ���}\���b����:o��ɗ���fb���\�茆�ژ!��Y�x�������P��?8����nch�i"���շP�Άh�'eP{��̻����{8i�wa^�b�qw�vt gls~n�����@�7�JƸգH�_!�����t3�V��Ȏ��T���|������� $ ��r!�8����Y�X��;�7�2W"*���+]�Ի���2������o�P%����C���ҍO���6v��V�)�	����X�$��w�<�l�/�}��h2ǟ����ӛ}�K���	��Ҷ���]�(Wgf������Ѓ�	�zmmu�%T(����F�sY1n�O�+hb$�$Yon�w\2��Y0��r�9������=m��������h$���Ğ+}���ǭk�z�Y��Y�+Ĺ&5P:���H`�%r�|��%�sݛ�t�gw�i㊗��]S�t�B�A�g^M@�'��@T^$�_�l� �x8=�"=M���w�%Z�2�Y/��O۩�'u�:V�2�U8֊���c�v��C[Y���:����0�����Xшo_�������Q��<���Lhܦ$ad�{&���w��E�<��*�!H�u�|�^��M%AH��7gk�8��%{�� �o�̸�)�����	��O�	���	����)���@�����A��A��kD��>�t�m �D��8�A*�m&e�J���<��c��U�I�p'<��]�+�Y.ܤp+����MB��~���=�cN�3�������m\�lkB����W]�ǩ�P`ӼC�gЈVֽ�&���b��p��.�<ߟa�/ۣ�6a� q�L�o�A�L�^t��y~��e���������?B���:��?#;
_NS4{��/)N׫��Sl�f�'M�2�X����<!���ݻ�{�F�W���n�'6՟�����6�̤N��t1h����e�j���^�d�"r`xC=By��K��L|?s�����卟�h�xPuR��r�}��nc�0;Y�m�	!8�A����&���O�ߜ�)x��!2�:������=���7{P-h����bШ�h@41+��	`���}4WF�I��k�!WhS�L���}�9��"v�[��m���Q�6IU�m�gY\CT���ǥ�ĬG�)B�Gs-�D%���єj7������/>a��/�:��uA��
��Y�3`%��Rc_�x�3{��d�Щ�r��p�i�XV,�L�ڨ.�[�n�r0TS���$�'�x�����]�	O��w�\v!�FFDx�^�͂l���|X&N��3���P��^|��؅��:ϑ�\ ������ �Yq���-����q��C�J�z�@�7�+&mk<�e0��~��t!�b.�OY����R�[̘z��p�&}RUm/��ҿh���ߟ��/I��_p3$��#��Z��&'p���ɴz��o�s"�X2�)q��z"O�)�.GP��X)m_+����'G�u*Tŝ�kHҭ��.�mȶ�nX
�gg�P|���,�%:i�.�"����i ���3��qS�W����4�R� �v���esCd�~��w�.��u"�=s��bv�NC�  �s�0e��h��˙g�h�� ���8x*���Ծ	���R׊�5��᭦�{1g�jֿ����_�{�Ǥ'lRc�z�#0-���Q�4�41~��-���)��.��������jFZ}RJuq�L�*`G����Ҫ�Վ���r�J���9�ի�h�������m)b�/u��.�<��6��2�BM��-������s�O���U���~��͙/�dyd-����[�Kq�mXM{Z�/�] 52�"�T��-f�\����J�k�V�k���U ��C88/u�H�Ġ�@��y��n�/��(�Hq�"���ȗY��ea1B�4lOeu�g�kJ����s��͡�8��"�5D�{�����+05�L>M@��Dy�e�l�I
�ȶzw�����A�����a��{o	�=@U'���Sd�^�����ytz_�_����u>̷Iw��mћ��܅
�l9O�sF�����|5�:���	{V豝�A9Z]Pg�{��~�C�Ƴ*������1����3!��(>��S<WcQ+q��c�վ.Cy�qP4.�x��ǈeh^qU��w��Ƀ�a�rN�d\�%�3�D��]��	� �4��fv��E�c��6�^1E��v�	��_�
�@���r��l~��h��{�Ag RP�~'�r��p���1*�W-�/
�(<Ȅ�ʐ~�Bu�켓� ��hx'S��A��6;F�q6�E��>տ�fUZd?z� ���H�E�9,�GE��S��$]/�Wd]z�{��¹��Ju�1�|�9>���U#��E�����?��R!v��%�
ٜ
�hE�"n�漱����5T�-�ٖم�ݮ,)J�ܨ:n��$�A����h������vK��z�GS��+&�J)������z�H�T-�Dج�4��3�LN9�u��`�y�
�>^P<�I&7��/��%:��F#���oɒ#N氎��d�۹Zs>o&�4�#�'A���)�f�*���#<�Ͷ�m�w����?d[���8��ƻ�U�ET��L6�J�D�:go����&��[����(�� �D�E����7�y�P��;�Ks��kn�m�*��r[Q�Q�"dH� ՙ��t�_2*(�:��z�n���B�Qi�N-�;B}�ژ� l0ZVnD)���
ǐ�2����[�;[�E�E�,D�Õr��,�%ܸUx%��&�H��:�e굉������'#�X<�7B2�����R����K�Xoo��&,�T�1(s�<�hM������+W!R�g.:�O���";#o�~ˎ���a<\�{�iP��ś��<3;�:�=��nzg8l�aC8%Z�*�ŠÂ���o�����4�&�·��X�*�㢶B����츉�˧��lo�a:�3 ����T�;�)w��C������R������y���Wg����.�n�&<�u�^���rr���zȕk�8�|S���/�� <�w�L�Y�;ӛZL�)D���k�V�����\������]�I��ӹ0a�t(��\�j!̾��\�x�?�G�i1d�T+(K�<I�,�i��w}���k&G&���P%�D�Z	��5˘�����g4c�<�۔c�;0)S&�K�;�����<���Q��ϻ��ZTt�]j��J���l�}|��\��UC�y�Z[�Kժ!�E�Xhucw4%\2#"Al|��ƀժ�.{���q�L�/E.TC�oI�Z�x�b:UQ�1�!�)�5����DšR�*��_�z��$[�)���M��1n������cbP��4��
h�����V��"ǜ�?}Ǜ���߷ߨb���Ԇ)#���j/�����ٹ.��>�����t����Ƌ���M��V$k։�$[8�#�7YYX�z��q�n��L��Ɵ��.�?��>B���s�8l\ϧX���ZBb�$�]�8T�nLm��'|~?�ʝ�K�����-��������u[�X�6�Y����[��K�m�$)��Ȧ[�'��c��cɬ8f�7A�W^�|��p����?"�WՈ[I�$�2�w3s��a.Xl�u���CPl鍍�[���͂Lf�����Px�Z�������;�4<q(m�o����+��%�w����:T��=�9J�4�[v���@M���Z�<+��#	�Y�\gzj���;��%W�7���v���Z�����gaG
&��o������uo��\�*�Ci�Sd�齅�X�K�x]~�k[Ä�������pa8��'���;����J]`�}pF�$k�aӿ�]�b&j��ZHJ����[�Nj[��{u{����m�s���N�Y��&ݙ��qw���x�2�Ѭ)��W���g1`KzI�-nzX���_N���-�#�?7j`��r�/[�D���\>�u��L�Z�13�o�B�9.���h�4�$i2Y���"�����,C�؉Υ�-"� ����u��p���ꢁ���g@�������۱�`�=I;���&j"����NmJ��am٢�2WP�&gr��#�2�D<j H�(W���B=]��?���Nf����/N;t�"���t�}�tOF`��S�+jRԸ���d��G�����i�H$= %Z�}u{c	M�0];RJzD�<S���u�v�Q~)gʎ`B$��Hf!��+Ֆ^���̠���_=��8ABL���Bq��zb���R�W�rImK��� �WpK �=��c��I$��3��	�Q��_���z5ʥ�4辉@�:,J��'&bY�A`�xr�s��sm�hD�&�+9�O����tk����q����Wr��`~��� X`������֛KS��������������)��ő�x/eV�C+,v� ���*S��yW��<~ �4� ?�$�i�C���V��w��`�����Ub�`������Y�%��}	H6��P����B,"�G6��xW�C����'x�H�T�����e��W�<7T�GN�����'[�caE~Ks�3�JGN��t9���3M�_Ռ�-�y�;o�S�������zC�c"k�%���6� �b�e��x\#�� �q�|��9�s�]��eM�fV�E�/��ą?&s��:U%0Q	e���F'�ڇ��U';�C:+��wބyMy����*Y��|ǫU{L�e�,�9e&�n��«4h�&�4Rݴ��&�K�N.�%�Z2����\،�z4G����lk/V�E��e�s;�
U�����du�`g�sҾ�$�9	\�������beJ�P;ߣ�aml�P�y[�#��������_�a� ��ƶ�s���� ���n�
��	���nҠYD�OY�aM����y���u���>��f<ݽ	N��Y�&�����eq���{���9O����(���&~M�� �Ѓ!��?����*��!Ѷ#��!Q����V�C,H6�7���0]���ϭh�h�c��9���{N����?�����h� �z:57Bb�Dy�D_%�8HB���Ys���ęS[JsY���@A��O�^&�9�+�k���e��(�n߹De!*���-�a��58��:�C�~��p�fiF�1�1�1Cn�������DJ�m!лTWN'�,����8�>���A�
1����c��񥧧��f2����e��I��������"���=��!�� H���=c����rj��,����|6m۰�8!\˱��Zo$�;G9����mmy�cm�^�QgHTxIƕ���N�8	����˭�Uܐ=�N�>le>�|�i�̀�ާtt�x�7�u�<�o�es���"C5>��h�c1"Vo�l|M*��q��wk`Q /-���$�y�w1�@�����Y+��]w/+�� ,��s�׺5)�}5~T�a��i�o��hH����?�b6;���OL��5�|C�i7X�<��Ϩ��<���+?7�kao�`D�)@Խ�ː��l�?׿��G��_֎�A�PAD��Hj�#-��-�xi��3 �'�H�H�Y�-�"b6�y9@��=��zW�A[O����P{f�)���*¯h����3�B٦_)�4/�E2m	?�M2�h�#d♍�L3�����G�7㏕2P~.�3N	E����������ܝ�B�y����yO�TA��z�/&���BP�d���u�;`v_7]|B�I�]8��Xn�2h�87�{݀�%�]#��;�����ʈ�0bA�� ����#i�a���D}?Gћ*ɻ>q4_j��^q!��?n8x;WR�@!o��(��B�Z��hh���_�|��§r�/Y�(\���i|���S#M��5��O#m�@} 
ܠ���E5�������'x��\���'�y��̅y�Ɠ�ѧ��d�>��*���&�Q��tI�_1���3�`;������B(�:Y�P��`�<[�NŘ#Ή(��op��Ѥ�y��M�M%�j�w�Xۘ7֬`����R,���/Uk��0z��?���wD�0�V�~i>�"���/W�S[�?V�DHBzs!��5�(v����\������fDh�PG �������xۙ�����
�WR�+�j ����x�Tt��p/�$���������ĉ��;	j���j �⎸���ƊweI����	��k�X�13�\��ݓ}�
�_w_�����=���HO��m�v-�S�-�U���8I�N�����Ln�
ɭ�s\d�ɸi��`;`�Y[�Gji��ґ5�*��o�!�C��)�������p��a�z�Jز^%ʔ� �� �.��;�X�I�Q`�G
�y*�xf�3B��C��@���%"�<>ܜ���7��MƮ��b]���o�m₌O�<�A�@�g�Z.�u1z�����D�΍�u�S�fo2-���I^�R��t��0��M����8����H��h�ff�8��<�M���"v��Tؠ���f�����z�՘C��Dٟ�xɡ�oe�����paRD��W��1m�����* �k��<�.� �wo��.+03�W���[���bUQ�g��,����T����џ��l�-�+P�	�x�Ar1ЀBc��1���ˏ�wJ�� p�oN9+:@���8��RKbBN7�N+ӿ�crrO��[�=.�w��d(/fj�lV��&X�;�ϱ��ຉ±��@�;�D3Y�bCY�L�)��@Pa��6*�S��[d=#�["���R74�����&�֦$I��1S�d��[7�;t�]t�^��7B ����q��u�N0,KS�\�X�(�8��C�q14�*!�B�^Ϧ�������ę^I�~\,ߦ�Sǀ |,l���[��!��z��[ɲ��JS2��Ԩ���L�x�����6>	;�cYX�S,od�HK�0�i��ᓎ���o�m�Z/�ӻO-f�U�F�c�7m�����	����;YXj�̓(�$���H17���x�ӻG�.��Y_y�vv�	�tww���mrTRFq�+ι��nY�tj�?Ŗ���uY�{砑y�o��6�1��"��5�7#��1Yʴ�	��ϙL�x��+Q��&+��Z���Y�=�3�֖q�K]�*:I�����$!���t�Z(q�oXI�jdB]t�0 "ÛKΊQ߅��	jɐ�>�!Tz���}b�d)�`3�]��m�Łs\��=��=��e��m슧ў�  ��vM��*�Jҧ���'C�y\F��F�*?r9;�uM��I -v��R?Zy�">�IY�s�ʍR�=�-A�<�?ݓ���)�P��vX����{��1x̤j��Z�c&��O��{�j ��c>�4wp����Db�w]~��"�;j4�^��r7W���t:�0@����;y�o�/�xzX«��J�3b�v?�
��Q�^n���8��8  �y作���5H�TT��\U��XNym�3�����k~��ƏwC��J�H�Ny����|�l᪑)�=����'V������ ��^7cI�ǧ#[e��̜�O���!98p� ���欕�`eF��E�Y��z���b7�(�)���1Ż������ԥ�~4�� ��$21{P�[��_=��V_8�������%����#
����b�����3?��.�Ow@�^���H��t�޶��/L
dW���_��I�:��J�.pG�}��`�eQ~3>�/��A���:Y9��a��5q�Lpr��;&U�a�6*����.����a.C	��u�ջ"$3"0�2F Y(.R�^*��;��+�E�h�|��7϶��]-��\y5Iư,O��2F5���"oڶ����P�/����=Ah>�j%��9��
ճ�����T�����C1�31�w����L!�����
l�ɚ&��s��c����R��D�<RS��:�wc������W}�Z�ꊲ�ȁ��>���T���1_�~�w�Db��޹A�v!<TA�,^<E��BF�>ZX5�k�~Cd�Y$�
wÎs
f��&��@v���v��s�� �:�+�Β��,��yw�5�xr��G�a*+.�pZ:�B��/�?"��Ⱥ�F�ۋI�,���xs(�0_J�v��;W�3w�-Y��\����������Opr�Ao����5�čM+�ѯ׵�P�^�i|�puc��VϪ� gd���������-�9��ɗU��0|Co+�b�o�2Avn��ʱ�H�$p���5�w?Ұ�����+�
%3�B�q\i�>�8�@��ꒈ�q��G�N�sYA��5�(�"�Hy��l��Dc������9�b����>b&fT��Ȧ2�C �(��g�	�
%�$�襒��QU��Sد
���K[�a���p(2�gr1 (��z�=�9�Ш��&�H��D1�������-��(�".�ءF�� ˋ�و��S�W�P��������m��N����<u��Wu�x����H��S8D�܏�q�;f6�4�v��հ�uA��%�4%5H"���= y�1���������*����Eo\���uә����I�F4�"�#b�k���,��g�f6?�;U}�j{-�W�� /	�x�P�nĠ�
��n'�+���\J��OQ���q$"��$�S�J�8ƳD���C�. ~�o��$8F#��/r>󞆫�ſ�A��>E�~K�;���&����Q�ꛡ?hq_�~&s$�V��Y�|Q%u�i�B��hM0ۆ��"/Ɛ�O�'=��Եa�I����J�������e��%�ҀH���EM��,/S�?�D���O'�AO��g�h˔4�A�\����Y�b�:'͎����'Lc~�3^�D���G_�����$�v�OC��-�����?���@]"��J��<��A�����q�Ue)s	p�HbԽ��w>Wćf�/�u`�JA[w�o��u�����4�%�#�4�.�RJg�-\/��g�Q��{�|�gTN��[�)�
�MҫA�9	���c�W�zӎڽq'�E;HG01���-���+p{
6$����Wo�:��MF���fv��f�4»Őh!�s�g�A�p�IL���c-u�N�����)X'k�ȖYQ�N����7������7��B���R0z��	�:�8F�o���ԕ�)��keO��ӱ�MV�S>po�/M�J��mJ	(U�ӎi�V�A P�N_i{ �H!A����s�;ć_t<!��ƥJ�3��_.�$����E��:����s>�S��<��+��)�/Ma��{qX�1���e���ڧ��G���.S�>&j"��~[�´L��onYu�n˺SG�0����jG_����+��#����ی��N��t�9����X����k���g�ĳU�we,�ڥ��tM�ӾV�{;+ks`�h�K	?��[�U"u��#| z>6m�}��z�]������)��ltĉ�O��I+t\ac&_W���4��-U/cO�pܜ��U���J��ݸog#=��s�Bh-�(�TyuyS�@��{����BES�l0�9OBPqO�B?���5Kh�n�3��B��Ry���ѴX	�
/���w�VB��"��SY�e���t�8'�UG�I��W
ζ��H������#v%3*�k}n�coO�j�g�*ptTN��"n,�W4_��;bª80������[�D\�$�:��Q0����S w"i�x������]������X�-um �}Ko�P�b7�~�3QY6U���P�z��R����<�U� �)\/K��w�L[}1A��9JM����y����=3������_,�[�#�w�Lm��H�wEiV�8W^	;�2�ն�GN臚f��a�>��(چ	�������'���r��~��I?++����<K>j���O�B}iW&�ڶo)$�|�4�۩�;Š)dc�!�j}�vs����W�U2�=܋$ooL��4��+TΡ,݇eC���|Į�:k�5�I�?���Q��o�� ��ٯi�������g�u�&��՝���cL4���{ն��.n��Z�P�䉨�$�P��vzK�r�D�%��U�f�=�Ps�~0H�?�ԙY�����Ȝ>��#|nh3u)�'u\ד3lr̽��g�n�Z~k� �mrXWtߤg�0�xH�z�w;�7)�+ pIJ��: �e�ypG��޽OI׫�H�\(�'���Ua�S9L����] ��J�o@��
]'��ꊆ��Ǐ�b-D9��~�)
쯝!�D�XM�o�����`o� �b_K�_��=�������NQ/�ڰ��ķ�T*�WS�0�s� |@���Q��T�kTJ�$Tcq�?�����=����S9�Z]�[Ə�����?q�.�%����?�Dwǎ�裏&#�p�F�(_Ck֖R�����9ulv>?��Dh�J*�ї��VBy��>8k��2�N�|���5sf�|���>ӊ�U�.�� >f�u�LW^y9u�O3N��2�F| �"5�a�z��gì7H55u��2������?�T���/���������C�a��.����A��.a�ʕ�F�U����w�Ü�
t�Q���ߓ���./��t�J���~��ʶ�;s?�0d�զA���=���1*�#�1�
�����i(p����������ߗ�)e��c��~�q*-]Cy>����0��Ր�)�z�L�8�y�B���T�R��ǐ��<p5)�*���i��/����P߾}��4z��_��W<�x���P���V]�VZ�t%�0 w�o}M	D3��`fa��ul�[_���<�\�p�$����@�^�CѰJ#��B��Q��������~���|�̥р�}��%ũ���f�z��<��^�֮[Eu5���ϟO�7m���uDF-/�D�FO��/���n]����x�*����Abp|>8v�}�������$(���|p�Y����}��E�6��үi�UL[yL/��w�U�6��y�Q$lq�#p��}z�,Rn����䂿��Rԃ/�U�v��m�/嬟�d-� 6e%b��E�ԱS<�
��x+u�`�r��d�9_�IlH���?�<��xz	�q�i�����oyQ@>T��.@\ȁ	��W]u;s�>7��i�TX؅/YĻ$�#%+��d�jJZ^ڶ��:u)�+����� m޴�����iM��j��ch�"|��5k֌��%%	�*/���ϙ	����M�\{���*]J��EG~F�֮-�Ꚑ]l9@U�:*[W�Lⴶ���4�P�+;Ā���9�1 ��G ���'��'�� �����6��;Z��m��+)T���nZK�C����p�x�h��-4w�����A�!CQ�>�U������j���z���?����W��Fz�����30(���ѣa�E�xS80�z|A2<�o��CǮ�.�3y��(�08�4=L��,�mٲ�����8�^�o�2oPC���1�%�/�0��0 ��\D��y�ƏF�:���ҕ|m���(&-_��j됴.E��A���N��������իv�m]�w N��JQ����W��9�|n޴�^{�E:��)�>Y�a-{ư!(�e�__���	�-���#���C�zı���]���.��
P���JgMǃ���Ac�r�F�֮YF��WR,VE>R�&ȃt��o�<o���~D�5	��۱�0�#0aT4���j�.��K=�#����?�����G���V��+nG��䥗�kdz�s�"�t�T[g�דφU[Q��8�$�[n���)�{��٠[YY�.\��Q�F��(���о�m]t�>˖|I��7?[�N�hU�reo���D�)Z���o;ڴ1D	�K7�p+���y�>���|��t�L?�}l�#p�WΙ9�QW�Ϡ}�G�z�^}�?�����)�{��tđ�r����5�LD�A�QUU-���@���ʫh�I� h�>�(h�6<�r�<��s,y�a��T�38��sU,AL��+3n A^���i$��IR<
�~,~���h���޼�i{e�?����O�K��u�_�=�Ye.@q�Yԛ�C���#x�k��o��ϋ��a;�@:��Q�1��ø��&�
GԾ}7�2�H�D=���6�����2k�!ھ}���;��4v�g�}�����w� u�������|����u�d]s�5�[زq=�{�%<�7u+�H�W,���6;�;*�%h�7�(�C�_������^�3N��y�OӺ5k�8�����r��!�Z?�Pv.��%]L�J����?��:��R�n;U�l�bҜ���i�hݺ
*��Fյ�}ޅ����{���w����d�>x�W^y��}��!0����@rA��u����LI�C��6�	~�@�$D�'�Q�C�(C�> ���K��oSUu��� !=:\���7�J$��������i�?�۴v��'N؟ƌ:H��'b�1�<�����d�Cy��dz�9:���q��H��g猷�z+��C�5ft������4�#���nc��*�B���4�d"BK����D-�UUo�H���>�c	2� ���Bk�ld�m�Y���I��'�y��ѳ�=G���6� ��Fh�$ZG��O��舩G�9g�I5U���I2'�u�z�Ek(/_��HY^
��Q����P^�*9�l�!�4�����p}��]v�et�����T^^��@;�� " ��. �C܋#�2�[층C��WD
zUvB����:� =OЖ���ʸ�����S�~�bfgVt�_�>�Y�q��i��8��<�ݾ��:w�gy�5T1o@����H$T1x�l�k�Oe��y�*� �:�;�<*�ѝz�!��1���#/8}`�=��C.L��O<��:�(���5�T^V��!�����C��C�E/-Y���7�8�|ew�i���胏?�pK��>�x�6��7��ɼQ<�d�w��t�Yg�AÆP,RK�U[��r��8"Q+�d�^Г0�F��H�G�������/���x 9^��	��#!�����R��X���D����M�雯>���j
�}*7�O���─px|D^?8��L���c��/W�w�t_��8`��7�?%���[����U�D�Y!Ês�GdL�rN/x���ٷ� α��T��OU�CN}�ʉ9��g_PM5损~��0�í;|�P'��|0���do���v��`��F�j�����G��W�i�F�rĀM6�~��!�P��9�D����#�������z�x���4���l�>`�lauG�M�<�N;�T�ٳ;��VQ2���3G������CAC8�î۷��	�@�g�[(��u xб#�� T]�u��JE/|�����2�2В�g���i���H�8}-��y��L��iS����T����={��h���>�d�@8)�'ڎ�$H�I�'6��Y�(��2qm��R�Cg$�|�53i�hX�6�PR{�N���R�G���<<�˚�W�ʕ��r]�̰XK��
l�f<�D�Ka�+m�}%�0�2&^)�g��� ��&��NU��ţ!WOD� n��#*�ߏ$��j:��{��, &g�M ��eRׂB:��cXY�=��Gh^)hc�n������!�O;�:u*u�܁�-�џ��L��s���^�U�V����`�׏��Z�1���i᢯�w��[���1��T �G��:��?�A,���S�$vk����*C�eu��WL�,��փ����C��q��m�����x[��o� F�!���oLd�|����|�s޹��c�q�8 �A0 J&����^ �-^�m߾�>s��d\mg�yLQ���@ｿ��a$*A�i���z��co����D{x�n���[��7��&/��A[�L}�	���:�Sg� Ε8e�Ef�.y�)�+I�dao0�C�����p�ް�����"�8O���[{ђ�幄�D�ޭ �,��G�^Y�2�������	��l#3J�F����R; ���<d�a�MR^~'�<�p�/Š(�|\���\1̲8h�w��s�,��j�5���!+�|�|��ǻ�5d�`���0)�>E��	�1�H�_,`�eH�P�����4�7��G��)� �	w�ѣG�ĉӞ8�M�3�H�~�U�Ѕ�ϋ��%D"|=p}��G��(�+��������.��w���3�������z&h��iC�J%��1�DurMP?y�v�F�;�S��Kp��xRe�D\��bٚ�����Y`c����r_�/�#�s�^��8�3W|'Z����8�8Ydd!�׽+�,���@�%ͷ$��;��v�eW�FԂ'�+�"���) �c��[v���󥾄 ��&� iJ�E@[ȿԻ@_�x����kQ�I�O�w�}��_J>3E�D2�>#)�� %y����Qu�h;�б�<� ��GT��~��ڸ��~w�oc+�?��G��]��c��ǜ9s�D��_"��%0����!�"E�eG�>GL�E�@�{,ؒ.�	��
������vR"w�ഖ�6����$��a0 �m�F� gܸ���v���D͐ÿ�b��z+}�����/2^���g��#G�y�����Z��cၫ'4�>"�ҧioJQ�f;��B�(�f?�R���������>��:�*����ۧ��L�j�}t�Z�P�|�  �F.�s�'1r�}��/@+�X��~�i�jc�$x�#�
-����E��sJ2.NyN]C籱�H�~�|J�|�� ��� ���Y}7%�,��]zۤo�|��ޘ빂�|?�To��c���CGR
	�L"V� �RA��ku�\@E�=9
�5}�"N��r���!��&v����O�;�z ����pA�0�y睼c�Dh3�;�v��(�`d�1[�h>X� �ʐ���?\XTpe��i%�������a�hDe~T@Z�dᓉ*�������<0T&����@�2R�"�
�P���q�����s��>���O*߾��"���@����j�"ڼ���*D�f�Fzo�'�d�챐��Ճ���k���K�]c�	}&�4�
`�J&�l�dLu�_^�e�B�H�Ut@����:��6�_�r�����
l��,$2�B�0�E��.� Y�t�^��m���N�Rr�>)D$�+�Q��Y(	}.I���`G����+�0hp�	����G�+���@G�7pu+�G^�H!/��F�n�����;v�	����{��x�ͷ�G�|���#.�����v����(ʉ,��C��O�%d ���� �%��HLͿ�c�\�^�I&\&���ŕ�`�֪��)��,&%2�q����ė��q�G�|��CI�!�i��G�d��8�A2RaZ�v)�Z��k��^Z�v͝�1��*�����5�\ku�d��'ͽ+%� @���g�E ����`ӵ^L^	�G_bl�ѩI�����'=d_
wX�s�w𿠦p}�nF�`<ڀk�}E9�3
 $���e"�c�w�L�_��SG��<�h�����˞���~�/���P�}w����x�V1�Ȅ�X��=���~4��IdQs!Y[�s�X�9p�>���y�F�����@�����[hђ��������@�z!�3(]��t-� n������@d�q�$�t�v?��

��5k��m��9mz��U���f��(���D��\�.����f��Ź�q��`�|�ǵ�L��~�v �>Ĉ�E��^����P���6Њe_S<���@�JK7л�>J�����r�	�plk<��L��"�Z�k�a��h��������ݔ�1������ୁ������v2V� }�<� ��y�E�Ƃ$;H</�{8�%���0�b?��1��)���� &;F�%��*#��L��DD)<��(4rd;O(h3�Aa��]��c��㑘���a�d�v E>�z�J�HE��&��7n�rD���C&<�z�N�(�x�����|ҢD
6b��kp,j���+�p�1��9�}�)]����B�!��E��cA�� :�J�CY�kd�(��nW��1.���"�4�6��5|ݧq��G��k�2x�Q�V_���߲ʋ�&a��	m� �#x?�t��P�����~���?L7�����Q�I(Բn�&zw�'\��4����O��;x��V�G; ~�?�8�O�X���� _{��B�SO=œOvm22Q��Ȯ�>F�$�ɵtZ�Q{�^` Zl��Q�M]�������N���0��er�f'FTD}��w~>����4�u0?�s�[ ��믳���_b��/�g���}�a�~��/~� Bd����K�&��v�(ϔ�=� 8j�6�#����H��b��b�^����P"�����JZ0b�TVM.�J���y~���p+J����g��;{�%R<�.��5�,��GqE����x�]�Г���c�1 S��w��߲����;���`3�ْ��)�.���	��B&���̚� &2���|:_=G�(��|/m�\F>���&����B0ОV�*�y|F�*�컌�?}���&��ښ��<s�L�P�\QO^�LLq)6��	��l��0�Ђ�r����x��y�B mF7,$�uY��#*Z��a�9��LP�"`�äǳ~���gM���y�~�I�&�_D��,���]`����{Pp.�{�M��rr,vx6��xθ&+ v�9�ոq��Ya��������B�+�'��Xu���h��)%�{1���t��jN�fQ2UG�L�'�"�7��OI��ӀA#�������@�s�@6�r?��@�讶>�M<v��s�����D���:N	���j�Yz`ZI�_C�ʋ��>lԁU�vݒ�!��354���y.@9��|�h����w)���D˗~�Y=M�Q���Z���U������k��b1(�8���j�hъ�m}��7�A�`Q���1�-0��Ȑ�K.I�'�Z�,��t(��Ď��������f`��O~����#�0��?b ���3�h x}�_Z!*���\W�S*Z�Î�B�Wp���N`� 9�v�L���n�İ8��x1DPǊh��B9��7�a����]w/��=��=�=�-���P�K�����1���$vK$�h��h"�t�㬷�t��`�R��]8���A���ߟg�tFb7esB�8�9��͝�믲3���z&;  �k�uA0E�[l��ؤ�z�����'m��w�2�]�a�.�������$��t�]u:(� �3�Mhcp	e��j�	Z�b1��[N>�E~o��Q���'��|;���TFY���Ę�4�?s��=�@h��U� S��16���x�@� 8A�������>~�\�VB��K/����cq.���(�@��Y���������_.��_q��)������}�g����TԮh�h@���{���
��BH�,B(����X�d�õ�;Eܐ+�`��n �� �yj�̺�)�@�����Z�\�?���v�x��<i,E�8�c�R�&�׿.gWϣ�:���	�n��~C1�_�{����>����_BpAD��E3�>�3ĉ��XY�Equ��
�~2g��'2��9|�%G�\�	�E��#����%�.=�K��m�����Ȁ6�����	��@�d���b$h��o(T�|��f���]!���\����y�C����O$�5�N %�֚iDO#H�4*�q�k;���KJ� $�;$�B�t�E�@��?!�4=?��#�W>��w��~;����?�1�eq�<�{�w HaW�����ڴi������T���x ��1�(&LH{��>�"�	�h<�	8���L9�98��-�]���s.B.�+D���u`�s�y���E�w4���!�0vM�:�,� ���
�t���	\u���'R4nq�^s����#�3(�?�r��������8�]z]��y���ϐaQ:uW�F4�p�iO�BU�d�}t#��ً6���� ����x��; '~YY~��;�` ��Zj�o�����27    IDAT�(���ƊFԾC7Z_���.+��0"|���߷O۝�u�t�xa ��I18
� @��M��c)�iUF�����uA�����y��ǩg�^�9#�hZ�׿���TPX��x�hh��^�S���c�� ȣ��,V��@����5cG��K ��\�7���6j�Е��5���of�4Y�s�-C�c�wh��E`����i��c��;�B"FmQ��ZN�;~��zVO��f���NЏLJ�$bI�s�.��#�Q )C��<^������b0�/]�2c//ڤ�� �sYGd|:G����~N�aQ��g??��mP�o����P=bm��
t�1�g癑�Y���89'�^U�ro�l����-j�b�0����!�9H��Q�<������˧X"ɉ��O={(͂�����Ř�P
�/솤��h�H�'5@р�����c� ��9@������y�^��c���`���7���� p�\�]Py�߇~�;�@
P�1c�a! �ʽ8��&�馛ҁ� g|�Pa�B�kKIP^Ai�3��#�7d�G���>��)Y$|C6�},hX\�N�+�K���E��}�$^�I�w�﹂��硔!���R��ԑ��d��~��?Ծ]g6�r��]��J��rTSU���s�EC�|�wI:8Ѿ�0"�� �3[�n�'��􀓟�l�d��X(L(�x�`� `�K�-�X�w�q�_�^�8�'&�cnJ�ʕ�i�ܷ�&���~���~;�Y=��mՒϛ��%܏z�(TG��Z/�Ȑ�H�J�ᢿ�cE;�/���>c��!T�ѷX�la=x�Hv�D�\ �C�@Rn�H������q<�����������<�'�P��*<_Q>����Ba1B;�o_\[E�p/����!��RAN�y�� Ա�by�[�v�W_}�89_vI�����F��kz'����sp��D-u��P���k)�qv[D�#�-�z"���ǞH�����s����<~P�w���ڎ�$��9��f��3;�Ocm�!�9�W��u�7I�늑�@��ud�\=ۮ�C��l�d[��~�cF��ɇM��p��l��2�!�xSL	��N��|ݗW�� b��DRɫ�k�Sgٲo��l5�=d%c�1*H�={��\]A�|�5UVE8�F���Ѐ��Ͽ�k����q � ��N:��W=�I4T�%:�b��X4` �5j11ax=�i���L�`��w5vH&���ջ7�
 ��~���.���i��;���ޡEc\Q����y�B������d`�Q]����?��ϋk'vH���(hY���C&���}�;p�0�"�0��XH$L��+�
	@�	H�*�7�<�&����)i�q��.�\V�*e/+�ѣ�҄	�ϓ�?�����~�~k�}ߗtB����� #�ҝaT@@ �E��8��1&�0Bt=���â��d�I��{-�W�V뭻��|���[��Mխ�y[��=�Ou������<���<�͟��T��FƊ6o�b�����X���I2�����=wr"�ց7Y���D,��zW���;�|���^�}_(��yԺ{{�g$Pd(��e�d�+�V�#&)zF<�����k^�j��h��3aae��3�Kֈ��8R鏍��:`���W���F(�`<=�i~29��F��UO�!T�x�N�d�h�\���(|3��Z�r��{�x��6R�K:���z�+(�E���qu���(a��r84�g���\t��y`>_�!��0G6Z�={\�%��G�eB���#�g������B���8�	��^�{�ġ��ݻ����QQ�0i���c��*<'J��SJ
�;4yNA�%��,�Q�<��r���;&B=�p�"dyw| r�J��u���p��5�o �չ��g�^�5�������`==��÷^�͛�{y�L��Ț�綶�V��P�YG�l���W�x��{9���fQ�4{
�~�w��<31/�(>Y��}2���ԟ�w��VB�5�f�:W*�-[�,�xa��T��*���l�����s{)�R���)�q3�f�@,�f������wO��'">���k�m"���m[��*L����X�`�KkU�c�a6/�	�S,�ȨdQ=���D�;^�[�z�N��ju��Y�~��^-Z�����y�sx����6:V�F�bfk׭��+����]ҙM��I�}��#"'\�C?���f2��į����#�F��ɣ�C���@D4��v]�M�0�c����;~��qo�q��C�&@
 ��ً�Z@])E�KX�S�XZ��}Շ�"�uP���(�1��@����n��5{�!͟5��A�4Ԑ�p3���<�G���z���|&a��y۹�^�-�(Y:Y��n��Z��iu�9���q��24Hi�X!����Ü������uA�l,s�k��f�w(a�;�B�e��((���n��;za�cHpO��:���6�4��������mOJ�6��ͥ�^��/���0]3%h�yX�t�z�+��>�D�N�:a<�]ג\���m���U��\�ȑv7á&��DGH��h��Ֆ����p|��Oʢ������n;3�P��\�;��2���}���6:ְF*��TճQ'R�Ǘ�T�̉F�ɘ�zPYߠq�b��`s6������Fи�����/|�A�Z��U>�s�\���ż��������)@���8v�r]���'��7�r�SWh��L����G�#�'a҇
QE�P*�wı�D;()KB�{f�S��¢�^��L�?Z+q�X�X���c�<����>���͋��7_w��_��V�^i54Vr*u�ow�g����~���y���˦)�@?�e��{������b��ɢ��p�ʅ!��S��#���ظ��x�����v�?|�P~��2Q���?�8͙�e�LچG��g����M��K��ƍW��;<�R��U��̳OM�8	:l��z�>�5���w*�_�4k��K읿�v��l�T�a}G{o�J�d�Lڵ���CL[�i�������y\ D� �4
�cҵQ �"I����w���hf����<9筷�;u�ی��H���;`8���q`�[�Ɩ/���|�����7��K^k��y]�	�Xiˊ�bnЖѬ���7�D�G;&��_ו������	�����?����^����-�ͺ����l��:d��r\�[
�h�0��A(.c�x@|�3���'����J
��p��1�x������c	��@���IL�
�M���� ?�O�u�[V��T3���<q�>���5sI%�Z��nW��F/�ݺuvͳ��|�l���dl%��C�8ξ��x~���?��I����eng��f�XC�x�T@ɲc~8�d�ŋ8M{��I{��'m�L��ǜV�g۬X�x�E�����l��%�\����V�Xa�Q�X���i�={�xhh�����dO|��׿��v�O]���~;u�=�k�ϟ�S'�˲�H�ldp���Z笥����c�S�cO��dN���N1�_~4�OZ���:�)�3���#g-�L[&�a==��U��86��&������ݏ-�Ϙ@��1�R��B�㌖̢��������LlEca��b9��7{��; �X�YE-���͋�G��x�?�2�gh�>�`��gº����7���;o������ODٽ�i�7k�����)18�y^����ONe'#9�6 �� �!G�
����B�`)�
�F� ��/��K��M��ۮ�-�iX�D+G�ի7ؚ��Xjxm�l6�a�����yFm���(l�&Nw��F�}"m��G졇�^����J@맪't��uyn�
�U�kTG��w�����J�UR�V-��[�a6^(��c�v����7���$��_��_��u�Ȣf�'.�v�����/6��O|���=�������&����Ä��}���|�b�U��o��/m붫lt����?�ٰ,5AJ劝<~ʆF+6p�lo��o�9@�Z99O�c�������R�?��Y�<f�d�Μ9b�=k��l��Y��?mc�����������㣈*7���`��%rg��s P6'��E3f�J�D��QCu�K��ht<�?�g���#��2��ٖ�[=�h�O�s��#��ޫp�2��١c�����J�'|O��BOhМ�c�	*JH�� @IF���}�"@H�C  ����]@(@��	T��8��|��O*Y��������K�Imݚ�m���,���*�`=_B8�;:]��5�8|Q* ��z�(��o}���X;U�|G()��k��<��J���=k�ʈ5�e�;�g��H,sK2�fǏ��b�aǎ�[��N۾�j��=��<H�G��d�ό�[���������J��{����ۿ�V�n�j�?�h�]���"���b1r �r����<6`��,;|d�6l��)Z%� ڀI��Y3�ACCӜULG��^�÷2^���\�a=={���V#q(�m��� �i�B�2�>�l��e�F�9��h�܌;>8ru�b���,B�(@���d�Q=�lp�)�+ |��;��/��"��=�:B�G����@�a]P3�?4�# �5Ƚ h-B1�.��8�cD9�
e��\�*�rh�q�����p�N���`9p}�'h�XXD�`A�(�(i��fM��B����i��E�D����\�m�Ԯ޵���%��m�u�Zd�_q�Y��J���HeL��'�X�Fl|�>���@1����o���Zd��Ԕ"� _!����c8~h�����l�ڥN=��+ǭ���}
�Z���=쾉ѱ��Z�����wXG�l;yj��z��S��[v�ghx�C�4Қ�+�W?�^/��ݳ���7��y�c�{�4N(5M�mhpغ�{�����c[�&�I�X���h�T=#��DLl68q�ԅ<�ٜ���p���IT=sq�8lgN���[+�[ �筯�k�����sV_ �_�3o��4'8{���Q�)�q%�B�=�*����P. ��������誉
�g� ��C�q�j�ε8O�;�& .JJ�E�9�/�%�&��r�u��T�kI �x�St���C�����uT��5۸����|3��KY�e\�#
�$,a�PO�8��������_*[.�r�/��յҮܴ�2�v��	�C@5��8~|rQ����sv�0A�1��94|�֔2���r�X "ð��������|�6o�`����w����b���B�n�=w�2��v��/7�S�|�
��7R����۩��x����u�݃�C�>��=�6�j����T�f���}��u����^�����6>Vp��d�l���9r�R�Y����bӎ	�gS�� W����H�4�8�S�Ntc�l�yq����D�j'���=�X�FB���Ȓ = ���z���J���X�("�y15-�8z��[�x�d2���_߻�4Τ�,��TV�����k�������Щ�s���y�����M��Rք�		��1���ֈ�wx|�<�YϦ���u�q�[���Tb�����*߅��`_�g:���/Xow�����l��Wx��<�u������k�o���h�r۵�Z��Ky�Wwx{;Ԇ�������D� ������U�ư�H�D��̄�B��88�}��_�(�9sf��C�}L�wTm߾nK����Q+V������jG�#�K�qԺ����En���}�|bhh�7��=&���������w��_����~�N8}�J�b�O��P,ّ��66^���5��ҫܳ���I6�q��MQl/�+���(,���*��'~�^�h��>���O=lgΞ�������:M�H[6�n}GO۷�����,��l���d�ǛX\<�o3� (�T���&i��p	����څ]\"A�^��N�y�ֵqB�-v�K�I�&���h�uX��.V�tr��}	E�85F�v���,l���8��^=ח�YA�r��zg:p��y���m�%�b���'�k���C͈���ވ���uA���n	+Z�Z�(�T��͌U�)�5�~��W[��o�6+�	���x\����#�4�^4���}L�oYc8�J×D>�|'�D�#�����)����b��-����?y̪��[��2/�O&�e�N���K���?d��s���1�����+�_�p��fjI����gQΞ�i�|��l��%�ޖ���_�+�Z�6�_L?�;��Œ�����Ƭ�t����w�㌍I�6&E����LD �S�� ���jT�W+��h�,sm�<qB�9`'Ou��\)xUO�Rx/��}z�>i��,7:�f�r��?tBJR���M���P|����Pb!�zC�V@h;��&�^Cm\�ǉ+�Ix~��f�s��4��u�P#��s����9�/IJ���P�,�����	�PP��-�f�L�j(�4�\;l��K��b��Y�{����3~��8�{����|.e�zɮ�b��ܹ�s`���wȵ�{M���k	[�z�U=�&�}/��I|��>g��/����;��N{�k~ƅyDt1O�����N��O��r�>��}�ha��S	;5pʊ�1�1� �z����q������7~�k](}��G=˻T�|�/��$���w����Ї'���j%�F�[n�����6V�F�h���sV��G!X4s��e��6tn�N��5Kvٛ�����<B�T��E ȓ~Ы�
�:�Y({���I$B�	gQ���*�P��>Lzil�Ν;c�:����Y:8�̒�W��И������k����k�y�8�E�}BS?����� �ٔ5GY��k~*�����E�7�����e�:�����t�/KA>	���-�
QNa$����)ԶC�Z,�@W���JX{du�,�4���JP7[*/U�!�/��kVZ�&�?��7��O9�R�9]Y�;���uG�xT�����Ȗ�x�t�KĹ�X |::���@�D��������O��!��R����������ر�����;2|�
�v�d���7Jʹ��:�y�IK����s{�E�?�V[�d������w����po�
b�^�ɝ�n�����M	���Ă^�|���]�b�ͷbaԆG��#�|����D#2)�eʽ���c��̳k����L2�rl Ջ�!�VzQ�S<p�lZ8B��r�h���6�&����5��g��=K'1�Փ��|QS�0�k��B�H�Y�v�z3��	���"!.�� ���7���4�f�#&ː��<iѡ�>ḇ�G ;-���}�Ly����.��9�C/C�<�eB���Ofq�<�q�Ӹ���BJ(����T�<%��f�n�g�Q�����-�({�Wi|��u5�Q�e"��b�b�sl��^�'s���p$����V-����)��p�b1�Z���C6:%�(#��(!�����[�*6p��>t�N�������6K4�^_��Jf슍[l��U^���@�,�p�M6v�Fc��h�x��TEB\�u�ַ���Fm��.;sf���N�BR�}�Nۺ}�D��K�B���u�?� p|�m���P/��<0�	�ęL($Rǽ�b*��'�}�8���Þ^�j�ly��b��6^�������M ��������{��Es�����oH?4[�=�/� i�D�6-�?3QP:Oc��!@���|�eYH��y�V��]�#��� Y�u��K��*,�&�3�4����v+������m����L����E�H@�X����,YBmh��F��XH�@�.��a����z�T��W�	��I�ܰ�J��[�yKPJ�����w�    IDATa�1�>0p�>��>g�Ҹ+R�Qf�*�K�w%��P���	�ݳ�+�
֖�X__�=���=4���âF�+V���o���̙��B�9��E9tz��gF��n������_�J�WU�Z��Y,�{ӊ��Fn���I;E�0o�Y���p����=���Q�(&���:���P%,TZ�7����T��@�ؖ���5m6ɲ 8@ǿ�~�N��X��=q{:�p���{���=f�c��f�^%��[�bu$$�+�x�>���GH��+c�����;�R���m�N%<D{|��K���t/Γ�PXg���<��s��9�<r�N��J
�yo�y�B���C��g���ZD )�?�~B�*O�
?�'�����][�P��7P��J�D��U��j�T#�?����Ջ�}�e��͖�G�I���w(������1��"�oo���>h�����y�����w� ����16�C�w�hb?��
7V�U��`���J�IgG�G���%'%0%�����xN�9h�o~���v,��%�Qѹ�>3�o�s���{%�D����.�ȭ[7{���~����{z�%HĿ>���.��nB�S-5�&,�E� `A�!J�Ϳ{��y�E�ڏ��T~tޟ�rq@�U���,۾��@�/�z�liZ?&���s��i���R�膜7���K�)�-.nIg9 
9cƀM�u���D?1��Y�*Q�xJ �2��/ R�fb��p"��P�G`c�q<�AT�^c����9��p׆� #ƞg&v���]�~d��X(�D�l5�x�,lz	M6� �g�W�%����[��{�X��D�����pMţ��Y��	���?W���M%
��g,�G�J��%ͼqnX�q$�AIz/]������	O�"ڇz��,А�y^}�&+Ǽ��$v5��'i�5{�]�e�G Q�n^hހ?-�3������w���ٟ?��M���\@��G���}����Ԍ��E����[}	%oԫ�k˻J��7�I%��D}��oG�qw�tTl���,����i��1������+lێ�v�����Ʉ�g�r`ч�t���A�%ٚ$uQ3���L���OD��6��#����[5s����#�m�T��k%��F-���B Q���}}�v���c�굤�]�>���{�.�CI[�j1�� �f �qz!`�v�V$)������a���G13	U�Yuo(�FF%�qŜ�: !ay��l<
�~+͘��l	��������͍�M���4�H ��zTڤ\��}�A�l\(��F.�$�OB��|��'�G�Y�Ō�Z6�.܃�PuX�EX�=nٲş�h
"@�*V$�+�'������Qh��'�źe�B?��Bk�8� Y`<Ϗ��5�j��U�P�0�{'�����&�.��	���Q=���m��N����^�皫7��)ژNd�TnX�m���3w�OC��:��6��j�Q����g����w�����n��V��#ܓcM�?B����߉R�>q�w���Q�Q@j'��")���ɧ��y@�Jd��]��'��L�󟺼CӨi@e�+CVC�c1���dܵxMJ=������I�' P��?�A��{|)S� �0Z�����j���9}�z?g�҈�57sm]v��xTۇ�΀������3/ry�K���j	���Q@���#��	�c��ËEŘQs���%@�	� 4(�����E�y��G�MŘ�`G���G  Ҙ�gxX
�Q����� U�m�|��ا?�ihr4e">���fF � P9���F+$������^]��C  Y�J�`� ̈�WD�.��@E��]��A�I,�Y#�1`iV����r8l��y#f��C�I�����Ġ&e#�;�G�ERm���<�04ɅX-���� ��$�"��*��9����g��zz[6ٰjm̶m��v��̊��FK-a�L���Zn�6l��IZ��Jw�jO�?<;�V�
��}�3 P1o{���C�kpg<QX(�G�&(�ЂcND)�*7�NtR@O�'�1�¨�h��o�u�g���?�#Gd���Z��u՛9_E�4K_-��-@`�g�e��� h��[����W�j�d]�.��������iTk^ҹ��ɉ�nQ3�FT������.3� '�ECcs��Y��� �G?�Q{�k^��-��L�� F�B[D@0/l@�z��Z�	Z�� 	@��Jm ��4rd����c4��kM�b�U���<� �l� �(�v-.B:g>@(����;k�͏@C�N�0@���Z@�G���'
�!T~4��ތ-��&H��d]!����ð`X�|�*���I_c��cҌ	sûBePH��5<7�KDy��"4��v�!�0@h�>܏�X�|Tj�#'���J:������@TϿ��r)�re�vn�ܶo��C����<.���XǬ�6>^�j\ٓ`	�ѕ�j9�ԫ^6����
���}�{<��g�b	a��֩�
�KM	X�5s�5��q�~���w�5�x�}Z,�j���XͿeU�x�B���P (��9�Z1�!'�̿q�����j���aΫQ�%�ܻ�����e��O����Nؓ������rVk�����#66vk��bY�����{�}������VҏLd�l��y�&
�r���D��� � ���1��$�Q�8x�cs"\��;�U?y>,1�h�9�ȓ���Ei�*;V����$n\��h� *-3P�� k �x���������]w�����@�g=�BQ	"@��L�6M�i����]ԑ�5� f���tPj\���E�	���L l�������a�b��bC��@�1N���xƇ���ȉ�����'̎n�W�6О]�$�����L\�?�ߊ����k��+��}�Wk�^j+�\i�:%*���4�N����LD�`&�t�A<V(x�^��GuPذ:��+S�RZ{�#��X(B4��/֏�����G2�5�[v�~Q�\����hIi�k���P�H�7��\
�G��;�1�, ���%��l��ג�M�^AC�ٹ���'�F�>�ԸOؑ�1��MN3��zRҙ���3�p����d��w��0XGP2l*U�d�Uvm ��PѪ��DB�;>|  ;�8�0�k3)���C@��riV�g��M-M�gCp��w�s�� �?��s"��]3��n���~Ο��������D���Y�\��P\��<��E�@��z��"� ��yg���̀���JQG_,,31��5�c�b�7��1�Z���`e�<ļ3�h�X#<��1Y9��J�\ɩ�B���������|�T;�k�F۾�rK����9��z�[��*�6�V�'�A��Z�����#~�<�b���r�|�9ғ���wG�S_|ƞ�fܨ.���|�~��0�K�-�I��!� ��hi����o1N����wF�����#��T!�#�r���Q6���ߘI�\hQ*��h��X
��h���k��7,�6;kǎ����yR�s����3�?�����������F� � ��)9 d��!�D�������C�x @�#xo��c��E�b̠'�ș b +� ;ԉ����� XC�\_�	�q�H�h68���������@��9~�"���t܃ka)��o�[����g�Fk�Fh��:2�� �j��
Nj��x���NW�AG��}�N�O�ϸpm			F���X.�(��@���c2�|x&(N,+Q��������&�d*Z�����q��1���*�^<����F�*6�R[�f�͞���;$29KT�zD�e,��ɦ]������>_�zT���c��T�9U�g�{	נhq�a��K�F0�\Kʢ"�Z�����n���}n�whh�=Sq�tih��Zf��t�Ĥ9M5��|Y ���hB�)'����A��7��ꓨZ�6j��!;s昝8�cV�!�_	�Kz��Ѩ���>4��G������@�KfY; �$�V\04`�JX�M7��9�GÇfPC�8�~E��^6��0�8�c�9�s�����8D���<#߳�)ԇ6�?�v��X�Zͩ�	x�ݰj��p�h�8����K�X��@ A�`=�}�4d=���7�e�@s�R �yg�1��yXT�3�$~���&4 ŸBc��2�9��	�*����!|��4R�C� �emx�z��~48q����2�p✃pVn��k̉O�S���9��Ba7���{���Q+�V����d�ƸY��c�,a��$;q��<���ͷy�;��h�T����;�z�h���P*<4�ֻ��Q�G�:o�@	;�£C�AX���J9l43W�e����{*�,���w�Tܿ��Pp��C�˹����5YD���s4$L~�^���0KT���G�T�eSu��j�&���NB=�����oT�?k��<� ������4PQ5
d18E����� Z'�1c�E�3�aB�) 8R����	x"Դ]4���
d���V���������w<�V�/4�k��b�p=��`m�vۻ��?BI B�{Q����Hy�6c�?�*�8[�l�J��G0����;����F���?A�T���gM3X<�/��cqM���r,ϧh"�Hh�r�ù�0h$�3��
���'��O3��[OOTҹn�y�Z����I��`Z&=�GJ6g�����a)��I���l��g\	#��λ��9ͷS!7:��yY�
"�~������؇�������l���-Xxیl�8�K�ntw�0�q�prB�j�2Y^2��[��8�l<b���h�o�bO?y�x�?qι4�a�nƶ��0���o����ڻl�P����g)�����S	.Z�DHP�Q22��R�o���3����^�"���dI�����cj-M��C�h��+sqmy9�B�D@������~���uq�P*PC�,��D!�y��XD� ����=Ѥ�%ᫌ�Ve�� �;��b�f�xVU��$r=��wFH��ܛkb0g֢��/���a�w#��5˹ⶹ&τ��傠��X��"��S!C���/њ��D�Oe��/Xo�a��?:v֮�z���S�l�0�;�L֪��n�:V�,���WY*M[Ժ��qͭ{�{��G�c��Oi��eh���B!�5�R�C�����R_g�
��֘07��ߕ��
[�y+����U`�s��ܥ}6[�'��,*�k��Z��1���N����A� �w����W-Q/��fuം�,�b%K1��ځ���Ǟ����'}���r����b5s�F�C�$�Yc	8C�����@���Q�ތ!�E�	�7��ax�"M�0И���$ņ|� ж�x�T�.�A̛�6�^f;@Z#<a|j̃���%�Z� �ϵe١y�
�û���������]є��.PK\ޝwCx�[ ��&?m+�֋�5�D�qo�K�1�r@h��:NYuSh��W�.�$j�ga�3P]�{��	�����Ԯ����=�MĚ�y�5� Z�w�*��^�vݼ�&8��+⪞�"9|)��qGj���M�m��+,��z�o�ޒtK���Za�dU/�\�|[�;~=�2���pl�+|��&ٓ<���\�Q�F�	�sQcr��]�5\g���p�$E�_�F�Z���,\����җ��������i��3�,X����Z�)TO&1�b�i*�xX��X��o�y�%幷��l��Bi6�j���h��IFo٪%
WQ�6�`_�elp�`�D�ʕ�,q�˗-�����0�a.tލ�6?!��s -�b��@	`@q��Frt�'����� T�7 e�����+�G<`�#�EH	\4�2�����hL9^��O���1�z�C[���%�U���yމw D�l~�#�����>Pp�D��`�6M�)`������P.��揟 ��Z�̬]�%|%aƅq@�p<�
M�{a����0��<B�s�P�^�R���A�u�_~Q'-@��\<�g�
/�|��D��Mٓ��kE��H��Ymf����)����@�'V�&��HY���\�͊�(@�8>�}F%�P�%ӕ����(2֒
���Pȅ�(�kM��0��f�*��Y����o��o�����ӄzJ"��*�]��f`s�  �]Z�jvȡ�w �4���S�!�P�tp�:F�)a�`���CV),�m�yu�(EͿTI�h�j����3:-_F���.nw9
%д	xW���`C! T�5 ��ln~'�@�)��#��i�r�|4t�08�*<6�~� x.�A~��&����>D�i��W+B-\�7�E�p}�(izh��MJ�뉱A;�U�F�O<�:�j�+34
�B!��/��%�9Z������� 0��DQpO��\0'�cM2����X�#Qb��S~"�p8�ySY
���r�<>#�V Z��h.�d� �~X4��XOO�u�wX�4b�d��U�4<J[��h���g�Ξ��6n�f	�zE���1��eU/��"n�駟}��|ܰڇg�0�����1d����h3�Z�̍���a����1dO�\�l�߳珇�o���+�����ĝ�Q�d^n�^���t%"�́F��l��
ȧ�Ρ���-\2��*ɋ�'��������Z��Z�D լAU�l����g��R#�n�/Yk+�/���HR��q�Ffч�Ei��5#�_��4om
EN��F����Fi�:�ߡ(�#E\pOi[�V�����

-/��d��y|�dѦ���ϵ���s�4QMat����QD��$�Bk��d���T�A��,S���hL�!ϫ,w���3+��Q��9��q_�%��k��Ƶ5��;O�o.�����cL�8�S���s˹�(چu���K�X�:�e��(y��i��;��x�n�V�}��N_�"h�h|3n�}�'#|h4\@Wc+k�C��;�
�C9\�1W=)�%�f�0D`C���A("4�(7~�20�OD{
���Ok���f0����%����:�� *�y4=8LņK L�
56�xa��{�c!���I&jv��S6����esIKԫ��ʣ-:���}灇md���x������5��bT�x்.��ؠŰ��=���yKi�l,�IZNH�79w%�Gi�y���X���ϩ�' �Uǵ��#%ABBڜ�Eq�l��tM"kI� DJ�~���7O���Z���9�g���y<oi��IWֹ�+t�A�r@r��Y'��X1ךC�'Q������ʟZ�Mt��:]�l&a�ڸ��v��tnT"���m�7��-�=�����:w�9��Yq�lt�i�Ko��;~�-���7�4AI���� 1���"k�c�
&V"V��=QG�&(�'(B�>�Kx%`*v�e�o��3	�+76��8��Xf��&4�"M�c�˄�z��8��H��{Q"'ؼd�NI�$��w�#6<|��U4\VQ�p����a����~�
cKg��J8��{��b���N�"�i�r�3C8��j৸T��j�(|�kl�fB�I�� �����p=6����k���mq���G�&��E �@��8_Z��$��>�X��:N�������B@E��}��r_{�IK0!Ƞĸ�4x����(���}=C(�$����$���CKq* �{Pҹ^����aˤ���!�r�z۹�*K6"��)�\�P��l��e�e�.+V�6,��{�&���F�-�?���>h���֬��N�=e������C �J�#c�>Ƿ���^�Z��QLQ4�����/�����>��>�B�>7���v㍯�&<I)�aw>���޼����_h[�l��wy��5�IDy`�� e*����A��c( �*ԓ�t�3v��a;}����/    IDATU�c���(���\~����?e�Σ�Б)�&��K�{}.V��(i���%8F��%zi�i��t!�0�3��K�4���e���I[�!(�u�*�%���s�kB�c�f,����OBCt����9*�gܸ�'�{*��"ǤK��K )�M�U�c��)�� ��Ѹs=	EJ5BY`�B~ 	E�I��&�?/ ������D�oV�M�а7Z&E�fT\.��]�,�d�lպKl���f��&b��'
�������OM�d(�K��d,�ې�Cd��Y��ɾｷ[[[��mY/�|��q{�{߷����o`Ū��;���a�t���Pw�����o�/h�/�����S��K�w���p�l�D�������Ν0h��� �U��⥫�k^i��Q�)�q�L��~E���ӂ���Q{<9�ظ�>��V��&�����f�L�Ϟ�Ç��b��k�C�g+9v���S���;ԓI^5����o^��¢;H��Zn��n|��@Z&?�'p�w�G�d�:�j����- ����F`���l��d�9N���Ӑ��=��7�D\O�o��hQ$�^xvmx	{i�>F��k~�ֈ�AE�	h$T[�~j���� ��.�z&���%�{zڧT�m[/��;6y���r�b�d�.{�.�5w�e3m��ztl�#���z�j5��l�C���Oz�s�LFY�a���5�ߎ+B]�Xw�2BUٕ+�Y�R�Ju�~���l���V��-�H�u��>�.�|�m�~��)A�L�����O#k�g �V��=����F�x	�¼��֭o��
�C66|�N���޽6Vt�ϻ��='�v����+I�;o����q��r�<�f$�[���Ą��O#
ca�
 Ĉ��*�� �Q:e����ؑ笧�+���\&c�|�uw������6�sA& ��F�L�A�����H��}fuF��DE���V�(c#�(cE�	ILQ��W�6E8'@U�i��[�7	ݛ���*��n���s ��Һe��9
r�[�{Y���k&�ώӏ1����y�$넱iV�uC��z���Um�����q�'r���m���M��b�F�/]mk.�ʒ�v+V�^�'�J{/���X�)K�纎2��Iu|�Ɍ;g�KE��z�����{���g���;�����ș�G��{�<�φG�hR��
R���F+���]��M��	+���hѾ�կ{QH��~�VY�/gny��J:k�9O�_�h���i��?��-Y:���<u��e4����ㅪ=�o��������.�p���夝J��-��c��6�8T�>$<v-7w#m�T�����Hة�����,����$g�ݪ��&x~a7�FKs�����'~��S*VX��ЎD��8�\T�����U�� watl������Bg��q�lB2Y	uĤ�C$���$�!JK�ҶC��{`��k���;D�8%�qo���x��Y�8p��O�h�ٯL�� �N�	��O���d.�?Ɓ�2j"ϼ�S�p�a��/O�U�|�R�Nh�����?��zy��;7Z>mV$,�Ҷ᲍�pɥ��tZ�R��D�9���9���s�t2�@Nm'������=���y�X(z	�H��LrY���?�����z�F�O��O���Ҹ;���Kh����6pf�j������b��^����}��H�iB�_�I�t�\�of�aK/�z%��R���'v�+��$M�{�[�i����cG��V����C�e�.O>Bsd�PGF&�f�_��8[4?�<�Wm�B��>��U+	�fR�˖���C���I�T�L۱���f./,��O���0�����O ��fc�H�v-���������C����p�#:I �Xq��0����>e�)����x^�&d]s�� �ʼV�l�"2b���z>6*N8������%�9aA"�W6̝�"	LDl��u��I��Z��#��x���A[�j�+!X'T�Ĺ��#������Ci�G4�L�LK����C3�-�.�]�l�|�zѬZ��K����vX:�?8��Rz��>$|�͒Q ��4��mDh�];=�\�H�#Ɏ5E2�Ah������.��w����_�����C����s>�POc����{�::�ّ��v�ƭ�����^��pw����:u©ח5�Iv�-{��l�X�W<Bf�ʕ�[��[�j��ࡽ��w��j�g�8��&�D=i�#E;q���>=G���;<}���Ԣ�
�(��d����pO��� A{�yal-�z��&��l�'{��@��=s܋Y	Eu�W�OU����1���S�S��r˥���Xp���h9�È�j6象<���pp��.�(�' ��LZ���'��0��"��|
��tE�.��JHK�秢v�`��D5���`�����/x6�9��<6w��-A��P�L��\_���A����~e"�MO$��:�*�#~r�>ƃ���ь�������j�yrc\Փ6�1��s	��kǕv�5��j��UzZ����m��E���T�?�ō[-f#'>%! tJ�D4e5Ŝ��F�&un#󙪬R�Kb�c��.�?5��Wl��ˬ���{�.���3Y2���S,�j��g�-����;u��M�pj���!�
�̥}��d�F�%[�z�}���3�(��O����W_����w�5��d"c�C;v�U*i�>�?Z��o��J��|���J3FC����/�뿣ɲ��rQw��k�^.���3���g���&�!��N�[w�@Tҹ���Z�Z�}�����Lg"39t���+����dI�h�	GlowNt��elr�)�S� L�LS�js��M��B�@��	L������|<;N;@\8s��]Ř�;����u�������Z|8��9�g���|hͷB?�t��Vu=5�x'��8`��6

�$�D� "N���-���pή��*۱s���-���IZ��0Kϲ��V���Kl����9&��F"�0S	s�k4�.ؙk����	س~Y��]��Z�R@�,��s���y���X.��cǎ����HФ�ܡ�G����ђ}��`���V��Mh���
��8c�8NG��,��d�:�������u��/~���~��2;ܽ��Q�=��C�#v��	�V3�w|Զn��5 �^�E#'��@���h������{7'�ςB�g���� ��M�$��lh�%%�g^��z$��������X�Ƒ�nk��ˋ����
� J}�G�$�86�\��X8/��:G�XDu�0�Rܚ���<�� :�%���c<�7?
J�P��&��͇&L������A�����q��=T���/D8V��!U'+�9���ޔ��܇�D$�p9�~Rl�|#����(�-�$�Ph���z��Λ�q�;
��}�9��7�у��
�]�H��
��$jhZڇ�==n��#v��+lێ+�Ny�l5/�l�U�d���]`۶�Z�J�9�T�lg�J���|��]wOXz�e�4��p��)�֨ΊR��l�)|Sp�(}}{��o�/��ʵ.zz��Z�!�����Xɞ}%`����Y���5��5�N��v������T�`����f.�3|�!��-g����ys�X�������֯_i�cC6<�OF�����;f����l�n~ÿuPB�S
�pO@�C��P,V��͌_Gi�L.jD.���E��M�qPKT���'�H�~k�S�d�3}]�E�I�[O7���9�����Y��<_��W-�kw�zʣi�_�-Y��n�G&Q|7��MC���p���h'~2n}��@��]�M!�F�6 ,�	�Bgr�+�J4WsC.�6s#*Fs�d(9�$�(d��z:j���J��C�b�K����8yk���߻��.�8ʹ�����.�}>@��%��`�'�7�}��1��_�mۖKm�+<�'A�;B=3yk��l�P�9�ث^�+)~����~b�� ��wMT��C2( ��)�>�$��K��`�}�"a�(
��=��7��3ms�̲��38m��y���#�ldt��O���ڛ�g^{�7�yv�>/��E,+�e�o�
�U�L��J���M7��n���f��k�#�$h�,K�?[�9WΟ�S�m���������S>�Z`�q�UE8A�
y9���'��aѱ8�j[��U+E�7��P�8bV/Fez)��ى���s�mx��>�锭\�ܖ-_9�����_�� ��r�~�~�ߏŷ|�R���W��Lԯ��"�І� �z~�w~�#��}����&���f�`m�	�6�h� +?Q>h�,|��\���&��1/8e��XlR����1�jnx6Υ.��k hb|$4$,ࢱ��D��I��d��q�a����PH�Ї�}�O�����w�r5xq+%Vx?�k��1�k�߈�Q<7�w�>����V�h�t�๰4�o���PP�;���M�>�a�C�#Ը?����Z
��x�� ʵ'�L�v���lTҙz�����_��.�b�7=�륚�sY+��R���ZmX�FV��Q �RX8��t
�>N�5���N�@7���ظ+����cL3醝���s'm��Y�JH������1��=f#�{ǯ���`����}��}Oa�Lc�-X��/���|�L��9u'�F�J�Zd��Kv���/���6����s��SO��J�FTK"E�� �,�]���;V�dTT���Z�1�p���lf���" �=�7��b8�y�RqI�L1���U\@5j�*{�?B�\%3��,w����96^"d�b��|��X��
�޴���}b�R�ģ~�	���t�Zf��t����h��i�X�� �u����ȣ�� (m@J��!c��� 8����В�3�X���&��y�&>;Pо8_t�TH�iL��9<#�}�K_�,����0f�a9`��� �`��B@vZ.�l��=�Ԧ�	�L	`ʈ`Ma8��J�v��: J�φ�2�D�!�yg������.X���˚�3�Y�Șk��z�|x�3���5��FR��Nh#��yg�@�E��q
�yE��T�a�^��d����d�$�����V�|J2ac�g-�M[��4��z"��(K��-�J�*�/{�$<q��dv��T����xG�Sy:�8S�R�(41�˹0d�iPT��[W{�|�z���(�uKeӖMe�\%���i۸y��[{�c4�_�K�7���Tz��;s�����}ph�]2��xs��HZ%n�<>:�����z{���R������������������a�V��׾�&K��zł����U'���bƹ�4���'N�t�s�� :6��<�q�8M��mu�?q܎�v�?�%��:��L��600l�t���B�
��X��J��:c+�'��;�t$!pQ�����fuL4� \٬$_1ԭ��"d�D��%2�1@�ط�9S(>*��;0�h4"���k<_���ƕ1Ҹ�a��3��x�d��0[��b�)�E�C��*j&`I�c�I`�d/4Hx`@��[h�p�1T�7���������h��8����XB����.�hu�s�?����ܯ",5y8�G��p-|Mh�{� `�����u m�lƁ�&8l� jd4Z�\�5�����>��D�0F��%P憹b-  ����IP������V}��k�9s;�R������V'E��t�=�6o�f�k�v�Xs)��	�60?�G>�)�(�x�b����%HY袁yO�x�޵Ò����{�g�'�ǎۙsg<�c��Ev٥���l��n��Dʾ�������}��E=^�IF`:����|AΛ=+���|s]w�5�������>�4�����uk-QoX�3~�644�?4�o��f��h�y�r�ı���h"^����ب��	��ھ瞴3T�L�,��Y�R�Q���t��C'�������^��s�-[���5#��Bm������,b�n"�`D''�l��e3�b����Ip��Izcs#h ����3O=�&36r��9��	P#�µxv	�x������2��46-V
�E�/Z4��D�V�GQ�G�]�[�/�����y��Ra�� �x���&ƀ����# T�z�k@��X^��>�4��LX_<'�������1h����'?� @#��C�@� �8�Ʉv��������Zg�c�Ag�8?� gm�[�_��`�P��(@�o|��'�SZE�fj����P��>�4���2|�N�@��֟���x��/Xb7��j#i��:���eg|[<t&���½h�B�19�qd3��#ㄦ��\'�(w�wݾu��!��(<pp�����  W�Zg�]�622f�]�큇h��W~�H�L�3��۪�{�0�h"Ж	�$������WU�^6��ѱ1���v���kAl��,Jܒ��F�q|��؀���������`)@�xDJKͿb��>j���d��5~*�B��l��=���=aC�t����YV����ޭ48����Dҙ��>���'lvx�
`ġ���O�k_�:s���׿�5��W^���F������.n���ccqc(�l,
�b�� ���>�FT�]���VZ/�B�)�/�e�h]���Q��SҘ�8t?~z</c�,nE��,<?�����C <�ll| Dƒ{2�h��?����k ё�aJ��̀P�3�!<?���&c�u��6�;� J����F9��`y�����8Xdj􂠅��:P�Xm����{� ?]�L������"�Zh���t_j_U��^����Y&I^J�Ն%3Y�d�FƊ6{�|���<0�.x(:XfШ�?�K��p_�v�ڭ�[@�yG��S�>���������׽��8j���A��j7�(a�"s�\�H��������w��Q$*�MHw�O��(�\🦍#`Ƅ���h���h�L�Wl�-���Ƥ�_D�@E� �*�M���j`�"�p�hЄ=)a���Xm~�v��ΗҎqJڧbGz���'���4�Q�!w�&��p�){��O��%�;�Z��V�p�GV�T�?�@ |�cI{g��n�J���=������G�,Z;|�-������Zԓ�?1�)��q��c P�u@T%m�t�����"���wm8�ņ��A�0�r��@��.aYO�<��q�D�@�BQ>ʁ�'�O�K�s \z�AK���|���s�m���#��oG��G�=���Z�ǃ����f�l�a��5�X�PwX�� �h���g�0( �\���u�څ�йV�� �=��P�Ϛ�jb,v��I�'��xX>Z��͍����f��;��{�r٤U��z�z۱k�%�eW�Ru =m�ɜG�\�y�ժIKeڼZ�C����G���}��_�E��G>2��b|�g,w���*ժ��,T栽c�]q�+�b^�v��x��G�`V�Ç{���r
S��N�
��gl��t�>��,2@�	Ne��F�*e�1Z8v���j�}#��бǩK��Y���9j "�z�$XR��?Q�BB%�[q����lxp�FGO���i�}(E��s�Ġ}�[߷ᡒ�ۢ"j ��UK]�F�i��cݐ�Ef#-���/~8e�Xo_�or4B4M VM�т�� 6���骫� �	�-	m<�m��;(��h�|�8��8��^e���f���]������N�7�6�W%P��`g�a�+GA�E�T\�(#9|�;�׀��g�~�%�)*��b�������}��|:
c	��Ppli<*�O
��u�������r����sq_���ZQ�@�J���zrT+(��eMqM��g�r��8^TG���O��Zͽ~j>� ��)3|[��v�����
۱sS��e\#�?a]]�mΜ%��5�/Yn�z����?�L�ӗ+��>�G���E@~�w����)J C�bY����)6R��1    IDAT�gfnU�;��f�%B�#b�����K/qg��X��A7��SKD��{ǭWy&/:���?s���;��/Ȓ����'���ظ�e�У�^�s/��p
K)Ւ4���b6�������ܤ~�m��T��tf!Q�`J�oDF_[&�)�=m�O1_'���#>n?�d��H[�T�K.Ygk�E叧4�X�{ m���F�n�3.�0��~�X�[Ex�A�Y�߷ϳzh9,l�� F@���G����E�1D}��|������A�I!P,a�Q	�ph> j�N,5Ȁ�����>����.�ڝ|xfq���tM����a�����W�ʩ-��+?s� exVh�2��zr����"����uO�����&|P�z��»�""�k=N����h}��� <�ƃ}��%�����; ��<�s4��/^Ѥ���h���)+m˖vݵ���;!��x�ƆKw��+�^��;��A���{�tųR܍����r�{��`3� (���r�χ��KOF9@h��e�q~'�8B���3I�����"��C��7�֚d�f.��t�Ʋ4�x�ġ�?��g�b�4C���D9hCiSPd�@5@6/+��s�펅%z�Ο�:U��H#JZ:��.^�D���{��g��+Ke�Xo�I{��ld���Od@�l�b��}����X;:�"!��c����B��[�0�<!nJ�
5}Ox�{Ȇ�����������T�V�-����t�{7PÇ�P����59_�V������\�MO�)`h*��s��
 6�j&XQE����_�U6�m��6��::8Xq,����/��}�����d��<q�>��(×���d�9j�� )�IYq�d�/��V��l�R�uJ_e����q�6I�����]�=Y3�j$0���Q9q4�tsnTc���3��?O��1g�k�{p��-{n�����`���y�����y�'6������U(  ������
����� ��V��  	N��h��4�G�U[.e4j:v�:�Uk�3���}���>j#cD-D%�q��\N8be��Sq����.���=����*m�����݉R�g����N��V�2^i���xL N�WtL�M�gCX�D_ hy �)�ĵp�J���j� /Z8<59��f���¢t\_�S?��'���%�-����Z 2
��jG7�waX_3�s���]iU
�ў1�
��ϛ����q�Į�f�%K%jV+���ˮ���7Z�Ay��[���(�V�|�#8{�O�O�uwT�5��=���DAE&)���Y?-�gk#0�YPJG���r|�N���Kj���{�ǳ��<ON硝�x ��O@��������ln�"�Z/덨�U˦y��uz�z�z/�l�͝�ǎ���<�Hk��zfŲ�����2�3n�ieq�}�t ��C/8��Ǌ��Xw�j���CZd�I���55�ԊQ��6���e��qܪ�W�O4x��AX�i�xm��F���vQ/� @j
�ć�Q�ZΓ6�spO��p�S��X�PS�<�P�#P>|G�?�1 b�1;��$!p��_�z�mW����N^���-���s�c�ev�u[�V-X�Q�J�jK���U�l����6^�z���N�d���8%ӨW�?������#���M�ɨ��9�J� �&-�����?�9�?���5��[&�:U&B0���⣨Y�1��)Z�`�B ��p���BH��o� ַ`c#gll쌝�?aC�#�6�JS5Ǝ�L�?U>�5����eQ�H�M��3�ȑXuax6��lt>ߩ&>�X��H�
Xm(ƀ(�ƈ�_Xn��f;P��G2!�d��A�uE����	��P�#A��ɠ%f��!�SA7q圏��kh�xo板au����;B��@Ӈ7��z��Kr�	Łkആ�x1�J?�B����ի�z�o������`==�Q���]��J۹�
�L:a�j�R�v[��޽Q�\M�jn@����I�әk8�H�'��"��d�b��6�<Z&�|�=�|�%��.�{wk�֙��/!p���:�VB<�ł���'��3)� 4�?_�����R? ��؉���@�Ɔ���G%_R�6;�7`߾��Z�����4�˗��ZםJ��Z �@,*%0�|h�Ӂ/K5R�m�iu>����ب	�H�Nw�l��ę�6���G�����P���gW�>�V�6�=t�J���S��r�</s�ld���Y x�Y�sg<%��.�v�۸/V � �Q��t��O"�_ Z����45p��9y��7�|��X#�s�e�u˥V��{�b�����*ik��U=���*��oo��J������׵�����r�7�H)�\���i�_�������6p���!�4���F�hB#�nr�'�جh�a�n����q��4K�-�"Sr��������8j�Ҙe3˥��]�;�w̱#����S�BUh�+����ΪY��C3BP >��je��8N�p I9V�ĮPs
AZ!��C�C�V��i��DA���y���ID*a ���E�*�F��(,������~;��k����s���������_/�!�}Ё!�F�^����?����ʃ�k�`~�����\��������f��A۵�J���͖JT�FD1�n�u��x�f͚g�]�j-�-��p��{�R�'��:�%I����)�p�7��LE�|&���[S>��(��S8|��帝��A�C�h�>��Xlbi~�z�@��V��^{Ķ��mլK�g��Jy������j%��LZ[{��}��~�)�4)V�I�'��B�Oʣ�������y~�a�TdC�Zn�y*�G �	7�+Q�l�i$����xEIp�q�M�Lo�O<t�4q<����&��$_ׄz�2�Г%#�E� �*�;��է`)�@�yF`p}��*Ĕ��0���r��B	��@l���.8|U�'������s4pﵜ[ӣ��o߶��ch�J8��Ixe�f�����M�Z�Y"�v�8U]��'�G=�{/�]ȘJ�z��T�P$T@��iGd����i�}��}�����00��(�	���&�\0	/c�jz�5e9��kG��d�h��h:m��wl�*�#F��$��g�R6{����B��J�l6��˩'ν0�������J�*��c�㈆�����w�C�1/p��7p� z�(+��8���y*#	���&�Fq�Y(Jl��⚊D�#Y��r$��g�A&6�|���0�H���r�9��W9�0�D������h��=�x��(r-j���h�{?�E�,���Y���,�oV+Y�2�Y�:,��rw��/V�\JX���L�ݪ��er9+�"���~~0j����z�S����d�˼`�[����jg4�O�O&_��f����K��f�vv���8<<��ZWW�'Zș'`�����W�� /i��AܫUy?-{��{�"�4j$$%��5��.�'��L�#3e�j�8Y%���w`���ݿO����
��^@4�v���4v� E,)��r%1�/JbGCb���K���`��wfgg��������~��eؙ!�/��s]{�Ιs��y��������4�dh:wx��܇���K��s��P����9�D���}�)��H֬\�bi�RP�UK��̯Y5V���M-�m��,;P�Z,i�x�^ۇ�<�\32���*cS�L���W��/t"4`��ɣ:�.0���
:=��9��������Z���}F��?�����2|�s %-%_{{���'�oނ��h�bkjn�b�`'QX�����>셖��Z��mJ#`�ʙ��D��~�]1�p�Q����G���?������Xv���ɘ�ke��b:�����%;|�۲y4#:=Ǽ�ϼ���/����E�PE�g}�$�h<<H A�?yF�=z���q��#f���>5/�]�	�36y�Xˤ(�V��Y�,f�B��?�.��f�B3���h���O����G��?~ꖺ�&�!�o~�o��@���������&3]rT���j����cC����Δ�o�׎>f�==~��Jf7π�?|.�?yʤ�x�?=t���f.$q�������
d�-[�£+H�bQ�z�=�ڹB*�&�v��qkۿ����7<2m=��"�H�!,��pp�*� �?8OTI�7}�fC^��}ʶkףv�s���ojL8�{נXʒ�&۹����v;q�ߒ�Fw`�@�3;������q��#N'���E��f�Q:�
N�@[I8�
���
�g���
�7=Ŀ�ᛈ�l����v�RkH�;|I��KY�T�ɓf؆�[��D�56��8�b��e�X���S��)E��:F�i��!AHTAx.o)�''>�/k�3?c�L��!������d>�
�B�f��zh�}��o�B`�ވ����G+�f͂������R{�e/{��$9�6V�y�R�d���8���9,�xZ���X��O</U��%�0d�ǆ�4.��i�z���ݹ���>dU��J��V��KZ:�b:���������[��٩�ٳ��O{J	�����U�S��M�ld���#����B��X�N��u��7aȹ�>Gg�4���RD���5�ym3���c�u�e&��S}�y�_d�
��)��i�4y��=4��t`8�u���J,@��<���=���(�¿r��J����`-#jzz�F���������>�;u*�&�yt�����G+�K:"Mq�^��^��ߴ�&
d嬘�z�*Ijjij�~!�7�_o�c�Y�q�;R�i��z7����&Fm_lJ�aB�9��C� 0�}�$�{��>��������:h��)��oHc�P,Y:�jm{=%ɋ����-��>8|�?R�/B���Ĵ��8�t�OC�ۢQ;Q�����}��Ϲa�7��S��$��F��ty���+�T�ui��5�wcV,e��u�57�؊U�,f��Oo(�G�m�稱��~��?��p�(@�ƴ'e����Om��Paޣ���D}g���%���T �����jժ-\�ȦO�i�M�J7xe�}m쓟�����Y�q�uV�>[�m�����Z�
�8aV������������y;�^{��?��J�R�FsC�]�b��^w����$�P7 T�=��s#D�j�rS㇘a�ˡ����|caRu2Z�-/|ڱJѱ���tٱcv�H��v����Z,D, ��=�e��+���T���s��
#�w`c)5D/����y�_�.~_a�}E��2Z��#�����xN��������>/�y�J+��M'�&mN-=�V��d�w�
eknj�dH�:d�!�1V���GA��د��Z��l��	����G��?�yg�r-��|[6��B~����:w����}���㌍�0�^��ټ�����Ŋ��=�ȣv��
�CB��.�?i��t�m�������xOo�ug��B�Rɸ���/�+.����Az觶{ד�L%,�ΈU���ռ�ґ�ݶh�{�^7�%J�I��ۭ�B곐�T�;������g�d|l��r�$��/@����U*v��k߷ݣH�u���{��6�CcOz�r���>Ϥ��(6>�����ƣ�Ȅ	�|N��Tq���F>/:8j	����C���b�97�g��v��\�_m�<`kW�g7���d�j�l��O�j�nt��n2��3C"��D@!��By�������
�l�r[�q��� ��@�6
UpaB&|���|�j�(��jκ�qő���sߙ�6;r䘭]���ѓ���n��K_��=��9�i_^�u���oV	�ل���}�-[z��
v�}w۬����T�:�a�R�q�%�iJ��;U�W��k��/>��� �$qू#� :,�Ph����8�}Ī)K�O5k�N򪞅b�'�466[[�A�����=A��@�ޣ�����o�z��$y1.�K'�W��;�E4u��te��2�yM�bcC�\�9{�e����h��%���=6X�9�ۜ�X��6oZm�*��kV+Vm��%6k�*+V�V.��Z����ӂ�G�� ���G�b�[�ƌku*�� �3�u!���T�_�?e?8�rΎ����`:;;,I+�xh��Y=|����g-�/����fϙg�x���;�5(���>g��m��zz�����[�O�<���G�q���������9z��zp����w[��#�y$kK��R��Z��7�<�4C�P��B��ҡ�����]��<l$6E�p��覧�l�z��b�͚�v�H������}��W,a�;�����S{��X���i��U��x�Ё�+_��]r�e~ppӺ񢋶�&�l���/�9�a��&�.=CY�r����-�0�c�S���+���˸�r.��Z~*�B�V�a-���/�t4F[y
��U����������*�Aa���>����4�Ud-���I�ɀ��i�pMeG�*(�.c>�x����E!ߌ�M~�9�����-ާ�E)K����՞Pb��
���p�O/���f�b۲e�U�}�L&,^1�>k��Y��*��b���:=s= ��Y苡�B�����2&���y[�]�W�������N$��O'?U��_�����'��&Nh�	�Z��=���Y�6Y6W��;;�RK�ɓ��v����rNM�O�3�x�VXt�G��,�}F�PՒE�?w�]�u���>�����]v�k=R���C����fX2��S������i��q�V������R�'�:��fs���OO������'�����r Y�7kH&,��Y�������;݁��4���uڽ�?d�\���Й����z���ꆍJF�a���osС�O6��m��^@G/V�OMz� ��9P��<(<T�) ��-0侀���h"m|���(�34�@ 
K5v�q+��ļh��V�ͅP�ƨ�`	�A�Q�ƭ�b͇~�<J H��Ґ?�s0^�c� ��:�� ��
�1N֌9�s\�N��t�%��4]���ֽ���u��C���D��*�%�,0"�O�흼���7sQ'���%��X��+ϳ͛WY��o���e?a��]��;y�����/��͵r������~��)g��⋼�<?
g�fCP��৒��g����}������ov�sm⤱�c�ϭR����l�v�9`k�����\���B�x�����=%S=j���Y���>���[���v��U��@�}�߰�/�`�X�����p���Y;r�U*��v�5L96:�ޮ�_�MMo>� @�����}׭��8��u UR*��%gt��J�����}����SGͪ��h0��X۳'8|��g.�����!�s�h(��h'����c��<c�={���;<�B~�֕$�ѺR�BQmz(�I��(xHs�ʀ��F#�� �� �!��Um 	"��Lt�+�O���{�nc0	��J{H *������q�"� �p��B�u��2~=�,�cM�^�F[����?�HT�%��c�\SV��������e�N8��p���u����+��P�!��6�X�p����o�8�4i>��x�ɚ�L�ISfz#u2���N�C��g7̅yt������-1�G��G�O�'���g�+�K�X��ڳ�q{��o�ʕ�l��V۽g��$��Rͪ��=���4���'\���
�U�yٮ={�'����G2Z��Po1X�{�����?�^�ɪ��>�����L}���'��[.�#]�A�G��ѡ��,"�J
�PP��8|��l43q�j���<b�o�`:~f�OX�T�LC4�x���i��費�}����&�T 5�3O�����P�\�4s���6���^�!�P9\�k�6����0c#���)o,�|G7�6�4h��@F�q�'j�*�,��QPR䖛�ޗ9lE*�vQ�d���
n����S��PU�b�    IDAT ƳH;}$@�΅��h.���q�
�|J�������o�;���X��yn�8lֆ=�ƪ����T9������2�%$������{�{G�uGC�����z�۴q��q$��|�X"�%�s��G�<�"�z�,I"g-D��kh��]]��=�Wu@��8;�[@YC�!H�f��e��٥p=����<��~������ĉ���m��KE�R��lޏ��w���2������A�����mFֽ��9��w�?�GkK����&O��η�n�S��Nul��D���T�:1`��d��/��^�җ:xP����o���'u����$�:����k�7��m�ڑ��<h����&;S��//��'�#��,�Y*�|$�D�G�9��I^ݧr�L�X�Z���9�3�|��_���_��_ٛ��&[�|���b��Ǒ��9��	~e/+�M�T4ę�( �
�J���h��p@�4K��z��4z(��c�gS�(W/*Jܺ@?��.!%zHt��*����BF 
�3o�>�����{�y�% ��2�����.�2�c�ŵ٫p�\KN%D͝Nn,��O ���Y@Q?E�ϴF<�z\h=�N�g��O�{�f�qo�N��WY<^�r)��=e�c��/k�c&��/~��*���O�;�D�P�+����i*���Y"�A��F�'��g��|,<�����8��}�~t�]6}�8ki�XGg�ˑ�PW(�~�C��ȱS���o/x���+�\j'Or���/|�N��v��|�V�YL�����&�P�xʶn��^|٥��sº�:�����8y�ʕ�%q+{S���c);~�{���&�_��5N�pҹ��ˁ���~���XhWl2{��A�_u���=Z��r6ƦM�BM��7<C$y��8j�	�$k�JIgw8�c�δ؎���;��;g�t�K��S�'1�#w�Ղ�O�UW]��� @���w���C{��"��j���E]��1����-��0�QJCܺ�n6���Ґ��^`!MYZ��q�9�w�;E��q�v���ʚ�`":F<u��$Ǯ��k���`�~Y%|�W�bQ;r���FAC�X��`3$��0c�,9��ή]�|��@�{I(���[ȱ�Ϩ7��G�,YC�LtMt]~
�7/��:�|:"��×f.O�}��_��Ų���CSC�J�|�y��Y������V/�\)ǩ�˜�7n�;~�~����zg�@߲�?�я:��<+����}h��h�����u���u�ú���l�+������	;��k:�X_o�^�����f�2v���; ��*hρ�(�݈v�I3���׿�Z�Ҿ:�ڮ�OZo�)KRʙ�o޹'i�J�j��󗬶+��!��D�s�{�8�}� ő�/��O��/��n��&w&�Y�!g�{��(�U����W�R�Y:�D2f�b�R�F+Wv�D���5wX[,f��p`f>��>h+��7�!lj����r�']�|�;��!��gy@���A�C[=r9(ꔅ	ˋM�5ѐY>��h�(�A���|>�;c D!�!�9�X�+g��|0���5U���" Y'����Su��S*Ғ�{��)J�uHj͹�"���s-�s͘��s4K5|ѳȂ���]�z���&\�R"��s��PEX���H�p]�IT����v(9o͙�>��Ng�)A��D��(E!���8�-K��J`�4E��.�8�O���~)�L��榘�C�D�O���|�i��U��(�@Ѵ�eZ\�O{�>��+���A�_��Я���(+KJ�g���I<���jլ���i���Y6G���G�Bɚ[-�/{��qc'��������;��A��3ٔf6jU�xh�H]Up��ۅm�9�j�����O~�#;��a�b�-�;ޖ/_a��l�Y�X_߀o��[�V�?8|�q�I����?���]w���x<l��f�\(���G�;�k���Y���T�fU��d��h?GtO�,��д"�$V%���U=�|F�d<�&Z?4����N>�ʳ~�S��tTϏ��\2� �Ќ �K@�"��B`��}��ph�'�y8�&�$� ,�.-|$��0�9��LBp��"hq���c�)��cf��G)cz��\�3�G �<��3���Ҁ&���V}���K^����p/��K#`"K.v�ʘ��ʕ+]��pD������sM9b�����d���5t$��{�;�\��9���5`mn|�y�����x������e�l�B���`�����݊�8|�	��˖0�Eђ���b�X�
Ţ+J�Z�&O�i˖��J~?�%�I���Wc#M[ʮ����u@�'�����W5n	tYV�=B��[�E��ﲥK���wn�n��~;~�;�)�BH�̙sl�ʵ^h2F��Z��o_��/��t��s��!0Z=6�Lu~�u��i�F����Bo�́�����k�X�&L�ds��3/�M$~,�& ��X���ȍh�lG�I�r/�o��o�q*�tp�}v=�����I�Y�R�)B��ԩ�=��V��_f��˂�l��V.#��8��WB	�fӽ�5�sڈ��9�����;�0ǯ�إ_��W�Y8�D(���@���>g�|�+�
 ӵk�:� ��CMH�A�O^UNB�+�xrσ%G����kD�5k�g��0gPvX)j�~�m�����6w��hx$��A�%�C�@C� \\��B����"��p=���q}� ��? ��e O(@+ׄ˿���z���گ9@�RB��<@�#��Bp���[n���F�+���A(�,W, ��A,� ��]����g��,��3��E���������}rMX#� ���`��=4[��ૈ�D�)�oO�2|G���[8o�-]�Ъ%:��=I���R�f3gͷ+.�;W�����)錒�X����=uʱ��y�E���u���/�gy�����\�
�8C	y�k_m��u��\(�Ѯ�v�P�𠱡�.\lc�O򂊍MM��?�/�v�ϕ�h�轢��^�4����$+��~P.��W��!�6��M�ߟ�����������?~Jq�lT6?}aqS1�
�\���_�ʠ�)� ��X`��\|z���_�O<hǺ�[KC�J���ͦ�Ix�۾}�=��G<f�B�C�jη���
����C����׿Ձ�g��׾fO<�sOhan���@q��!����t8�� _��v��)�2�4y@Q��p,�\��ܓ���'�=�y�s� ��.�`ܙ�\�w�֭x �	5B��9����T�y��b�/�uh0ƈ?��lXH 4���S L�}XX '�A���l�F�'���	��!8s�<#τpŢ �����ٯP��9����y�#�*G�o��o�}X։�@�s/�k�6�����,����1�&�N�}Ü�̿���ꂛy欈Fb��'�)����f�G��h��v4���Ϫ��m�ƕN��I_��j�wĬ�e��]�Ɋ%B&���|ɝ��7�C�;��n�[��H�?a�$Wz��ST${�3L�?���Žy�W��J�9a�Xߋ�Jy��Q(S��[=���;��g�5g=��h�6W������ji��0O��!�K���D�������^�>��x*�>��'o;w��~��v����2�i�p�ho�xh��o��MZ �D����}?�
��hh�̑���l���Б���Ү%KŃ�_���j���{~�����=�B E����B��ac��‿�s����::� P|ի^b�=�<�����h� 0g^8$r2����a����G ˈ�Vh�h��6 
��ÆF����%�!�   <րC��"Дo�sO�t@��v�o4~�eВ0P0��� P�V��r`�,��5f�h�h̀>ό���	B >�3�@�4N��5��'�)$F� ��AX"�����Cb1�>�����D�p},&����A�#�{"`���9�^��.�'����#9��� b�y&4c��Dp` h�OΎ"�$ ���;|)�P,���5K<cߪy���Z�a'�P�z���u[,�i�r��u'�' ����?�1����,�ٳ�z�7�6���|�c�R�ϣ\$@�yϿ�.ܼ��iTidM�p��v%�$Mŭ�ʺ�w&!pVW��b�����y�p�O��Or>�is�Nu�9cƌ�C���lX���~Sf�Y��ϡ��&����CE���� ���Pa��4��p�n�R�֒9oP�]���x� �}8�2��,^|�M�>���G��PB[�N���k|�2'X��O��2�(���������{ #a��|̫,$@����3�I��������Ƽ1���
���so��f
�:tȅ��ڱ�rJs]@���1���9�p#���c�q�C�kG���P"$������=� �'����~ m��S��Oh�B����F�h�PiD�(D���[).�`yp=��8q�<��ڡ�h�X8�)��E�@��B8 �/��s!�z���j��=Þ�o�`�Z@X#@x&�-
7)oӦΪG��9ڇ�ΔQ�$����R�Z��W5|l)��B��1c'�KVX2�h��R�Wt���op���|��.(YC����}���d�27��!�."���f���`��R����B��X����ΰ�E���Z<a}�Hk�^g5�_~�����j8�?�$�v�"M<�B!;�~����t�oEˤ��TZ��B��_��_��Dy��C��h�����-�q"z-�x����U=���Wky+�؞}O؉c�,ӀI�������j�,�ޤ�+$y-�3��V��h�?�q�$y�I�1 �}�� D��PCc( Q�Y/Om����������I����Y��]�Ce�2��e�?�C�p� �	x�
#�@c:s���4n@P�|O��1&��[�L�#��z ���@`��h��A	N\�ﲏ?ό Ch�>��2V���%��7�G��X�D�H��3
I�E� <PMF@]{T,4�dyvE�)Z�9�|ȷ�ȗ(��'�s�gB�����{�L�nY����O�����5��zl��e�y�*���Z�jD�4�،����ɳ����C����k�t���y�5��S�7��>*���<ɡ�{�_�A� �a>�'='ק�K�ۛ���!D���+,s�9E���r�����2���=|�]񩞞�7�nB����Oo4B:}����K[?8�нG���f�)'���q���9�8���X@1���5�{���G�R�Ǣ����s���ai	�fh��n��v��S������>ف��b�:�/�&R	����11^LN�����(h�������"��?h/4>Q��h��1�����%=��b�a��
	�o
)0E�ֈ��'�(��Xt��U�d�H�(�C�T+�� `|Ou\��>�Z��\GQR$����r=��M֤"�؛\K�+t�g��*���r�!���e�!D���h�|NJ��#d���?`�gEI��<p-��n���:��b%p�}��i����y����}�+�АIX!�m�/�u�.���_�ڤI��${*=�jP<��;�G��@�<ɋ�?
������8�U	���U���B��u���@���38���8��h>���i���@Q��4�)�&_{��f�������I�����fU̓<�0s��җP1����7eZ���wP�OA�
�xk4A8Mi8�������>��G>2�@h���*�v&��"a)KZ���L�b]'xI�b)�<���?l���'^�ڧR�;(�R��p�����p�vc����b>p�AO *  �Qx
��ϡBbJ����7�����[U�l\��aN�	3~Ɔ���@B���u|�4~w��+|
��;��X�@��*?@Bٰ��W������)M�����ݮ��{K8z_龾A_��q�����T��br�	�
G2t����N��!����G�Gs%��s�̫���{�4����SF5SM!Q�Q�$���[��8^`k�,�t�jTM�C���KmּU��W���d2�)-$t��hL{G0��sS��O����� e_�w�5�Y��`-�|� <j�� �J�=���u���zC�
�J���B)���z�s��f��m�>�����3j�5����^���
~BX.FA������]*�tS�8yN�IT�d� Lp�*(Հ���o�;~0U����UճZ���=Cq7�>5J0c2;z�ö?��� ��2����{?[�D�����/tǫk6�vc�\�y�X4�F�I|���s�� � Z<�,��CX��@ �
�s/zB�%��i�:P�'�4DJ�LS~���e�&d�E�1i_|A��4Ƭ���"��rUn�������wyN�/��Z�l��D�B��A�/E���" x�Q8���e �������J���a˜��+!-Ag���|f(x�<����tV��Z�B�������B��p���S$'g�-�իϳT�j�R�
��-\����_c�J�2���C�Fē�z��Ԩr>��W/G(Z=��,Z��!�'�H�#��u��ϧS��T=��s���)�����M'�<�s��030�'b�$n�
�w+�/�ԁ{+�U�6�{��O&��4�W��{�ő&�CqzA��E��u���ٗJƬ�����s�>q�k�P��H���G��w�o�Y��]F�9#��� �5�����s�n��R������C��� �04�Q���H?��<#��sv�P:�kp �� ��f�=_A��m�T���z)dt@��ӜųhW�\h[6�6����)U-�j�9�۬��󗢇�r���p,|����`�̠q�T�,�`�?���*��n��di5fBR�W�> i�I�=�B��C�����ʭ����y�p��B�	� n�bg����!rE�* ;!��<�B�������H&��c6 �?�hrI��a^����:���O�c�d/�J��il����=���
�PŇ����_d�f�䅹;r���ND�?��NJ]*�ϸ���,����m �_ڰ��у�\�g�5��'����/�n~6?�pc{��O�R��{�nظ�jeJ9Sч�кcl�����:ަL�a��YS�8/�\Ĳ��W�lx@������9T`�4{�9�S�Ƈ�#�NTD�<gIB9��"r�T>���Z
V�5����OX�<��?i�|��>;t.��s���?^�`�U}�tTN�`~�<��S�.y%P��K�e�e�G�;�F�Y��l�-( 'Ǐ�P�UG�v�P���u�I��Q�J՚[&؞������C=�	Vb68�PO|u�p$�!$��5�\��Q矿���0�I�����""H�h��Eل����^��p�b=Ȁ;�q�z4ƿ����* I^O�����C3�zd�mӆl�����ސ�X�HDƊ嘍i�`7]h�<�C��*UK%3�h@��$�|��A�od�K(��ɏ�)�Q���N)5�y�B('Ih!h!j$�ǕM|�жi�Џ�7p?K�$��J<���3A�NXA�w��\� ��0�j$�}���$�37�k#̐�I��Åz�����G�\���7�-V/�[�O�l��'��{�%�S�&.�g͘�tV�p�����f�����t�+��ꡉ8��w��ͳ@-��I�l���<�8;�� 9N�{�����ϥy*�?��C �vklHY6�m�V/���ά��(
"� �X��Ŋ�3Ѷ\x���!L
�'I^|	�-�s�\�5��;���9O�����ij�e��+��R*{���	-G4}�ߛ0�&�:�O�2�/����{�i��D�T��o�+�����'/� ~P���N�B�#a!� J�@��G�'`K4�����B�CT$o�    IDAT=��5f8��'Z�����UK���֫Ikk?b?r��z�I�}p�͟;��1�	�EG�F���ybŊP'��@<8B�������AU/�+��{.��sm��טkY�RZ��ϵg��2���O=,r����CU�T�,ޒ-^0Ӗ-_d��P�Y2��`
��?�2��l����b��/& V ���_��C�dE��E�I�Q��a��b�!(T%����G
������������ng�O=���n���:���$/xp�RK�)�Q��G�"qy)|���(� Z@��(���Ђ밍�Y)"M�Q/�ŦË�
��[�Zo�I/�L�(�&V�ZKZS�D��/x�z�@%[�p�͟7+d�B�h�K8y\�<�-�08^�|@�':ģ�Ik
��B�P�gb=���2fEJ�Sʌ�tT���2��8Nk�Q�9���:���Z�2��%S+�<d���P���Lc�%S���<�*U��:�� �zb� /�y��Y⥈,�a���5�.U��AqW����x(9%"���g���K0傥����O�4����G+�P����h�l�F��S�jH���-t�pnii�E�e��,�;�vR�66��uF�5��Q�o�j�x�I]���v's��}m�����>K��?Md���d�}y�1�'��Λ�%��//�k8�G\����o
܉���\����X1��p4ro����}�=���ϊ��"�c~Jy��U3�O�����>��t�Ϥ�V*g��9f-�)�2�+18�A��ĩ�f�z���cA�S�z
0τ�=�aťpVi�Hi��E�D�Jm(d�L��ǒ��CkS��\�ԦN�l���>Ι��<�4�87	���{��4N�R���U���b��v���`��fO�m��_�9�f�E���MJ��kRH������?�I�#�H�����iq��+��n�,�pm�6Q��?b��<i�l�e�^�ө�QJ�'v�c]����gΜn��~�3F�	��|.�WQp�����_q�K9���@��p��B�3�����g����w�OQi���?3�s>���:E�-=��Z���� �C5Oj����9k�]z鋽�o2I&P�p���!ڇr�p�(e仼���p�3�T�q�?����G��	�$'f��6�lkl�0���X�ʢ{���?�'�[���B�D����Io9+9��K:WC&/N�J(�If���+^�r�0n�s}D��S�N��\2�0Ƕo��}l	o��%�dh�
� ~�EI�UGvM�̹t���JV�^��b%۽�!��M�Ȃ��|�7N�f�ut���&%~��U��G (!e$�׭e�~&?E�Q|%J��Z��
@8ʔU���� ��Q2���
�hR
�>�@�E���~r�X�6�(��CNa�<��!�\���F����I�o9�d��}�C�+�\t"�a���C��d9�"HX#Y����"K�<������h�g.f�]�|*��퓴B�7�wX�ܬ��n+W,��X-�h�bŒ���[(a!�����;`�&ݟu���6Dӕ�^���W؟�ٟ�Y�B�zq~ɘ�ҭjT)L�(��m��\��Ək�=��'�0c%8�����;�)���`��fa+4t����Z����ꎢX�3M~�_do|�묥�1X�>|�v<��u>hM�F�=w��w��:e�KUK�3��J-6
�!P�v=un���S%�M�g�?��O�#�xp�>��{��ah_�x�v�z�N�8`�B֒�%c���IKc�x۳��{߃6�������i>2����hN!*~�vv�u�ɆV�3�B��E	I@ոK��(� �����åB����G�5%PD��k1&e�J�]	/�[��響�
�IX*ƛ��B�{�:�k�\OUe��7����s�R��e)Ei���sܛ�Y��ҳ�7����SB����5�	�_O��~�O��P�t*f�B�mް��o\a�b�ҙ8ͳ<ο/�9�Z[�ٺ�<ڇ��yXl,P���Tۇ�Y{���k�[�盽�P�-@(P��o��"�٦t���Y�\�\��k����<��,��#X�����^!V�>�
�P�`}O�'M�r�Y�u�֛�{z�=S���$��y\�)S�7_�*����V-Yϩ���#?�'�|�Nv���f���/�bp�]�l��^��#` �������
�S_���ԽA�!���fΞ�%��4
�C� 7R�'����	�9u�N�<l�~zc�V�X�XC�kk;����Bm�~(��}��3X��Z�lF6;σp �pg�R߈�a�J�^�q�?'�U�+����Ł�����Ɛud>)��f�9c�GF��!sH����q]擒J����z|���N�Q�D �_�� �}d���&L|�^�ʳ�ٽ�AV�E�����B�j��{��� �oX�� sĵm|Iܟ�9撹C9�w�&*/j�L�2�+�j�x�$.�mP�_�Ϟ�<�G�����S�e�r[�a�U����$�����i6a���I�@��垓!䓤O/R*�y�k��G)�����y6�d��A������#�@Nb)3�I���K����{�b��{m����s�c�굶v�&���%�Le�;��fh���BEÿ��ugga��[?���s�3|��aH� ݛ�'o|�l����kk�i?{�^���MQ�b�jI�!�j��_�%KWٺ���9����}����)�P�p��+��~͵oqI ��<hm�G���zmr�U�=�޶ݎ>�!��$2�&ۻ�34sɖ�ݤ�ϬuW����q �ď?��mkmE����u��9�S8(<֍�u@�������=���T����>�`��6�8�i��e� ~��O:�p㾔� �ɑ@s�z����cԴᙼ�s<X`���Yփ}��!�(W�㟱"����������C�s;�^MI���O>Z!�{�Y�ʝ�	z=pO�hQJ��_��"�3.������X�p�wXc�\��&h �%�����5#y��O-�b��3|�}⵼��x�fM-m���6v�T��˚�.�֡�C2c���,}~9��\������;n�Az#�����9�;��B��#���<��`A�R�q�i{�ч��'wG�1�K���z�5���V*�l` g���?��Q3�a�
��{����m���~8�w����Z�Z�7��Ͱj�h�>���������`��KK���w>W���S��_��lŮz�[h �]9�2���� ��y�k�>��O;� ro��M�D�i�=(���?Z��Uc�I&,�(Y���־o��j%�P��\��G���)�?!��_�X-�FJ��� 	��j��@?�Y^��KD��h�<� g�	 ����e��?��?�k|��?�/�@�i:z���ŢMQ�N�� ��V��F��É��`.Y�@G.�=�3`]L�:Ʌ%�)����\��hX.T'eLX>T[���vN�̯��9�K�y���?�k����;4|@��`�ױ�G��P�Mj!!d�/h@ ����{D�QdA�r�
?t"�E��BbL������g�UF�}���)�`���Z��֭_j����9#0n��l����a�Q!��]h��D�F1���:0f�����Vk<eͭ-���WzIg�?���X��a�{�ö�\>�O2Q�#��m�欄<u�{C�|��kv���,�����~�-Xx�o��|ͅ>��|RZ�(�svk���?� �i��ٟ�ɻ��a��}��ٺ˭Z�Z[�.���]��Y���v����f�tۖ���9|�2aY�K_[�G( 	��}�{���ń�۶�,@��06�\ФG�},n�Z�j�y��v�X��k{�
���
�����q����M� -6�G4?ټ<�f6���ƾ�-Fh�@�2ln9����̛@t��j)@{�'?�@e�5Lj5�ȸ/��T��µ��i<���+!r��E�s��d��C��-娱�кyV��5�y��_�6���ͅ@���u~��<��'w� �U����b>���p=,�xz#�Rv���c��+Wz�4�{
���PE�!X<(X!������e/1G졨������ь��?���D�V.[`�6,��J/x�����Y�-o�V��{�s��sJ�y=�9m'=������s~ޒ�}��wT�,`����+�	�|��{��߶���)T�N���o,�Z��}V*Ǭ�x��ʥ/�K.y��3����ӳ�i�r���=��붭���a8��DC�9m��p���J��:q�~��o��e�������ug��R�ӝ����l����6w�b�r��g��jY|�EW�q�U���e 0���"� �5����DȌ�Ex&E���:����y�
�~�E��D������i�_����
�D�'��.~_��&��w�.PD���`i^�3���IVh�h����g�xa#<�3 >��(�CA3Ѷ��];��� ���}����چ��h� ����}$˫\)�8xa�߸?��3X*_�Hx�G�((��K_�VԞ��#�lX(T<廔�� ��Iz%�	j@����}�.όe�����)8�y߳k��=#�g>��\ ���G�T�'�Wq��zU�P�'I!�ꀭ]u��߰�҉�F#��Y���u�H4[�d0�Xܳ� tѢ�&g�g~���>Ŋ͘5ӕ��v�g�Q|��P|�s��_؋�S�'��c?�x�-_��&�c;v�E%�$䥬�7k��t���v�D����`���w{%�#�N:%�s{h�?^��?��������y��m7�`�I۷�q��[_����V.�Yǁ=�M�S����Z��C��ڎ��KVx�T �k�Q���w%�GQ��b��C�븃D����>�P�3 "pJV�����Nkk{Ҋ�^knL{)j�留�}Z_��`i��l��YV�~$�a�W\?T�ҥ��8>����^��Q�]8oh4_�X>80�<��&�"(&N��3�	���C� � f��C �e_s�N��v��2� &����ϐ�?��$3��j�O�<���������G�:S��b]� о�7_��^1����h�?/�A�#��cg~^��K��_��S��茙�&X!(<B Z뭩�ѝ��
A�傰Ta����������B�Y�*���N^T�ݸn�mش�j��OTi��V��9K��������4y5\b�CE�������hwkݣ},a�}�����7��)^�q,a�S�	5��X~"�9�(��{����a�2�8q����J�Q�L�-�-��]m^|��'g=}y����ߚ[�Y.[��|�c�Ѿo���9��O/�r�Gz�{�:��_�7
Y8���Ʒ��g���v�7���������|X�j%i}�y��+���w���e���Fʣ��������B��h� #��Vv����v���@�T��/9w��y��;rp���V��Rλ6���X�ہC��{�L�LC�
Xϛ7'���k����+�ꪩ�%����'������n�Mp�j<�g����;��w�P���] ���,%4o�V�Z"�`'�1 ,C�i�p�{�X�y��o��8��>%�X#iϬ-�`�<�Ȝ�7Y�'�{X>�=����>��<3���������+��F�0G(���w�� �N��Rr��ޔ^{I���B�OE�9R�آԠr:Ȣ B(�i�U	��8�D���c�#fӽ�?�\���(���O���[�fm�ʅ�y�*K'jV,����V($��a���0�����uʜתa�]!����٩>4�P2� ~ᅛ}MX�T�jemI�"�G�����??w�z�~t�7lŊ�6}�T{��G�Z�'/h���,�h��G���d�'n�L�����ܳg��&���ׯC���_����~�<�d��Fx������w��55��Z�ٿ��?�E�-m�W����!y���~��~�ʵ�=^��.�
�L6a]8�?��X�K.��M4/�M��p-]��7����nΣQ@���Wԑ�{T�|�������U�$%��*W�6n�4{��6��COZ_o1����m��6w������r�у��P̊� j��U恟�gW��*��h�\W	[��G��F���j��\ �\��o�D%W)�_��Z����
��}�[���9�џ�R�38e�)7@m�J@SG�~݋uT8��y�3��5ŕG�A֏��T)�?��b�?p�T��	�g!c�9�H$���O�mUP�/�BC׋�c��14���H,,�:y͝��N^�5���Ջm��%��o����:M�ן�1�&��~�R���{��J=�'a1����[�p�Z�I�я~�[�2.|?(������s*kN������g��g����1}�577Z{�^��(��T�1{�g;-�i��ǻmݺ�쥿��Ǝ�d�v����S�N�?���[g/��F�`�1aM��r�6[�v��,���ʀuu:���]����J7ہ���y脝8U�����\�����)�8����H���щ���ܻ��ݩ*f�/��hn�t���Ås�}�N�Q��s�
�>76���L|�����x؎�pb��Ϝ19�i�*pÃ?�*�#�s���f-j`E3�=Z�Rq *��<)��M���P�: #Z/��?@(�s}����=s����氢a�!�=�/�&��X
<#���+ˁ{�ys}�+��s�;�Sy�ų�󀇚�3V�����%$��3�¼���{pO�Y;w˴�V�,��ʭ���7��2��J�����ESro������i�E�:�Z�(���~	����?w�i��U<�w��́���W,؆u���-k���'E���%l�l���j�/Xn�\Ś[�?�Y�����[��Af���!jg�	��Z��BAOr�yvĬ7c���p��+���'-��B1�:�3ꊱ�-�c��?o?��Þ�՛�����S��w�|F����l@��Q�&O��K�����N�b�8�P<ekW���\s�UJ9+���c�#��Ȟ�ŇO��	ո�eK�(���.X������㧲K�����+�� �N��p��׹�@4�����pM����f6���-�g�'��b�ϓ�0)S�9�{o�=�}��lt��l���6s�3JZ�� ��p�0Y�d�8q�/���9p�lv�`����������9<�CB� �t��	��3C����4Y�(������*x2��a�������<BN<�����rc\|�5b�rƁPC�#�/������@ �(�7~|!̓'dM��kϸ���S��d�TB�H�W�>�a~� "�D@/��f�j�0�`��٫Ap�7et�������b��,C	,��>�KSԂ��W�N��ГV++Hc~
��4�o��L��^[�`�-[���P�������y���<j�B��O�����ʁ��k���k�Tj;g��r�-!(�=�S�e��Q��3�l��U�}�־�������',CK�B?��ez��6o���n�fkjn�����˭_�g��%dߟ�Uo�r����+>������8O�f�KUZj�<���T�����~��ֶw�e�h	w�,�`��۰��;���,.�@4HT{��%��F� ��c��M�1݋E�� ��!���>�i؃A5���=�i�|����!b�b�s�X���V,�(ڢ��'���5�>h�42�q��
-��w�r�g(0E���n����K4Q4~g���l�� a�1�e�XHD�`#�=959��4s��7�a0�����D�0��:"��y;D��	��B���p����0v7B�8k��e�#܈���K4 �{�
 �m���5'��H/�V���A� ��׮Q!5��8h��J��u�Þ�E�;�'_�T��@;���ח��U��5foHj�D���	0G�}$��\��=b    IDATG�ߟ1mz��{���������T�p���^��S�*�����z�2��6~�Tki�h�}Yo�B�x�O����H�T��Q�z��#��"�e@ԗ(4YF(6��Z�`Ǐ�����ܹ�:vX:�r��YҦO�iny�-Z��b�����/~�KFU"�Fz���?ra7B�b�@��@s������:�?g�d{h�`'O��G:�6q�T�>m���0�
� �qڢՉ{�@�9d ����w~�@�8��� p�1�f��gpͬ}�>{�G�����U�9�N��Œ�u"g���x��*U"�ʶh��={�����5���c�U��o��Vki��I���p��Y �Z᪀. �Q�A��{r��	r� ��L��;L�� �ѦBݓfP"bEEf1���y��Qr��/͔�� >�q�L|r-7���C# ̱$�=������N4"< |�|��)��%�M��~��pX�V���yf��1��x��rҨ����s�8\W&�0峚	)-eq�Q�_�蜨�XV��Y~}G�CV\0�0	Y.<{��s�����P��7�v<Q���36ab�ūeKg���L�<O�P*ٔi���/���4��>�XҊ����T"��n�5��jj����'c�p�����|D��(�2��o�iӧXKK�u�:aǎ���9y��Ek���lμ��L|���;v�W��ekko�Ʀ��p����+F,�������F�m��������
[�t���9-^E����꤀S��O#Z�*5ʉ���&�Xt�.g`А(���녺�.p y��H��fO>��>��V�D�f2�Gi"���\���{к{�Pn�g�3g�͙=}��	��4���Bp�]]�|��PG�k�dx�MJ�����? bM �p��������NT��ׅ���a�p1.���4l~b����.f6�:V �6��pFx`�Y�ϸ� �p����j��u$�@���s*�-���`a<<'�\�
Q_�����-%�ː=��QA8��9a��o9��KQ�;�ы�����×����t~2�*�w&�"�)?�׿�w��`���'F�[J���p ���,
�u�{3f̪w�:s=��\�ٚU�m�U�<x��$Z��^7a�]��_�^M�c��A��),2�����@_���;�|=�?�>�x�;˺D��x֐u�|�+��+�!(����l��M[[�z�Fj��FX�߼�۱�I����G�p���)��;+�}Fn悃,t��@�ĭ��j�9k�4��.��6n\ocƵ���d/c��'�w�s�k�Q�5�Iy��k��B:|0�OM��W��8sB=���u}��V��;~f'�z;G��	�DXa2����~���!��@ uP��ϡ�H�l^�3P&���}�k_qpE�E��	��xf��d0��M����{�s���3��X U ��2P$� n~"��_���9��\��.L�Do0� >Z5c"��sPX ��'z�g����7�@p���\!w�5�8�@�E�>'���Rh����>� �b`��;�[�M�	��H/�.�0@��v�sF�xi�cBԌ�'��Ⱥ�x�τP�rGi��>e,������ʘk���sO���@��B���I{e(D�?�$�,
B�4iJ��^�?�N��n��ev�5���Z*�L"c�r��u]�w6v��Z��� F!�Y:�`U��jN�p^?����A��NJFdh��V2�{��nͣ,){P��]�K�㖑Q��]I?X1w~�N;x�@(��sX��b���j�Z�2i�gea���8R�#����K�ZM��%�Ny	 b�d?y�7���{,]o����,8��& ���������h��f`S����7Ra7�:�&>}�����FS���������?��T�
�!�J:��q�9G+��a'�u��� �E��3*MV5  ��\xm �a�E����y�&��� ���=�@�= D�����YE�p-�V��=s��m�{@�0���	���,kD�Q2�@�]����@P��C �yc�h�(? !��"���hrMb��h�0i�\��M"�9�惤D%�y< s�P&"�u�>\ۭ�tz����9o��~/�c����S�eNX�B�����J��ҳ�I � Z�5�%��q�?�f.���[�������X������R5�i+T����-8υ���i�BD�"�����7�)��66X���^����U��^�0?��^��b��;��Y�g��:8�<�´������Dw��U�EK%C2�sWü��[�ʒ����C<�)�t}ʋ��J)$	ł��� ��kj�;:,J:�	p���x�l���z�'k�U�������$�z̳�?��R��d����;R� ��4s�8
�s�eL�P���b�n�*iH�N �h��zդgNWϼ�.�Xڧ�4F��84�����gĽ2~Ơh �3�7��6�h�pW��r�	+��9S�-�仌��Sa��}$�枊����O8a,H����9�F)���h?��C�� �&;���yQq!���^e}��e���~��{�}�s/|-�e�K��B`" �h7o?�:%X��	+,�#�	�G`�Z`/Θ>�����!bi(��鞵5+��u�\9Jz�k"��է��isl���ij���B�l�J���S�롞��>p��Y���&R)+�r�V�/��5V������"��(b�>7D#y�!�h�4��M��j}\X�����b�����}����
fR�%;���j{��zCo���A
>��,H����^r�Ձ֏���D��P�#��'�[>4OBBh�7O�<�����{n��y��r�R�c���p��u�k���g�?��q��(ِ��IA���<��m��1f7��|q�q�r^lz�I�աW��(��p99��:5�L9�&����j��:�-�V��Ys>/�Ut
ϫ{i��$%����D"m�46�����N}nDo(�����XO��G�W���}�;4Hi�DXae<���^��1 HZXS�?�+�Nܓy��}�53��דlV ����ʇ`]��_���,�:8ЙX}�M��O�0Ux(�+����^�2�X�X�Z(�i�C�W�����ﭽ��~���v�4ѨkV)V��e�-Y��2c=��.^iώ�z
����	sa���ߛ��S��\�W�d͘/�rg:���9��N���+8X ^&\��H4�Z�{^<h>�P���(�;��=�L�� u͟�^�����Hl0�������F�_�%^��A��g8DD�l��B��Y" ������ 	������w���Y��S�*a��G��͜5���B�؀����w� /LH�=���V4:>�Ӕ�D�h�p�p4H9���B��h)�(� 0��VH"��eP&h�P9�Q�T��{P2h�h�P��JEà���g���c� Uċ(\?��c��l8kq�)����$��1C��S���U/��% �B@�F�Eĥ�S_��9�/�{(�ZV�@_�������#掝�����_[*�v|��I��E/r��ń��9��<?Bp0��r(i��ի9�%��4�	Ʌ�S�5�2��$�h0�/�!�G�k!�
-���Â?�/��Y.{�6mZn7� _��&�*��]a��-�l�l���Rҙ��U"D�Q�Y�����ł��
)4n�+�����S�J~]��{�H[]���[ �
_E�Rb����>�����3k��^v?��CæB�?U�L:���o�����$V]�ߞ���۝�� &�qSۣ��{��1���y
��Ъ�{�d�VJ�`:�����'�!�\
�Ā>�ihy2>��������"�	�c���w�#4X��8�8`|0g 	�K2���g�Q:T�D��!L��Ǣ"j&Q7X]|W���h� �N�(�%�b�B���1_�7@d�h��;�	�?�G\�U�q){��8]��'m�>J$����hd�?���_�h�]����O*�27�?J/�$��o��{q��g�x�R��pt{�{�A��G2�`f.��TL?���Ǉ�~�~.��%N^Ԣ�!/���b.�k(I���6uZ��sZ�W�o��C���/jum��/���J�d�r���/�CQ�������k�p����`�>)/�m��� {�hG�Z(��K�'�Gđ�9$1h�`�����?�_q����t��ax�B�Y��/
8/S�τ$�@w�0(��
�BY4`�)�C�Aw��������А��0�5F���@"̀��y܎�g�r�A�fko��K��J:W-4s��l4�_�9��V}�e��1���o�fO�����I�*��.��E2�J@��U�	`��4����@  ���P�8 �d Ѐ�*��|�*Aa5����c�!��.�
����3s-��  
�@�po��8H8�X/�<'U������/�3�����%? �$�ƺ#���!�g]�2UrӾ������lf�q
������Z.�����!�%��ĺ!�A+A%`�ܱ�]�/���|=��L����^w�y�3��ZN��
�cF0c�!DP0X;	��t����N���ok�.q�'Uݮ*��
��ҍ�_�zMj�s���רµ�C�p�cu��c%Z(�U��:�pܑ�߱�V��7f	�r��C�Qh(Q�N&�5pf�0Bԋ�&O��t�nݶ���==�?#�ӭǝ�1��s���>8xc!
Ӌ`�D�������%�@��()�;� ��h<����9|)���1^���v��n;y�Ò�rp�Vj�H5Y[�Q�羇O�%��?}����f�h�`0�n�r�cf^���ޅ  �s -<?`Kr?q ��7MH�͠�-��`B� ����E�>?4��5 }�w��� �.s!�8�l���z�j   �3r����h�|������R ��x&ƅ3ap	 �e H?����H��b P�)!�b2>r>��u����c8w����A���Љ��n!q}�A�s(�J��Y��,XM>������M����S�3{��W��khl�<ւ����{���G�����SXŬ#g��V��8�6p'�+��Wm�t"n�j�V�Z�߄�-��Y�Hᴄ5��n���Vs���Eע`����{0;��\{�gF���r�d[�l�$?��9�Bs�$�%�	qbSB���P\���$!�⊻-K��fT�h$M߳�>���=�myfd$�����5�=_���y�zֳ���փ���V�T�-TCX���gT�O��H �;FX���k��]r�O-�/"6 ���Q=����ܲ��==ݿ=2�G:��+�y�j���@�x$��[�lSo��2�'+�>�>��8m�U���ΟI0j�7V�C�vX{�~��=f��R*V),�Գ���n���������o�h1��gW��@ �D���-�' �{>t���j�i&�B��` �X�o�� ���%`�#��^2� �=��my6� ��� e (�}��z��K�P  ǳ�;W ���� ذL�2ѯciC}@��?1�U�eL� 	m�c�i�6�jG*.Yi���:�����^oL�PY�˟g�j�Pb��.�ω�	�b��b���al�� zyg,*�w������챋6m�׿�j_t�&j4�+��Ip�X�;�U�s��Ρ5��zO�w�����b�}y�x]��9��G4��iy��3��ʝ�Z֊�-\��.^�ROh�z�c�< ��w�>��	1�x�p`~�+��@��lO W�cx�����%@����޳����0'��6}�uw�z��O����G]S����+7o�FOo�F,d^��C���A��� �Z�c!1f�R�Z&I��t�^�SBQJ}���A"��5X ,e�q�'�`��g���^��XC�E*��G�7��]?��r��54R
~v��uf�
`F��k��ď>��SX� )�\�pŽ1��$��X�����R�@W���X�⻙����o �����Yx�G�`����c����B8�TAE<--tx,&PB����|���|��=��k��N:�X�B'�����bժt�(=��(2�O~	%��p�\�!��}��]�Prܧ,�����m�\ v����x2�#o��1�Yp��x�|�G��:V1��vIlǥ����546:��x���L��њc��1�v�{��Xg�#��! E�ܹ�O��}��O)f#��_�ފ�~�t:k�r��_J6n�$��%�Y�P���x���\�Q��$fG�/������|�j�:v�0j&�l�H��w��H-;�~Ľ��/`M�'#�y�hL����4�O	V����O`T�g��C�\(\�B!��{�sN�v�MwW,M�5��bV.Pf��_���f�^>/+¥m(��J�*H'~�c`�B[ <E/&wb�v�c((D��'�T��6s��`����G���~�|�q�>Fk"\I�y�Y���>:�x�G��������P��{Խ���s�9@u�X�܋��`�K������<;�����m$���`���^������ه�� &��]��K����]`aSo ��V����X�ܧ�`5����R}�����|�uJɽH�X|����"��y<�2�B��NUD��2:(+!�G&�;�
���/�Z���b��Y�y�P~|�u ̞��N�9�'xx%ހ��g�������ؑa͢������~g�w�9��g�s^΅7�K�ϙ�	�ּr�	ڧųy-V���,��kVZ"R�����K����[��l��(�� ��k�A2�����Ywoh�ٟ�YC*���?�Y����ƻ�~��+X�q��T�b����p9���?��;��1���>�Bry���UJ�S����ӯ���ۿq�Y���>f>��������I��Ix����CB
3�$��E��
�(Z�e�B���=�����h�W���p�'Mg�Jɚ���)cbx�-���v��[gW�����q�6f͜�Kny����Ț�Z�p]!X���y2���r?�G� �~��@�y"���z��"��ZM�	�D$�H�TJ4��$��p�s��¦������R�<�)�NV>����<₹GY{R�pn%�q/Ҷ�K��O%��̉�p���xMx)xP��TO���[��?��g��X��t�L�����c��b}:��#q�Jc�w}��>|/�������,�Jy5U�Z����� ����dB�(�J�8xW���+?���*��s�8~����=�W���6yJ��k�>��@\�x}���{m _�δP�d�¼L�k#�u����.������7_�ޗޫ�5׍���Ҽ����Պ��q��/���C"#�9*5�ϱ25�*~̐�w"?`���c��vr1eAk�c��p��sw=�t2�I�:���e"���y���
*k���$9�8MMf�����V���aY���:X̎v���V+��Y�Z�bs��O0y܄�6P(Z#�,zXT��/�ksg��C��h��`�t�LƯ�������
P��1 ���Ƶ�>���'H�*�zЕ�㗼)q٢K4Yd-�2Q� xn���6r���i��z�N�,�kl�V�����{l+jMV��1����_sl�A��������D�������Ρ�J\ �
�'����*��#N�	����,f���pn-bl/���#!�/�E�k�Vc;t�X��˟�2�C�"���7׌5;�F<K��<*�w$�oȦ-_豄ap�,����2����%2Y�4�;����N�����U+�iCRk��ݻ���@��\�x�I    IDATt�E��>��Ϻ�#��K��]=�%.�-�m��ܠQ�o���E_�~P���m�q0���ij�X$�6�yG�Dj�k�{�m�Y���}"0�e�9h��e˫��=�iC�,/�� ����yйm�|� ���-�1x .Y��r�ha�� ���@�i�X����n--��ˤ=��#.Q��g�Z����{i2�I�d���ϛm"Ji$��m���+� ��T)�p<Y��U!�wՕ��U�&�����_]� �_�qh����\T���������-eYr�L��D5Z��S�|��k�z�K+s/J���U���[�eK֠�x- <S��v�8�<C DupD;r-��� d@��>X������N��I8�Ȇ�������u�ߺ�)���ϖ�П���w�x�AV���<h3f�t�b-��L-Z\;�t�p��"������}�!�����G�8O�:#J��,��v�U=�.�i+V,0�-���܍��GgL�n���ם�)�B��x���/�r���h����-�_�ީ�o��g�3�����_≃��/hl8��lC:�S��J��?z����$>��9�*������?�Ο`�T�o �믻��]�B��\���bu�o�ץvP��;d�q�A�z��]�jչN��8TO�>��q��yˮY��Cf�iY�X������c�w?�%����)ƶ��_J.D�aGfB*8�X�ҭ;���{����e�>D��,]�O&e-^�ʗ�{�uC UqY�ҀkR`�����5�-��N �`. �w�EO�k$�C�9��L.��J�d�s<b$��4��c��*�>x����y(%���Ȋ��X����5h�g�q�d�s\���E��hav�2R��χ*��Q򉡼�
��=���r���=���s�<�V�ȸN&��HB��3����1u�+��s���i�?�i�S�Ѕ��r��p�5�x.	���)�0<��S�k���Vڅ�s��{�� �$V�Ž�������K�a�W�������@<�"���&��1�������[�t�0����cbC����pA����d���t���93��<���E�u�ڈqv׏dw��c���b2u�4��?��$y�V�b���NϘ6�9t&���|�2���O����x89
�o-Ł���y�L�@��Ǫ"�&:���@B��A���B�`;w�ԺzY�B����>�����ms���^�9�o�J��}O��W,d��:�Fp�[Z��D:��2�wJ2 �h�YXP��FÄF�$���Ft饗xP���}��>� n0�8X$ @*Or,�E�)E���J�.��a2�h��"�Ċ�o�&19�2��*��;�����-�<=p������Ce�M��Y9/|0E�xތ��	 �x�я�t5Ǉ.Q|����F &c�w�@8cL���`�h��x�=��� �\Ƕ���R�s�����B��9��do ˟�� 7Ή��kg_��k"������c�?��յ"ϲ~���=�l�?b�;рıh�T_ۇX��z�{m��e��5���v�o��J5n�R�Ə�l6n�r%�u~��{�0�w�g`���_��7���j�f�t�����"��2��x�4|g?1��1����@��qD:s���y��<[�>�e2$�%����=_��sx�!X>f��N���@�	N�>���o��V�<�]�|�߶m�x�>;���z��2$-�M�.����3s�"SU|6���4�L8L\H2 ���f�Q�< �Ԯ^�[��b�wv�ֶ�V��F�5_�5��%�wo�=��v��F��h���7o�!۱�h��y���C\�	�\'���@� 90�lQ��< ���H��&�{��# �dâ�\,,,"�+��)��YЋcb9�|Ѣ�3�X�XX)�`Cͱ� �(^H b�}�+Ã�<o
�2Ӹ~����ɽ��&.��<�7����ޟ㑸�+ә�)S ೨�����=� �����G��F���2�E3��L���ճc�O��O�y>��V ���?���?���YE�?��sƻ�9S��g�"I5 �3�(����wd� ���q����T<ԓ��k���˸`Fyĵ����YWح�����X�V����;$�H�$%�B�����l��ɶp�
Kgm0_v#�󧼇u���4��9d/O�1������w�B�\�2.	N���sc�+��{���x�믶���pgg{�=�����S[���7j����k���um��3�Z�y�����{DQ����=}u�[F��|�)�b�6n<�^�ZR�y�kn�k=|���U����)���Ҩ;oG���ŗ\��\}���I��Z�b�P���L�s�� �﬉	0a%���j�hR��ԋU,?pܞ����
��Ɇ�Ka��UϿb�X�-�P��U�f�(�P��)H��|Os��

���ʱԙ�ߋ�@����ŁkYu�yVX�,�,xz������aq� K��,(���� ��U�p�u�Pٖ�3�Ylx)�6,8�EZ��]�=ۯ
	���\�!����,"\ 1�����0tV4�b��d	�+d�+נ��|�'��C]���b
Xq� sWO�{9�a�0f9.ϗ�Xt� �� c��v|xWlG�>j�o�y�8�Œ�(�8k.Ԃ%p�ߙW�'ȳH�����1�����_��������v�R۰�����K��l��6}�|�0~���|C�8/��s�_԰�+���}��N����*6y��B�x~����R���7�)��*��n��6��?j��6n|���Z��>5{�寰Y3�z����vo'�{S<��8�7����nX�����k^s���a�%beoܞ�Ĭ����=�2J�R
���{��y��b®������L,'��QCrԣ�k_�]@-�D �Ky��'�?n�Z��F&`��e��n���\*����=d�����w0wsm���,(�H��������d�2��` hi���bun�`u�`�tx�,�,?��9�� �����>@V�,,HJG�i`U1��o��(րE�D0��(�@k��%p?瞻�3}ѕ�;�Z���k`q���Y�w}V�g�ǀ��҅��?���y�O�p�Tw�= ��
� �Kޢ���G��R*	L�N�g$�'�<��}d]C�K��s���ȣ�X�޹>���'�%ZJq����}�x(|`����y�#.�{Q@�,�������3�k#�>��_���y���J��n՘M�:�V�y�������c晐��F!�9i�|Ǽ��_}��LG��l�Θ�)p/�:�Zq<��^���&����֪��m�Σ���v�Z;�d���Eڑ�.+C2��|�M�8�b�?����n��.=WŉN��>�7s!����N9���=�o�tܲ��v��mͪ������u;ׇ
������:�TN���.���_�T8@�)`	������2�\l,?TG�v�$��W� �Wy��
�Ճ�J�j�׬��նm}�ʕ�gf���}�?��J����"/��?�#����\3Vu6��4�@������p\,y����m��� :�29��������"l <�?�����e�1�U�sJX� @̢�����n�kp��_q����{-N�3�[���11���\/ �W�g�f%� �b��xlâ(�7V?�f��9.�ͳe��&2��3U��.�lx7�[ �Y����<S��8d9��c9��J��$�,2�I-��s�/�c�O%τg�"ʹ�r@�f�xx�.��=��5��X$��)��:��Q���@
,�ݜ����;Pw���\�qKe�֬Yj/8�b������N�l���h�:+�Vȗ���?���{Tq4zG�I�P�ǎw�_�t��� �����^�;�`Jf��k�^�f�C��'�s��J���wYC֬�1c��^�� �:�I۵��i;x�î��[v��K,�����[n��C��zE`=tZ����C��>Κ1����m�R�;c����.�� Q�:��A����~;x��
Ť=^��3�z�D& /k_*^
r9^:�@%K +x��+\Ѡ@�`�:`r�^Փ��[��X��a{wo�d*XU�.����'�)���ޖrΜ�/��~��w�&^�g���w�4LN�^Ԅ�f�� � 7 �}�Sn�����-]�@��W2S�K9�&�hY�R�̤��z?��z�����-����{��e��j{ (1N��Иj��9�ԓ�e;%[j�^χ�=�
���?��8���zO����;������ ���H;B����kd_�)T(q � �Y�J��}���x��w�޾�6]|��Gx'�>X<�b�|����g5����jW4u;�x{Jv`1�	P&��P���%s��;)�����Jm�V�^b�?�;y�����'m���6k�Y�m�b�A�Ū'|�H���Z����j�x�c7�ڇ�>u�L����s��0�0Jx&�R��ϒD�K:l����lŊy6u�$�����BE�*I�q����=��6�i�����u����.>p�e��[ Nk�߼e�{z�Ӏ�1d=ׂ�ꬕ+�k�bM�������wϝ�i]�r�==]��SM�u��:b�r�����.r��������I�t�r*2��v�%�A��h��i"^�R��v�x̺��z	
� Z����t6z�Vk�h�"�3w�s��:��_)� ���I�A�,T~�"����lϳ�X!�: ��.e@*�\���\+�	@5����� �&%?9�~��nط~A�5�'p�3Wb��Zt�VO���X�ܯ��h��4.��K�(J�d�k�X
 �3���g�������pmx-����XR���Y�Q9�!��>ʑP�-4���1c��9'@�5J��R@����� 8cZ���?~�����&��H��Ϙ,
����h���N^��_��=p�,��VZ2�j_�z<&N�yα	�g: �C.	��D��D�% �?�2	�֗��dhlø#���Ž��c�|b���!����c�����b^��ҙ��ݷ��w�_*F�J���iu�����U��� %�@�홝;�ٌd�������_���~$�'��@]�t���~�*�A��;f���U���-�(��C�^��C��y���Z�Z���g����6zEJ&�� "V�^:?���I�$���䤙|���0A�(�������jǏ���������K��V�V2�4��t$�t�Yͻ�-��_��{*��k�v�zB�Aq���J��W� ��7�&)��ǩ�(IJܴ&���kW�W�e(p�'V1ϟg+�M��.���7ā�� �R�7�=��^ �u ���s~�'���iw}����u���&�/%�AaQ�=q��C��/���
���g�;��' U�`�B�Op�hX\�<���Pw,4,.3����q-HCG��Y���P2caN��;���KGa{��?���\7�� ��{�_�����i��Ӟ�5`��.�u�V���Z0�bi7q�e'Z63��.\l�Dƻy�H��:�hL��;��En��a����~���Q��������;O�4����-����]v׿��F&����{�b��Z�P���n���$;�v��{�?�J$�r@/�ݿo��3#����~�-'��t��9:�G2���'؟��y-�L&fw��5[��L����4�Vн�VM[_o�Z[�Y_�:��v���}5g��+c!��y�v���p�X����#L�%˖�%Ǥ����'���k��y�+���[��m��K�,c��7j�qaSm��N���G��)� �Zd���hI^Rp=^_<�:�Q�A�l .�τUr��tU?���J}kC�� 3�����A0y�K �v��n���@&zH�E.�ߎ��f{BD��[y&m�L���ST	���y�,�sX d��3����8�8}QW�^-,</>���#cDIO�PP�= ��P=�G�t�{#hK��uk�V�<<��<c/}��\����ze��3�ga�������o�UW��v ��?ng�\��@_�_������PG���3�S�$ׅ���_F�F����?j�dS1/�p����a��V)S�'��3$<��Kem\�D�p�ž ���&"����X�c4��'<N��/�ߺ��.@`� �g<d�~%��%:`�C�}�uw���i�N��q	g�}��/=a[��D�юu�lٲ���o|�Wm?��ϲ�H�s�� <�
�}N[��rOo�5#Y���2Y������k�s���-�(Y>�c�����e���LZ{�1k9�a���]�~�Ox&�*�r� �,� V��) ų���z�5��f"�J�+`�`%ԫ}F��#͖��,�1��u��ke�;����;N��e��/=|�J��fd�g��A�@8��]���� `���}q,I�ا�W��z�XT�J7��?E��L$a���(��}�p���H��[uQ�e-(|�8�hyql�~,`��⟵���!�h��`�����t�1��la�S��\��L��3Bm�3c�I1r�w<L�	),V+�`qs�LxD��.q�ߑ�@����}<+%)�W"�}��@��(����9�#��|���'�u�E��	�s�:?Q\1WD�`(��G�?���p��IXn��6n<�.8��}.�z&�]��U�)ˤ�s�Eό�{�^껇�����n�����qp�����]>G%&��ȳ��"�Q���=r��j%o�>m���HV����/b�4%-kv�h�5h��#���׽��]�֟ŝw��^�H�^������vǭw|����O��F������s�J{ӛ�h�j�*ł5��}{wz5O:��=�#��r�j=}�6}�"������PP�0�Eo����pR��A��2q�wדg��T\B$�N�T����	���
Sg春�p�Tm+�O&	�M�&[��#�u�;ޝ�Z?��f۲���*.$����җ�4��s/Ǿ��<���Tő��JR\���x,I,�ƢW�5��Q������U�< �X�Pyj�V��%/�-���5�/����i.spc,�47��.�l�_5� @Q5���m��F=D�`�J�����򈤢��&�a�g������έ��/����L��e��\���[s�7;�Y:��{��)��Z>_��	�-��X��={f�{�Y����<��cV�e0���e/}�{4ܣbP,N�w�������� 7�Z)X��xd�7EJ��
0x�i��K���k�T�]v�+���,���v�w=&�4~¨/�����?r'/+�X(���dMM��7�ٖ-[�u�a\�~j�g�>x��ʅA�t�B[�f�-;k�uu��D�7+�8I��ݨ�8���bB�
���:�k��+�í�:��y+7e���C��eqf�@Y@��i���5�B�xͥq����Ŋ:�c����_�Q Ɓ�J�~�,}��Jn+M��U}(Qr�)�p����+�l o��@ � B����j��n��nbN@�a�@7�v�;�AX�쫚F�2�M&�
}���L�;�ʊ����y*���o4�w�'��b1gMM	ה�� �{2���Ǜ9e�91h�Z�-j�`�s���Q��8S��jN�U����_��1<}�J��ŋ�Y�R���G�g�v��<J�'����Xn��]`��&o���Νv�Wi�EU��˿蜧5�o޲��{z^?���A���6A�3��3,��Oˁ����a�r��Qyoά�6k�\+US�8n�[Gdh�ؖ�@���ѷ�V  9'.9|,�����p��s�d+�7���ܼ���v��ak���L�EI�1c��+�c�e]�F!������ٳ�����\�,�_h���A���׌Sh@�PG0� l� �
Œ�Øb�3�P����L�|���Ǌ���)!��Ʊ��}�    IDATd��3( ��İ��U<�le<���ù�sa��	��"�˜!&�, �$u�D�wά���'(�V��8�}K&ʖL�l07�q�b��U�����d�r��ͯ�T��K(P��A8j��"������e����K�͛�h.�u���dA�3���빱p2�7����	�m��&��hs�Tow���y��p�*X �v�-c���_[{�W
�Li�<�Nk�r˕�����G��w�R��8m���nx�M�2q��T:�rp��8�b�W�����\+_�=q���FH~�}�IU>���KC�OQ����/�=��ּo��ckjL�@H)GFa�={ۮ����������,���&U����_�q�}d�364���+ �$hȮ`3c��R9 '���n�ɍ�N5�H������C����!@����>�+�CX��`�X�ϖ)ٹc���5�qCG�m)���I1?�@)fS�aQ]R�)����Ϝc�z����n��B�l���v��K�j�ު�bE =��gΘo���׽�s,Ny��d= �M�
�>G�����R�7_�V{٥���"o�k�:QAAeW�9�]_�}Ӧ��W��M�8ޚ��=������;�=��*�g���]{��-u���V��
ӧN{�i��9�埈k�I�Ʉ���7a�xzQ ŭ��D1Şsv׏�vK�~�,�X����[IxA�̠Ɗ���2�ؼp�1b��8J=�������ÛTSԍ��Ɔ�[X(V����~�����4�F�������w�������w4�7�lKD��ĪG#KRk�)����θ����PQ&v>jdþ,���>�O���� ���9�Z��k�W�q��^T�T�q��it�*����?�w�aI��
A�#`��QI�[�ϭ�Op7?�kk�[a�6��Ze�j�UJ9$<V��l��i�f���ן��x<.J>S��8�;��٧����3����߱��\ڍ����9F!:h6���ޕ��w������gKsY�	�%�Ugj�������:ފ2�k:ʍ��QhdS"�ͩ��
Or���x�R_�\�[xJ�����U���^�X�r5>�w��f����/�8~�%Q��!����~ ������]��Ԑ�d����Z�&O�a�w�;|���2^�%Ȃ��NYc���Ͽܽђ>@A� �C)�\X��we3��A��Po��Fߗ��#� f�U�o�Cy�Mݤ'�x������Ko�tz�H����]��M�<GEtǠ�%	I��E��C�t�2�z{{���O�
�# [Dȣ1�؎E�Le��� z5s)נG�����e�ןe]x��}������U�I+�)�7��n��-��>b��������K6��9-����ɖ-Y�^W�ҌA�*����爸$��y���z����&M��m���m���~�۾��t����à���{�0u���{�m_;y��:�o����a$ڇ��In�/���χ��^ld��ł�=n|hP�T��g���g�a�A��EF�/^8ٗL&0A3,;t�X|(%+�a8�?�붣GZWW��u
�T������.����>cV,T��3�r��NA�i��>�\�G���� ��3�c��&"��J�%H�$ aٓ�Ż���[(E�( zz����F���L#C���F���#m���,]�؟8���N����u���f��Xx�7d�/@!�9�^��zw�(ܛ��p���}�h�o���]�ܥ�I�?m˥�%��mʴ�6q�6u�l�x�Ű��U$�<W��p���_�B腲m�t�]w�[\�D�B�c��k����T]&)��d�޸=HxQ��B��,޾�^����8NC6����YG����X�V�O�>��;n���s>�=��ӨŇ�������+��O |�{h���Ui��cM�	�y�*�'����PJo{��<Y�	"����8zsg���K.۳w�l�ci��5ҵ+f�-�v���@�!��4v\R��5*�h�_,<�r��{V� �]C4���
P5R�0�@�` ���ᝳ?��{d�����V6��ˌ���Q�A�@]Я�r~���&su���A���m����!����9�z�=�}Y����#*U�^ݓ��|�袋�f.Á���s�]bm\�%�)�H�V:3�.>צ͜�u�JU�� �Hy"�'yEy,T�$�듟��Z���0���?�C�Kt��xv�R�@��˳�=`4��;������a1�ܳʐC�])�ĩa2\v�� ����Sq�/h�8��Fo�`�EE�"-���x�dM2y���O�#� ��=Ǻ��Ο	�d���YC*i�b�R�=vؚ�m��`�/T��7�������T,A�o-�nՓ�<��>�k��Ac�?i#�O�7��L����"D% �ÄfxY t�P<:�<	�m۷{�0�' ��l��>ۏ�}��ӄĵ��2����#���k�������V�^�F���G�g�>x&j��v2���`�?��J����͘�6��[��x�b���[��9w��SU/���x�Y�h�Z˗0�2f���d
'���)�h�nN�,��������k|��dqkjhp��8��uq�м,�F.�� 	��àO,h��GH<�>p�ӦO�����O���WC��?XQ-���>'�?�(E��cM��S�f@��M�H&��Vw&21QV0iFj�k)�,�IXS6fmͶw�V���9H`iii����r���' �MM������g�M�集
�R�@���ˇ�i�9��rI�b%3��� Q5O7�zD��*�xa�3V��?��%xw�I ��A�'��A��5r}���#g?U����b"��}@k@y��T
פ�o5�q��lq��^؍���f�zB���yk����˽��}@ۅ�δ�γB9$m�jP>)W�d���[�fNd}ui�O}�Ӯ�w=?%�*�ސ���l�G��u�<���,D;ɲ�1�^�e�{{z^7��_�h�jH��S��:�w���y�b��X`\`�9$e�äQ���n=�:&�Aޚ��{��J���"���J:?d���	�f.�梪 �<F���������󢪍� &F����82��� b��f���j�˂�*�e�Ŋ�q��1�����R�c��/-���5��kb��9�x
[�|�&F%�|��O�Խ����	>��I�+���E^F
s��(~W�!�9s��U�<�Ua�lM�[�֮4��:�SΘm˖o�L���-Rޝ���ۆ���%T,��{�ֶC�ٿ�,��bL<�P�d���r�(F#�&>G��O�8�� j!;�9Nw��;==��}a�����q��G-�ݯ�h�l3a�S���	,��ކ��U��D�z{�[_�u��Xww��#��-��v/�ݢf.���cD��⎁����5۠�/���2���]��ϻ5�A�hJy���Ϙ�8.��sw^���<	�r\��0�j����� {�(�r-c[Mdؗ�p�x'�cK�/V=�\��U�f?ߑ�����:ߋ#�~� �[��o�?��:Q��|�]x�9v���Z����x����>c�M�6߲��4N�B������s*����v��_}�
Q������K�+�K�bj�=*3S/�74���TOp��_��� �#�8,	ύ��~�Gp�Qd�);W�
c�KcA�Ť�����H=�X�i���f/�L[8�QjU�L������9m���#�왡�`T�v����?a�_=�cq׃?�E@I!ۡ��~�; %�q�ō���
Ń��lT�)���u�b1��(v���B�*�5J^T/�"�����!�W�R�;*�W)��Iu�D ��y~G�I��\�ߓ���������S6��a�
۰�\�T,���Ӻ�h�����V�m�}��P%���뱱Z�z�����?�s/��s�e$*�������Y��Kp��8��:y[���~M<�8#��u��~�7��O�	����?/��	�	��9y��M�ădo��*����:�8dmx�#}be��4:�V+)��l2d����0�Z��]���W�VP��?�\/]�����ON]�z�5M=�C숚0d�:hᡂX�
�dT�w��'?�I��_UQ�i�"�KZJ-@��2b|J�L�d�q��|Ϣ��,>��1�@U�gScP��XD���Ăǵ��S�d��x�������[����U+��mݚ��s��a"Q��W�	/�R��m℩v�K^扑P?(�<W���Я�q���J*��� ����<s� )|FYw=#�-C���Q^G0>��"8�;n����Qi��_��
�ؓ���xl����Rɪ�U ��B�8��� `��j��J�L��R��j%�V󖌺a�g2m�f�����l�R1���^�(8c���	�����>�B��,jh�C��G=�g\�DH��Ģ3�yM�9s�G?��� ��t��\��e؇r�xxT�e�����g�{�g(���8 ���F�-�	E�ꇅd0�?$v�����im����4�q��\gϜ�
�� �TUO���&V��m͹Km��gӧ�ɚ�g0���\��,Y��ZjF 8����[���|�;߶� �er����Ӟ�v�~G�GGY'�.�8��<�>����0����N�~�wo���O�濽���|�K�Ї(�@������Z[�ڑ�W���;��L��R�y�ZD���D3Ed�{�1 ?g�֘IX�4�HH�'R���ޢ=��6�Xƕ�R�-Yl�����Β�����&�#g�� /T6/�.�'W.�A�( ��Ή:��/2QJ%3�<}j�6���>�5��h��泟�ĳ�	�B���'@�<�*����8@�)>`�J��liJ?s�|��͟��,Z�9ǎ���-Y��ҍ��:	�C� ��c�P�͚��s��k ��j�����p�;k��P�V��,�t.��۝v�����~D��'��'���=P���l��[-z��x��>�/��)��܋�BA�u��[&��� �L����+7o�VOo���|�V��54f,ח�j�&��uM'3�
��i��fuB�����ِXLLJE��sTkE��+�<U*T��x�6����'��9f���V)�)`Ԝ�,W�)�,NF �A-n�.��s�vq�S|���:$9Tp���r�)J�׬d�_Mh�տ* F�H� �s��l���7Nd)��T^	�C�|�!���`��}��c�(���7��M�|�9�dYTH.���Ch�hu�W��NU攬��J��C�������?�����"+�������k�xUO,�Pճ��[�f?@���V)3��r������M�5T��S�[n��ٌ?��ɤ�ko�굽h����\�/u��� ���}�S���� ��5G<_.xŀr��� �΢LǼ��;�rȪU����`(I�ChH3�紶�GO�%��j^��R �d<e�]�R�;g͚��D�]R���b����� <���pl���冻����RkA&�5���C=�t"�T��;����l�\o�%1KE�Y��L���~���4�f�'l޼C5R�����I^����=�3������>��Ɉ�x�_}��սB%�i��JU�D*�ႊ/Z�e��y�O<���a�w��.6 Q�3���M�8��А�_)�d�B}�������F�-�xy�{�;$��PB� ��Y.�Г�8�k�
�˸Vj�qȠ`,O�:���s��	���P#��ڄ	Y;c�xKF�J�B��b%���[`/{��f�z�X
��q&�F����t� ���T&��	�x0ڔנX�EmK�Y�P�!es�Rq�l;�앎3fd�!���7`;w����l6m�R��r}��~#Nk�r˖Q���p��usή����y����'O����ϼ�C�����(����i���z�������D��FI^���5�k$��'|�l{vo��{�ZB�M9����T�|f�>{��m��M㖬��;g�-Z�0���b$����M�uY�xp��p�yNyB��ū�>/�	8������s��P�����ࣨDIe���ܵ���n鲅������;�UvA9c�����[�h$,S�%X�x��G>2T �kW�k;�:�Cc�{Q�,�(��w��]�HhA#>k�[�p~���퓌�N^_Tm��œ%[y�"[�z�{�rɒ� �4aǘ�4i�m��+㖈g��o2jd�blE��찏�|�{|�����k��z1�H
ʜ��G4\}�r	.��R���mΜ�^��Z-{��kjj
yh>X`����8�U(���T9*�=� ;����ͷ�t��i$�-jw'�Y*�����W��[:2�r��^%�h�;����O%A�ep�t�'�����A4iy�������+eȜ�J�����^�:.���������'��6�f� )��2��Fk9p���!���[&KY�͝7�� �.X5�s����������n�C�!X��5�d��A^4��;�6���+�:E����=`-�d���J��������c���a�(XI�h��D�W�,U;�Ia�����իz?�C�� �9�K,W΁�c:�V�7d�3�Pq>-Ķ��\%OX�Tϟ�>sf���z��r��֯[i]�֬�w�'�(�X� 64N��7\��o��P�Y�3��vx��ԧl0?���^L���8�X�'`�G4�(-l��+^��v�K/�d�R,dq����~2�T��=r=�rr���1=��\!gY�Y��?�W]��+��=o1�KE��)o�r��+�寸�z��z��c�;���O?��4M���sV���o�q&{���R��LQ;��XT
�s�Ԁ?�1Oaokuݶt�X������;P��С�ֲ�U���(nc�ۻ�m��O*M ��<���#p	�U���e�SٝJ�g0�z+d�X$FRA��x�3�:�S@ �PGG��h�W�,��� ��w��k��G=�K��:(�DUZ�	�sϪxn��f� :�?��O|���:������+�Я���b�@f���y�{���.��8 j%Ā?qU�9�S���D'�@�b��X�{�!����q[��L۸q�����W=�Z�ĬTIZ���I����.�rm?}|�ޛt�-�,�RZ�����+(m����K/���Z���ډͰp1Wd$�w��K.��z�o���J���ჶ{�km=d{����x�2[�t�-X�ĦN�IPK�����py���S���:�����v$�'��I��5kV�u׾��zl\cʛ��w��F�L��'��JO�\�
%���앶x�
�\H�ԜEY�L`$Ȑ���CC�[n�ś8��-o�^��eM`�SO��H�hW��9ܺϊ�ǭ����./�J5���mv���Ya��/���m��%6�l�Jb	��4�*p�:!����� rq喳���LX���G������f<�A�99�+��h
�!��{��?�f{G�, 	��$� x�y��\�V����Զ'}�R���BQ3$�\=��0d��/@H	
��P�;�g[>�}�˸b�q}����%m6c���|O�H�J%)��kk׮���W�%9+�l�3�-�Lv��3M6c�\,Z�`p,�^�i� ?���t�v�H{�;���hx)\���h��s�])�':�wB<d��q��gv��n��ͪEK7d�!��\>����	S�׮x�M�1�E���Wo��:;)�w*˿Z�>u���e���-�����s�H�IC��7�卶t�|ˤ��Ҽ�J圵j���nO��S"��.Y��{,W0L�;���>�$�Pޕ�����?��ݪbB�!�]�U|��x�r&&ނ,�z����h\�l"c�Z�b�۳o�:�-I]F�������m0t�( �9�C��e���^|-
�LLx\]^
�62��    IDAT)�~>��[^��ƌ�� 2H=�(� {���3^X��,7�|�?T,�_� cE�)�鱦q���0��Sr�cqn�	 �o.�.�?��<lG2�T;�6~�lG�K�$rn	*�RK��@�cɰ��Nr��^�YI^!˶��$��D���3g�V-�������Oٔ)Sfۜ�l��Y�;��К��\�`�����B���s}��G}�p�Ϛ��$Ç8���L(�{���X�R��Zﳖ�v����k�X�\�*�:��*��3`�J�~�^ms��̦bw|�{���ĩ��-�jq��iם�U=7o�bOo����}�M�b���7ؔIM�L���߿��\��K&:�<�-&D���6�׬�Xɮ���p�&����ʇ����qH�-��ʾ��/����E�B&�it�gܬ�kZ��l�� ]@��a���Y�<��Fk����1���@��X"fK�-�ӧX�B�PO|4�_*�MLZx]�E�� �	��k��?@C*�1�O �!���W�@�<C!z������\<���, �&���/�=���|q(��3��L�c����;��qh
�V�����".�^J5z�b���s}�A�ߡ��XCn�)����e��"2v$�4�<�-�)���騼�WC�
���r�f�2���s�F"d<��Y��L���<��-_��E�]���"�z�s�>������&���?q�,��' ��w�.��?�q��p�)X���m{�^K���>|�r�3 ���í�֟+��`ͮ��7m�y-��؃?}�n���!I�H#,j�~����+����{ð�O8�lz�2{���n�b�Y�h�����K.���B�k��:�&����m�uX�����}�h�
w�x�j��B3��Q3������2���Y|�!��1X̸��h� ���Qy�ᥞqK[��ʃ�M��%����`��R�X��w�p-��%K��i��Z�I$#�?��kf�cyj1�u� �[Dfn��H��ol��'��d|1f	��H.[� ��6xdu��c�d�m��$��.ՖȌe���� �l��N W	d=�U`��9����A�qY8(E���������op�d�K3Ͻ{eT�_����F��T�_�تs�؅���E�Vڂ%묯��|��QD�0�jV3J��	ć�|������
���44��ʜ��	p�k,d�Y ����v���k������w�[�l���h�-���<{��W�kw���nhN�6׮�������<������7�w�g%*p�G�X-��,^do���J9gG:�O���]t�:ˤc�ܼϺ����N5Z{{��,�h{���k/p���!���Sn!/��c1`v����,g^��s	(U��p�O%_��q)�{l_�6;ұכ��h41n���y���	�Ƭ\�[�Ry��5�KU�$����j-�&$�- �1��/n�I���ǳTޅ��#�@��ի�k �xW�?���G��]%�i!����'�!�?5�1t�E�w�=�`_��j��,V|ǘ��e�3 #���^ƍ(%�˼`�S������v;��ɤV)����K��ɂ�x3h�E��;�S*�J�l�������
R�[�\�_�xc �Z������#�g��'/�6�������@E<)��]��kw���v��sl�����������;h;w�l�dk=|�*��}�C��K|�o>c{�����ؕ�Y��)U.����J�~;��a��/�`/\g�B�;��	L��%����n���m��|�*��UW�}�{ߐBCV>3�f�r�X8X>߾�;���HT�� ���p2��|�FI�����юfk��g��#8U.��4Xs�ѡ�/��ր�,/ i�W��(	�[t~BC�09�������H#�?������L� `�2� fx}������E���w˾�U�vޥ�����{}�R�����'s��{?��@/�P �ԩ��`,b�
�]�{M!�
Y4���!�,����ˁNT�<��Py�(���o"^�b��֭;�6]��9�|+����ON�e�W�5�ĳKZ*�`�\�
v�P���'>����V�<ө7����@"��C���K�Ƶ1���b�o�������s�^lS�N����T��d!_��{Z�\IX�^�TR�я��������ܼ�KL(��>��l�o'��e�L�2�>��?�Rq�R���v�7l��U�y��փ^���?�tο����Ÿ�i9f�6]����kM@V�5�U7���7�n��@D�`yPPj��[Ա�57?cm���ԓ�.�(Y�"�Z$i;p��ԓ ����A�|*�'�%Ǌ��U@˟=E#���(����� �����qw>���ƫ�3�/e��r�ԱFh@���>���fl�p�, +`��z����?� �j�����[�@
G��)����˳y��}�f�6@kB�
�#��sqN5p�����4~J�gSc�����V�E�y�ԓ��J-m�M��i�d;���V(�,fiK$�<���ϸR�8������7W������%�Ur��ϝE<�tv���?�|�\k�fl���n8�����\�v��o�x֎w،Y���kǛ���:p��-��8O�����n��m�}���߾�ە�7���皑�>h�����h�_�-�?�j��=��}6�����`_xў�D���l9h�����]w]�����C�#���G��d��gR�s&�{��׹��-�?,(	8�H%���쩧���foW�M'���Ja��	z�v���<hǻ����=���z��8��8QG��:	�"Їw*�s#�`� :�Dy��~���=	EX�H/���*�ޱ�6�S d��R��&���]���O�'�:��O7.���E��wj5�1X$X��s P�]��(s���i�GM�J%cV��_{�'yŬ`U�7$wR�N��K_a�Z��unt�X��ڇ�\�Go��3qy.h x��_�5b)�7�����~N��G�w�0�bǺ�Q[T`qj=�i�]��~���k�`�7\�E�ܺ;��o<'�o�A�?}��n���[N?��r������e$��lX���]�Mv�k_k}�]� h�mmV*Z&s�����~/�0q����W�����V(E���o�;n6�~Ǫ�A�U�� �.#:a���z���E��re����b��sO!1e����b�<��-*b&̛� ��%�p�r�#���)��U����*E��$Y�����g�i8�
t�/�MI� �(�>@�"�o��+I^�Y$��*����0N����2FQ��v�w��E���)�E����N�`'�㆘eh<�c>@��!p^<%��1^��s�Z�	w,Q���Zb�֞c�t�*ł%��n��9e�6s�W�T+�ư�Qǅ�8���˾���9�so�L�ʰ�s�����S�#۰�bPʥ�#v��>��hsj���R%����H5X�T�;�Y2�`�����S�{ىo~�[�ӟ>4��)�v�������t�y$�@�/�\qk捿�z�3w�M�`--{m�Χ�ۭ��{(U�K�Y�m�s-�j�����N��Kd3 x�b�o�8��������@F�dU+<�QGh�^v�*�56em|R��%"���$���Y�N��Q�ki�|2|�zEQ�ꑤ��3��=�p����τ�?��Á?�*�1h��-����1E���0��'��z�� ٗE�W�I��%����3�n���߹�[N�`�(X,%��������@[��)��?�#��8��L���;�4*�2�K
�z;�9�ς���ȅ�&Mj��&{UO/�Xt*��05����T&�4Y���c�]In0���Ɛ����3���:���-���	�f���Rgh\6iG:Z�8���;�����^8C=�����%�^fM�B������/���	���- ���mw�z�WO?���>^ځ�?��^�y筱�_�?��?���zmǎ�]�s��O��d�̚� �R̃��H��%��ÝE����o}k��?�4z����?��?��L&ܠ�����?\�77�k��X�T�$��(Z��)�ʖ�d�>�%�F�^������j�Q����_��M�ZU%�>
62�Ƥ�?������v�n�±������^x?P����{
��E� +@�g�ƍC�d��J`c1�P�*���n���;h#�9 �𦼁<Z����������Ϙq��ba9C�2W 9�sB�: |����I%�CU�t*���>������:}W�%~=.�%K�yrd� �<�RԎ�gt��a��_�eμپ�>��%ܻ!��c�!ཽ���y�HZD=zĽ�'�|��Cpl�˯Y���=w�M�8œL)�����ǝ���t=aQ�$�1�$M
�8���T�/�d��f�&M�	��Z|����n��
�H�����>ॺ8r��ċb03�xXE�_�YX�d��
ϯ���`��m�3��b��~�R����
�Wl�S;�)�b��*D�����$��(�� I�	񏴃�B��`5�� {��6��O@�Z@Ř�l����h�js9o�5�v�\�9- �D�
�R��*�'ޞ�]��Ї>�/Zs>��Cm�c<��p�,
@ �x��P�?�$I�i�H�/c
��j$�
�k�܇J���Ϟ17�}�'qkkk?��1i��?g�$[�p�UJ�fR�P�͛�{����W���L�T�L���.X�Qt-�W�5&Bc�8��x2�B���/�`	�=�1O$��MQ���\�%j<�����$�
100�`WO�3�|X�K���7�s������-�e3Pqu	� {�ej��w:�,2q,fl+��Fݐ��=�)4�*U���X;z&��%����ޡV�];�c��<�Db
@R�/�g�a{��^���>��͎���9O����
p���ͽ��[�'���;T5��0��?���ͻ'Y D��0�G<3���w��|�� 8�� ˛y�1�'��Up�xrP�Gq<��}�W��@P���W�wE�n��ÜQ�"2��:��Mg@s�>G�mBL�RW�y8��k|�6h�Zf�_mF�R�X"��$ǁ���k�lm�Ԭ��B	�Z��嚢��2��_�����Qo�y}��/�o�>扏0���
/H
 ����3\��c`NJA�*�2Hهg�������JMwZ���-������Ƒ�J<�1Ȕ.���dnP&/������->�^kؓ��2�M�'��ŢW�� �%�TUO��F����3+ێg���P*��Y&��~�P���Q/�Lc5���._�$<Y��OF���k��^|X���\7�/W&E�d���y��7������ċ�nx��HOJ�y���&y%t%�_�+�|��R���U�Y'=� 0���1��X�(�THF��J�
Us�1$�Bu�6� |�L�W*��E�%�W}!�����چ,�����β��g�b>��wN���Ujq7�[{�7�
�@������y<^�Q,:<G����s���<&�8���Y��>�яz��W�A�<+B<8�����3��𼠿XP�����d�c�?
F�
�UISJ)%���jG��s*���ZH���AY�|��h�نA�W@�Z�u�	��*�'��Xaox���4�8ٵ;ةZWW���{z:��U:��������w�O�y��b��-^��fϙZ�UF���LV=i�%'T"�\�z�y��' �V�, ȭϺ�������"eч��pT�$8q (G@� c%�L>�ˈ#0�⃪�0��4�G���ƈ
�i�H&�W�.�"���o|�ϋ�EP`9]ŠU��/�|^�W�7��%�CUφlҊyJ�������Z]�>V1yz�O�4�Θ:�/^:y�)�q��>$-66f=��2����н��w�*j')9��j� �澸O����IU�ERυg� .�=F�:��^��H
���P��JӧN��4�z���K@%i#��˲R�h���|��>�C��,��n��i!�K�Ë��L�b�xSVw4�cB�`�H�y���\*�-V+Z__�<�ú�[-�E�@�Ѥ:�e?��a��H����-�g�fOwz(^K�j�s��X5xUp��&`�*�� դ?�e��A����eA,�n�
���$�D�;�� ���Bg����{�2/�`̊Ҕg��\΍�1������,M
����;D���3��x%|8��Ca�V�N^�U=U�٬X����t�rܪ��%bY�5�L�4y�54��L��
%4��~PBC�[Ro<ݛo�Kf�ӷ��Z�0i�'�a���H���ûG����_�Ǭ���L���^f��,m%~1�����j����������#�<|�i�Ղ ��� �@�`��~y���$��!@�Ń�G�n3����眀?n#�q��[�qo�ސa ����Xs�6��h������;CU�\�b� ��ϵ9s�[ie���*�~Z�4�����;��k��P>����C�/�%�幊g,�D����AF��V�!N����ƽ��Z�%ٔU�1D����ǖ�,�EsPF�"���b�x6m�<T�M�ζ
rj���=Q��,OEU=CI��4%ɻ��ϱ��?Ǫ����9�;g�^`����Tz�W�-�V$^���{�*������O9��
������|�	�X�h�U�n�h;C�.�AϙsS�D���/�N����2�O��W���)e��B�W�/\�.^�"��Lhd�������Y˒���-�4�xMx=h�D��;����IKO�[oO������>�S��w����'��b�x谵t�"�3w�U������g�
xVr�5����+��|�O�J>�
���>��{��� HW?��g��ƶ ���q���b�y����U�K��~
��#/�G�D�Z�W�2�D%�k�˜k����Hj29�P=�J)�}NJ:��a���a�ٖL�Ӄ�l�|�*�:s���d�s����H� ��<����3_[�a���}th�s}����
��QZ�1�Ƚ@�To�K�g�g�©F:||���UKގ�������M�z���?EwM���������{��]������ٚm)�R�Bh�iIDEE@D=��S�v��;˝�������"-	M@J	%=�������g~����g��eg7!	p�/^����Oy��y+
/?��4[nHic�nt]j'��Uf5��aM�N9�\@�� w:@l:!k������+�d ��;�c��L˺\�@��ƣ�-EG�Yˮ���?bd�U��D��W�o_��&��q�1P���������\9�����K��AZ�\RH��z�=�G�,;eq�:��\~<֛�#���La�tMi�^���w5�rƿ�y��|7��9�����!˘�ƌ0m�1���H��4Ǝ��c&��D7�`"���L���η.>�hU��c���+ĭ@�����r�����%4�����+��!���z�o�Ĺ���_�O�s���b��kim�����g��_B����
�� �ߵ�\ʙ�d�b^K�T�F͞��c0}���$0��Lw�:y�N��G � `qa�{'�/�+��ͨ�9�#�X�~��e�ǳV"�g=��7n����n��O�lZ/|~�����C7�+��G?F�<�2�Hu�J�R��7o�|��	�.��8q���-��;����m�ē��r���g2�T�Z:t��7�+�c왑6b7�Dp��(�,����� �����u�x���0�F` ��4-2���T�沎���5��w�)�OO���D���`�UW]�g��>����زy�ݻ�ݽ����Ne՘�葿Z'�@0
zy�Aq�V�Z�Jf,��9��Q8ɿ*��/�3�F�Ў����-��M�g�-r�PUgvЏ�3��S1�e:1c���1�D!��.�E�4"V݈��&6�    IDAT1�(+���l�p<��+s�y��i޹RKU����,k��x����R.������P�/5p|�n�zj����+-_�kZ���埓�HDҚ��f��ڠ�!��Kn�~�ݐÆ���m�J�}�D
ȧ�uTU7`��Mx��g���ΰ-]�ʍ�EC)9����R|>��[�v�]mh^��څ�
_��&Rq�T'`nݺ�������E6݁3'�S���O��"/�;}A�
Q�3E44�⤙���u�+M)�ƸX���mZ&�=͖^�[ɋ  *|����O�'�F�P<D��4�!�/�2�����|�L�S����ez	��wU�������_T�qoLA�C��XA��Cy�K�����|%kS�2	���g�ƭV�L��9�I�X�v�Pd�����ӳ�z����,�s�F�P�@߱#?�k�a��V����g��������i��=���'��O�fl�(0��3��"��aX�p+�"
�(3�`+��n$q1K��\�$�:ȏ�y�6V��4o5�SXB` �oni�~p��/���3jk-2oZ�I�B���r��l�
�޹�<_ח�Gn%	 Å�@/K�)������?�ً�h !���2�Y�C����6nي'�z��$Ba���p���1f�XdҎ(�ii,ء�G�
��:}h��v�Џi15*�����ػ7n�?ӧ��I��ǍǉӧXrD8��c*r��,�ٜz��5��+����c�f(ȇ�A��`v����H�6��x ^/^�{����'YR:KTV�>PПn�A����+e�w�V~6.,C�)3%�W1
�L4��*�#)�;p,3RE;��s"{��2�'p�e�_�p�u1�U��#�w��|���j$��رk7�T�Y�R`�Xv�:
�T�hXiL9��<��޹ۇt]lh�c�W?"!Ge�HvPkl���k�oτ@����$��#hjn@.������ѳ�s驝�Rɜ�|(���'];Ѩ#g����`��b?^��!JQ���tv5D�Λ�"W���4�
#p�e����"/i�^
N��i���J[J`e��xj�fJ��o���6y�
�tM�k�tHiJ�R���S)~��?)����N&��N�F�
WYos[�� �H!V"���#hjj���G�豣1��s0bD�-b�&�@G�������7~S`�����%1O�����r�e�oP>eA^��ٜ�1�Ҏn�����|��cu�ً�Q�8sYa[�q�- ���:
� � >�w�gT����}O�K�\b	�D��*{/�����`���x�����N��[
W&�᭭8��3��:�t��+-�i`X6L��u$n�D�P��ތ!	����{L�����a@�]]��gFO�˸ TU$�t�?\L)�"4o�SE:����k�{fΘn)r
R�`��,Z���v�!��"+��O��%�,K�x�����%ȿX阞�;R;��[�>�j��x�K�;�t�"38x��딿�wޏ�+��5��3��Vz�W_w��������RN��}l��4����Ǿ�ml�Ej�|�|i*Ϣާ�x�/���ۘ��|�����t��c<s{�g]�[��7��,�h�z�����wߋb!`����(��DCat'2�j����t�"�[�]��j�c����k��I�����5�� 8��;X<��q���G	���~N����>��!�����b�ݟE^�-�7J��܋L�t�����(䄾�k0m�q�1P�3��}o�ހM^���b-�T������|ģ��r�x}��e�9���(��ln���<�1�&q%���D����5�*�����{����ꫯ�s�������h-��4���f@2�s�������o,J>�6��������]>�t��b3�ѕ��3N�[=�'uD >��7(��u1h�̸#D�~��]3o~`�!��?l�� P(&m3�Ǎ&R1����#9ʡ�;��H#�A��n���Q�,��:�*<O�ŏb!_ dϗ�q���E����X�
pj����ek��Ϗ"��C�_4�y�	���2W�sW���S���Q��A�g��@��5*�2�.�r��vr�}�qN�
�f��h7?n�
șu����}d��d���B
���(�Jb�I
�5k��?]��_˥oz��t_ݟ�{��ʲeϛO���G��$`�u���<�����������u�7p�N�gL���^ U��woL�g��{Nq���8��_@??c�n��P���TWע;���K�3�i�%@K��>AG���5҃��?��������\����p���"��D0����²�F�le�y���	3����)S1|�([l�,�]�|�M
?�{��Pr����j��U%�O~�S��\ ��4P���'ٙ
*�i[���Ի`D~CUHrQ�r���]XR��~_+�+R+�
sA�cˋ�H&�6�Q�E�y f.8���,V/P0.j�N���Q��[��aaN��l��,'��;>��ʆ7��;>�}j����̆�.Y�
l6��X�h�)�%���6z(2�iS�dQ���&P��p�B��}���s��2�>���RiLl1�$`��������i��tPd!R>ւ�|V��/WcB���B1�N�0���=8ͱ�w���~nŜ�)�.�bP���kɕ�ci�X<���_����w�{�:��c	jn�l�*d�7��dZ5}Y�
���W�p̵_��A�We�]����u�x`*~׻�X���	��.{o(&�z ��^���fR���O௩�K9���w���a��عk��SScƏ���3N�~�������sK���O������:�ނy?��;n���,���8G�>��C���LC۲e�|�Q�;���0�����ο�ǉ3Nø�l�R@��G?*7s (35졇�x��i_�U>w�\9�L�,�O�� %�kA{ϯ�a5�8��6H�Ks����ٳվ��B*܆�a����5��!g-n �Ԇ��#	
�S{$�dm�>ט��:�l|SH r��M;��A;߹-r(�]@�.��.�Ի��&
�a�%����	rL�%�����/?r)���!�r-q|d�p,,�C?p0�xe
E
K�E�\|��ˢ�,�Hԏ|��K�_��~��s`��Y9� >Q�	U~���06W�sI:�Ɓ�E&�:�����
~�r�oB�ד
�s~ow������(���|�w�C�	�r-վ�/A!�GkQ�@�W�C��*��Ԟ�P9u�)Fa�����Q�����2�g�����g���n��I�Mwa붍xq�2�]�Y�c-��s�4kƑG���M�X]$���7��'�3}5��_0�����gZ��ITǪp���ٳ�J'��Վ�;6a�ڕ�XҜ%v����ޑDC����ך�g����g�d�YH3�.!���z �+'����ȇ��\���'��``��kj�Vֿ�x���M��9��,�ȣ������hf&����ȕ���g�,ɥ$�1A��1wF �l΁-�P0Rr�el3�	v��c	�sHf҈	�A��	������cڤ ��|�H0T�hx�Q d�����~ݿ$t|�����YՏ*ӈ�'��I�܉hU�	��6|���m�Fb�:��Y��C�e`�-����y}Z]�R�!��v���>��6�����|_�o�~:>G՜-�.����.}���o�G�����/o~(ʆ�xȚ���ۓ��������X�E�l
��*g�����4˂+Q�H����)�bj-���B��/�Ӂ��ͣ���ǐ�¢���g>��F�F��R5Y)Oz�����>S>?���5e>�B.G���ذn��چ*r�\&�5��b���v�L�s�F�Θ�/�+��)=Ͼ���1�����ߏw�o���S�rݼj����$��a4�U�ww�S��d"���6��&����۶�D2�Î])\r�[q�Ygوs�٨�����G$p���[���Z;"�Y ��w���hCie�@�/ ��UN����t����H�ՍƦZD��X~n�u����[�)u�+~�3��O],�@Е�s��s�s��;���Q����(Z��I'�� �pO�����\�֚�F��Ӊd"��a���]�W@�#Lh�K&��8] 4�0���sYz�z���6�;�C�lٺ�R[Z�͔D?���_&ldb<���	�g*�A$\���v�wU�0������%�3�``n!]
9���v���)�ڣ��khmѰ�P������u���;�mn5���F��b$�j�N���o��xI(Ïp��d�w�Ecc���e�0Ǎ�fKZ?���\�,�0v��_ l���xD�Ae%E)�Rp�n�Z?X�_�Ϸ��(��8��5Z4	>7��I'��/����g?kV�R��\<��<r�n��ғ�2��y�F��1���-�͛v"ѝFWg�]~f�<�((�)��寑+d�)B�m�q�n�_�����U_!h��Q�F�s�������v�0��S���ֶ��7�`��lټ�`5V�ۍ�Ǟ��~��f����]�(���G>�[lq�zR(�˿��� >����~��D*gn\o��P�}�9�����|s�<'�e�П�!�u>��[�@�B۷�㩿����{pͻ�j�'���R�r�_je��H����K�੿>�a��8��3Q[C��TbOp)�-L�n����~[6n�I�gb��1�{b_�B���{�X��R˪�d�YhF��T9�aAD����]���>�V��g�Css#�:�4C�
`�8�A:�3Mه4�LWdp�
�x��'�Pi⤣q���/cq(���A��OR� �q[ :;�x�'�Λ;��KY#ΏO!@߹��KMxؐ���������SO��L���5wV�*��P���}x~�Kv��SN��)cM ��a�@�IQ�_)S.��aǮ��랽����X<����8��	���o���;z?,����5F�C���s}�k_���>����Y�ϦM<�^����FMT��ɿ�c�D;���?b��ᨭ�F�Ƶ���0���JᕗW!k@[�5v>�w��^�;v첖�[�mvsPR�z5��_0�{������E��TL8f<>����V�Z�g��N<a��v�؆T�u��ՙD[�&���qL�|<>������I���B!S&ӹ����'�P0����C�Z���Be���J�/]��WҾ��M�.-���@��-"�9�~��Im�\6��/��IG �ڃb.m�j_>l�`A�b�B�y�`;vv��G�!���/��p��@�im�&�F�`�|h2S���kVo�#�=�au�p�[/E>w�}�8�R>f�d���?��#X���q��:�(�3=�{�=��.��L*��}��q\�΋P]4�`UU�4g��JUz�e_۷����?��#G��K�"_ �e-�)�r�&�g9dr��b@�����59n��v�t$��P`��#닙h08ZL�62�B��r���9gOGsK����Dssn�S*��*I>G�y�V�}ϟp�)'cƌL1��ǥ�z}�.5�M!�!��%�-�O<�3�:S���v H� A?_�b*�|ϴ��c��v,Z�8�	��yfS#�Z\����^% � �� +����-1� �����d	�%��#F��v�l��n^��L����-Ƨ����OE��?kּ�'�N�6MMðr�ˮ��AgWk�lB&�N|�����_Cu���.������+ʬ�ڻ�̟!���>Ǖ}��q���o4M�ޭ��Ow��9�M�ݲ��DW��#�Ύ֭k3�߰1�	��7-^��� ��M�� ����ċ;� � ��A�3!�23�߁}��\���Ո�ʄ���_�/�8��Y�8�� ��c<D���M�C0�3�~[�ua�%Ȥ�����Q��ȹwf:�e��4Sr�(׬m�c�=���:̟w1�$KrJ�����ӓF��j<��X�b5��9�?�l�U{�h�tG������,��YtttᲷ���z�I�O*�	�ְ���lX�>�c��/:��=�D�˅�D2�@$
�$�r�0��V<��X�v=��0	g�5��N��R�9b��~?��\���6�����~�aÚpڜ��:�� �RK��y�Ɲ��_1>�c6mڂ����8�sp��Lw�Ͼ/��K��{'��!�z,_�
�?��<�TL;a<ry���A��qə��4��wo
-z��.k=
��rZA�V��>�����Q�>�W�J%�����X)ۇ��~T�W�5�D��/Z[M�a;����wYV��X/�y�[�����N�3@W��5+���s��!d3�\��l ]�Y��E|埾�`�ʺ����?�굫LY�{�/�������@d���#F��|��e\��n��4�8 ����TPƢ����[�+D�qs��x
n��F����n/�2������6,\��x����9g��{�5��m�L+@���[�l���c�+8?�@)n�]���Z�3�8�=g6��X,�7��#�4ͬ�1�7RÆ�Y�ޓ£���T2��_~b�r�����ϥ�Q2߶T+^Y���|��:\�ˬ�]u. O͛�T
�]J��F��ú�m�5�$?}�{}�s'���'�s�JK>C|o����i\z�h���=�����/C6�|�e�h۰�-�*��r��"�NWe�u�.����g�o7���X��q�_�f.�c��|�k�1�KQ�b1��N��f:+5�?���w���0�1�r�-K�.'
�_v�"	 �>֮Y�|��~�N�Z��;����Rx�o�G�2�=�|�
K��h�������cǘ_��DP�G�>�y�|��?Sx���ٓ��E�ބ�e0��;�̨W����װ�����J�+�{*��
��J�KqM�'�?�f�2w�ҥK�eFk��t٩����i����	ذa�~�^�7�����/ K~.�zC�wc��G�c[5����'>���aX�n#~{�-�M���R��b�����A��e �`J�>������z��]x���8rT���]�{M������љ�捛�i��j/����5r�Pkb^��f�?>^y�#l���W��c�a��ٸ��������M �8L�
�-i�}��p���bx��U��3�.�ɓ�@0�u�UV.����o �?ņ�x�ѥ�z�;.B4l��������X�ڳӹ(~0E�P����.A(\�K.��/�p���L��.64<�ebVK��۫�x�_�~�F��'Ok���"M"/�P[_�\&��D���5�"�L��������s�%� VC-�Yg�nT�� ��a�0RE��*{��X���3;����ٵ˄K0A6�<�����ۑ�&QS]o.��x�<�֬^�Y��a��V���teutbյ��l7������*��;���=6�����OPW?��2�v�4����~��]���?`ƌ�s�$:��]�1���z�5$)+��T�a�O��4������ǌBw��(��6!���+�D��h�hG
�0v�N��+���E.�L(�]q_��G�sޥ��@�k�B��ʖ7[HnQ���������R;ŧ�=̿�׮]kץ��Һ�3�O}]�~�>�.��`ێ-�%M7�ջ�CX��{�ص���}�1���Z�v�e����^�=o��/5J3�|>\r�[p�y� �����e�b������2��>�5u���@ۖ����_�N���~��X掸��կb���fR�8����$��1����shp�H�e��.�/ҫ����`��-XH��gҤ1Ȧ]Jlk��6����G�Y��w�!W̠:V��;�X��Id3�u�y�U�H�hEZ��Z1z�K�?�^�;�	�PUU��k���Ï���W]�6�	�|Y�=b�}�Q�ݳq�F�m���mZT8T���[�5k�aΙ�b��#-x�L ��Mhmn�豣-��qs6nX_���~�b��O��@����CJ8A���    IDAT�������l��=;�m�f�X��b�Mx��'��P�K.���_,�b�w��13z��֯{�V�������I�m؄�'LŌ����k���c�����Ƙb�q����B(�@���������a�Y3��\gV�)�5c��񨮪Ǯ]۱e�Z���.�T�~�I1k��Y�`ֵ�y�9��˦����-��=Q��]V���Ą�c�򣻫Ú��6��@g�[�m�Ν��L'	נ=��,B<�,k�ƛS*D�AyU�W���ڂ��H����}����?|_i��!�s�e���[�j�^V��|��!�
N?�t�T�g:�n�Kصs��@���Hg3�ҫ�fV�K/�6���W����܉��.,\�PO�Y���P�oni��������1�A��uj����x�ϓ���ш�n� ���ȫ=��>�4^X��Ip"���>� N�}:&N>U�l����I+A�L�d03D���>6u��0b�H�[�� h@����ޟ\DFJ��~>ܜX�:m�����X��l���w�-s���I��M��L<u�����8ַ����]����)�w�"��_�֋�P��a��5b�䩨�kp�7�70f�<�ϊWV�i�}�jq��������Ǝ3�j��Tr�Y�ʺ��I�i�},��U�0��,;)[�"�ǔ��[u'��\N�֬Ya��-�:;�x聧lc�����\�8��駝�|�o�[ca�%��3O����m�_�����!�O�=Z�����Fw"oEl�\�����+m�؋a��Eذn=fΚ��'M7৛�����8�����b):�v#��Buu=~��[��쬳g�e�0d30�9u��o��@8��ӆ�<i�Z���W�5n���'L7Z�L>�qG���e�3Q�*ڸa-6o]i� �b/,{�=�8�;�\L�t����Ģ�8y*��u.���GWW�7;:��ol.|�l����c�1ۗ�1�_�ֳ��c�o��,)b^k��\KS�Y����T\��ϸ�<�v*�&����F��شq=�a	6mjC!�A�u�˙�Hkw���8��3�٦r�=��w��]�v�ǧ��?����"���l�5uHuw�8���p�EZ��ݝX��9�̙����S�Zpgډ3�3���n�����ؼys��YY���������"�b�Y��O�w���\D��SS؟�}��I*Me����ތ �s�������QG�1�3���N9���
w�옝ǚ�+L㣏���E�6��[�z	jc�( �#F�ńc�������*dy�]���=F����ex������dc˴A�-��`�6ړD%ScGb/���æI�U7�~���u�}�Id#�5���N2_��9f�6+W���V��Dx���gA̿�\��ģ"N:�TD���,hcЕDy��6�>��ۆ����g�Gĳi��@um���#�M�,_�ľ�Фe�K/c�ɳp�qS-B��ة���[���֬{ъ�BA����n�bU8�hh"wL#F�������+���M'���{v�et�btIΜ9�O8��+hI� qԨ#��A�H8�]�����9 ��^Y�Gys,�j2��4Z��q��i���?B.��/����L(�^��>�{v�j���z�`���_��_���Z�5n��3���֯ ��?�9ۧ�����I�?+������bP����n�E*k֬r�D��{��ZP��9s�c���1�-��H$q��oǣ�>�)�Km��A��@�@>��?v�����;�\ǟR*n!�15 ��ј-�Ԁ;w�4ʆ�^z��wS..��'L�����7e���5�QV
NБ/Q!�����ӹZ��)!3��4o��g��|s瞅Y3N,q��L�oji��ˏ��V%�k�V�?����Y�=�l=�HG��Bc�(TU�ώ���S(����c1m7�{���G�Ōf��u����BC�00W���8R(sh߻�,��K^�Ë�9���̓���n��I4Է���,1��Mw�5�hߍ��^k�I@۾5�+��#��3�c?u���kh1����WU��u[����2�}̽�|�9�]{m\he�@2�t�w�EZ��oCw�?��ο�0a�DTW� ��Y�OK�&�
E�2L�d�;en#V���;�c[.�w	F��6�U8X���ᨎ58�K��H,׍ή=�h��K/��SO=m�o޼y���2¶P���Z˰���u�T�,���N��)�w�h۸��c�%f�dShj�Z�2;���YDcUH&��s��3	�}���a�fd�yK�e�?W����wߌ#������Be�y}��3%RhP�E�u��FL�"�Db��(����V�y睇�有h�4�R�o7� �G���R>I���Ltw㩿>a�E,2WR�׸�J������7���OM"��t�3�	J�?�S�֙��,���0�E��1N	ݨ��}��f�o,�Rր5����rQ0����9MEf�9��/e��g���(��L�C�|&n
ˮ�pՕW����@w�����K>Q�.�?�����"���M��M7b��H���e�����;j�Q�2�̾����sK�����_8��0�����d-��M3E.gi�N�8Ͷ�{���m�މ�-Ɨ��O�h�oFu55_f� ��U�1��&�Gx��'��_�����U��,!�\��L��0��-%0_�r���
��w?��O8��Ӎ��2_��1�ч`�u�rM;�&���g?�)V�Y���w-&M9�h�K�D��'��j*(X��	��꘽c&�ړ#F� �l�s�C,,еBM<C-�� 
�<>���z�U��{fO�n�,��9��S���4r��ձ�(���o`��Mx���c��wOյ5�˰��DB��,��*�4���;��o�4Z#�DM(H�z��yy����ތ�5��M��%���ܫ���-���ζ�<���x.����*c��!Z�sΞ��g�RBp�%����?T���1�F��G{�^hB��6���"��ń[r�z�5���T�~��@.�\�}�J��Hu'��@��#�iy��H�B]��n�fA�%K��ɕo^t�ܨ��\X��9������^z)���
�F�lق���[#��G���V�'`k�_����T�.����@�wް����ry\~����>�qJ��aʣ�8�'�p���6[�KKK�}�{1bdS)>�F����N�s��r���x啗��}����y�7o�c�$�u5+����L�|2���p����w[�ͧ?��3
���8��
8*
Z�Jv�>�X˖?�[n��=i|�_G��<�d(�ppEZ�7[�TM����p�w��{�ԩ���>`<F2jst�T�/�\�b������ ���obÆux���o-6	�|_'����	���eEV�`���}�߬0�C� �Zb�V��#���F,G�P$%C�����L%3֓��ʀ廮yg	 E]"��3��T�Θ�
�mNw�܍y�.��g�m��9����UE1˭�.|�_0��B|?Ο���[kwO/�����@� �G�2)OR����`���c	�7\w=�=�XK���c���5��Y�O���B���U[[o�>y�dL�t&M�d������L�,e���|�)l޲�h������
sO��7���6s鳙��L�&��<S�"�*�U'�{���䗮.�<�6,w��=V���=��w��]��f�� �3������q�@�[�8�>��{�\^��3��mWX���9�b�JI�GkJ��|7f8�}p�u�YIw�l��Vk�n�Oƍ�ϲ����o��/�%��s�W}�@��>��������+�.�m��vwZ��EpV���Kˍ�+�̚�B���j�g̜%��	aG����\�Ɍ�p��Ԟ%�պ��b�����������1���q��e���]�������|�Q�Z]���C�z(�'Y���*3o�k��S�rt����OBC6N��Hi�^0�k�87]ݝ��׿n�T�gS�S��"�ý��<^~ �oޗA]���7�lV(Ӻ�}*��r�������q�l>}.�G����ɬu� ��i.g�K�?:W�cj���|�u�p����-U�
�mQ�g��"���MWcN�?��?`Ŋ��;0q�D|�S��2m�iS�I��r�G=L�mj.Ϋ�~��x���ֳ�y�6І��o|Ê\�r:z���p��ӜB�*�a��͂\��R߄J������c�Y����3�\ݻ�F��X����.!��\Ι�Ȕ�}�=����fw��ח����	Ǣ���^承���5�	��ZR%�/p�W��SL���8{�7���\s>yi��p��'�ۇ
�2U*���;�k��`3�>[~WIx����S���]��z���>��h^��Ũ�A��aP�B���O��O��3œn^
5�mR0+�G�}�kMy�0SkC�$כ�޵��$ �����n�����������p�X������<����޻��x9�,��O�Q:���X��O~?��O��SO�F�R���9ܸ�ٕ������fk���ݍ�����J�����GW"� �]�����C�5�����0p!�s�y��>�7�s��Z��2��k�E���6��s��eQ�gq75�)U��[g��q����,S榛n*[w^��2}J\�|>+7�O�Ss��M�Vp���y���l�|^*�&�k��XI��k��(tLP��Ҝ�7�T|f��_ti��#KV��+i��%�3��?�߁������@��>��WZ��?Z����g̭C�g̎���ts�QY���s��ˊ�Kq�
Y�"y�>�?�'&X��N�﷍�~�Cop�?4��c5��4�}ьg�We�X�/�R�����4N��J��1�!^��z\�W_��JD�'�A�K.
�?�;Ǉ���$p]{��S`���ečB<���E4�p"ë4 �ݧ)N���}�ƍ+��qC����H��y�	��ɭ�}n�� �����bޗ�?��,i���:+Ҳ��$���
��j�^W�B�"AR)�J๪ %�����r���T��S�j���eM�	{^�;��	׃,!��[�x��i��)P�Q��?;����˕ƹR�W
��k����ה�s|��x�	k�Ƚa�%>�]�F���ԓf�U~dux��!���h�aY =-��&m�m����F$['9��`�� B��w�X�e!�}��ɟo��?�ϟ`Lp��T�s��I2���N���DN�����G���l�C!z��� ;P7[������U_U�����X�?�~��_ۦ%��%����njC͟�d�,�� .2�ļ����PY�CAI��c���3��4Tj�^�qf��`�K�}��Oa���,��֟���1.fi=��~��aM�XZ���������{���l�e��ɱ&s's�Y��:��)��b�.!�w~�N�JH��Y��_�u�[��������i��X�g8���?�b�0��H>����%U/�MB��� �<=���^ӫ����ͮ�+�Y�\���,t��(��뀚i���$�q�8�Y%*��1��]�a,���{��/~Ѵ4�T��Wr2�-G��[���	qik�*cD�A�=5�z�i�H
��n.��el��.����O�����e9h2t7�閠��?��Σ�e@� F0�Ї>�Oo�Jc��p'��y�FL%Gn����z!�݀�g�u�i<^�Z=�i�󹔦���5ſq�8�|g�>�@�8	2�Ko7��u貚z ^kDs�U<��z���޷T�{��������������$ؗ�X���:�O_2����4.
Uj�	�<N��?hr�?�k�߻�}B��]���]�8��N	�D�f�]�L��ޚ?��c�l+1��tKP�_J�/95p�ɾ�8���ÏW���ڠ��㩽3�[�L#R����I��k��V��S�3�ր����o��4L��ILŀ<0������7O<����]և��g���g�	c+�w�
����TO�+��FA�Ɨ�Qh0���)Gj�{��eE����_��=��y����j�e���d�p�6�;� �  -J�,еT]O���'MS8#�����/,p-y*���#����;��������.kS��ڽ7��w��˔���X  AN��Û�9�f��	��
�)�h��)��{z�!����� <� ����W�}�9�=�I�A	������[np
 �'��&�O�;��;��\��'�+��c$���}	� ��Z��b�6Xa�M���!��@�^�KS�'S>ǅk�V����/�嫴Β�q �+~�ؐ��v����x+��9�Z���)�%O�'!�w�6�h�Z���s ����pK�'ô!�D���+�Sօ6�ib%��-��e�-�|���8-N<���� @@��`/^ %ׁ�&z�M8������;�_�`����C'�D��Sȹ�G����0G�����	D�M
�@�a�����5���xǍ�4i�;�8N�|x�� �%Ùw����j��O�^vdJ�q������'��&L���H�Ф�4���Y�}h�|@#0�4\�+�b�=M|P:�,EU��v�.���T��J�r���6��L-���W�Cg�qo�NU�e�Τ'P3pK�?�2Y��L��1����5}Q�������a�)x�
�x�J��\�C=4C#``�(�}/�v� ���<NBA^�O��z]���zPk��R:����'Y�7ρ�Ţ8�9V� �	�B�-غu;�[�Ě�����M�''�Z�R�zg�ȊP�N�ƿs�9���|��ch��#P)���׊�oJɕ�/OS��3L`�8@a�:��޲�z\�.�Hx1�����r�m����W�]��C{�O7P'�t��'������3&FNYɛ�((Ĭ���>���◿�\r~Om��}s)E�o� �<�N�1���+��Ga�
C#04o�(LռJ�^��8a�8��!y��*Ͻi���1]�B����Ć�ͨ��`/��^{<��J>�P�eeĢ�_��y��s�8[�������	bfN9���햮&>
o~/'�����=�R\4��L�!�#���=�F�Ў �CY@��`vi0�2�|������V�R^�J�
짟~��՛��lP������nG{�#���2诧����_lz-M��7m�|���Y:#'���	��g�2.wJ_�U2��Yy*�~
^�a<��y�����GB7Ѿz��eedV�e:t��������U+ �Y���8�����U�KE��_��f:,DzH'���Xu-�i�4�J#0o���������3�k��Ϩ>����4�]��h����O?�-�6��C���c��)�����z���D�NV�R2쯺�*+���?h�b� ����}R<f�7o�;5~��Z\�P����8�#0P���7
�*������pԘ��
ho߃��_���/�9�$4�c��4u
N�>�N�2X���F&�c��{v��;��U�b����>_|!�?���GG�.lټ+W,C���+״�]��/��a��=hj��_��r�.��S*��6"�<�<I�JA@:���;����Yu$�>��
)�W��C�d���f�J��ߦ����o����ys�	�T��=���d��*b|�ᇍ+I-���,���=�C�,V���z\'������L��p(�DW�v�1i�4�{�\�&�F���� 	#��b��f'����y�e�+��6K�[�p��cxk3�a/�#G�!ѵ;wnF"�i���c��{W'��rؾ'���0>Jb6V�_�B�yK���ok���3 i�#�7}�C�."c%3�xi�io�3�t:C��#vx�W���2�L��� ���q�����yZ���v�a�
;�>NN+z��n�_���N��X�a!��g�KN6�ö�q$ytv�p���4������� V?��R:iI^�7�������s�W�y    IDATq��{�����
�|�tn���s�I�6)������=�شq;
�0�m�c�)s���Et���R N�.R�ra0����[p�h��j����xQD��t�!���n�7�Շ���5+^��N�\�l\3��#ͺ��ץ�;*rO�Y�7��Q9���?���[:gW�<���3��uQ�X�"
�����](ॗס��	�mÉ�N�o�d�ܼu�%�l۲���{�J.�\sK�����m��o������!��z�أ�~���nj[���g�9�|7�n_�L*iڸ?@n�6�����6�cܸ�֞Q��_���)[L�z�[�b@O���"sz��E�����:(�;yq���(��\��o�i����5��`P6�ܲT����O>e��dOe"��(���iՋ?�$}TIHw�S�ߋ���ں6mZ��nrd�ΐD2��ϯB0P�ݻ��|���~�2|�E?��f�Y���D^E���������f{{���}�l�Q��cƖ��W��p�ٳ�Iw`���Hg%��:;��~�&�|�X�������C�`o�(jt��[]T�Ϲe���i���L���RJ�����������P(�����P=�`��hY�1N\<ܣl���6�ai��ʑ���I��fNl]��Mvu�����˟��܃N����jlܸ�{��J��o+WmD6�Ggg;v����/C�%�o��k�������#�Jc��1����4��R�N�~��p֜���Ѷq5�.͓����q�m؂L&�u�:p�)g�{��y���;��'�D3��6w����L�`�L��9*4Sw�����{���{��4������¡r���_��/��]~�=Nk�,����~���]�� ��><f��x|�]�4i4ZZ�a��W�˧��`c�4��+���Ua���5���n�����;�������imn���n�y����������-�i>��`dK3��<^� F�jB�Ѝ�{�!���y}~?��3ؾmv�N`��$\�vK�$�3��\4�.�"q���ӭC�9�	�����;	�n��~�LM>���c��^�(��}�ڱQ��.��7~�������;�q�W�ޥb���g�q����E�̚�`i�3`���]X��"�TPc�捌��G���;;�ص�\x	�=�D�bx��p�-�X:���+e�Z��/ۇk��<A6
a޼K,�3�Ma�m��ٻ{��B��k��<�gG�6lC8ڈ��q�;'��o�TOQ=|�k_3�gF�z2ݓ�AGaB���~`1 /{���6���A�zd�܇�y�ߐ� ,�_���"�̦3�\bꕀPU.��ty��M7�d�B�5l۲{vmEGG;�9�����l�p��֬݀t*�+���ǌ����nK!��������o�����?P�o��#�3a�x��w!	��&���������Ĉ������Z1�ē���	��g������ގ���:�������N�nQ{V������K�ސU���uoٹ����j@��U�C�痦"�h/Į��^'KJǊ�[)�bB��\����MT0���(�v��y������y}��N[��Z�I[Ԇ��[���?�2AҎ�W�H(��TO+D�5��i�0F���K�E(��3a
O�/�@L����;��{Cc�&6�{;�ʚ�R�����uEE�)�j�#�@֬�-���zy8��_����g�{S{ϻ�1��w�m��T\T��I��S3"V�~���<��/�͛6��/����ծ�u*�A8�$S̘q2�u����mہ��zK3�{�R����y��?���R�7��ۀs���ݍk��N\tх��E0�����F�����{�PX���b�'a��3W����R5YuG��6	]=��ԧ,��_�2��f�i�`ж��|Ŭ��������ڜ��`�^���q1�	U`L�`p�L��t}��4����м.c*e8H#���ܔ]t\3���@J B�,��+}O�ϟJ���Ϟ=��*�CA}�(K���^>�hx{[r��#�c����	�us��GY�p��[Q>��_i���t�h<ԉ�?���ΝkkQ���i}�ƍ��̵*^)i�<O���֐�U�\o-���i��IF6Ї�s�g��SO-�K՜j\U��yb�<��wT��~��`��E�G�/�������'5s�?���bʔ)`;L�'A�}�9�=ʣ�c�����D�f�j���{�j�
[�&p�>���KQ_7d#(|����Z��b��c�����h�hR6g)V�lʢ�'N�n�܈�H��,��0�� ��"",��Հs۶mX�x�i��(h+ �����җ�d������Y���H���j=��{��*Ս ��w�۞�@��'P��gg��-p<�
��g�8Â�
��$�%W��o��o6�2��o�G$�]w�mD�e��w�	�����a��s$�x�)���i�eG3��T�Y)ܴ|Ư��e롯���~̸��n�^��nu�i~>�����M���c�# w�R$�2��*�'����-�%�sK�X�I�����2��J�*�4Shm{�y9�V����&��@��~�T 4�R~x-u�b^�O<a>u�[i��`�`�x��kM��t�R�df�=�̳x��l���
�����[��_��_mdAr<�'��'L��"�t⬝R��'.f���/��K+�;�S(�����/�ws<�q}%�_Ҝ�C!ׄ��/���/�	<j�X+��ĤS�=��ng�Z�Ҹz�z�ro�>���M���}C��Y=�<�pT��i��]o��4�ú���4<��;��P�������*�Z
L��XȦM���8�K����c��/8.�P�|�[߲":�6��κ�����y��n���sx��|�,
�����YL,ܡ�ƹ�Vʟ�'���P�'����:Ӧ5!W�c�����'>�ѣ� ݝt�鴍g>Wj���~�,zx12� ��"��&���4�\c}��$׮_��~�����3�
	�a�?�S����Ϳ��q�1��nPo�y_뀱�5ZT�����߼�M�b�}T����*;�DkF��K�Fp_�z��w�'�t*z,� `��:�ݏϨ����;�-�<y2����@��2�@��d&��h���x�������y���*��d�m�w���?�wį���<�M��/���b	���aĈQ&�#W��c�m�b�H\\�r���2k�,�`����	&4��{���{����a ���X��k��|j!��%���9K}-��	[�)]e%u��i����oV��y�j�/^���{���J_ڧ�Ҕ)|9����%
�4�e�!����q�Hx	�5��X 3�.����b4�K^��||^��8j��}w/��9�т��z;Ə��ꪘi�Ŝ�1A�߬�l��N��~�%K���b96����80퐂����y]�?߉���_X�̲�<<_��֯\�\���ϟ���>�ƕ��j>��y���J»�:��B�2d8��I(��k�YY@�5 k�d�RYܡ��^UV�u׾����rl���%v����*� ���SӦ��jL�:3N�i����Z�\�(�
ؽ{�Y�_|˖/�`�Yxp��IH�ߧX,f�[Zo���^6�����W�` l����h;%-?2���}���b�č� 087�|y\�
Ԋ�� C�+]�r��Փ��:s�L+�b�@n-�}�C=4K���"?�Lpj`|~� ��ǟ\���h�`z%�g������ K��UV�5k
��AG�$�;��I��97��xg�mJ����^ם�W�����1�t������T\O�J��}!�PЇ�G�D,Ze׬��3��s���Z�w2�l=���� 	���"1#���lr����u(5>r7�
'6$Rq��Fg/�*�D����1�y�ǖ ���WZyA��N��8����\^|^^��*/[��x���Z��ť�����.Ɯ9s��X������~r�0�DE���U# ˓���pMM-fgry
��)���q�;�]��/ 
�?�p�T_�Kk�����{��_d�h���v6n�w��:l��6`�~̂�a�	|4u��5�F޹���h\,��c0�~UnP��e��dpL����IVgi[�78d�3���M��Lݔ����H3���+�?e-�R��@����~�^KMA`>���	�y�,+l���u��y׊e����r!�{�����5�.���u�}|��<�"Zʱs�Nz|���[��Cw:�T&mY�W�;m��#����!!dq-�)�l�("UQ*~'A�FD;�#���Z�^7��-ŀ�:Ї�?݈��y��'��\^��)6����-�,^�1�Ә�8a�Cʅ�C9�P�"�����82�ɖ�,�8]|ʝ����&L�0wkIY�4�C�_I�/2G��l	���}6�����28_A �w� ~�}9�o�<��XNjE�C�'5f|����P������O��@��p}/_����ƔF#w��@��m�k�C��8�jb�ո�	�x/�W���'���=�Q�,�L��|yms[T����+뽏6�4P��xm���_
Z(���x�Q�o?y}9㓊R������w3Ѐ�(|�XЕL"�ݍ��%BB>�57|F>��G�{��=��Wf�U��?�nP�}Ya��������;�0J���T�Lk��O�TP_{�{}	cY\����|?zo)�^+���|q�r��w���|���:�ڰ���,Θ���w�Wpk���ܰ�C�8>-�XUM)�9�B�Y���ks�u����@n��>���Uޏ_q%߾>��O����j>.�o~�.�\^��b�t�wmmm��HM�	�|z�q�ۥ�b����w>������c�F���8&qӊ�n|����&PB�2���9����
��	��1�j�����	_�ц�������]6P_�� �E#`?	�;ݎ��,A�� ��է2�}��V�[��|pL-1@<��2�4~���ZEWy�5�׼{�Mq�}
��ރ�Y�W�e-����y���t��Zpoփ�8�R�O��SƞR_��y�A���[0�g�xǵ�|�}�������k�k���11��c��w �G�r��R��w����'�&��f���iԇ�k���m����*ȕ4z�p��#����������Q;��W�ل�G �{�B	�$ zP��i7�_6�����{+��9���WC�����aN��{�B���L!fŰBPy��'�Ng|mK�������b�U��S�0���@�����;�C��k����iT����*��c=އ!Ϳ�ٚ�`�/�����^�/W�4x�b�?X
ZQ�C�!�]�J���K�0y}d�݆����}�f=�s�ұ\��E2�EE��"X6Iݜ���S^�}	�y]� �==ǻ�D>�5��o<�~Me��_�����p�L���h{�Y���8��K�;�w�Cm^��R�@~�ײ��!�?����>N���t���b)�3�C� ���>�`	&�B5����|�S!69���A�?�~_�P�˗�*X�0�$ �R�	�S�2�5��e_4����!�?|��/*��}z�?��l���3�K�O#������p.������e�x����W
��J@����A��3o@Ϳ�p9��.�n�G� C����uL_i}"�� P���ؕ�/����^�UX�C����:ʜ�ޚ����3��f���r�i�o�n9�{[O<z>����{�!�<���_(��1��7����qzh�;I�$	 �M)�._7d.Vs*7��+����a��}\@]�CK����+�?}��Z:�?h�>ݩ��;P�t�!�?p�}�a½�z����U1�� ��-����[���om��`��-X���x��*���A��9_�:���W1o��0&�������h
�L.�M��������G#~�@��+Ư"Q7�U���U,���7j(e�0E���������"P�~��������ZB���R�?��q�|t�Z<��*�Qі\i,2�Y6W��Ze����y.�->�ݔ���1�G�����0�^�z-C�S E�9s�(�O�U9����nx�p�d7�錍m&�~P	QV�����|V�6���J�9Q"��p��*k��s<ʬ��b�bU^
�ǎ���X�� �k<�TZSz{+�5��ޞ���Y�益=�{C�Z�'�jo�^Q���G�\�-aV\>_N�渲��\=~ �h����=v�+N̻b�e˞7�qWp6��?��y�"���������q�?W��E.m?F�����zm���>V�=�B!���&-�j`�&K��k�8��*�i���#��?��% T0t8��\�L	�ci���w������n,��R+T��Whv�L�6���U9����K'皙x+O�!is�oW8�tm`iS(�"/���=^��J�������E�+$^���������r�����@��)巪^�hir�Q�H��.9��8q���lh̩�X�TI��
�%�����sz]���~����|g��8�t�QPp���sq�xoS�I��kk]��������)o�s/�'��Ϥ�=�i�ڐ��U��.\GV�۝Fsc�1�2|ذ$Sd�u䆉�k��V�$�[���9\�\M<�p���/��m,G�Jt9���g�y.�{>��r�O:�4nFiuiv_�۷�4C
m i*� "��F!�	���w/�x�B�`��F"�i�RW�~��/�1I�Tۻ��	��	V��x��}P���N�J�7 ���#F�w��W��ss.�R)mb�8���;����x
x�Yc-�d667�S��ל���_ȣ:Ve�.���pu �Q4��
"�c���Y.���������:3-��E�,&	6�#��(���	N	X�{�ݏs�{h�Er�k�;����Ha�߇�E��,-	j��Ƿ��ގ�=^
/��'��s%���g���0�Z���ӊ>aډ�����W�.�h4�ؾ�:s���T�zV�X���q�Q��-�@�ɞ���/����x��>�>$v�3kcU��e�I3��oKS#2���X��Yk�F�-.��ԩS1i���k���.l�B�a.|.n�#�<�ƍ3ӍVB���M$-�C�?�:��~ ��MWGg���h��_<�V�	ۻ����{r3�1������ �U�oV��m�L1	g��ZB��TE@o�W�KSK�Ϳ�CZ��xe�\�Qy���w|G�]���Z���ޝ�_Ȥ��҄=#���]���=w����!��RG����f-!���Xr\ml
���:+a*ˇ���J�)	yZd^b;���8n|w�I�=	��LyǕ�	]�	bY�K�P�{o�Y�)���:֫��~N�:�����~�s����r��9%(�F���q�U{đ�DB�fRض};�y�i�w��Z�Ţ��;|�H{�h�Ŀ�?��'k�h�i n�A����a<�qc�oմ����q��ދ�G����(���c�`˖Mf��������Gy��v2b���nH�L�~�7qQ���<�_c�@n"i�2����5�v�����˟1o�E��H���|�I<��2[%��ߩu^xᅶ���
8R+	@���&�Q�)���x��)�i���8q�]OZ�W�P�}�=�II���^b.�#�l�C�^j���e��r�xP�����;y�P��B-͍��c�8��+7倾�]1�<y�]w݅�/�����F&H��ƙk��#8_����[��yK_x�>�h��D+�q�e��36GlIK^S�7ޗ�p�w�y�)Di�_��O9���J4^��uE�C6���l�Ə,$�}8FrG��ټEc��,Y�[n��L�,�X<F���1a�8�
i��	,~)^Y���&0�!\g��L���3g[G&<��_����j��F^\�7�s���?h��?�'�S�.����w酸���+f�N%�f��xa��,(GL�O-lW{J��s    IDAT��������r�����F�L'����6�}�Y�[��� �!7�c�=f���J�����;�k{�K�5Ea�9�6��K�$���{���\m�����5�\c��X�x�cC3�{��6m�\�*�F�v+-��8y�d�i�r+�Y�.
�qd�1���K�N�/�7�bw,cW,���s����c�<�쬪��N���IH!	%4�]P��2"��"
D�*���S��\D)6H �t, ��i�L&m2s��~������̙3%���'�̜����~������Q���ި a��}6��{�=���FΪ�j�p�~����4Z>��#�;�����f���Bs�8���2^��/Y�T[.ug��Y�|G�\g�64���˵��|3~uS��ڧ��ֲ�Ro��#���4S�Y����9R��q{)��T�E<�|����i�(Bt�y;J��J>�!y�'���u��qo(�\p��Cy�S��?����V��{
��"�3�.���mr��G��%y��X��t��Z	8���e$��� �l�Pe�w�o&��^q��2k��2]��c�� i@���Δ��6Y�r��tw���<��w&,�ΐ�9�<6��p�X�[@�Əf��~�i�%Lb����!|m�r�є�i�����y�W�blsr���qPbl�{u_ɺ1��5`��f7���D�E	��ۢ+��h�ԼV��i��9�����g��5��� �W~�����C�h۠F{�6|(���i9h� �O`�`lX�?��������t���K/��ӧ�����k�W� *��oֱ�/���	L���s�Ygi�l���1�e�*T��9��́�N�lNۏ�X9�kZ��0��DkHU���|�u�i���|��k�T�� �Fu۫~�k�g�ش{�=���|E׽�]�y��=~?��hw{>�=~�}③ll^,�T�������˜#�X�(/��5M�$���u媫>&3g�.�lA�x�or�=�H,��}n};#]��~[2��J�j�O�� ���ڨ�}�r�����r�rI��f-�M�NGd��9��cK}h�������	�S����Р��CM��S���3��r�����8E��̵r���1c�>����#o�q��hO �i{h~F�������K��u�P7���q�  |��6W�k��J1�b�?�^54f�Q������yJ4E��q��&(��Z�v���_j�E����瞳w�/�P��t����E8��Tł������ G�q^�*��;�MPs ���35�ߴ}s�+�Qp�6��)SJ��	_w�y�j��h��Dw���t6�6׀?=|�^0��7ø�m��+��_���9��W���UysچR���i���ӟ�eie�yN�w��Hn�g�zHƍ�˸	�d����U��tN�-]-�\X:�S�����sϒQc��ˋ^����_��͙;��ɶ�+�?�3,�ٻ�&W_�!���ic�<���r�GK>�%MkWIgW�ĢԨ��斤4�k�l6&���d���Ҳ����җ���'�E�hٴ,$۴��'NP�0-�4EӺ�Kܞ��s����cƨ�vb �wM�t�E��pԨ�ȖIH�ײV���h�f�"�\ )���`416\_Z�?�/�B�'�d=�����E��s~��|l�an�]��/��8-LШjh �1�t���CF��o�k��8�]��q2f�o�ͥY<G��9}���ic�o��8KN�~�X���J�w��-��x�W��u{��W��c���uO�ߡ�� ;��{��gk羦&GU�u��O|B��|�+�'#���3F�,}��ڰ'��c����"�iiMI,Q/����$D�I.�ma0{��l���G��?g��&����G��s���#WX"�����By�O�!��-�XA֬]�m1�
��l��.�6�O�F^^�V=�(�B�(,P8bQ$��pL�����Xx�Y4A5����4__s5A��-n�O7��1�	Rv^�����67	b�e���>��kn}�ôG]��xWz�:��1���� b�c�����>����S>���'��ρ%,q�\�:��U>��/�?��aB����� >���O�z�{3Kz{��Ӭu��>�\N#�h�������{�.8}�~��l}A�]q�J�-_��<��{�G�'Ə����)Ţ�ĥ�+/˗5)�l��)�Z;��o�Pԅ��䎟Ȋe�J}�s[�����j�Oz5u�NS��k>.�b^��.��m��c�L�]6nZ+�=�.����d�4��$�y�ؒ��{�E���*~4>�i4`�J�^8M8P�p���;��1���Ȩ��6y{.�j�f��Z�@�`*�8L�y��}��7�EE��iަ���>3���=�����;����Aɿ�	=�,�����ܒ���(�&����k�v.��]���+ 6���o�3��M �
�	�Jc���߿��*�����s�������2����� ������Ϗh(�2���X�PfX(��׭�'{P޲�,i�8ZV�y]2� ?#��lFd�+�K$Z/�YIeC��]'��Uo��fY�b����R�Ap�������i��}��1r��?*�u52nL�,��Sy�>�J����u���ۥ�G�	i� �[��+#k�&��S標�Åޙ?~ɁH��SN9E��Ǎ�R��[nѰP��\t�F[����j��&f,o4�������L0��i���f��`?_�5'���K�F<�}4��9���h����(�Uic��H����l�|6�v�6�c�='��} �4�V�Uc��߿����)��l��������}'�/��y�fY�M���j�f�� ����9��w,,z_��X|��ΎM��ӏ�N�GI"�ի_�Tڕ�A{OO^^|a�D�d���r�ۏ�y��֤?��w/���������3�gvĂ�i�7~��-yU%ڇ�Y��Qrּyr�[����VI&7�����"�0 �➡~��Y׼Q�6o�T:$W|�*}`<�[o�U����׿��=1�h�\r���%�m���.�C��k	_��,zc�x8�/�\��4/_����/[���[>0�Z5�� ��7 �/��|喏��]������<>�җUe��K8�}k������J��ӷ<�}_Y�����6��/��p�z��Z�׵G~��7_�~"��?�|����͊�Ә��@���j����ѾQ2�N��R��C�����BL򹰼��5iK���^";�<SCA~�a���%��T��w��u�=w�}{����/���xC�=ye%�ϓ��T�n��v�X$������MR�Nm���K!�x�N�;�p�m�=�D7�勉ǂ��K������w����%���A9j��x㍚d�S_���y0���Q9�].��V3�r-��r@,�0 ���%`/&tʩ!Ӽ����W�����������2��}��\�3��e�F9��[ff��c����W����TK4�ݗou���r_�9�4}�����$`����Ja��l��K�'���p?����K.��2I��*���חȚ����t9k�#TN$��ttfd�Y��A���@$:.��^eFՎ���77�a�e��Ͽmā�$/�_#k�9�t֙g�	�'�I��Eem�Jy��G�E�4��E���C<DN8�d�0q���&����s>��'1���Q��	���-Ġ_w�u�v]�j˖-�gc��e��+4��6������26g_Ԑi���� �\s���G����1����s�F]�w}�5|����[�3��)��@����?._A(�r��`�mǚ 1N��90������1�[}��h?b�W ����XC�w�;\ߊ��Ӭs�s���WK�K�dlD�� ��<���}�{�+�|��c��j��_�����4�]��� ��g��M�9��s�}$�/j��G{T��կt�`�/pM����M��p����dā�����f���*���k�/��޲�d�i�0�����.kׯ�H$�^���Q�'���x�F�v{�-�76 ��,��,:�a4��{�q�>,6?m~��w�߷LO�2��6�m�j������V�7ЄmL�¡ڵ�|>�����7�-_p�S��P�Y۹lN�D2~8����1�9-⬿5�h�Z���i���ߟ�r���{���)�}�A���5���kв����w��cʬL���a��E5���:���.3w�x$*�|J�I(]�\-�J��<C����Db���勲x�k��L:���Ek)���;�~������)h	�?$17gyW���c�	z�n3R,��ڶ�X��H\6lؤ�(�`8{��q�<c
�>?1�"�.]*].�Ӿc��@o8����w�\����\��U��>ܱ�����w���	Z��\)�u[i>�\>������KHM8p.~�4q��}�9��{Hm]��pF�Ơ�s���W���ߟ����w�a�}/����
`���T؍	r�TzB�ϸ����d�ӴD ��<$.��W˚5k4-�� �Gc8�st!|�ߔw��r�W��C�_��7!�?����0��l���\~��-^~�9c��(�.�n�3���1��3P�ӱX |ƌ�g�$.�x�����߯`mt��[��:;z�V>��#d֮��J��m<�%�)����/��ؼ~�
����:�{�
��Xο��kRa�]c�b�uM@��3g�t��ٔ
2��E ��n�KI7��'�"c��D�|�T���p��iZ������V��b|4���YMPq�JiB���m5���1�n3`����ӸSj�S����Z�T�%�+�}OUU�^@�6|��h9�F���)Sd�3�&Ӓdv�x}�J� l�����ߜ���\�ol�)ٞ��R��{(��n�� ЇM���+�f�?U+�j�HfK�e�=��h��=���t ,�`���{�Z��~D~��ȢE�Jac`���l�d5�,�6����T���lc�{ ��ߎ�7��~f�PoW"���ֱ�O=�TU��A�ɜ��`��?�h��|�8w-��)���}��8��	ܾS�x9��jUϑ��6sa.�9����s�Ľ{ci�����a��s�2~��7��Q>�yv�Z�.b�����'�"ف<d���z�qu���ʬs��E�7i\���6�q��ގ�w�j��MX0C���Z�r������O�'�?��u3�9W�y�1\3 ^vL$���G��� ���w�+�F��?w���d���4<��SIO�>�$�o�]X[X ��kSP���9UM�дa���Z�2�V��pJ>x�AB"Na�},���!}����i�&��~�-.,�-��������������3��g_X2�%l�!��\����J)=y���{���U�H6�@�I8fmb�*KmM�*\q�Ǚ�^��M;�#B��#����xK�=yI%��|>� O{�z�Eh◭T��{�("�|o-u����� ��_ViM���a�QŐ���'�/�o�m�X��p��%�X}|?���E2X�J���p���;f��},`¢x�ꯖ=nܻM��('����5�q���Vp>�f:�v�D��������Wp/��\��B���,��3�4�������8�*�O�n,��F D� ~H�0���F�
���j�Y�u�c��'�.�����c�@����]�\��Ec��p7����#�4ݓ�s�Q?�EE(p,��M��Ꭳ��{�՜&D���1#��}y�m��a�zO)ʡ �bX����tc�z<7֓����	u��w���T�����g�r%,"N�{�iڼ i��^�Z�
7
��7�Is��G��d�?tE���\�4��
��.�;�R��Pi&�����c
"L�N2 ⺨9M\�GhX�
 ^V����
)dz%�����m�2�/+�ZB�{�k����Z�6���4�+>t����Pi)���L^���9��SUU_4�5Kry�21*E���D����x4��H��Hb���9��3���MH�<�Ũz���ϲ��֞�H��	�hB�Ǣa����ϥ�~�K졭g��o�˜�VEV�� yʀ�֥�_�)��o���xn�G�>2���
Ղ2S�d�}��P>4��!3�%�0.	���}O�\�v��sP�G6�W��#!��b��$1�,�6��� �Y�]X�E��D
���F�����-��s���?f�I'�K�w�y������ӱ�5	m��|J��X �>������n2�`&��8Z2y���$�1	�3�tHM�[:�֋d���HݨIR��%��c"9"������ϰ�Q	SS�%ߛ���l�N
Q�LT�y�Q+�ܲ^6nZ��^5-�C���~��d�`��VdN�.�ϱ+�3�����7!�X,��>��-�ʔ9W&ȸ�j���;����p��l�Y��`���9����0]��J�*�|���?�aҥ#��Ϗڒ��*i�L:@��C����a�e2���������g6�.Y�����r��6�Z�v�g�;K�O+8�
y��@�i��o���f��_��u����/
�c)�$ �m� u6��SN9I�<{���Qb##�IL2�uHw�
y��dݚ5���mǾSƌ�(�bA�E<�0�XC �<�
��Diբt��k$'��8I�k$��H1&ɶ6y�OԒ݉�:�Td���/p��̙��YT�$�Ȣ�,�k����O�����DùJ��	'����{�Z.e�s�b��}�����e>=��h��M(���zA�%��{4H�T+.PB��2A����_-��'~�i���k�FMM�F�(؇c[4Y/E�� �B�F���˼���n���P�M�I�Nш��e`<�̢��;��=)��Iy��h�#l��\;�l��Xb���!���*�l��J�G
R�I$�*��:���Ț�Kd����ݍg�����y���6�m��d�*Z�)���J6:^�?C�z���i�I�������vB��'�r�c�� @ȳ:�3�$	�>t�	&@��}[so���$f�(�ǀ�$
�q��aaS�B��������؀0N^��P= /�5��C�R?fQ���2�SJ�?��[]�o�4��YҹZUOʹ�)�ȡ���ۅ[9n������b��L������+�V�i�,Q*%�˨��F]�Z ��S)�ɤU��L�H���t���-5��&"�#t(
Ю	����{�±Z܊��D� �\���I"�"�^p�lްF� O>�Q����G�F���ry=����c�}$"�P��#�$/����-H}�hy�EjE�ui�x�s��{�� {Y�y��2�47'�>3���g�f ��Y�Ͼ�i�n��O"��XY��7�կ�ϱ��@ྍRV��r�Vp�ņr��ou����J#	8��ܵ���c����;��dۇ*�>,>�4��:�ҮA3�#�6���w�}4������
h"h&hZ<L4��1���M|���|�v��U���%�؈�	G$_�jr�Y/�x��82���wu���qN`C�`��c�f=|�J���*d�.���P��:W�}w�"��keڔ�2g��R;a���Tt�`�/�׹�)�~V�DX#��IE�J66Vr����b�F��H��I:�s�x�|U��P�7��8�h�Dv�\Y�4�ӟ������cL�5���&�:�,�����k������?�W�u8���-�����d���RS�ڻ����h�
���~�D\B&�SkE��׈�j�����N4�|XT�pL::�d��3��w��͘Q���1Rp��ާ�|w�,>�i4�%����Oߏ@���Q*��%w�_�K,'s&eD�D��gs8<��Y%C;@�0�H���p����3��)��&��i�f;%�k�����n���52i�$y׻eB�N��I�)��I<�W�@�O\�֑��|1,�P\ґ1��-    IDAT����Lx�d���
jRc��7|O��Z�B��r,�2��G{Qd2
 &<�֦�����G}���e�����G�{${�,n��u�ܹ��'��)K�B�ׯ�iJ�P�����Q=%� ��!��|��r�1����SU1����ē�* ��]J��T{�#��5p'�V�,׏�M���#o{�12��4M��f{4�C��_A('��P(��1��'�����vg��o�|���a����z��|Njh�I�i��pF�|�'`�!�i$'E�hS�lЧ ��n����@ ����,�^�7~�g��F!-�BJŤHO��������2m�t9餹�0e�tt[xja����POH�BB��h�9�	�M�j$����z�>C�߰a��薛�E/�0@�V�۞ c9! �瞫�}ӊx�-&h�ϛ��|� (�ƽX3h
�)��Q�*f{=#��L�(:m��ɹ眧U=�����&�F՗rn ����0�A::����ğ�T����j�/��dD�>��������G+�>x���h������|@b���]'==���+�i�Ji�h�D̳=��Kf�ds$m�f�7�t�.V���o}?���4����[5I�c~=�<��-�J��R���-?Q�?����Ȼ�}ݜ ~�����$���4�����w{�?��X]7��#��vi�u-ᨙ.��%^h�pz�ܿ��Ҳ�I�N�*'�|�����d�]D$L@��7�gP?�����? �/D%��tt�d��[/�P�&|��ٞ��������R�\���@��̔+��s���a�DЖO9�Ufx�[���<s�G��5i�ja�>�VC������k�[	��4t:pN�x��ަ�N3���e���I��J(pN�)@�˚�����YH�ͭ��ZP���=r,����#{��C-r�N�;Zeٲ%���0y��m�=eԘ��Jgg(�L��ؔG�Z.�F4��il�v�=��J����l&/ӧN���u���mw3v��\�T^~�yy�����E�A�%@gƴ�e�}���;Z(���z��'���]�t��g��P<���L^� <m��kl����a��5�7Ż��U	�K����$�RISP�����XM��p��%W�v���I1�)5�#��&��*���Ҳa�����O��:�cͻ0ϡ�4r)� ��>�� Ӝ�I&2�9|#��KǶX,!=]���?��!I�9�a8�>>�E��U�X8"d�J$�O���0��#�=��$�
eb˾cc亥���w;�ʐ�&K�4(,�p�PO4� }�#?��?��pn���_�Ĭ{�@Y�2������n�:�h��y���?��J;�C5�1�M��e��瞑�uM�A��tugd�]f�G-�춇��.��GV�m���9��w�?����B#jf��lZ
��,ym���ҳR(f�.�~�$�HWGJ:;3�����G��
��w��]u�(؄���g��?��j.<0u�i������g�yF��玚��x���P���L$H�l������m������s��(��P�S��Pf���[�e�j����j�)�?�揀��Z�B��֬Dk�P�JN�%������	��p�v�wȝ?��<�ğ�TW����۠% ����I�����wb�)*� D��c�t_����+Y`
ʶ�~�������������}�$Q��c��|���dJA�B�/0�J1�W'k&S����䢋��C�=�~g�)�����ַt�~tc����_�4l�����^��^]$�m%�^'��:I�����#�~�z��݋P��]?W_ k����0i�#2�s��9�J&�?^I�g�y_{����.�fH,"����"�F'��e��l^/==��$��rE�ܒ��%3r��)S�(x[M��i
\�f�Gu�nD��X��K��అl�}�-��K�`J����$�$ �A�
��)���}
P��JZl/��UMG���4v��%����������e'h�������0��|�o!\�"Ų$_�s�ђz�6qٸ~��z�O��?�4�m��e c`n`=����k����g�r�Ъ�<+V�(Պ1+´c�?h�"4��-4gֿi�f���l��QF	��Ϛ5���D׻��V>�����Y�k�>X����(c�D0�P�$��{�{�k_�����8���.�HA���p��4��/�X9�I�tHrs���6˺uM
�(A�C�>���^�^:���K�a�Nz����k�#�}�'ߑ�z���%���l~^�N����5��6�{���v���e��W��#��_$��u�7K�ڍR��,[�^�9��ڸ�M�"�����d�����f8���|�C�/}�K��iM)k�q�8���CY��!��d���z-E��8οv��
��2�k���u�����餝�{�	�L;%Z�,��*���M��NS�?N�'c'L�t7��f���߬\��a�0GaM��b.�%%��d���ʈD��i���G?�%˖J��m�/�P�`�_�������X)�A�Y_����΍ՊF9m�4}ˀj��9�ǚ��?������6 h��Y066�T�S&�	]�N�6V�p^&P̪�s��u�]'+�-�4�cY��%���|�;
�P@|n>����o!-}��2u�x�PN^}�F���¡���s��2v�N�t�j9�'ɻO��x�Ң�jo�,ݻ��_O;���/�s3��,���c"��l��$���r���b�G6�4K{{��c%.�iY�n��sY��]v�uO�n?��M��/|��ݢ�������8�8|>�я
-�xX��o�߰�]�~�W<�ޠ������Z �_5�=�/�w����U6KK���c]���'�3�����e�r�#�|U�'��������t�<3q��)��eu��3;Dy��D]M]��Ʉj�G�K6<J2E���g�f�*��?��Mͮ�S�(7��_�y}[�?y&֏��8��;�	 �~XVn[�&\��� 5����8�aj~��9�� ��bV�YF��=7� �?zf��뚀5*�_��<��g�^��Nj,z�(=�Qj�~�U�Ę�@��n^/O>z���,;�N���AW�?&ٌ��Eˤ�v�4��$u���ǯ�V��FIgw�^kŊ�zn~�����h�l�0�k���CW^!�pQV�\*?�k9��äP��VKWW�s��jd��ViZ�IB�zY�z���!�)g&�5�\SZ�,z{8ַ�
��ޟ$R��8�m�9}�`���s>��� V����5�	p�u���o��匇�EI��֑���
:�!
B-f$�k�Da��3����&�}��ɪ�O�?$!AcZ�?�H�\J���7,�bL���;!���_�1 v��%Z�aS[�UE%t����mƀ&b/Ӝ�Й��|�R�P�7��zt������$8z˜�s����\�	�q� �����H;�()s��}[�:�F�"�L�.9�i�t��gȧ>�)u�ҫ��k�U`��K�B��&�h�x��e��k/���J�<r_i�4V����1���l떥˚%-׷KgwV��m�caٴ�EE�.ݲ_���Vf�h(4�=gϖ�\}�Ĵ�C�����;�y���]�~�jimkQ隈�K��NY�z��r1y}M��e߃T�ǼE�n�Q�>X��ӊS���Ik(���g	/��@7�v�cK�qmAT?����\2W��?�}�� JNi����^�+ڡC�������?�q�u��LN<��D�K������|�.��?~��h4RD"�!j�Nϗ��d%$4 ������}����#	��(1��|G�l��5Do�������M��F� �ti@���}�!��1^>?�uW~,�e�o�I����_�m��˵�"0G��6?�o%�IO��í�i�Ҵ}_0r?8|���<��#�<R-�;�C�.]�S��g�(�����<����̖q�G�kK��K��D��saye�r���ٕ�L6,���:=j�tv���C��0&?:�����n���5�5������~L�j*f����ˡ�'�b��Z�B
���i��M����뫤�#/k��ȱǟ��?���8�j4R1G�q�<,6+&�]w�UJ��}����M��^��m?k:R�R�4.��k`rSBAk�����x�C��崺'��2�
�E��ˠ����Z��K��#WKD���f%�k�p�E��M�o��u�d��i��O��JW� ��GjS�;res���Y<9��\l���%-=��C5�'��W_����/k}�����WU��d���b�ͱ�),�}_\������[Pۦ���%
ڒ�ݞ/�K@���S��,��^������Fa��^��P�,��PV���8� �gs�Z����(k��a��iz]:�h�p8"�]=�|�jIeD6o�:\�8���+�_[.w-�/�5�m6���ܹ��L�]]���]�F�{�{������ukVJwOR�6��\�Gyr�$ź��U�o��Y���רs�ŀ���4v��v�J�{�WZ���A{D`��㎅R��s\s�j�O;.��JN Zd,���u�>���xc�����Ւ��q�:)3D�E���u�jA�l6%�t�$�Ih�g�Hj�<xϝҺa�L�� '��Q�O�.�T�GE����{�i���	z5��aL.2Z
�1Z�!-5"�z�<����_��������C���F�;��sh���r���A�<���a�>5����l�}��6����oK>M��K��l�K֭}U2=mZͶe�&���n�hm]��^�$[���ʵr��W�����p�N~��?�/�KF�%����m��8���m��+���ƙTJ�._���$P��d媥�|��QL*,�t��5������3%��V�1swV$?mq�qN�iF�C��x�%n�E�B�s˜J��ETqkT a�泙��:���db�5;1W�=�5�kj��'%�Z7��U��?�u~��-k��1�[�y��w ���F�eR��vK,��!�l����r��ۥ�y�4L/���4��O��H������<���2�4²q�a)(��B�^r�1*z
1	'F�g�)��w�-���Ev�?�����/�}i��Q@��?��X8u�@���9�9���/��ژ�3�����M��A	%�GK8�q���7ȸ���N)Ƥ�'#>�;��?�s��~��ɫJUϠ�b>���cG�YgΓ�;X�]�m��i���7JG[Ri�P!$�h\�L�*���Qv�6K+C"�)��׿�����x8�}48U� � ���4�����kU��*�O��q����Z0*��%�i�OKWG�߸�E����$	�Õd#;���@�/���S��f.��{�w��х|F����%%�L����_�*�Vj�ƹ�d���E���lZ�ZVZ�IT{���/��/���I12Jr�Z�)F%�-�L^�Q��ǷH"�V�v���b���,D��2F��GI�)�����w�h�믿^�=`N��7�B&5��x,,�L�<��S���OHw��E�g����Ւ��s̱�����3V��^�Q_KJ���������++i�tɱH���0I�s�<y�[���DL��Z6o�H��+V�����HmM��7^r���?�L���ø@�RY$h�˖-�Tp�r%j��vq왃W��ΰ��_� s�r��O>Y#���:"�Y�+�fZ|�UWT�z�5�O�1��<�v8���N�����*g�{��I!��P!-�ѼD�ݒ�l��~�lni��;M���q�$�FK���Dj���ϕF8�5��/Z<>�0��:)D�$NH�>��:���R����)��H��ڧ�2�w��ه~�nԜ�D�QR�`�|nV?�d��Ib�߽�ҋe��	l5��sҶy�,Z���\�R�'64(1z�X]�������=��qB>��_��?w����+*�?tN	�pxf���w�q���{�)��u����%� �ߵ�u��IgSZm�����-�>Rn-��+��� "p�P��/�+�A����í����ꩧ
U�Jt�g�����|�s��д,�?��I�=�y}���~*�%�&M��ft�m⡜�r)I�Ҳ�y�!p���S����K��ه��O5h��<��#T �HB��I���ȑmIm�M�em�j O���Ù�ߡ�7[o{p��c>9����M�+�y����^�����l��o�8�!� ��sl6�ў�T�em�_9.��+��������Sa��1�uw�q����46ޔlO^^	���IM����Ak�\CC�w�}�|��%��C(�鲓��K�_��,~���q�\�߉r �k�]w������H j��3����@�[4�j�A�ᆪq.�K��h��VD�B�}�1b���E�S�`�M�X9�� �j�ѨjN�\A{&S<-��Z^
�n���G�R[C7��� U"q���?Q���$��Ȃ���91�XH�X����G&�W�N)�"�R	�X�n��/�},J�֩	�сo��/L @�@����~s}�].��6N�i�2(��f�TAA�US����fy������N�����r��i���8����HX,��.$+���̓�8q��;Fv�4YƎ'�LQZ[��ҲY6on��x��f|FA�h���O>���illT��駟Bİ
 ( �~�����G/m`n�DS����@�NA��k]i�����s�nL���D#��N1��
��pQ��٣ɴh���ҔF����fc�*�e�xI�Y�G4Ɯ>�Ez�F�bk4^��c��3��(��ZKH��[�C��ܕs{i���\@ohhJ5`�*{��k�.�{([w�y���`_�P�~�����t�"�&V�J�n���"��YY�v��X�\�֮�J���Je8�S.���z'�[�gNc�-���%�4�^�ؚ��"�J@K@� +@`��"���ʩZh��l~��Ԇ�BVl�c�.���`IahF�{ktMY7��(����B���-�6���)�ઍ��E1��r���"EpÚ�[Q���h������x�P�P@e!����I|ύ��U*a�`�--����`q�V��O������'�Y��	|�����Lk-�vMS��������5�<[�4i?1��k�߯Y�ܧi�(Y�� ��Z�~�i����I�$w���to�M��?�>�����̿u]3!���YG+\�a���^T_#�g����Ȏ�N^CE��j�P��ҕ9��<@��tJ�o���n&Ο�Ë��;�s4������Jv��	zr�i�Gi����F� ��Z>����| �WH��m���!� %�+p/}��n��p^.z� 	������%V/ޢN|�|�1XL��s~9 ��FeP�pŅ ���=h$��mnݢ"��Kz,�B.�^B΄{�롅㿢�N�����˪�Z9
n5���z�)���u����_�@m�@f��,q�G�PG�:��h�֢p�X������2��:��]�����ޖ�����ی�i��)�
�1���p1@ӌ� �@���O'Q?<|8?٢p�֤�<�[h^��]��Uz ���瀻W�@_-�-^[&ܠǀ+��ZVV��IT�e-�$z_N������c����7��'�O�:a}�R��i���[-״{��
h�\ֵ�t����,b�Y��+_<�ׅ�|���z_`��û���,�J�P[�(W��qƫ 3kz��a1�~��&J�T�=|���A�?�A9�c��K/U@�o�x8A��"G�h�Czq��r0ƔI���}�`D��@i5�Kt�o�M;���(�JZ�3�\sj��X�l(8@�l67�  O��
�ق��P�[]4�7��0���5|[ݴ�ܒ�\��`ӻ�x	���m�KTSp�����?98�X7Dy����~&����5��E�JQ;[�oL)��>��iHBt�����n��Ÿ�H�p��j���:�4�H    IDAT^6�����2�+�5�K�'9�zDd��b��c�ҺY��j�X�{3��"�'d᳧���Ju�Z}.:���#��t�9x�G��6�6Wt��+; ��`�=[�}|�|;��_�K���7.��V`����n'��3Yՙ��d����fZ�{u�Z��>ڲU[��>�?X�zەuc�����7x'h���m�WI�!ʧwc��p��1�w[��J���T^Vc��%�k��_恵u�ŗh�M>���&	���
�Ma�3a@EJ4U�	pn�QiBd@�Fnf������)��oq/�X�:��t����S���1�����o�� 0��>y��'T`�z��h����"�����E�Q{<C+�`֎�OF��C�I/]��:sQy�·o�c�>[������ι9�l��o��  ���X���p �x����X,�.O?�^~��׭ҡ�c@0��g�}s���������ӁƯ1��a�Q��������"��G���;�('�P��pf������b@�o��
��'��¾l��Y�uiA�Cz����}�l ��?�x	p��d��p֟�S�'%��G������W��͌lo��Qg��4wb�*X 4�D�'���R���_�}�����@@���9��}� v@��G���ZtE��� �~���V� ���<��C=u�IL�s&�h�����O����eԉ/ }��Ea�ꄘ�"8,��L��/��m�;�;�T���
4P�Y̹:,:�D��:�0V;�؂�q�����cJ�O4`ͽ����;�*�"
(� �D����o�� �w`���h����?�.��q5˭��ӈ(p�B5RR���&�O82�o �y-'d8�i`��O�:���&*f��U}���n_����e��$�@���k�6�̀�5��B7�۲�}F@��7��+&<��nA�8G��=VYw�y�Sm���f.�&y��O����������MJ�b�3������a��LR�ke!�>�lQ[g�;�/�7���J����~| >�n�(e�z��Q5��¬%��Q�1��s�å�]t�}�o����}I\  ��唺/�pm���������ș���?�����_3A�s�2<�4�<V5λ�/ � D���0�(+NL: ��z���� ����4\	i���V2
�ǜ�|��?���J�H��!��A�x��O�Sy��ϕ�f����5��R	���uNc�k����RþeW
�E����?т������RN�����Bä�.���-�@i��h�ij7�l�:��6�����@S��z���s�/�dN5{�&�M�0��ie�)�f!kV�m8���n������r�>���pL碆�=���%[�J8A�4����0"�BX
9�/$R��L�Dc	�*/mW��_*'���B?{�y��8.?���8����KNK[8�c��I?���eo6�EI� �|��@ͨ�lxr m�g�]�����a�a�s�lH�9�#HL�<;~�_Z\�{!�s�� �K�,�I��Ϲ�[��3Ӳ`�Ͱ�Z�e���s����d7�d�������{F�1ɦ��Щ5��Q����̿c��y��:Zp�ߪ��¤ɓ.Zpׂ;��q�)Ù��w�6�ؖL~�R�'fN"~])ˠK8 �q��a��ٿ�]�͇fO,���k�+������Y�0�!��6��5Sq[��@c6*��}b�)o}Ѹ�t�d#͔%k6�I(z	S3(KW.%�xL��^��6Q�VsQ4�ׂ89��3ʩ�.kkH�rBݜ{�xUt �͒�*<D���^[� �  �Y�+%Rm|>���-j���c�Um0��/~�EȬ*%�t�Ȕ��B�t��̱���Z'�jWe����Y攥�.��Z�|��֪]�,�r��k?��1A\$�]���ح��+	�\М������`�_�F�;����4�JUOJ�(_t%�'D�g�M�2MC��؝"o�����^�|�K^iO�F��c�Μfl2�M�}5���˂�Xk3K�a��U[�&�q���������E1w��VN<���6�̉d;3RK(�Y��$U�H�X��E�%�l��Tid������u�����й���F�VQ�8�m��Tm�������Ǝ[�!��	�4zh �V�U��������)>����D?B��¬v/}}�=��A�;���>��7�!�W�����#6'��Bm|��9Pko[���y�@��+,�#1a�+f�k�� R��y�{�5#�a� $<��%�Y��VUJ5K8Lq�ٜ�(e�WT.F��?gn?��iܑ+�dS����շ�dRZ���C��8P�O���@��8��^xi�����Z�ro���ݚj��y��dr�jf6��a�Y�C9f8�����gt�J!㣥4!~�	0*�����͇%F�|`!+��uP��Ϡ�@��_*�a����p){[D�k���ԓ�V�֦t\ȅ�moڠ�|0a�٬C^�	E�0%b�V�l��O��F#ڇ2$��n����%�O�ܼ)A?����2����]ˌ�,��?^3�V�����h-۷v/%N?k��9�� ��w�]��{�}���N����K{{��{��e��Œͺ^��TֱA�J��

�]4��;�R�:������ɫH���l*źb�Tr�a�hݝ���S+���,6߲	y�񚄴%;d�UkBR[\��mE��/Eܨ���c�ir�J�/	_ֻ��6����K�υ\�����.W�'�L����3Q*#񀟌�Dr���t�R���|1T��C��Sh�oξ��B=K!���&\��;�Nf��R2�ZD� �q ��0����Yw�%��Y�J��+b/+����/9��O��yC��_�B�q�R\�똓�|ù?C��ZG��w(g���N��\�=�9��bn8�	H�S�_���޴��#��|*<���}�q:��	���K�6.�tZ�@&��g��U~�Qio�T�ɯ5������No�^{[�>9�F�Y,JM<!��V�={7�䒋�e`&�a����SO��5�����{�m#���J6_�g�yFc�-ӏ�/��6������A���~�3uH��+����d��@Y$�Ql�u;�SW�P<�j��#����	Eb��B�I��IM� ��aɤ�$^�L!+�X��c����A��6*�AK���� ��j�J �2g\Oڅ�U�AM�f\Tyd=�X�o%��B��k�s��À������Q�?k���,4r�܉'*��7fv/�`ʧ��	&��#)���.�0�����=k�Z3������_��SOy�~�!:T�m�j��e�/��!3f�R*ߘ*�_������haT�LGt�W5��9�Ǝ-��8]<h_�(U(d���<%�$�6l��-�ƍ3Zv���t�2e�n2f�x}0����I����9I�[����EL5)����~�#��6-�8Zs�j%V9x[V�t���|ø�J#�;^K �0��X��ĊiɈ�:����W��nA*v�[e��骍Ȕ�M���[`�tە�_^x�����'K�~�9Wˆ� �-��X�o�X�<C�A�`=0椯z6}]���A�@�ˢָo�Ws.�{�t���1״y��1׼�s-���<�߫��P�����|ǯ����|��=��x�;$��X,$˖.�GDk9%;�5󺶾Nv�<UN>�4�y�LIC�f���C��o������=�h�3w��$�mWW��!T��#�K.�PR�.)�R�ʫ�ŋ$�s�(�X�����1ǟ$3f�f	���A`a�7Z�O<���{D&P��/��7߬ܧ��i�Cs�����W��j�_߸^&�oP��D���D$+�LR��V��rӍ�	e�x��g�#;7�(�Z�,%����JqMV3�W�O�GKw|�d£�yY�k哟��$�W�����b� �8���"�|筽g4���Eq>�j�6&����9�~���ܿE�Yč�*�;��<{��A�ܱPp�c�0�F��Aik*���D%���+�ʋ/>/�������b�����%��%'�����Y�����mwܮרV�b���<`R��!�/�lJ^[�P�lX�$�74�:^�Ԥ!ʆ��;���TH����j�Z��#�<��$��D�G ` ��Oa��ú�DYT���+,΋���b,Յ�^{P��x^_șF��& #�M�0n�\����œ�	�%&]͵J��"�L�����K.OrRX�4ΓS���h�q��_��Co��~U A��B��;�����l^���~�����߮�0+��
~���`�E�Yh�i�vߦ)݈������ޤ������n�F	0�ǀ�w�o�Է��<��E�*{�֬�t���.��Ȕ����L�SR��e�ڕ�a�:Y�����N('�C[7wʆ��RW;V�zϹ2k������������s���P���&7\<"���̝��d��#�45�����U2��F$��_��^����%��U�WH6�rE�����eg���D��w��o;^{��`q4A� �l(6)�>�Na$:B뀈"��"��h�9�q0��Zp�ݶp9����1OY������Z�F5���)��/I�8zIB����N�����&���ߓ\�[�Ѹ�i<K�M�-�|t�௢�^yu��[��u�����L�Fƕ
�1? ߂{�|p�U-�
��=���QHe����{)�}�yM�X����	���P��Ox��vO&�8�w W��r�a@���57Ա�I��snj#A�|�+_ѐU�a��?�����ʻ�<��?�S���'7���>&���$Y�f���V�p.$�tNV,o�H�N6nL�1ǝ('��?���^��%��O�o���Gn'�*�O�B6'{�>[���5��꒮���}�rһ��b�G�4��Q@���I��KV�l�t."�W�ʁ�5�y��8���Э�;���A3@ۇ�4��6���
Vv�8},�e.���ð�B B���{���-�&�T�B�����w�!����$!�?��$V�h�E��n���}�����eΜy�ӌ�%O��W���ުm~7���.+�ՐK! ��=4C���R�4������]E�WP���]�#6e9	�4���O�X�A�'�0���<M�)ꏡ\[5�2aPm��ތ�7�f�0�i���s�Y��y���/jH)�$���sP�xAa��p�z�ed�����
��M��Ϗ�J��wW�0a�,]�DR=���LQ^Z�D��'JSS�4L�.W_�q�������X����-�����G,��vz�w�ے���+�
��n��U�R��>������C%����HGgR%,}f[6%��i��N��h��<T�z J����}�Ta�nB8By�L`u6��f�F��z�D�+Ui�V�Tw�F�u�Y��EW����� ��8d��xp��J��qh?G����-�~�
�jK�b!,�PN��E� �o�����wϝ'Sg�&Y/%~p���f�'�lU�i����[=k����W�������@ɞ�Qp��E +��h�*�O^�L�[��� ߄C�1V^v�rJ���E�ʩ���R�-�g��k�Q9����?�i�+ <�[Ț����<Z_�җ4ʏ}�g�}�҈�y���SO> ��L�0V�-_,�T���;�e��ՒN�ds[��������F�+������?����YC#��46~;ٞ�XE��Y3f�G���$�QiٸV�ӯ����p8%�ׯ��֍J1Dc5���)�[$����u�2}�n��O~R��L�u�]��ll&�Y͛7O31�������$n�\�b2��-�8�*��9v���{�:�D�X�����X% ���u���)�>+�ʲ(Gq�Z?�A1.���
�;Ϳ��N������Zy��g�ԝgI��;C��5���6�}���F�G��>������9 �hno����`�?XW<����)|+�5j����JM4Z���T�P��}��0�V( v���j�;������w�Y��'��	�TA�Pv��i4�F�S���6�oʔ)�-W�Z"���>��ݥa�hy}�2I�;u.�+J1&���H�^��9�������_�DM��(��?�ח/���✹s��L��/�W���ҢL���|���H<�h8/�T>ho)�es[����ꦉ��=���5�d��Y��SNx�)2w�\��l����'[l$�8�I���eQ���� �-����Dk��PIh$�;��R!�l�тF�M�O}J��7�������DC���v���$�����rىb���-7h=�p�^N��?���:�������k���Y���n!����X5�j�3�ʱh�PD���|�V5�&��	�ٳg��F4~˲-�N�Ž�ڻ��HM�����)(6vߧ�y�{&��V���*�p� >N_,gzPn��n�����3��g?��ww��SO�Fv�e�����U����Q'.AX�.	�H��69���e�Y�HM]��Q�z�J���y2�gräK�ϟ[���__ح����E]S'����-��!5�<���2vLTZ77K&ө��<�I��d�Ƥ�i�,m���+�Y4���n����o����6.)�d�ZV�ղ)����%nX�E�P�j�x��<����(��s^Uƅ	K�x�.��LP��f��a)�sr�)'No���OL�@$=��&�)��o�;o�A����i�g���H�8�Ԟr��^j����4���L��1�޴ȵ�u���/�Ɂ8�yA#P�� �4?+�փ k�5J^
�4� �|fl����~&�����m�������Z�q�o̲���e��ђ�X4��_���g��ǔ��N��%��l�[6�4���O�|(!�6u���kecK����d��p$"x�O�8��t4A�����_����k�q�G�|@ҩN	�Ҳb�bY۴LB����0ц��	��²is�L�eO9������Z�������i�?� ���E��ԤZ6<����M��$y�:O�R_W���7F��DB�r���fiK[�R�Ԍ��lA�����P$�)鍧�K��;S�uǥ�3R���-���;�'�ߩ3f�_2�i��6C�M��<���8uU�7���c�'���"�L���:媫�ڂK�@8�s�_t�E�\�SM3C�T�4p��N@���~�ܔTF�	�ZQ�G��xs����(<p?|�����%|Yة��T�d��l�{����\z?� 7���ɼZ$�|�C���l��j> ��;���
�Y��"�Բ^
���ջ�n�V
��,[�$;M�.�x�I"r�P�k�dR����'Mn�l�]~2�4�j_�,��y���������)�\V�z���<)���	B"�e�<i���]�!���S�5�
����o~�	o���_ %z��g��X���e�Z�5�bc���J��U�I	'�?�X����
�!g*����"!���:[�q%a��J�q�����~����K/���~�kFr����3.��?�W-�j�<��s���*9LK*����os(k�ݾz����o��,[[*��GT��M�lx�>?4dӢx>P`���_�܁�P�cn�u�*`�Z������`%� 0��iԈj>`e̕�c@��8��s�OV =�q^�!�,ɑ��mfB��"֞�� 2V+��t�2hå}l̾���p/���P����?�Q8�n?߳,`��L��1}����Xs+�.�t�GǬ�%^#uu�d�]��#ߪt���O���n��]�j�W���{�����2|��O�E�`�Q�	چ����>��j�(6���n�g8>���+��( �w���i�(����v�M���ok� �C�fX3�j�OooY�h{i��U1/�HDk�G�Š-ڹ�x)��AP����+�B�h��$H�
V��z��,ި�%���K�mG�Ux@��Mڹ�y��k��Dr�r�-�ӌ騂��2}癚<d���9T����0�PL��'>��>	hWW	.��-
�����@��>p�* �mp��    IDATk��&���7��u��h��#���/V��^Z�p����~��G�g����̾"J��s<[ȭ�B�%�k���?�#t�$S.^�Z)+8̧�|�߄)
������gF�|?sl�c|�#�Ep��1��fT	&��a��B�{3G=Y��~�3�j�ܴ����~�z�Eۣ��+��$��3�h����c,^k�d�Z��駟��k��4���� ���4 "X�x��u��jR��BAM�bT˰����G��Z$�m��R@A-�E������\Ahd?�O���_*Gu�V��������z���yN��M��p�$�����&��j/_�g-SX�4,M�"������ |��!��ZrbEdQo��Z�L������7ARm��ל��@?�1��/|A��=L('����� <��K��I�:Q#,��s��!b���D����b>+��wh�}�@����\rnY�����!���uڃD�g�P���<�W���=�����X�p�V���������ϗL^�\��ˊ�tP��zݖk��|Nj�Q-���~�.�K#-�)��`�B8T�����2��U�����S��4���4�7;�w�v��ш�� ��'N{SK�
�lp� �� �X��}H�k�������v��m|f��� �;��wܡֵ�a�<����r�[,,�
͟(����O5�`��Y����f��v��V<�=> � ZWR�Ǭ�� ��������:JKD�]�|�w��P�
�C��a���Ϳ�#���1�����2��Ĳ�X��e�Y�"�3�m��u�^ܯ�c��]q��p���,�j�8�~40�3�@,�El�j������6ܾ�����I����4&?Wt�xE��=�?�գ��}�A���ϣb�?��(�(�or����F�F�� ��@��}~�NZ4UA��������?c6�Ф��*Y�80�o�k�kXn��?B��g�ؗP��?`Z�6��傈�s�'؀�H����&�/��BIq�Z|�%`]�u�����1c�j���B�h>~���a�U:ۻ��������t�Ι;����k'��Y�.6̀��$eaqF�w��O:7���/	���-|�-��P�;X��@�-���>�C�@؄
p�QI�H�����.4w^�܄�����4�j௙����>�8G�>�������i4Ž��{�/�9|����g�h������_\��v��m|�4���t�w*M⃿s�;%��
6͟=�%C�ǣ�C���?�����/ �|&��M���m("�Ц��1v�V� ʤzJIZji�M���ʭ����b)�7�2*��N^#4ο��d{�r���s�ol��i&��AZ9�ɷ0N��i<��o��,�dq�!��ބ["�z���y���8���P�װ[l��4���?�q�h���p�M���������5ZY�h����\+� J�2��?������Qee�.��(h�O�~}Я�����?��1m�/���"�������1`6��2>ބ�Y�������-�������7�Z^6V�5�r�+ױ����ƹ�?jK&/��&�m���<��o��k����w{�v<��Y��%qY�-t~�>�[A��Q��ĩ�B�9�q�.^���M�/Pp_U���}x�,h��q����ڧ+:]��1�o���i�����RS|MD���$�ֈk�u���LR"���3Գ��7�Ǣ}��њɏA��e��r��ڱQ2P��	U���t�6����iS�6�xߺ�Y�$���ri�����m���9�y�ʼ���{�
V�k��_a�̝ss2�~i%�f�BA�0p�T�຦hT���^��_mCb�
̴R]_/y"��!J��x��L��X\2��d�"�0�D�.@�8�[A������ΔS�}���E�@���h��>��{6.n��z��WK(H�y#���'Ml����`��U+��'#�N��f���LHl���3��k��i5�xȤ����󀳼����m�vaw�]��A��A��A4R���&Acbc��I�Q�`��&%	b����ԥ���l�;;����{��s睻s�.;�J��������k�-�9�9Ϳ����!%�kF}�9>�|QHϿj޼�_�I�%����Fm��%�5á�N�ܔ�ɿ}S�?��6fa)Z@בE�@�,I(Q��H��Gs:�cZO�h�,喖���%ʫP*Z�R5�������Th6]��+������V�v�ε���\�/9|�}F@�n���M�(�v��~}Y�M4�a��Z��V��h� �Ƭ�F��|�
���袋<�h;!��C��j+�o&|xV�}h���F�����^� ��x�o4WR:]	{�4ք�s���;�����O@��Xf7��ȹ���6u�5����%�R�m&uX�Z�l.8�� ��p���eZ[lm�z��h�j��?_1�?�2�P�bs:ϱ����8|Pr��ܣ}����O�������<շ��� �������LE7L�?�>ǏF���u���B��{z�����%�ܾLʎ7��	%��Q\X����FC���9��������8�I��;z�	�����J>�s�x��~��i#��8�CŞ���yS�X���T�/4�UOq�\R��l%��$y�����Z�>K�zp	���A��������ߠue|�AAP��R�j�~S'�%��t�3\�
ȎMm�;֚���v `b��5Η�#�#��N4��*�������3.J��b�wliku�u��Ͽ���xĴ�"���hA�s9�3Np���|���M����#m&6�M@<�����,�ac�h�x�����-����I�!L5�#��*��[X5���+Y�J�}�m�����3�i�Bۉ3�8��r�EV��]�_p���C=�?�Xdn���_�MH�(�E��P�f/�'M>�jDT�X׏�n�{������Xo�C����
��cy�0�^�Sۭ�lh���'2��9��4��E���/�����V�o0��t��5{����ҠK�ġV��q���P~G��b�+�k<�(MχD9Gswm-�,^"�Z��ʹ�{6��įJ!�����]��L.���J�5��H�/UҞLv�)'�e�����3�-�"�'����"�������6���o�Ǎ�}���B�KȺ���M]��KqX*����v��I�Xv�B�u�l:���0�XWZ�)�c/�J���8��ⱎq=�SO�	W�Y6h����x���� "���O�6X�B�|5m���D9(�wSP3��뵃^�*;������L	��=ے��׮��]���߽���x�0k�h�T�|�	�ٕW\��>p�.<��q|yv#Գ��R��/�'��M/���2��V|~�p�1�"�?�"cZAʋK�/�����h�$�G�c�����5ݍ�JH`�C2}ϦS��M}�?�y����4��1���=��Ϝ5���o�����O���Ku��\RB�0;@����o�Cʈ���`1�/n4|
�Qȉ�Ʉ�@M@f<�F�?ׄ�)��v��ϲ9�����Vs�fq�fF���Yw�z�����z��{�����Y{�X�O�y��!;��W�UW_bϳِ!\-ZKe����J��s���iU���W�3�c���t.�B�� @A󧄂�q�#s�5������(�&;X��W_I֬(�p�\@�84�,��]2ӳ#l�7�c#�����*����>��@��G-�O�'l�$�������R0�s-�P	<�/`
�#h�0�ͪzVK3g�x���fq��c[[��f"r�
���a�v�y��C\���t�Ig�t3�����͛�l��LUi4 ��>�!|�{��@�j(e]��ߴ������F��JR<�1{�l���7y�>ז���j���3\qՕV*��b�h��p��d�z����r�Q���5=`�r��U�[� �f���v�yo+��V�T����A��0���Wӓm�u��KLOp�ui���5�`�j ��8�\o������̈�\2�4V��I<�l�/�3~��j��b ����<C��#A*��`�
��8��C<�u��h�D�� �)W��#���O<a+W-�r�j-�4�
ax)��G�q�-�jub����}���/*;Sj����zՁ6iR{�$
�ļ�y��/U���@���뮻|�dV�V5o�6<1�h&D� �|��ޡ�?	;���aƳ�Y���Ѵ��n�lB���>��������L��'���כZ ��
Dۭ\��L��J]I3�U�͛>����L�ٝ�ێ����?�a��L���nV�NVP�����~�%�U�g���0vZ߱,v�}�9}6ָ`�r�r���Z����EK�BG&�;{��9^�eŚ��R�8��c^k��q��M�p�Jh���6))8���k�y������B�`��ϴf�ђ,�$`+�'+fvg���=�kE�Դ�JH��q���/����5�b�`}��}r����͜i�����=�2hȿ��/] h�0�u@���c�Q����3�\��뼪'�%,b����Q����k"ph�'�P59�c-��P��Ѿ!�����nSuJ�ͪ�3+�Ղ��^Ye�b�}�Ϲ� M_�ﶓ+#�[�ol	lP�2#�9�����VjٶֿVB�
�$����,�3A."-?��a/J�b��aQd��5>�	篨(�Y�V6�����7	%�1�|	�gǲ+�{Q���9ԭ 1��׼�Zr���������f*c����,C:CK؜�E��O��Z�iߘ����Z�К�9�v~��;}#��}@�6�LV����㏵r�`��m����k��8y�n!���v�񯱝v��
�Р�ʄt��s]��G��u�8���?{�w1��5���as���FĢa'�X8��gu���6�O��]v�e��?Z�g�j�b�r�\��]�Q^e����͟�J���?{ι��n������V��ץIR�: ����.Vi��c.m�1�����V�t!.�\�k]+XB R�&i��˾�}�q(n������jo� ;�}O�q�o\L�Y4�>�o|�y�˦-C~M~�=�Я�_�<�T��ε�Ge��q��N/R���ݾs˷���V�X�q����z��74�R1^��:�����k��bi�2���X��~�z���V����S��p¤�מj��� ������pg0��'�OO,�R�Y 4p�q�<���G�g��g<�����(�+L	�s��$��IH��ў��
GWlֶ�ؿ|���:"O�5W�\����W��o�w�� �v;g��t�s�5���9�T{F�y�����
�l\�5���㙻?�s�*�k��M�Ԍ^ �Ϛ�?���8� @q,���ԱT����:�q��g����}�����}�q�{��l�vKW
�j�2{�
�5����!�r��'Y��SՌ���cg���aͲe��%	���	�1s�w�z�����O>ڧ�����ο��gҡ�+���;���-�.��yOY_��\�Ժ׮��g@�kw�Zg��e,d�]7��;�Y���ַ�A���B�w��S,, �9?��3������cNqS.�)KRB��#�,q�Ҷ8g��CSH�,�m�N����-�	!��R�Z�U�V{-W\g����߸���m�s:q������sd�R2�[Ç�s�HX͍��
�l���_A_������l ���j���O���O�aq7����D8Wt���P����3��~�;q�����?ֱ�p��ҬH��"�d*W���Ъ�O�V�(����~�"5g�;�Ӭ4�o�}kl�����m��.�e�����T���ݽ�v]���~v������6�c�}�;߱_����'�
�fw��9�����!��������v���K=�e*vם��1Gf}�����g\��j�[�.o,���ڲU�v��'�\��ˤ# ���ڦ�zϸ�hw�Ue�}��x�����{*�&֬�����X>��a�Z�)�-�O��uLF[Iy��ʖ�>˖�Y[e�Yq�}���Y���X���l����
�i���Ӹ�뱗�~�ӱ��Ib�{�i~R�:d>�V�}zZ��W>~2>���W��ǳ�F��Haoq��gu���-$���4z
�3�{�����k�j����7�[�����i`�_|ћ��4�a���3�K�=kJ%,xƏ�㾮��2��㿴�P�͜��=;�i[���{�
u��E�ʴ٪�n;�����ϲt��~��Cv�w��@o���hkuBk��tv�SOO�Ɔ�5��*��]��k�=����k��w�f�q���Ru�E�\_\���A[�d��*��pq����������Gc����8X,��;��}�+�WZ8���ŋ�O�bO��9�6u��<E+(tT��4�X+��Q�f �3,��ђ���Gl��휳��JѲ�!K�z����T�Ǿv���S� ��Yi��W�~ɴO<P�ų�ʈiJM������g��d�>���[���O�����'��-�y�3oФ
z�#��z�OIg8t-��3Xԛ#�^�Bk��b��
�_vɥ����}v����4�~��&��k�-�6Qqt\�b�=���۾��bS�L�矟�ډS�ٜ��y�b-ֽv�v�y��򫭭}�[7}�f[�d�V�o�@fϙ���|��������o�\{��Re[�����e��z��}�յ��z{���U����]��?X�EK��+�;������c�|����BF+�ē�'��{�mT6��O⋇��vl4��Q��{���U��P>�=e�4����Wmr[���!K��<�kš>+�)��\K��������v�G$6BbD�n ��,0��|b�Xf�+�v���RSt��h�/��'��3k��o}�7>G�˗��%�?~�����X�ƲҮ��Z;��|�1o����󛥜�����I��}��uk�zT�BTIY�?��}��i�@��g���{�q{��w��G�	��>���Z���Y�X��O����|�������g���]0|��_��_������HMh���9��?��������Nv�uW��t������)'g�L��?����>�����l��%V�v{qI���+݁��ô}���_Kؒ�/���ooG}��s�9�Ezǝ�s�@5��&����n���8&�%�9kC��p�'�(sV��j��բѰڥJx[&kE���]3�y�b��h����I9d#Rd8HkDZ�f7}9O���F&I:��Yk�e�6z4��6�XJ��v�o�.�x�Y�H��͟��3�я~�Aozӛ�W�j�*��>�яz����>����m��=��o큟�eG~�M���-\�B�0��
Q:�b�>���E��)�G>�	�2y�����׾�5���s#譭����sf$����F�O 6k�v����`�-4#)��}ێz��V�5kWY��5.$hX�b�J�^���dE�q䱮ɠ�,\��#~Xtj�ƽ�T� |��g?���{｡v~�����?��c��@�r�nC���%� �8�˰��L��28d9��V��{���� ��A���}�a���w �7��J���d}lrix<�k`ԉ���l#P�(X�P5dU�Ҋ�c�?~z���������� �F�O�s�y��Y�{���_��g��P�(r�]v�;�|?�����O�����U���w��{�lmm-�l����'!�<b�Z���t��s�}�ʫ��z����^�%'�JK��Ϛ1���n��k���'��L�omi���n����暫l�=w7��#�����Qجh]���W�T,�C<��s�z]��YW���~�����;�?��O4��tLS�s��n���������8�R�c�m�m�Qj����Kg���њ��gCW,GR�ӡcX1]���,%�	�䟁2���ޗ0H�x���@'p�c��lL��
(    IDAT�?�K��(IP58}��f���۴i��+�� �i�8^g��e
�D��p�^~�e��>��5�>�����C=�� �����<��`�|������ͯ���cOe=�z��d�
�Z���/��?�Ֆ˶;�t��_�tv��CMY*�<s֌+o����N@����ϤP��M�o��k��%m��?c^��&Y�R�����1�%˺l�=��#�<�@L0Q"�/���F �����O��a2zz�{�v���/Lڗ��I�Q^>!d�V�+��P�V
OQ�7�T&e�T�J��-�.g=s��?)�7raK�'{m�[�v/�:�B]% ������Fxr��(�F��;��ֈ�C�� �G�����-���W�"<�M������W�}~G��-Ͼ�� ����:�i����V�E�����˭l%k�d������)7c��csm�=��O>Ͳ�V��l��η=wH�ӈ�JJ:_uǭ�~e��ء�$y)
I~������ra�Vu-��}�y���?�×�a3��̘1�Nx͉����y�;��mh�Lc���=���k5u�5�M����s��Ga�,.%em�8�-��]8UCMO���:�4 w�d���0%����2�!]	UC�-���U��� Ц`3�x%��Y�>�^����7�w���h�?�n�Z9
�e������{�5׸U���8�������> w�ֶӦ{�t
5����ş�/��gS�~A��;ﴃeR%[��E����l� �@w���[�~�Pr%e���n��ez�m��Lo+:w�\��׿�B�YT�����O�{��n��KG��BU�C>8Ak�Y{G�
�6�3������h��Z<�v�a'g�;&Mqg��������}4�~����JO� m�����;(����3�BMSZ�c�+N�x�>���f�j�rմe�L�R�lE��+�%}z��L�J�@-\tʇۖ�!Z��X����q|�?�S��ڐ��8|�͛WK��8�4���]w��0_(\�3ڇ{�\[;����+.�k�X���G�M��߃F����[
����>$�N�h�\.c˖,�����}�����w�o�Wڱ�g��S���6~�B͠�R3Z�B�����n��扨�&��~g#�'��5�J��\��:�.��"kk%��6���`)0�CC�E��~�Y������MQ�C3!i���������'�͉G�$i�\��@ �s����e�� ;��sN��g��-!]8`d��cx<�f�kc��|��˄0OYX�ކ-��Sx<�����7Y+q�'mN�$И�Q��Q��X��v��w�Ã)ثh�(a8|k�S�u�a�0c�������l�#��Ѓ���q��5�чɞ'a��5�F��cO>�d;�3\9t�X.c==y���m7é�.ϱ��ߙ|#��p�w�(����5���sN����w4mve��7���W��N?�4�o�}|�x�\��0���g?�(����9*�8d�}�;���w�B�D� B��n�{đ�+��	5�N��6!B"u���8�{�>��zp��h�bn��]�A�(�{0�C�q�x���E��C5��y��������|�=
�9߬m�c�B4U(�~��b�ࠏ?�S�[�M���:1YS�t�]p��3N����˗���w�=����/ae��^�����l~�����ӿ̐�s@d@�f�{5ΤP$Q=$xQ�
�5a�� PQ�
�i���%��jqL��S�AN�Ϣ��f���f%��d&�Ae��H	#������R3��I�fB��_��q���7�x�GQ'\?���ˎ;�8��ǧ>�)�&eQ(���I���j�����{͝�WX7�^������K��i��B6��c�?�9��W�P"XZ&?E�H�H�h�7��?�X|�T��k�w�fD��b%�ȐEA��T%�ap���KfS'O���V(B���ڵ���z8w|�����w�?�������0gP:�~�pSwE��3X��@�?ɠ;�s�?ȸ`Q<�����\����, dBs��s:�Н�_Ӑ�I��2�Z�L�6�IP�1���D�9L��E��R������{,�!�����D;xꩧ�+$���U�g3��lsn�|ˎ�4j6�ֈX'�
bwGwRwF�z�IO-�=��r��H�DY:^חe����P�?�u��x�Մ/��!*����N���1|�����M|(� �Bӥ\k�gl�L/��a��R���P��U6�����w� ���W���܅	<K=hk�@�ȳ�?��FB: c�τ��sf���K�O����1���dVk3q\\S�8h8C�I��\ t&�s9����`
@����4:i�ٜ[�ݲ#�<K��Se�e����ޱ&)������� i��ט=�u�{�4O�?���xF���El��'�7 �Eϥ����R);�f�I
�Rb�^�ʞ� 䂕��A\K�B��<#�f��c��N^P?�>��k�P8��b:NV"��t����*�^o�qo	�۪���zgwv�G�'U#�_�Y�˱V���:���L���f�5_���ٛ��f�����X0�zg�y�Kw"pTq�"�bw<�s�[vb͌y��-��ZІw帎��i�zz��@����k��aL�H`p=S���@?J�ñ��艐 H<�8�`�q�(:=��%z�����e�och���I��TEb�h���/A���~'YiB̕�Z��,v�B�� ᭆJ� ����@�q�-��c�T����9�������|��F��+��A����8�J����-���\p����U��9oٲeN� �!�.Ƶ)���q�18�ڪ��,�X��Ġ\oQp��W�Xv-7)A�/kU��h��2؎k����^8S�����?9��e�d, ���N2Syf(�M3�SVl���%tmů����E#�ߟY���3�z�į"!.a,� ?��\����%@�@�1�<�����K44�+bc��j�R�5c�U4�s�����+�����$ˤ�yZ��Fc��i9G|?�7�o 2��<��^d�����Ƶ����t�s���L��?~js�4O=
�+������
����c7��c�����$\{C͸�Wq@��_�[5�O@[��="K�-�t.�P
NU*߃�	n���H�}�e�fp'�[a(���A�j�["��'��MLw���O�_�g�/xA��V�ϱ~�Jh�M�=�;��'�{�ܱf�9k�շ�r�M������9��Λ{��7�Xï�~bs-6W� P���4����z�������2�!��Ŝ�Kۖ[��C��@JA#��M�	L�f���a�|�$J� 䑲�7�.��2�Kg(^�=���@��R&��c�C��P*�|3k�3�y."Ɉ�"�&�l�X)�G�Z����˂�r�eE�;�b���.1:�g2D�T��	�-������U�����������a�$�Q&�%uJ��p�4w)�RP
�R*bZQX bc�Z�VgΚqՄ��sf%�﹬����I�b�I+��%�%�X�/�q}���LҖ:FZ�6�ứ��� ��5�`��e�b�S$[j�{]�Q��1H�;�����k�}��k�����o�|�����p�KQ2^ԣ�40׺�K줓Nr ���?�$3�9AԒ�o��,$� ��K/�ԭ	���.S$���p}�x�l��WG_�E��T YB�d.��2XE��Z=z�(DT�0#�.Z����fB^����ɐ�V�G�Y��=�St�ش�x׎Ώ�0�;j%D86���SF7	�f�w+������6��ɒi%@�F�F҄���8@ I��uo��ב	-gd�o��&�Hi2����^��I0ΓbPԥb�/��͌��o��o\;�j+N~4�v��������!�4.�2 ���_���[n���Ϗ���	'��?�>��>H� u���E� ���p�O�k�B%YƙZ7�?k�+�&�LLKĜ����α�pl�O{q?��P�)����$�>]�L���P��l]W�RI�j���V"O �V[���L����������>�q.�D�
ԳC� ��19��=�QH���o�1標���My�c�&K��)��n�$��H���Ц_AIk,8q�rR�f)��j�~��Ό�ų�ŕ�"��b�������B���ȣ���[G�Gk�}>'A�"f�iA�@Fc���/�Ў?�x��hŃ@��T傡���}��j�r@�0�\�gĪ �\�k�h掁�@�� �i��Z�B�2�����
1�N}��A��k�b�\R�����O�aKD*�%$ejs9B�O[K��9�J�leچf�ҫ�}(�b8�w��>7e=�t����E!庶�:�M��Jоe�H�7��'��ߌ�g�\�M)�C1�|�{r�2��M6�&De���MY4�����G3�5Y:��M��^Z���2XEn�`���_�4�XS��>����$���_�����������?� ^P6��������~F��: ��H�BB|�_p����x�8�K"!��x!<�}xA3Q�W~$i�γG�/��WrO��O �Bk�H 8��K�-Yh��͍Rj43��y����'0K!n�+�)�y��J�`�,��RVJ����)���Vk�%m���-�
���rnsC�s���hj�Y�(D��f�'�\&`a��Λ�=��7���1��] /
��/N��z �OR\[�!phf�5���~΂���#-8������^,t M\&�g�ӟ�4l����e�������C�w�ԃ�'�ZOh�O>������
��K�U���hd�}������՟�ٟ�` �n?�n�kB��~���=a�5�r��w������G<;U.���K�q�G��1���=��8���m��b���L�c!�fU�y��UI�80���2N	��%�[�q��L%k-�i+W
V�!KUKVv�?g�
I ��M��$�������]{�uȍDM)@@J�h�P�"D
���w�ڷ͒�"���?g�PO9[Ўpx[�qlB"7(� x��is0DV��c#��2ɘ�\�SE��h��=�G�}��~#���黥5YL�hƸP헱!����g,�k�Y���a��)����:��g� ܧ�z��J�_�0������q,V�b_�tVׄʁRB�#נ�V�@2�9�nR�@<� E�i��\-���W���شO=�C�S>p�Y|���U�k�Vm��w�=����V�B�bm�f��Y;%*I�*K�:�g��a�w(/���=g]��XO����2��;d�y�1+.�D  8?q��2va��M�3�q�C���O�	�GYh���~�8�B���0���L��Ϙ9�	�̥Y��(&II4H_6ٹ�ז� Px�����pP��<��.���¡x�E�L#8�-�x˄	�F���_^�/�;�28cΟ���
\��g�6�r�\1��5'�Ua3�����%*ǠBݯT� ��b�E5ȹ����|�r*� �i���7���Z�f�U���Z��O;��8�Dˤ����Ҷ�������3@\�;��mP'h�:q�А�,S����u����ڊ]�կ�j]+��Zmw�'§�D�T�X����Ж����c�r	氖���'�x�+�̹B`����Q؍a(��1}�hMh�oV�G`��
��s�:�N8�P��2���n�ZK���|�,��utLu��{���2��Ln3�̖>���駟��R, w��WOc�_�U�P��Sc/�L �����e,�{�t��
�Sē@_}�.�Q\��=�� 8K��zNC&�8BD��d�i�şK�������_�Z�c[��5�nf2U˦�V.��i'c�{�IV*�[*M�i�Ǟ���@��5�O��Rٜ�R-6T*�50�+�T�h�){��Y��+�h����k��?��m�]��J�^�)�9��4�VHyd�Lr<�p�y	N�W��?����;��k�S�T�U�,m�&4�7��$��*!��s;��o��P�![�b�����قE�\.��D�;��C�SN���lk�v�B��tcΎM$�_�_ٿ΅��A��sbPP�q3���P>g�vz��{�s���|�Z�W��}B��?�K
@����]*�������6�4j�6'?���:�F/͚��lTzAsͺ��(�4u�g���/����@kF��^ti���(�_�g$� A"Kgx�|=#�'h��n �{���٩'m�j?�>���l�v���<CJ�t��Z�m��1�Z�H-�ݷ��Y�n��"�m��Gm�o��RC�*g���h���w,ߛ���Z��=���J���-Mt���[�i�C��d���Bi��j�+�B����ʷ_a���a��y��.��ϡ�at����;V`�����#�w�Cה�P��'4�7��_�(��g߽�?��&Mn��U�����Gg��5�kQ1LJ�[�v��Î��:�'��&�0>%6q<�t��ALv'-��@m&mQ��EM!d����أ'�V:p�4,�x����	��T��c	2�
���" �!�/@�˺�8]WB�ϤM*�?��ba�k5��e��Z��H8�&�6���&`��1#��!�3�ϡ�U���~�s�k�ԓ^m�r�����mmڶ;��`ي��M���e�mV,T����1c�M������P���gh͵Y��gK�κ�.�j��ҩ�u��ؗo����X�rV&��7��g���X�g<'�G�[Y� �A�-`]��>�(��u�㼟5c;kɘ�p|rr�Z���Ckٌm��L{͉����z�C_p��9Y��Yi�����|���F�>���ʦ�6{��v�i����=��k���^m^x�z{{<b�D��F*e�Ww���C6u���_��ӎ	��~DgP���#D���	Ĺ��o~�I8����I�
����ϕ���S+������|ST�P��w�ѵ��w��a`�������@1S8fY��.Y /�'*�*�����
J�=�/��"
(~6	.�d�����xw���NT��e3��}�k����J��*Ռ��v�Y;�DҥlҤ)�΄օ8|{{��\�����v�P �{lh�ZrE�Z1���4�c)k��]f7}�[��b�T�U2P��T! 4t��=6��Y/�5�
�V^���}���3J�J�s�8�^RV���.[��{�鹶�7�t�?T,��@�֮[o�춧�~���ʹm=��[o�x XF�O'y��}b�z6�͔I���iӷ��2���w�=��+v�R��-z��}\S��ށA�Z�e�r�-�׽�ӳ5�8���-��ވ� �����pCy�������/x���!�|,ir,����j�c���Oc.���{hl>i��$��<v�BH���c*�O�P�S�0�"�!v��z�N��K� �yLO�7�*�/��{Z���;#g�$�3���<�4E�o�R�>{����I�=���>�fZ�c�^��nX[K��������R��P���´��&O�/�io)YO�E��/5+�[&�f+��K7�a��a��"�ԁ��y�u�A	c\Q���%������2��>����m�f�>�kKY�e�[�x�w9�500d�m�mɒ����V�Yo�\v�t�V,V����[n���h���&4�7��K�1lםw������X�w3�?�y����c\SX�|�5Pu�?���/\l}�f�W��~�b�z׻  z���Hh�LL6� �٘�9��u�U�\킀�!�nEn����8uƂ���?6�v��f�c�޹��6�w�99J�Ҧ 8�x��f��`9�b�&���u�����t��9c���Ɗ�QB1m#��A4�^]�T+���X�H�q�;�3�v�%{%Zt-����
���N������'a�r�U���.Gٔmw���oZ��B�J���th(OC����X�0��{��Y����׻�o�d+���7�ak֕\�SF�	�    IDAT�����_�>ߓg`�E0�\�`�PY�ˏ�dt3�(x0X�KϷ_?��}�����Y��s�u�;x��l�=�س��vؚ�}�������v�k�+W��<�ŋzm��"�W���s���lOw��F���Z.�>{�e�|�u�Mm�������c�y�ў��l�"����	�d�֓�%K�Y��j������~�����v !�����y����L����H<�y��>��x�v0�C�9��scC��[��r�4"J�F��{��>��̝�hb*@�W�t2_
	i�Ҩ9^��|��/��:�,��U��}E=��~=��Gk��R%(�N��_^1=U�p+%IЮ��Y �h�T�:�9�N<�(�z�Tm�=�:�Z�gY��/:��	`$w��������� ��YOOޓq�����Ֆ�-�j���{�k߸��v��b��MLmE�RԍVI<���d=u�Q��o��6/����C^y�^}�}��f�n%�Ս"8�����_�mGq�M�:ٞa��*EwDS�(��g/.Xj��$[ݵ�֬�O��=J�ZM���{���|<�-�a%`��o������c{���X.]�%K_�_��#;����R�ŋ�@G�˶8߿h���ڳ/���~�Wgd�����?\�h��ꪫ<��+�q~��pΟ"]J�  �(�J�l���q�V��ǠG4�Nr��$��o�� �l$H�o,�w�e����˚a��S�� ]O���|�)��m��@�?q�|VuZ��)�ɲ��� _����	�RB���[b!��#�w���W!�
��5�,U7�v��N�לp��J�VI����l��if���0�=X�sV����RgK�����2x����P/��
C�V�H\%m˖���[�ۖ-ﮁ����o�F�����b���_�c��O~��W�r8�x���|�#���z �������~�=;�l���J�h�\������-���Yת^�d��>�i++V)��ӟ��-\�|�*���X9���\�p�V1C�Y3���|��V)z&�7�q�w����UK�o}o����D^�p��*-�pi�~�1^G�����(�t��l6x`�Wac����Ss�=6��Hӓ8h۪�7����? ��;@2wp�l�_��מm)�Z!���UV��b����/�ιd��X����,rBD������B8��X��Q X[��v�\��ƽ�YOj��#Z��F����G���R��R�;o�T�,�1�Q��]��l������9�
C��ɶ۔�{Y*=9������\�t�ޝ���{�X9+���0���a�������
�P�ǭ��B��5��ׇ�|Ya����{��w�XSO	
������^W��f�c��"�W�Xh���ǎ�Î3l��'j��Ht˶�ܧ�Y�J��m��N�go�¦M�i]]��N^�腭��h
�L�J��I�f�d��Km��w��\������Ͼ{�`��]���4����x�R��Zo��%{Ӆou�`C0�ԭQ�8����cs:/�¹3��h��).��7��V�o��f�% H7��T�C=T�×FkYr�rGE�����
@0 ZD�!���zj�E`��gb>w�K�)�A�?k�{B'��  ��L���r"J@�kp�]w���p-��~yQ/�u�f+�(4{ u�_JX������W*���%����jf��b���#Z����ed)���@��U���r[�R��[*I����c�D�� 0N15w�Eفh�W嵳P ?����R���B́�&��ŖIlĽk�&������18:�l��նx�*��ڜ�7�QGo�t��>���緿S��}��U=u�J�&��3O�׿�4*���}���l�e���L*k�\���Zg+��m���|��j-����"�ŵN9���j��{�q��a�c�N��x��s����#(-Sa�lZJ{ �R!�����<�N�����bߍ��f��W	��:�ی ��Z9�ro9��q��g���# }��|�߬)�G�>פ�3k�sE��i+�D�EMd\�H��C�C�1]�G�����p�|�G+/�<>�R��M����J���H����B�E%�s ��f�3BI��uPM	�I"��$y�9GFio��G�n���<R�A@q����q�E�\��o�r+��.�[e�kW���-זAY�5k�=}�1y���^o]��-��oo~�%�݌�\J��w|�~����5Дc���������[�\�?�r������9�_����6�×����O�`���ˎv��o��ӦX�2d��=��Þ���i���l۩����w��;ʆ
%��@3d�C�F0��DBew٤�+N��墕�!���G����?����3��(hȊ�Q��;�K\U1���#iD1���hq��@������ơ m�K���h��%A=)	`�U�
�qM�����x�y���`�p" ��{�zR���� �zQ#	3W�+������'Y���ݳ5*��y�н�
hᐸ݆'
�L% �?k�U:C�^A�'1ܴ%� �u��ט�g}0�c,E�$OB�����c0�(x�;��x㍶��)�^�d�-x�9[�b���-ז�l*k�C�6y�6��:�;�H���N��jU��t�Ͷj�jǯ���`fwv~3ߓk�hB7����N���>�.��ki�X�z+�����'6�U�8x�A�ٱ��i礡�~;X�s���J�\B����4O{�����'_G�� [���S�WR�X�������U2��#�H��[���}x`�`�5��.?�/-PU,9� �@q,稜8�����Y[�8��(%\+Dk��*��{��f]J J���)��
urj��֨k�������Oi0�.Y�5���(Y����ܡ����h֠Jl]���U16�����7�D��+�(g�X� ���1���1c�Q
����lp`��Lj�+���w�e�}yW��:m��6u�t;���m�]����^f��q������En�F�?g��������S0C%�8��'���:�u6���z{�[kKp�6X6ko�_�Y_���P��~�;U�A�x*��BaC�,��niܿ�6�2/�H�M [��9�3�w�^�:Ná�V*��ŝ˪�󷦕FmE��7���}� �F�����UF'Bց�����u���@����7@3�:rfs�"~���q>���ǰ�P�$X}���.r�A.��i��qkP��AH{�ɰu�ţ����M\���o�;�� �[7RR�sr���Wj�FM�4X&��J�HI���t	�ׇ~�)�%@��B@��(��ߡ�O?�u64H�G�r-T~�vE��E��nc;ﴫ
���p�i�{��ahO�I[�H�k�WR�ab�>�;;���ɿ��.6}�v�h�y�v�i'������!U�g" 6�SO=�� ~O?O��)ڇ��?�����W�£X@d������
4I( 4:O|�V����<q��`ߏ��=+�s3�6���%�� ��ﰒ�S�$��|B �D�p/�s� 7���zA0�9��>` �1ψf	�@ @'r,4��s��\�Ǳ�[օ ]��m�X�xP2�څʀ�E&?	��9�j�2��ƥ��$�zR8w����	�>��B�}���������哀���� M���>hN!!,K�qf?3�8��8�o�� 3?*���>��{��z<(ԛ��z�ɧ���g;�8��|̳��|���}�1i�Sy��|�������Γpk�ʷ�C�'K18�B�謥� Tڴ�^g������Kd{xm�G����9�=�����#:�J�|1� <�lhLB6�/���������9�n��?�(ʹ*�K�s42�wM�R��ߥS��U`���%��a�3�̭Z�1�k����3� ���h�h�QQ�P�3����7�FP��$�?��5���M&J���V3��Ij��+!�)���q\g��c�<)����M��Ki��s�GO�I9�c9��4�kS�f��u��(��o��M4��$%�k��օ�O~��v�]w�~���+Y�{V����gM�A	P>�"�v�q{;��cm���9�-%�2tt��=��S^.~ͺ���*�vL	��dF7��gΚq���~S�q��s�t~�'��htͿ���R��b�r�!�'�=��͂$n�P�+�8������C(�����a���� �Kj7�=4�K.�������%{lb*�[aS�V�{�D�H&|�xw����"`�?��^�Xjr�h���������@փB|�+*��կU{L;q�k���N"����*�W�e���RX$|�'X<	�'�S��寪Y9��y�������0�k�W��^�`��0��2ou|-��F-�3�{l%�<f��|�U"�'^'�k2uk"~�v��; ��׾֕;4*��ЩJjd vS*>�
��P<4���|~�uw��|�$	��o�R[[(3aqo�Q�����C�XXmI|�����n�9fk�xQq��c�ɇ2@�3���dx>��N]s�5�9�}��j��7׊�!XDlLg@��������29�1�[m��ix��f�% d�|�S�rK�Yw�$?%�c��p��E}��qȋ�q�^��ω鎀�8�Ѓ!�������6�~|l
��>r�J��X��1��V��յ�@��f>��H�c�%��أ�:�kn!9�%P`В#�?���<QK�a��k�BeCoK�w�]F]\�}��KC�N���t������S�=����'���E�/�G�F��<jxѲs�׆j��˨�<��4�S �w欙WOH�������{.l���}#0LƆQ	A�	�b�VE|8Y�4�V$��=I��?�s/��v�2��Фah��Ѧ�
8��B;}���~����}�V�lGi����Р�0Nd�G[4��� x6At��8�3��˓���Q��J�s���$F��s��Xq�����߯��$�����f���b�������D��3vs.kF��a�0��^z|N�L�� �5Ф���y,(�^@>^�̔�4p�Ԭ�@Ŗ����)f��P�m���9�=��W���$5�j͉�1V@��/��-��ZK�
�|L��~�(���u�?�/��{Ml���%ߓSc�	>��l��R5�lD�Ol���i�M�?N36p~,���ȩ��� G�L{q����Eb
a���"�t4&(�[��-�������8xd�5Z�5z	E���B>c#�̜�<p�18�2!��)�'�G��<v��3L~��㇫e>��蚪���̋gB� (P�����<�� ��j��<E����B�9�lt*jJI�y��x&	]Yc���"�D=%eFV!�s�@"`�.���l�40��1|ox��Эk<�Ϲr�K�I�3ỏ,(~���o�A c��FBIyc��U�c|f��	���,�$�����w�ynRKsd���]M��9*-K� O�F��C{h�j�)Z��Y����{�:�+j���F}��^2�"P�[���E��O�<�|U"�K��><�B$�k��]V  �s���K��gNI(㧴a���9����"�T:��	8@�8��?I�=q�a"���z�B�)K��~�[���Nn��-�z%×h~P���Pn4�MDՉ�A`IS��r�+p��\�����O���Xh.CUP�:��Q*&�w5=���i7����+ƞ��	sc����x���6���k��fb�'0�"U��T��C�Ģ�糁y����)h]C�����1l�Z�i"h��67��Xm�,
QͿV#q��Y]�.�q/�+ A�:cD������.���g^T�pt�o6�cO/�7O�J�:J�����	o���d����Љ����Wq�����6�����B��f��y.��uyv :�s�.��_~i�Ϻ�'M�x�y��K�9�Mx�����j���P~g��x.��b�C�I�"��zI�F*ž��y����8]��>ße��Ev�-��s��4��p�&���ԯ����#+T4m}C�F����'�7���Fm��i�	���8�e����E68P�����j�-Pa�0@4%�H��8�
w��y�������/oX�Ζ�����$����d��Ҥ���pH����qrj��\[N]�<7��	ϕ0�W�) �f̵ J��$.Yrr��LkO݋��YJ�R�g	<���@�����}xO<;�������d�] �:Áy�A����ȓ�@�B�q.�o�w�8i�|/�Cd2š�Z�::s�G��"p��-�_*�C���}�(����3O�z\���W�%���4N
`.D5SNF 
5�^�~�
�1���wD��(�A����h�A&���K�!h�ld5��si�V��1��,l4=ř�@���V્΢��rP�D�/�7�m��N�F��ܺ�k��ъ����_��X����c��>�y�<�( �U�8D��&����̭曹��&�Gh�P9
��oU�Dx ᙹ'�����e��s:R*��15%+�u���R3���|b��L3�C��,7�A�<����^�7[�zUT	7D�[ �Q#Ifq�ŦM�nm�>��W��/��^*ݩ<��o��/�#���=}&z/����b!!�b�<c,0�	�f�~Bk�c��7�z]C)[� �5��Y��@�4|i��6��r�rY ǰ��81�R{��K� &��.�f�� ���t�fZ�,�!@	s>�	����|��4n�A�.m�EEc^x�>
I߇����?~�[J����o t�K������;2����X����,XB�S�>�g�����EY(�RJ �
�s�hA�N��O����`=���f���F�'` I�c>�`��#T�>=!�*�)8��Җ��l֬�m�?�Ψ����CJ0�D���t�8�'"�_B_�@���W�ޯ��	��[���sD���#��3g͸rb�z6)�6q��e-�ZN�@ҦT����X�\O{�簨��T�M���a6�;��@1�2'��M!}'͟��YX�i���኱�"EkH��Oir���U$��;]W�%�CTB�T�ȱ�N\�8%����Xm"}���T=�EK��E;4N\Ka|�uUs߿��Dhh��H�_Y�������xZ���3�|�s���y�=.��g ;B*	���yF5o��ǪDH�"+ �
���!�<3>�I���M��g��)�Ce�1��\b��GF,%O��޽��U��Ο}Ʋ�S4��a�n�������-_��È��?/�j*��p��֐�{	I	,�X�|m$ٕC���=*�r<�+�=���`�(	o��Em������v�Z@����`�y�v�I!:�J�k�V[Oo�ggs�����]� ����=Ĝ�&[�D�B� �-.���Х�iaJi��ڸ�X4A��:_Z����o�K�u=	�%=���_�a�kSmI�g\��3��c!!��g��������7��q����8t���ԙw��́"� w���#׵��3]	@�g�p��x�N��ܗ1�;�y\�.^�[�B3�;x>@��Pj���0� @�X��VD���
5��9�Ѓ�"o���5��D	8�6B�p������h���RY���5��/<��e8l�����<)r�'��%�N��qh��E�tl.�q���d<j�Ak��N���'�n,0�5�1K:�O��ϔ)!�pg`��AK;�������B�z�lhpО�;��1[�l�ku
��s&��?J��̣.���"b����\��h���c ��౳Y�4���-�A֎61 %kF1�S��H ļ��@�1�Z	��'�%�_�Z�w(������[C7�p|r�z��H 0l~QE\S@��XY<��=�9�q��:1�$�Psm>WY*�z    IDATG���{�
�^d������r�yzO�{��Eiq�rR���֐��|�;�i�|�V.�?��*[��n|����Y�~�lR�?~��n������~'���e݋��w�:s.g�[#IiW����X�d�c�M�����[���γ��	߇	��������������s;����_"G�4L-D��������4�a8��C��K�l)i�yY��i{q���/~�i��f�$�� 	��l^6*��hhp�t���'�$j��C�F��~i%��ka��9Oe$TZZT�֭�$�44rT�P��Q�]�s��X�m*�I�%�7��g���6�(�ሿ���2�f���ҸD�	����%�%,W�Y�þ��h ��<���`���@�7�Q�9�&s�0S�/�Pv|^�!���Hg:��k�tnSN;��3N���/a��J��(Mc�5nex�V!�Z���:��J�OL���)�-L�@N��E�*a�g�k�0�<� ��|��x�=QVX����9���;����K�ٝ��/W )c�أT��n���s;o�i��15&�EO���k�w���� �k�Hb^hlm�9+P�m���Z�}{��&d�����}�Cd��qt������I���
`�|�1�C(� uxӄ�Ȣ��8Wi��% `�'ϮD��;A�NDY+�4cA��&Y�L�"ekSIK��-�������L*8�Ѩ�bQ�A�4�ҋ���\BUVS���$ 4��?:���I�g�5M	%���<�E�i���!�_V�)O|���xM�9�N�_����GZqpȆ��e	�N}�j��p-�c�whiks�v�i~.�>p� g@��s�~���}$|e��j|�\%<�ȘB����y������,��T�M,L��BHպ��ح��ns�>�nO�k٪�7��:�t~�;�����ς����3N;�.����Q�`C�}�����?u3��6}�ǃ��Cl���I�C&�x	�㚢C(`�$#͗ʞPI4{x��_�E�ЬT$�x�����$-� �+��&���*G����Ǳ,T�?r�/�C�ݠ�dxg /��4�wBy):������f���{�]J���%i��1"��R
�$�%4e��/1� P�ঐI�ב��8�l�(M_օ�Be1�>��/IIF�3��
VF-���-?�,>�S����:V	d�{�Æ�/�u��3���.��?�iT��tu��=�(e��^Ƶ�oPl1奧YcJ�"�������z�2��;���D��ڿ�Jnd�xF��`~(��7_dS&wXGG��9���#�sK���
;�#m��l��P��>���ZWW�_��i2����3���|�Ս��X�l�]w�ٮ��Z�2u���d����<�+[�n��n���f���vԱ�ٌ�;��S���;�9~�T$��� �f�V �y������W�8�BZ��IҒ�*s\tE@�pB5�fA�*U�J2c��3�8�s��� @������Y���L[�c��Q�%pR2�l~� 'c��R�8�oi�G /�� ����ǪSct	'#�~��$��;q�S�=��+��se��)*��ay����D�`n%�@�DH3�Ж�Tm Y�(i��ro��i0���ޑ�QLX�N�̏��1�'��e%�]Y7D����;�_���w���e�"o�@�&��Y��).^�eoi�GQl��0��'ƛ�ZI�i)����m?s^=�Y��~���z����8�;�'�:�̳�^�T���h7��U_͒$'t�������{��6��-�gLJ����O�޽��=��\[�����`��q�-����U�l�̽���Z5	 �� ��(��g_�j�0�p�X �����E"ڠ�O(��Y��}Y4lp@P�,N4o>�"�cC
X ��h+���V	�(-�c�X��!�@)^�s���@ı,r��x>�%@����#��Cyj���A��{S�Ǽ6�(t# L?��H(�
!� 楱`��L���C��Q�r�ATcƘ2�*Ɔ�e�'�n�B���I�$�D�����q��K�zi�+	�f���X!��K�j���lHn+�J~����4��������ʅmʂc~�����Ip��!�G`̭, �7�Ǿ�={�����Z�E_�'�>�}A&Mj�� ���i��������v�gy�����q���zH�VͿ�̞3�������?�&ɤ�ɮ�Ϙ���������]w�e��l��EV(�ͧh�ۇU�cU[�v��=/��4��6��j�ڋ8r�E�_�$���~^r>k���=�� �?]����\� �hҮ�[� ���D�R!�A�@6 �6�|/��84��4{�� dXPb
��9;ƞ"� ^X�S[�����pGp�Mw�N^7��s�cm>�͙c�X ��+~zG�LƵDQ-�=��8�ZB�p��5�ye�r�1��!�$A]��;z�.���X��C�^� -
e��7�x��h��2#5b�t�Kb��\�ԓײ����y]�J�p]E�q���z��}]?��5�=뚦8L���/� ��Ų+�m����@����xɋVA�kZ�RM��E+��l��e���o����ו�{�C�6#�3ʺ�`���ȴ���OHh�]��?�{�*%�f*������t�1V.��E���\�i[���V�\g�b�.[gx�;rj������,�йP�3�I�������<�T�qj����7�KCf1�)�bt R� �~�3A4n�h@y@����;�	���U5ZK+���}i��>���3��{��#\�c�5[���ϳk�а��F�g\����b��������v���:4�l�XQ� �;Vt����M��jn��-?Ϡ"p��^ ��h�oE���s�K��N�g�o�%̽�L��M{�S+o �y_��~1t�
�y�.`d�# ���
�'%��[ ���Qx��|w,����σ:XÊ��3����}���`�ux��3ԟ�_��m�ݶ�i�;�g���"����\���y��*�zM���>��K.u*k��.o�l��Zص&����	M�t���\w>��F�?���g�W�{nx7K�.�g?���䓏�je�V�Zl�{�C͕T��u�ڲ�]68d�t���+��pL�����ᣄ���S� `Cv�a.���tg�Lhmti��4mD	iʘ� ��� 0c� ���f( �}�'��Nc��A��u�h��f)��}�B��0���1B0�q��b�Z�}b�I��-� ���(ʉ����k�D�W@�� ��;B� ߈�r�s)�|��=� c0�Z<'Y���.��� o���%�'�P�=��C���R�����o&b������{���w��?��2����p4�{��c�QV���>�яگ~����e�w� hտ�˿�� ��1��S��<�����;�C��Y�O�y����\���6�_�g�Y`����.��N�����������������hNa�U�o��Wv�y7{�{n�L�b^|�~�����c�R�׺V/����\��n]�-_F��6{a�:;�����x�ob6%�ڕYy�%�x/� �x�|h����O~�V��E�H!~ ���E�p=��j�9*��DE�<p��@y��@Bh�@(��P:�g@sAh���Z�|T����#@u�<��=��=TE��Z���O�TV�h8����|g��;D��S���`��F�W�NƇ�� Tm3QE�0WC>��������o�9繘/���،3�@x0�Xq�~�G�Y�ԍ����q/jN�Ys��P��=h��p4��p�ui��ǅ�t̖Y7�s��Ϙ����v�[|%���͚&G��o�����H��8����+���ڡ�c3fN�^���2�A2W�����-�r�Ŗ/�[�P��|쟼�iw�:���sYT�4��̪��c��/t���4�Jp2�������h��>km�ط�u�w�V.���e,�_k�����Z�Ζ.]iUk��K{m���eeX��,�h���7|SJ�C{@+���˜&��i�h�z���XXrk�� /�f� ^�L�C!�h���"U��o	�)�����������[|��Y[��u#�5��ⵡ"���~���M,���c��������\Cxa�J���-��y@H�G9n���x��k��V��Q���S�;j�uy�)kQ�g�y�x��!�'�h8͕H)&��-���	��	������ܷQ��%�K�"?��k���~�aW�k��C�A����(���J�͟�_��9{����C���۴�s���P��R��E֞|b�����_���d{׻�<��*��>�9[�d��q	>���c���ZҤI��w]o;n����`?���e��T���k=�~��,؋/,��]�mmw��?�-^	&$��~%K}�c��s�=�Ԣ��E�H��;��/[��ə�8�F_�`��I���|��L ���EI�i��t9ͅk�q	�Pf�d���Ikk-bHQ@�6����; �u��I�S<~[Z��{���=�??�S�9+UVL|��P����!h%��c(���z�}���a1��b���Z�2����\>S�#Ń��`�<��(0h���j�!�>t���H'	������׃�蟗r�M���;͹|=��1�>ڵ|.�h$���ކ��j I¥�3��V*�����ȦOk3��k�J�z�j �,�j�y�X_�Vuu��g̶SO=��i
eOo�֓���������[�\?^�tG~)C��?�Y�/�]�ٙg�n��>�z{�Zo�:[�f��^�Ԋ��X�
�P�����ޛ��]����Yg&$$B"�B�w"�Z��IP����ź�o�׶�����V\��KMX���(UPA@�%����6g2�Y��{?��̓Üs&���f�����[�����7R��n��$���]^���Z��c�5�h��[5�Ź�lX�9G�K(��}�r6i�*�`S�v�J<��^��xnv�h�C��܏�b�'�h��{	E#I��<�T��V��'����u	%�8�ǻ�X�����L� 
�8������	�J��w	͋�8H���w��%�]�KBw北�:�����d%j�c'&�AQ;ʚ�w�}4ǔ�@��Dsƻy"�~Z��0���N���(��yz���������/E-V�� ���Z��S�#ʕ��E֘�%]P	,ٺ�)۸i��ض�JղM��[-�����lp�j+�Zk[���eo}�͞}�U��~�;����l�#s�h�,��_���
��w4�} 6p�Cgۻ��v;䐩V���y���l��uT7������������C��N{�2����>�X�;�0��+�ʿ�Z��7����/���f��6��s�Øwf#+kT$�H��"�A��7����'ϣ�mi�Z�z�84��^�v���6)!$s_����eE+�~��������VA���&ca0�H��#�� ��3h���w���u�ݩԂ�c�'��X�`.8^�ɵu��+s�υ�������<��k=h����]�G�:��?~�;��W ��E3����������G��k\Q�����̄�rX6@�Y�YG�j+W-��+�yC�O2)UISV���u�y��c����`9���o�b�Q���V#�Ϝ>��ŋ_�8G��5�|��Px[3��dj1�ɋ^h/y�mBg���)[�z���w���k���-�-��ڬٳ�����{�M�p���¡B�P�MY}6�e����͆)Φ*��/�C�A�C+��6��ٷN�H�i%[`  ��x�7�V��.��K��I˽����J�����o��d���w���v�W�X�I8�z
���9�o��OE�$�~�Lڲ� e������" �oqss@�#�j�K�wZZ�Z?z�V��-�+Y\�x�Ю��s��Oi���9�_,9^����Z��U�,z�}4�d$���9w�(Ǘʡ�&3��L:G]����Ю&�p+�?������}Bg��c�s#��[��=��mdN����E]d^�r�V�^����,�e˖z1��g�9�y����̎:�y�7���w����Р�}=�}���;7_w�������P���f�/P�=U~�$���KmE���P�3��߱���cƌ�>�^�;���l����YX�~��}CSo?�'�E����rE��B=y>ORK���QYh�W���?���;�/?@��wh�X�y�X��CDE�rs��CWI��i��(��	�h�����|_�?�'n�g��Ϙ��V�Vi쌯Jr<mc%����s��BSS�Ɖ{ro���+��9
�9��^s�8�.�*	X渝e"�wAc幜���I�B�B*��y��Z	�X IK�����Z�\��|βD�O,������pP�J-��0�����)۷\Jh�&�ߘD��.<�T��h<��ݗ_� ؃zn�(� �v�*�%�O�l��vt۔��G`��#��b`����Z5�wt�����?�����B���'��?0�����.���)��w�PŇ�r����7�ѝb+4�����+&tǎmo��lHi�L:M+�� 
 ��[��V�U�`3�~������4�j���b�1�<<?��;�#ԏ���R���� Y���Ȋ xV��h�h� ���(�#\ �����w��g�TbB��8+�������e#K�f���bR�f=��k��}��)u\�1㠕ƈ�!��3��zH*zǆg-	LCƖ�b.9��C(sՐ��J��J� Z�"Ɓ
�D;�7��:4s��o~SO|��P���t�Ӻb�.������{�΂mZ��K��ё��M�b|�?�Z(��1ɦΘi���\���~���m��-�t�I�3����+h��+%G!��Zan�3{�t��"����c��;|/֟<�Q>x���e��X6�	�lGֺ:����R(��u&o�����?��;�Q<;:r������>c��nY��+��ߦ�c�[� kq�c�R����?����d�׿*&�����ʖ,y�^�%v��G|�]w��ݐؼ��ԅ��
��G�v�-A&�q��N���zQ�@�I ��ffa�0
��w�$#�k��.@Ģ&I�Qug ! _�HBR�H��
�8��1�t��3�q��V4Ҿ�}ėJ����:V�q�Xm���i�����T�&����g�4�'Y��	�)T�XT�[IZd�2~܏yc���/��a^G�S�Z;�Gt� n�e/{Y�i$��G�+k��^��C����%!�(%��sϱri��{�~�*���\&� �
��ZMp=��'b��Cմ�>�X�5k���6l�b_��{l�A覰,����#�u�%M���.�>s'kPY��Ε��P�s���<���ʎ:�9^I�=�N�c)�LV���ݕ�L6������ZP?��߮�;#m�IS�~�-�|���>@cp���*Ւ�\+S|q���I���|�	�I� 2|���x�� ��-FE ({Pe��w���� x��&͓{ΊL@!	Iڦ�F5o��`I ڪ������Pb�Ҍ��І%(��c�S<����Yisc��|��u��[���-򪬲H�)�ڌ��=O5c�Y+l|��f�'ƛ����an��5�B�C �@�ɪD�o���܊���=@���*�����P������������[b�u��V�Zi�6oXo}=֑!>�b�r�i4M;r����J[-3ѦϚm��j�j�
�}��k��ǟx�)��4���E	�� ֘񮪃$�]>1/���7�@F@��ɜ����#�������p-p�`��g�Ppq�[\�#O��m�f�*W��w�C�W(��UK���������B���>���F��
�;�x�5��    IDAT�B�g5YV_�R�/���2�/�i(����O�����^;Nk @$������rN㚊��Bi��(0�f/�Ţ�z"��De�*_E�x+��H�q�𾀓|	��POT�~W�6ׁ���2�5`�;C���{_���~�O�u%�>��@	2_rFs,Z�֔@a$��Ɗ��'|�o*�J��7��]&�c����r�s����]-�s��'�Q�xY	����?���=�[�@�M�r���w����趘���Q� �TyЬ<d�V���7[�Be��[��'/��CCUO�*��Us��9G۔��:�wz�_�p�=�d���!l2��.��b�Xrq`�LD�%�}�}�K_r˝r�u�]�E�"u�1��͘8U4y���o���PV^�*�?)��P�A�w�'���#��6�g���)�����=>��t�~ܙ��ģ+ X,�P��j�] ��OX��~��C��Omj 0a�Ӳ��f&���}��"o��3�i�5�U��X%�(�H}b�q�Qy5�V	e���`��,P����Uw82.� ϳbEȼ�;@�s�O}h?5$G� �|��/�k�\�Uc)*l_9|���i�K��&驿��#��
��8w4:�� p��\��^�U~�VI`Mh#�S���3�|�u&ڌ�#a�Ԏ�Q�'ϫPN �P2@|�ִ4����J�h�D��+���s���{,���Ƶ���c�ufҞ�J���~���8 תVM�l03��3�&M>���i�6��_���VZ'J]RZ=r�֚���|<ק?�i{��<�| ;�r.�k��}�<� d�3�Y
R�<d�X��4�D�|N�"~��}),�5�ã|�7B����Y	h���}*�g̼�L�j	��M��W/_$9,���31 VtO�P ���*�aP����������y�Q�i7oݭ�U��I!ڠ]��$L%TR �������� ����DkDp����y>��B&�@����;4Gq�,`��g��:��Q)��V�R܋��Se��K�_���g�]c��͏S#�q
%LT*�;|(�h�|���YT[�8�����P�*��5���fYc�J�MF�h�N\i���M��%��=�X��
�][%z�K�0N�Ԁm��rV�5�V��-����Ւ�,� ����TΪ�iv��ϵ��DK島e�v��k׻�c4�����?�'i1�j���O~�֬Zm���7����~ʂSߟ��1�Þ}}�k��D]ʊE�ↆBX1��I2����#���Jz�|�O�V�̘9��o���_k<�}����,*t.Q�'��	��K8�Ɨ�$c^�b�[ȥ�l�i��f��|i�, �8\����1�i���f�������s��sU�+�CX��N���1����E�v. �'@��@·
R�H��X�*7�3 ,q���� � (Y ��u�w���x
��DК��G ǽEY�V�C�Z�[\9U?U��Z(���������{	��h-1?qKF��|2��sJpKH�* �IDOi}J�ig9�{Qh��yN���i'�`��+C�~��c^�����ͤ�����A���?q�A���i�7m�k���=��S�'YJ�kY	�4Z͟{K@�;DΡ�S���N�(��0'�7��/��/�-Z�w�Y�A�Y򱐕BJ�N��)�(7R�5�T
ڧ���ߊ���-�I��a�g@��ed��ؑ�zh�f�6rp'�����l
�pπ�J5��]K�KE�p��.�f1�%\����z��,�&��k�+-��%
�N�)�x�[	1Q^zY>\[��! >��w�j�tہ��~��k��ߧ6.�)G�@V`�؈;����A|/ �z�
�JK���{�ΕI!�����R�RxX#G=S]�%]��.�x}����x.5�܃:Bg�q�k��r�i������W�N��.Tm�6�τ����߶�`_������K�ӹ �{��+�_�_
��]�� �1g�ׯH;|Z̟�nY�Z�4��A��9m���8vi���@5,�)Cs�j�[p�8O ��	bT �2����F@j�6��9)��'<���:�Mh	���L;�ԤM	|���:|/� ˃��9��:Ց��Ε�(^�Rڹ�M��Oi���j {����3~�����������v�Y����x��4F��"S~[e
�X��Kc+kP�1fXr
�%̹����@V�"��%4W$F����<�-��;�z� %��8�T�Ҁ��l��ֻs�u��CA=�\����;X��G?�&O9�JՊ;|���km��-MYD����h�I�/TJ{Y�1Zl5s��B�+|r��}:L�p�D��ĉ��aǡ�M`(��aއԑ��8���n�&�H�x�w��'�$uК[���~
��EݼM4yi�,8w6���ht6�6��G��1�h�I𝀸t]I,��2��'�]i�a�,:������������g�<���qכ���5��[�RG��(�4 |���d��=�y���%KB�p�rbK�yD`-p ŵ]�I��@?^��;vr{�H��²���Gkݶy�-�ԚC����gX�<d��۰v����p���X�])��C=�ռ~��6��Éذ-�wؿ��ڒ'���	�] ğ�̓�	u�g��-8hC�����+�H{/�S���Byaܓ(�B:���q*������<��7[��}�å��,�$��'��A�%����Z$o0�[�n�|E���<S�x,xb ��'��Sa�X[�5���y��Z��b�ǀ��γ
D���Lև�_����k�1xb�ƛA�I ��0�y&(�_�>�<�1��V�A�q���X�J+�/f5�r
�u� S�R $���� ֕����K1�wAP�+���V������4�����M|�YgZqh����n�`�};]3�=��}�zy�9N��6���6}�LO��oL:\�f�lϱd�j���)�Z�{SV����֘�Ա%1]Sub`!���+K�-�,�$A��l�q�g�U9a�8�����3�N9�6s��I-Z�9ߛ$X���]i��9�L��� TG(:=�|/�1��c��5�H��4�F��X�-Pӂ�~Ah��&-�V`�0��5��Jck|T\_QJ������#M<�}bMZ=~e�s�6z��^��K�Z!v;�hT$�֐Rc��<�^��敟��@9��)jH�C|s���ח/G�+%{:��x���8�=�7e��;�s�\����?�{$��p~���/�L;�&M����t&�͈z�	�{y�x]�oQd�?�B!�!<�)T�$V�4�u�<���%�v2I�"ǖ� �#k���Z�|vu�����g�w���74����h�6�_s3j��OU��i�!Ty��uV��qG��	-�����v�g?,��Q �w�7���s��cmN�/KC�F ��,J 8�2����%bm/�$F2y�1�Ij��D;�D���p��]}-#Y-<���B����I���S��4�=�UP�B0�!k[m	�T�:귣���+��w ��� �t,e/���;�Xo�7$r��wYd�����w�q�\�g�6�Xu�O�g��?����Li7V#}����֑�oϚ/-�U=т��"�R����rŲ��l��e;�Dh��YB��aa7)B̑�]މ1�
e�Uԑs�N�_�ּ�0��lG�[n$l�P��;r!����CuR���X.��a��V~��X�o]�!h�>95����7&o޼s��Shf�8�7*�*��v����,&Q�>ͦ�?����c���wo�Q/�&-J=�x��ħs��?QA�P�֢��(��ck MK�]G�[�}�����^���zҤ�;O�2�}M���K�$�s��]*$��*5�ԛ���n��;���@����_Q�� B���o�ݣ|h������������A�A��AV)돜2K�l~��_y�!�{��_�E�PD��d%��q�����T����	��Z�W��Z�����%�fRV���9��V�f%�}���Ý�MI�0GP�t�J���aI瘮��m��J��+E,Vd�/�r(Um�DҜs�Qv�s����&L���*p�|�
[�jm��9���wtUUh�ߦ�[:������zgʪ��o���E6��s|B���r专�R�y�Q������M�;�(F�W6�w�i_|��� n��f/�,���B���&Y
�}L�H;�ƌ���v�V��"���.��G��o�L�*$H%��]�P7)������J���4�%#� Bat�g"ڧ�;P�3�$��'���_���l"Q���44�v ��ݾ��o{���.��rX�4���_^_G�]w���34a\��^�'����?�����ČG����g����̥qݱ��B���̕j=i����[BC~�u͘q�W��;�8�y�t�|����{����k��ҥ���w��a����;���g��i�r�j�Z�>c�{oY����u����-4������P�L>lj�ܜԩ�_-��n�L�^��/8ߦL�T�����n%�~�͆d-Kel��^��^���1@S�����\k#&�l?��O�/x�oR����ы�Q�)iӇv�&;�H&c�s������Lp��( P.1>�`�w��OL�	���X3���{�񓟺P�v)�E�.�&1�M{!5���a*���E�A} (����J���??h�q�>�nD%��CH�������3n��F�S�r l`U��J(X	���Z�b$���7�#X�?J�����|��|�7����b]q��y���BG�&�\l5ǁ���������e>��H�ճ�/^�:[��'ͣ�"X�V,��Cfx��'�Xj�/�D�\G�	�'	�#����V��Y|�^B6oC��v޼��k_{�M��e�tնm�l+V,�%�?b��l�,����c'�x�}�s���ȍ�SA������/4 �۩�����}����Q��+��K�,�ו���
HY,&z�"@�8P'�W�d%����v�F�l^�W� �>��j�/0�3���[ns�U��w,�Z@���)��wн���)�����[֯��3|G#X��<�ǀ?7E�����}>��	�#�i�A) ���0(�} o�h�����6�( (%� ��J,�������}3YN#�5�w���Oh�.���_�}�dK9����U=|QT�O�-t>���4����VX/eֻ�y��m[69��!3���͵l.o��Xg�{j�*/'�z��?�h���j.��_��?
=�����3h,@*xN��f����J�1}�UJ}�}�f{����򧞰����iV�x��!���?��<{� 6����
C��_�����|�+�G#$=�]W\�<-ş����E��i�b�̵`�7�E�l�V�C�����_��o%)�`���i��Q�	�"�~l�[n���q�u�G���FZjD�#m�����?vFslɆX����G��\�5�wu.c�Ӵ@F ��W�(� ������d^o��G�G�W�.���_K�g���w�!����*Ҁ?��I�0N����D���O+��{���"�u��g�������÷���>�N�G9 ��Cq���g��H^c=#�����g}#�K�?�7�\�Ry�{�a��{�9�Dp��6�?ds�e�}�͞��x�G1��n��P
����9���M�r�8��T_�k���۲��-y�!{��-��zQ|fY�e�lgϠ���q'�j��z8ߗ��e�p��{�s����I�OU@z���	ƥ�H״-�F����"t ��5�q 	��f�NL-5�rů��*���B�i� ɢ�;��{�}�����K.�gD�yN��IS�ZV�,�}�9`�{�+���gV�Z�w~��c���9����p��O'1�D��{����h����5�s��� a��������s�T��5��;�cF��so9|��C���D(?�e8yk�>��p)#�1�ozӛ\������[xXq`��z%k���\���sө�elȖ.{̖=������i塢w��첁����؉'�f��y�z�,�,��f_3���4�����k�N�6Bg>o���]��c��T�h����6uY{�l��^��R�����l��-60h�ik�����y�?&�g?��kq��1� L�/~��&4ϸ�7���dS+$NL� ��9�|�T����88���� ��^롃q$�H�B�����1@?|4e�#�U�(���h	!m��8��m���?��'��GGçp��>����zVǩ���G5�YNz�/s����8��P GB�n lE}iޕ��#Q5�&c�H2��(tX�c��q�OE�R#�۽d��u�gl'5��u��CNH ~rB-L�o��?����������h*X�>�j��p�c@����f������8�k+�z��%��ښU+Bu�rj>7�֮�d�}CV���-o}�<m�<���d?���u!+ 큫����U\�3�����:<�䆯~���O�\�+��_dCfҝ6�_�IJن�v��'{�*@ʅ	_�0A6����*@,�0A�C[ToV6&�P�D���׼�����PWg�h��.\���V[�xbU��u�<1M�E��_�!��K������V���p�bR�$9���x'�h�h���sEg���
e�. �xʿ��}���.��r�_EH�Sf�d�i����u���h����^q�hȝ�P4}r}��a�vCͲu� ��m�\��5s��w|0�l�ga�`�C��/ Jڗ��%�A�p~����ۻ�CgL�I�'چuk�FQ�u��r�f+W��J5c��vۙg�k�{����k�-]��n���m�������T�s��q��?�c��Q�~۸a����;l޼S,�.���Ox�_b�k����m��V�u����l�	��#���&���|����	11�x �-�_����:�JQ�Y� �Z���(K0Q4\0@����<M�@��qBSi`������Y�ȝ�q���]}/��������D�ƅ�u��1�{�IJ������<��T�����d�ǚ�(A���c?.���j�����Bz1�-KNV�֔�Y���؃�����E����$vՂ �4�g�c���aܘ+�p� ��ĺO|���u��,p��"�/���l�#��_��N9�h�1�[�أ60��� |��@��u�u{�uvM�_�q�wM�����ƛlŊUu�����p��3�������o���>Գ�毥v�s�t �Z�V�z�~������n�T�֭_i�}=I�D��-ڪ�i�m�/�`'�r���M6�wh�C>�4z�^ >��?�&'�mTB�LR0L��E�z���d����q8����Z��Z����+�tx>�Ef2���P�lFۇ�G�W)�v`?ҳ ��>�J5ǆ��y���P|�`��)���� 4�틠m)�E�)	7Y��W��9�k�B��6�Iܞ����z�XP�^��i�~��n��KV��^�*[�x��k�c_@���o�i�J��;o���8�>x��Z�<�zz�0 e�=���Ga�v�����~β�N����o�b�r�	Qy}Y����?_ڬCg�'?�1+�,m%��o�h���ݶy�:��� S-c=�A[�j���Y۸��iej��ѫ�O�����L� q��lp���7;��������ϙ��)�ub�w��A|���3�n�k9RZb+��H�w,_zH1�#l�/>#�p|�a��d
)������s�|�|4�ǳ���c�Ɖ^��k�ɇ}�u@���k�|��������5����N��`lEi�]�u�N��'�G��6y�Tۺ�ە�U+V���	l��������w����1k������i�{���}�v�
+��i�N�mg^��v��m��m��ګ_�jN4    IDAT�z��=����N����F��w^�.����)ޜ�"
ɹ���8��e[���L��4g�� J:�xB�	x���?BVj>��Ku�#�>�x�!�G�/*N91����N���������=�C�8�g�b�;��{�#f�Y�kV�p �8���oK�\a����M������ezh���k��j�=����G��V��τN;h��v��U�Cֳc�mߺ��wo�Ri����%ˤ��/tÆͶb�FK�&�;�����~��1�h�$[a
����O,�,e������׻U��H��J�#�x\��}�
b���8rM� I��~��	��磈'ێ�!
��V|SK��n�������ڱ�{L����C�N��X���O�Mq�*CQX(~�;{�R����l˦��ݽ������}#,c]�{G�=��%ֳ��.���6k�l�T�v�O~j?��-����)��%cx�:|���QU�t-ms�εw�������[��=��a+�l�L�f���@����c�©6�9�8@������$ƟJ���DD�"5֮_��f��0��deӡ��H����?�m=~�31�p��V�+ �Xxj�  T(Q�s׭�����G�3!���c�1�X��V�]��ʏ}���O}ʁ���\'J��N�qQ���8�@	�_�q�h�V-�e˞t-ʇ��\�_���`�N:�t�{�)��uX���]��=� \j% �8�VU=�VO6D�,���)S�S����V��k�����k˗=�WS�5a��z�iv�9���鳼�@Ov%�J���D�/Z	�-���� ��N�V����J-s���7�5d�9�q��X�l�+�EV �1�OTq(t��1M�HłA����9���,h��<�x �XޓwW4�"|ؓ���<��x�c#G0>u{� }@��˟gR4?��=^t��T��Ѐ=��v����+�[�J^HH�<a��v�ة���5���<��gw�ү����s`W�lQ�_]��JE��5�bG�������Yg�n�Ҡ�je*؎�[��[��'|�t�T�e;�X���y�ų�0�lU�'��/�ω'���]D�ȩ�yh0,.�>o�1���h�fe�h���]���3kmK����=���TB��b�e��T�#�u���Z!����eK��iU��ݳ����Z�]�I8�	�&��g�P��������,E��	=����ՙ��ނu��ڵ���c��>X3gf�"��t�._f����~ *��Ƚ�g��o��Uw���(�J}��|_����/8ߛ,PB�hRJ�ԩVC��޾�����=U�/����W_�@�ǂ���+}�X����_yHQ
,���ĉ.��9�� �������0�S�-�]�z�gvS���P�b�W�H��0�U-�N۱�k�$B�<���z��р|�cT�	P�ު�p����+��Q��`�<��Hй��P�^������_w�[t,+��~����o�B��G}ܾ���Y���^5�\�~?�����
݅KGN�ҿ1��o�P+�F�&L�I}��W;mCyg>��eaB�l޼ս�j������1hj�v���A$;�ݮ����¦�|���f�����u��E/��pdƺ)Z� r�YH�m���RI�K~��a3C�ocl��Iy�V4��s�єw`̈��Z�ot�kG��hL�	5T�ߎ���l�ќo*9��7~/@�3�UnC�[��O�c��*˺1���F�&�4@�������Y:������<P"�s��@V*�uMԏ*�����^U�U����Ο��:"��G��t\��ڱ`b/S��w��l ��_Ia��vK�N^ټ���!�ε��&{73U�,�"���3"���==Ng��O�������3�?�{U�er�w ��9�|SQv�֊ ��kA�����z�^p�c��G�'�hB=�N \i��$���MD��JU�z�J�1h?�z���ΧV�C���0S%yQ�ᐩ�F��5K�P��| ��H���I-s6�j��o�AJ9��y�X9�v���PVl�Vr�	���v�h�}�{�kK�� 9�5*�9(*I���<�ϕ �2ʄf?�0�}�o��"⪣�KZ�?� ��GQ�\����C�k:�=y�s	�x���8Fu���
#�{���zdN��\=�����I'�uE��1.���}^��н3��gýR�`!��F�w;����߬\����!�������`;�Yw8�� R�l*d䖂êqQ�����'���� e`)���O~�K1P��k0���Ь�Z����uY������/��K<;��z���$�8r��w�'�2��1�uI��nu�������f;��X*!R��#�*!�ZD��9����ƒ{��۝��R�S_'I��:�\IJøގk�{��%PdQ�Y���M}�����E7V�˳���R*����7�(��8�X���r�����%y�w�q��ؒ�] ��v��|�a�8�9����&�KR���_ʹ`���Ă�n��(���;��2�j(՜��10��hh�����©q�aځ%1��W:�����& ,��iQG�k�$��(
M��.����n�4��q-� ����S�3Lnh�^L� %�<cA�CM��%%,Ne3rV	��B*Z�#-���H���i�����4��y󭷸�[%k%�)M��c���;���Jƀ��&�*�;�I<��6�~�r�&�����+n��F��I��=�w�y� �`Zq���)�����gkw�-��땠Z�$9�S���Ny �͟�J��/>88�'�h�=�H߫���Uq,悬b�Q��P'~R������:��4*�uKh'-i�T�d/�I���z�p��`�9t���c����[�a����:|��)�<�n�jA�G�
�t��b4�J�ĭ�r�w&NG/��D�o��w�Q�4p�	��4B)8~B�`�?=}��\RW��O���P�v��1�ƢVm�F�_�E
��@ʂ�7l,0�	��ӤƋ�Ն�����8|���t�Q?5~D[�n���$� -���/�_�\��o�y�V�֧�㿧�6�S\��)�d,��1��3>�C��D���1�ז����+�Hc0�wP䞔Q<�p#t>�񏏘������j�!���ZA$��t�M'�%����.��{/&��?��S4vj��9�ƨ~��0��̹j%r �p��TI���F팉Ŝ��o,s���v�]�a3�q��D#�����y�E���c�G�̹^��_���GE� mC�&	o��%���9|o��mN��;�GμUO�}|���ռ�, 61�<
�y�ERu�&}�1	�?Pn�~ 5�6�Nh !�^c���7���X0�bJ�k��%81VXI��sٝ���c��Z��<vXJ��6�ؖ���5��s-���}ޑ�Wt��>��{����M=���s	����#���[*%��L><Y�h�`����j�P�8(��c�lοE��k����HӚ��L#�j��PfA� �Cㅴεهs�h8��f���3�T�.�A6h�Ī��x�K_��_o��ݛ|���}ڙ�.���K(�H��_�����YG��ӈ7'�}�[�����Z�%�j����p��&��r��`����(��7�_�`ų���ʺֆ\H��Y��]Ig�� σ��:�hr�]�!a˽dep�7��u�[k�v�DϠL�՜�=���/���Z�7���/ņ[�ַ�o�(�MhY�g\v��۽����u|/�E ��Ou���]4
3)ij(q����^�B8y��� �]���B�'��F�g}�}�$�V��6(��������J9h"����kv.�E�*b3O� � Z���j*���U��lp	��h���z�����k�'�3s}@�{�N��h
�-	gv�Ӝ��J�½�������v��L�,��rSI��	-z�	��d�k�	,�m�=�>����
��y�K-�f��ˢE�p����ޚcͫ�|���3��:�_|�cu
E���<�p}���{�ܘ�z�K]KN/�����|
l5�;�m�Gćs��#k(���k� 5�w���5ͳ�}�� �@D�����}���,��U��4r����a�N�c�}��Ĺl	�f���]g�aV��%���ש� Z�j�qԹ,�봇4�X��$���ڔ�`k3K[��N	��G�^���":���7��ɤsP;�m�X̭>��X>ZԊr�i�+C�N��X�m�ϭ1ֳ�����Ƈ�cݐ�G�a�k���W�q>
oe^Y7$���_ �O�'��ց�ќ���F{���H�VS:᮫� �(d�1�K���G���{�ð��OJ�H�5d�"n߮��j�����5(�_ᥚ{Y$z.�����)+V�\:��[�:��0aP�p��q�R���bZi����Z�UfN���ŋ��5�I��z\��n8\(�Z�f3!<m?PA�
�d�<p1o�9d�2�����[2��P|���^��/ ���r���AlA��'`�l�*D��e��iNc`޳��c�T>��9d:k|��~��e����{�U�k:�~K�.��2������C���x:LUX��|��zA�v�/���g�9����E��e#ϥ������+�|߯��u�^X�-���W8�j!J��s�,)*��%�yX#t��3d�Ha�<�Zk�fَP�'��Tj�vM?X��/���l` 亠t��������fQ'�_�iH��gsA{��ET*A���	�삏/�dtuM���m�G�X��Y��5�"r$)����`���18�`k�O����o�������c˪����6
���v�?��ey0/ZC�B(���ؕ@˩����X��<�@D��Ɖ碥���|����xʊ�T8��=��كs�!��}+�_o-�.�ZPb�v�':_�[��["�CG������mw���g�a�C�JV�r�k�o�	C·"ɔ�r�c���OP:�Y�Dw��f�h,;�����eѢ�5��[��2�vH�pS*���<ҙH��#����zz��9��*k��2��7W�?G����i�P���c#$X���A9�c�kԲ��Z��z��3vJL_qSi����3n� V�\4�.n�'�I{$��a��r���D	<	t�ݓ�.}�.�5XG_�����+ϱ>{੓���[N�Ш=|����,���-T I�5�kX�D�L	����eB*�sR��E+A�č�[�#�	в���i5t�#�PX~ �O�?�"��-ʸ��Q
�|H|?�2�}*�O�4�'�@`��P�	��3�-4��#�wIݓ�u���{����I�ä��j����+��+_��L�4w8IY�h�ī��� E P�����P�Z�5H����t�Ӥ{���6w;�2Vڧ�{����힯����^f�45�9"����ii)7ɉx��7�R`�M��m6o�E�p} �� W��}^J�gQ�I4j�l�r���+�%A�t��(����^���{��QC�lҫ@'as׸��e�r{�q�^lq��aD�o��*�u��-<�,�o�%�޵�M�4��e�E�S�vJ���B�ּ�1��=���g̜����{�N^0<�=�Č�8a�k�z��k�>}�o.����pg"���r�
���d3�������S$'}�{�sm�c�S)��G13�Ac�yGF�D��]�����H�c�v�>���>#	����{����Ώ��;�M���T�t~�����Tkgo�"�ⵡȣ|�^AR�	?Q(�$�Y���a,c[n�3��ц+f�|�.�G�A��E����vy8���o�����w� ��h5�/zE��
��=Ĺ�o�g��	����,a���7��N�����3��a0��7�a}�\,��_����w�s�K֟�w����s`g�.���B��f�?���W��Ͽ���/�x|_�I�>�>��p#�-]�G}ԋ�!��X��$/!����!d�&�DkPן��4|�\���`m�FN�QP�u����p�÷Q���tO�c�v�����������d�b�1�lf=�z�{��^=�}��6����@��8�����J���k�j?Q���U��N�8-����9RO��:���^��:�SW(v�c�˾dL��ȇ�ͬX���	����n���d_��?��{�'��"�:�'|ods6y�A�y�6�ݸy�w�A��r��B#���m���5c�R��l޼y6�E^�&��o�f�
Ϛ���O:�4;��6g���2����#���7��<>���C���?����?���Ԑ4 ����E�&QO K��'5�ݱƺ�������C�'-p_ܿ�5�PX+hb�����x�����$�v�s4��2�&`"��}�)?��=V�����}/�Cs�s2Vʒvn��|
�#<�2�I(u��'��4y�Y?��T�z[�:�X�`1P�ΡW�%랂����~�m�C��W�%σ0�3��/���z��1����_�Z;���B����mt��rQ�4�����$�;\��Kig��8��3���[�F�$��Ϝ9�.y��v�)'Y�4h=;�ۃ������>!D��P�{�̙��9�γO<�r���o��v�Oux�I%J���ϸ��`��ٞHu�M7�BQ8� B`o�v��@��g�T�)vp>s���TH�Q����k��ۃ*2{�;�a'�=ޣ[{{lӆ5V跮���xJ�V���� �P7%���s���I���ȭ�
�쩕��uBI �	��s+�K|=���uS�����\P����~����Q�KKz(����g�A4��fO<�����_ن���EG�;����K_�J;�i�����3�����X�Ԟ|Mn5%�I�����=2gh�^���eo~����X�V����Gy �Х,mIĠÎ�ݶs�l�}�)�����d|�_p+�L�^ij�	��B@K 9�@	"\G�9ƪ9�������h����}������ڶ?%�N��J�^�nmw��|���:f|x^�8�qکf����{mӺ56�W0��)�x�\y��@瓊VLuج������X:�a�6o��v�=��ɤRR'��w�e�)���UI/|+�X�m�v����*��d[�s���N���?�K��m��'l��mǎm�ˇ���ض�������/p�'yq����5o ;�������G����f�?!��\Ʈ��]v�	�[�<d��M��a=�M�a#NU���P�6o�j�r�zz����y�{��o��>�
�BCIJ�FS�o���1�X�,�}�����4�i\��7C=�=�Cy��}"��Ya9��Z����[��P�m^�����[6U�t��QT~<�<4)��>ڮ��N�YGk��l�|�mܴվr�W폏>�+�N8ޅ�nr�%j���|�9�9���|��������+}��"��p��|�	�ʨ8�g}=�m���l˖��}�V+���O~�P�f����[�k��v���d�Ϛ�>GJ�C5������1��/�����U���#f٧?�I+ؤ�v����K_�+�ؚ�O�P1�Ϥ����o�W���!�������h�+W�ts�E�v�$oȞ�/QB����x!��(7I�g� P̡j(5���������)��=j
:P$k�}�{��u��V+Z�<`�6���m�,[��UܑN�r�g5�\��8�	�TƊ�)v�Q�ڄ�S,��t���7ڣ�?|4%v�ǘ��2�����g�����'?���wB�����>g���o��(~D"  �t�l���;��C��	9[�f�����~����mɓ+��s�-}r���%�_��I�z��-[���4�.92��`Ⴏw
ok�1�s�e������%۶}������i�t�֮{���{��e�����    IDAT�b�o�������csO8���	��/���o�' Iߑ��kV{$�LH�\�7�����G��J�ߛw���G@�}��Lo�P}6Γ�3��Ph�r;��ӬZ�L�d[֯���sT���x!!���:���9G[��If�[�q�]�MN��5�p��c3�PO%g�X[�k��N�o��o��ˇc��K5�T"�pN�İ[���_���v�I���i�l��%68je��R���\j��D�)XG���G>�e�=�._���ڨh$��f̜��3���7�oo��cY�l�a��UW}�2���Y��������ϰt�h+V>i��`����m���f�&K�'ز�[�O�+�����p�0���D�Ш�Xl��p-8@��r ���`e	s��8���z����N�V�K�z����1���Ͼ`ݣ��š�rѶ�_i;�n�|�h��̥�g=�W�x�������?�c�z�6a�:�_����ǖZ&��������/'� ]�^�erxN�{��]����T��}��\�(�|���=���7?��O?ΦM;Ȟ\����RC�\IY���Ǘ��J��ne�Q���������W��ei�z��
0�q�o���P��c���|�*������n��[���e��N��i�2����W�uk�8�j�v;�Գ|1�0�pH�R"���p�͋�uHn�{��_zM� ��Xi	q�X7����f�����5(�u�����1߯��S-�\�߲v���������<�����pNJ����MʩSژ�+�.;�����I9�a�6�{�I�>{����w)ɐDټ�U��K/y}=�����Ɗ'�+�6��|���n�Gp�Z��~����I'e3���_,FLeϜ��Wm����M�ի��f���_J���E��v�?s���,^����1hޅdls��9�=퓵��{���Gl�d��J���l��2��l����D��Sy��9`�W������ۼ�^��=1�E�VOU�X�Q���5k��0��;��]w��G�@ H�h�1~�����2�u����kd��x&�M[�0k^e���f���_.Yy��6�[e��[-�*:���s�?r��-D�0\2m�s��	��t6���W��	���h5�8zF���ڹ��m��]ٓƯ��4���>X���Ϗ|�#^�{�f{�ޟ�ԩ6m�[�&��j�O����-yb��Kۺ��N9�l{�%o�l��Ճ[�n��>�4���E��,DԠA��Mo�y�βJy�V>��OD��MV*S�+0qZ���wز�k�З���>��?�~*�+�-�_ř ~������淿e+V�p�W�Iu}�Q$������ZV�B��~�8�$�U�V�+ئ묷��&�3��]��fB�$J?�Pޡ��Z13�fqdh&di���o�����%K<)ʅ_�#@�Q(�(�W�J�ñ?�[��Ź������bG�9m5��F���gj�fգֻs����PiЊ��z��T���A{b�S�}G�]~����G[�����.[t�b����w8���uj��L�,X�B��n,��90�9�ܳ��^�5��|�=����z�2��-���UB�g&�����)���'�EA��?��?{B��_u>N?�tC`Q@��G> I:J�V���D�rm�6>��`��M��@M���ζro��};mݺ5�ӽ���L(�P){�j)�����[��pJ�lαϵ�3�r�fk׬�k���_�[�t���bv�m��b��GV/����|x��.��"O�BK��Q��i��fW\q���u[G�h+�z���1��3��8M^x���6ڑGg��=զr�z������
�Й�f+���)��Ќ�'kNN �-o~��ܼi��rY{쑇��?�gO=�ܵ
�M�2ɘ�SO9�;�X�0�5��~����U�a��kQ��E/z�O>���'�}�l��yZr�&ܳrW�?���bT�=���-��sfϱt��e��n�s��8��R&�v�5ۤ�����̆�;x�t���ٯ}��v����Kg3^<n,���Rv�BV�s�ᇻ�O�{��6n��A������ܕ<W�pL)���~�I��mp�����>۰a��{P�3���Km�aG��I[:�����{��7%� ���?}��?? ��/X�`qw���f௸{�e�v�An��>���b�y�F۸q�k�8c �9�g۔��Z���Jռ�%}�"����,t9�X8,~QM��n�A	 -�����Q���C�G`�G@>	��؇h��K�������i���JRO�`;��7�{�dC� ��syotB��2Q.y,�P^Y �[��f/��#�K}�TЯ�kO��
@�Wƾ�J���[.���'٤�]6��ok֭��[6Y�@�G;utu�o����������sg��46l�d]��R�|���h�\CA&�:�d�⬁�g�,jF�Y���-W�w�������ކ��rI�Z�B�������� �-��1�ݻǘ3~�d�� �>�F8�N�T��x~��E���?OS~� ���b3�\����/��k륤�m��nr�q��#y@�=��I�1��:�����_o(٠�`a�D!,:)�X�0V8f����^!����S�W��6�Z�����Qb�4y�$��N=��<�v&v��8�H�K9�t���v�]��D-R�	��#mGf��'���\n��Vw��!��}����kk����
�=K���c���n��ִ�Ls]V��U-nըf.O�2��}��| ��<��$d�f|o��q�!��)��B�k���.�GA��=��c}c��@_g�	�N������>˻{�96i�D�˱��W�xwa�=��?�w�����������颜�E��¥M����E��rJ=`�Qga@�I'�d�6+D��.e�n�:{rٓ�uTke?��^����|���������Iǜ�$���/}�^�{�g�������Ox�F�9�:�Gh݇it�x6g>��TÊgv�(�\:X��%}�^a�����pކ���z�*�M��aһ���b�Ja�h�T椌QK�ݶ���H��[n���<x(�SԮe��1Ӟw�q�QC���ֺ����I��� ��Z2��g����i��l���-�wh�B�K,��*�)$ӏl���W�&Y�.���+�K�I}�At!�$�aʱxT/����Z�*?�7���l���z��T���(?�o�G���V�F:sU)��M��Ϯ�<�(����@��Thv��tٓ���t���l�T�Mq�q����.��K�ѽ���5�y�G��H>�},���>V�s�\.o�	���A�� 4h3h����i�jq����=P��Z:|ہԮK��z�g6U�V�d�0� h�w�����/�ܣ}p�7 �_i�m��6����ydA�:_�$��03�}g��3�v���iQw��=I�zvvҌCᇲ�d;�c��c͓�"q"���n~������s�]H ����[�s��J�(t����9��\�<��Q�~���Iڵ��8nMg��Ww�ۃ P���H����8�"N<k��W�pfL��������t�v+��N�'�^h�� ��&�|�6�I�Rr����gqxƐ���
�5{�Z� ���\(t_Ҍ�i�hw�4�H�HׂD�F8�QC&#�i�${�(Xh�p��?�� Q�8mt9��=��,�F�R`���H��I{�������ꫪY9�Te3N}%�qR��"����ZXm ��3�;�Y�A�|b*�N4�D(Ś����8b%^+í��÷��0�`�?���`j�T�H��r+�|>�A3ޟ���1���F��q���u�b�|��i�E���@0r�E�m$�4�a]�8Gxb�oT6C�]��� ���[
݅�5�Ȭ�al0����ݵ�P�C��&l܀lB�b��y� H�ูs��_����G� ��|����ځ7k'��c�s4�����"��H���6����|�p�5J���F4��Q	u��Fo��s.s&
A׌��Aɛ	��g���]@0))�b ` 2����
�9K~�z�9=����]�曗@������/З(��I�S�%
�5��`sW���� ܓ�I�fb	Z=�����@���v�q�Ջ�)��y���k��U[�8�!�����hB� ��ڰ�$4^��a��*��:̀?~�x�Ŗ � ����b���;��š�qmX����M.����7��4���f�Цiw��o�}sd��j�Q������
i�~�H#��$:�g?��Gy��G�^"�D�i�wը?잼a;���w���e/�g!_I��Hӗ��"�#����<)%Nt�~��H���zaTJ��y�4�yXL�7n��S)XJ�ЇW�SFN-�^EK�okĺ�?�,�?��<h)��g�����������w A�5�@2v�{�����o���/�0��X��'�ä�$d��7"rX�h�Тb��Do5�rI�m#!�nc����O�n�d~�k��'y�]v��#�S����6��V~g�5�׽��노诊3��)ϭ�h�Q	�=��9</�Bx
��1S?��K.q ��C�(nY<�֦�T�?�C���~�v�d����� �IɆ䨘�ј��\���`l�I�fi��.�b�^`� Ƣpȕ�В5m�����beLc������0eLe0�g��Ɋњt��,��c�. | �u���8�9o�[���mh�с�������<�MT&�DX�p�C�x���x�Bk�)�����8�+�h�l��*i�!��NDD&�z�}����uɌ���{�J���ҾΫ��"(ش*�G�Y1���ַz��O��]�W`�����2�5XK��r������}�c@V)���F��H0��#Ǣ4} ��������=w�W�����Dah/����� �m;��Ԧ������O��ݿ�m�C��<�( ͵�K��i`}�=��z���X��t`�f�i$�W)_	�0t)��`ķ���8��bǵs����G��kk��%��1	!�D��eq�~� �`���h	���e4�M8���&�o|�;��m5L��Ip�o��q��(�y��۳�c�����$+�ͩ�
�CV�Ýު��/j.Q�Ma�d�V8����g+A�O������$�(,Z
�9Gq墴(6ȹ|�(�z�?���τE�j�b��-�,}�CH'�a�/8�����]�v��X�$�R�4��ź��[5�J2�+��#h_+Z,�V1��E�P�%��1pBkС=�C�sW�u'n�^
�<��$�HB���{��>M�R���Q�X�������^�W,�i����6|aW*aMS-����r�4�7���A,�4��c�\s�5u��V-$�<�?��@S���Vϱ��٘�?�,�GqB�G�d��%4��[h�1u�9n��G�ٷ�v�����_����Ų t�	�(�9�:�/�_>Ɓ�~��փ�����pD����빗Ʈ�4���@K��%��"��=�&9!�z�g���0Q���[o[;	����FzW������*9���`Q��^ba*�w�Iiq�I��	��  ��
H�s�o8����U��g��[-�z�q�V^�_�G1!Lrp&��X,{�	���PC��s��`��g��!�h��ڀ7�i;N]����5r˼����'��x�R��OPS����$υ���UO9���M�vϾ���%�{wzI]4���6&sR.���&��8i�Gċ4�Gy�#4H�{����2̳��4ƌ=��C��/}���������;�0w6�p�����w(,E��x��~|��O���1�� bE��p8�'��P@x'~g=b!���3���|���e;�Ph���)�(;�	�q$�F�_L�2�ڇ��~��J��E�J�c�j�;�9�5�����go����6���˓!\�s"Z����!<�����۔t&Ҋ�r�'"FJ�PցZ>C�%Ky"FH� ���&�����L�R�Y4L;͢FHk�f�x�21�)���SO�%�i���������/: �>�E�
`����6I�wؗߏ�1���	E�0?�6m�wN�]xw
�Q�	�j ��Z][��\@IQG
���s����������w��T<�a�5G=V���U�6�d<��z?E��"��(�����d��iR���Md��L�X 9���=���Xʖnų�7�F�  �<Y�R��(Q��bv}�Iu�l�f�:��BL���'����o�g�e�j5/���nj|@��k.�vO��&-.��Ҩj� ɏ�3�K1�9&d�i;�?�6W� k�5��/X
C#BD=V�XQ)--J�G~i.֕�;@qJh���Q@��&����m���x��Jh|d%p<�+�z#��kd�����w�6w��	�JCܟ�'���?��d]�����|�󰁪0K�ħA�1Q��X�_@��KE1�5[�����+SV�q�s�����$�+P��8���z&t�_U69�DU�a�Y��,+1�z6����`A��C(���<�1Yj��O��u��'�d�7���}VhKz����P�֮]��@��t��%���'�����5��o
=�5���i	�_u���PaS)��c�����;;;|a �;�&�@ ��O}�S����|w���b�V%�BT�P�0єp��PBVB+�'II���Ɛ��p*�P���'@�;�/Ĵ�H���Q��9�Je�����@,����yVE^�&y6Y~Ҋc�E`]�I4W��8=UW�x����@�gx뾚�v�'ZNjY�. �!�MTǒ3��;�·R�>����{��)Q]�J�:���	?D{��V,���yq�c˹����c�'�k^=�GN=h�K�^��z>�jmE��AQ!/��$�9�Ƹ؆�@�?p{�.\��B����?]S���>�>t�,��9ȗJ�t*�<hK��o����cB1�f�~�kV,g-�MIF/�a����;�vXDT�r�Lf���|:�쳝n�)�8	�j����P)8Y耇��:�
�m�}�}+���%s�<� R�x%�(>����Gs]=�"������tc���6lp��:{�E+��*���=���q'�^�0)p�gfM���;�Qk�[`C�a�H���`1T��o�����$��������;�$K
��X��O�AEO|K��z�~����y�B�}	ʕ�=���x��9a�u��N���s����~��۶�p��k���7
=�l��Z�ڏ9�h���WY��édS�`۶l�%K���֯[W�+���	�og�=Ϟs�qf�഑FF	g&P ?^��� ��b�U&??L_��|��\�S%P��]W��fϱ*���<�Ѱ1���}wa�h��� پ8���Kt�������AQ�SY2�c-V���~��� �.�v7cރ�NxQ]{��㋢Ě�'A���)�/F��ͧ?��\P��}R�.�)'i;�G�]T�:��3�K�����T�Q�W��(�/�fmA�~������;v�w�̛7�#���k/��^z���O^lV�X&]�'�\b�V���Զwo��`����{��v�igء�fCŲA��w�u���e���.���Pxw3�VC�c�:ʮ|߻�R�l�҂%[�~����{<�'�	�#^,��P���*6�������rV�~�eJ��� Ŏ?�|(�a���.�Q���h�8�����Ƅ;��,�����Ak��׿�NQ�nc��o��h�_c�@��;�ck�x�V�_�-�-V������>h�$�)}op�Ҁ�����:'%p@\8��'�Ē��西�ۿUVk���4x9dꣵ�e��4*ψ����x�b����ݲ�#��+�^�w�(B����A䟀�j��Wi s��W;ː��l������ۭT���N�J�N����vX��������3gz�2�/}�Z�0��8�7�\�](�yS�'ڬ�=�������:�+���G�\�f[6��m۶��Ѐ���&��d�;z�ڂd    IDAT��3`���]����ɇ�����!M�@&��w��Zil���\��_���9�D�Q�5
�=tl� #4�$q���}Ќ�Iʂ�F�_ ���}����[�h7���z?�񖦪��
9m�c�pH8�.ມ}�M�7�_�'
��E�ٗ���z�s;p��g��1s�L����.�3}b_M;k�s��wQ/�۟�2�4j|"������]���wgw�}�7jU*�? �/�B(�.������3U+�6ԷնlXc+V.��[^�D��l6o����y�����\iO��x?�������:���]��bw���f�_K��G�9�>�����@�M����n��.��� ֮Ya۷o�\��:�]�u�[�n�Y���o��N8Ů��
7�]�Z _� my�ƍ��H�yի^� �{*zB��g����*}��z�ȗ�ǚd��T_ ��
�����w6 �Ɔ��;���X�o��}H����w�+�BY�� T�h��rG]+����D�z�Nq��G?�dAU�P�E��u��FT�	�ڇ��Z��������o�AH�r=�&��g��%�g̘�5���|ͺ#T�dAA��X8c)��	��ՙ�O-�AC#�3FPP#3���07�&NX4&�q����d"b"Q.	J�F�^�`��@7�s1�xM��#q�Q�iA��޻����WOq(��k�jY���t�W_���<��>�rP�x�Y��M�Jc�����׭5~�ayy�ik��wW�o�˫͇��7�1�w�W�A���u�Ŏ-M(�i��H���<d��u�d���_�5eʯb��݂?�燆�������M7�p�|���<������Gc�MC�G��9f7L4Ti6|LPg�Ix�f����QGO�- ?�E����8Ё�<�P54 {��G��ի�Xx��J��^fF
�;�?��?}�o���Z~����[���Y�%��:�d�fu䘳>p���� T�8w�~0J.@�9h"�S���"X�6�M�EO�%
ȋ�"@1q���yꩧl �@u��$��3 ��/�Iu<=�("��RC����0�a'ث.��0����7W��>5f}çf�A�������~����ֽo�����bQ[�ߚ:��-��K��<�Lq���/2ш1�]e�������cL<�l>��cӴe�Ow�+LӖ6��ǟ����yo�f3��/��.���0l*�@J����ۇKI:"`y��[-=|�p3c������8���,m�S���R�A�C�台�.����JM7�dG���k]�G����g&���M�TI!�"�'��-�.�5� _un��<
q�|�X�d���Y� �|����_wQ>�f+�y�ր{��,��^ u��M56����9r�5 �V���QG�6���}�|P�.�$a�zM�ii��-M���%n~>w����kk���^�j���g[�IS&��m�$�����u�Af楗������d=�����<�$����47��`h(j�������ΐ���Ō8� ��N��\s�]t4�ܹs-/�;L�>�Eê��&��c�)�:@P����\௳ v�
�l�����MK��ϢH*��1��m%�FA�����V����hH��	2�~�Q�Z]Z��a�����~��t���C�˳᧒8�X��2y�9�G���;{Z�s4�C��|��]��3G�=���>f�wM{'����6�xȼ������N�HF̜��7Ѳ*Ӵ��zZ�Ye�?��UԖ��)S��/��P���G�0�~t�ikm6}*#�ŏ��i���f��LssS�(��ټ��ԯ�Ĵ�yf]}�w�?��*�}p�(��h��1cl��,����F�0dlD5�Rj�
Tz�i�/ �2�0Ȳ
��eec�0d|�,l
�y���}7�ߵ����Oh��;��Ϻ�R1�}�]̅hy�<X�Z��]@6S�Em�C`��N��@_���&�y�1��c�W��۾� ����Ƽ��-�67��_z�x�P3`@�z�*�mNUl�������۫L$��l�3�c�8�_L�>5�ݕ������?>h��/Z�����s�zZΟl�2���!f�W�f�;oϴ����+�j'�j~Sf������6��Έ9���e��T�e~'�kN�'5��xW�/]��*e(��\bU"��r��)p.���
��B�jN=�T�{饗� ����L�w�cU�?�%��^��N�F���_)��.\h���gk���m�R5�Kɳu��s���=7���+��Wz-s��o��k;v��������%ւR�<���iv��u��0��m:y[{��:&u6���'����]mZ[�滧�iFr����k���^��C�t�a�Ǉ|Amm�}E���LY�5����������ϛ��C�d�;[�����7�3ﾻ�������ܞ����io��ƦN3쀃�q�Oܦ/��Y��<��ݨT2rF���*
c��	E--�=��rnfDO�?�������W���(��{l�Z��(�02
�10 #
��5R�]�$'I����V ��G�=���v?`��;Nl���nO�
	��||,g/�g���b��b?ślX��Gٲ�Q�jAk
2���V�����u+͇~`�;�MUE�54�imQ��xɈY���f���jL��l�����y����r����Wjݱ�/Z�h�=���'?�;3�Ӷ��:�/�O7t�����g>��`ֽ�����?���z��N�
E��Qc̸/kF|�M�b��T����c�*Iכ�'k%�e �/!S��Z�͛2�}��kv����g`������m����ݢ�l��a�_Q�����R��B�?�F~?Z.�>���2(���X��(Y�
����qXQo��,�G��œ��>���Q����I��)�FԨj3x�D���7&�n�Z���_�����^5��wXs��:ZU��|��c��8ҔU��:���j���{MWW�Z���2h�E���w#�?�;=��O"x�3<�\p�~��6SQI5/�.v���&[�a��>��4π�M(L�0����8}6���S�G)�Hq#�p�|�@_���������y���!�s��P�}uV��J�T���ϗk����@���J�
HRTUc^�o	��S��8ܞ��M��U6�/�`S�|jW@}��/��v����Z,0�o2�ԟ����~ �?cٝW�-�L�K��U� P*R�M`�ޢ�T$�B55�S���Y�<� ˥I�$ݓ�l�w�3��N22��0~"}er��*󅹄��ء�m�Y�V�N���$9=�Z!�x��}��+�@�t��d��P晲s�ռ��u��4�4���I���|����oжй7�p�Ut�r�<yW�T�Ϝ��Czx�J:��x|���wW���B!�|�!>������U���o[ϊq�zy��4x��ŋ�Ut�����EA�Sy����T��iXm~��L�l(����k�͙��A8�� nZҲxO?���JQlmb��ֳ��ci۾(�d� o] +��o�l�w�y�n82����¸d�Ӧ�	 �߷��4�8Nm>�	��N�� �%����Lj��	��1Gw��{��ލ��� ��\�YʖM+�W��������)���.��gP(l�p�m�ؼiQ��ś3^��s�̖R��e� �|�?���i�(i�.G
�"< [�3�Ea�1�ָ [���@V�1'F�t�_����A��}��-��J�=�5/R��Q�F�8cE��9��T�=k��>�2{Q���x����I��}��r�`/
��!7_2�Z�Ƚ�KH'�I	�=��y�P��u��9)e>�{)л��@3n�eW���d{y^29dА鵵�w�O�2��Xl�iYi���^r�%i�P���2�u��p�b&GY�dA�B#+��E>���m M�g!N���D�p_���{�9��]ֆ�g����V��:�'VY���o��;����,O&���%o�k��l[��WXA����[o5����=�@�a	o��
�@���)�٤,X'Z:c�1mf��OA-Oϥ6���U�/`�����R����n�=2!0���f������<�J����?� �?�ܒ��u?���+��s<2���;��sm!# i��3�5���� BN~5�����IgO������H����)����d�k�0�k���y�f���4L�N�b-�Ħlz~�Y޶�8�:s�J�3g���@>���yF}�����K?��/�j`
Ɣ��xd���<�U��~;>�	�i��HnZ�<d����u�.>�8��b����2�m(ֵ�N�,~iu*��,"`ON?�}�m,hr�9T�ŕe�=%�,�[\"�c��h6n1�Bl*�q��������m2��ҳO�4�o斲�mO��
�;u
����S�>m��WUT����y��l&)-�k���x��h���r�=�	�]*�g����q����7�^��\��Qq��ѥ�v�`�x��z�H�\����SbN @��w_R�Re�} 2d�,�=�.�(�~���chqrޙg��>7Z�>K\�b�-�1�Ϥ�d���[6����c2��s�O��g��{}{�F)ɪ�QCCq*#@ԩ�J~b����w�� pƃGKJ7��Fź�]�}������C�e
Ƙ3)>�xP d��ٯ(�[/Y���d�Ew�O��(��N6�P��&�_ZWՋ�����4��>�$��92a ���
S�xJ���j�An�� (
E�k�IG�*j�T	cM ���u���J�rS0ڂN"nA�GQ����d|x"<'9�|�R۸�@UHV��R�6������*�Y��&��
�G�bL��8����]�Ck!��뤸v%��'�LjL�����di�&s�����҆��|����7�W<+� ���E7OR}�1�wJpd� �6m���3-��d	���'�p���/Y�ʣWF�֒�g�jf(�M��?8��,���3�z�V�T�2�}O��`��KT{�q�x�������^a_��`�^c�6U��Ŀ�E�fƈh_�oK��simm����)S�b��og�d�Xx-� �u�]Nյ�e�sf�YH�G��ʱT����D\�xg�ϱ�\���?��u��a{k��`|?���|��M���?�����pc��bG/rL���	@]�������������B���y�~ �>�:[�L���}{��~}}�H
R���񂠜Di���������"�2t�;�ȋ���Yw����nv����3�N��q���F@F�*��z(}_YW�||�Z��|?^�&t�,X))�����:�w��7X�^s�g��W�j�	䛗xz�${�1��Dɸq %> ��)) "�^Jo������/E��3�%Ydb�0�k֬�^s X�c.�,���7M5)�[ލp@^�"�H{^�\�EJ�>��-�������ű��)��_���@�)��N.g,�ׂi)3A��I�
�[�wJ�k�
tt��o}%ҁ%��r�c9� �Ud,���J�g��R XԎ��x|��tM�����/ZŢ͐���O���>���
��e�5�@���f���l�o���<3|�a�2���gPX��Z�?�Q��8k���ڂ�9����z�QGٸ��5�*��}tϋ҆:ԚBy�(AY��R�2p�K � |�M��K<��ISK����r�
�?�D�7�H�~�<���=��+�����9k��e}\�'��ε��KE�6��c��갺y�|])��xc�l<�ﴷ��(�[�F:��N����b���g~?����Am?s���a�R4�.nHaK!
oDm2���d e�=�Sy�:s�E�*>�2��X�qj6�( ��L����ܝ8�dIZ,�A��U�h)��7�{��J��od�5�CX ���{ �@��թB.m�*�Y?�ļ���nu8d�w6��!!�6c�!��象� �x"����������,}ι��=����$_���e+�U��`3纲A�lN?�ck�[��c���UJ������������V��D� J�C �~D��PV�A�+D`��3Go�����!N|S�f��D��p�}Cn>�$0��(*�/Y�X��/Xʌ᪟α�*'����d��k��"� ���������s.M+c�k�RgϞ�ND`O�	�-ݚ��d^dy���Y9��h<cP���衇ڸ�G���R%�̢.?�Y���\cEϡl#)���Z���amm�m%�O�����d�?�kd �X��d[ @���� ��ȹ��z:��H�:�`�m(��Q�6֩
L ��+Ț�Z6�F��~b���2b�� d_�m�@�����o�_)����Y	xc��I ������Y�� .:��� i��Rb�����X۠5b�?�я�gB�(
O)�xU�.2$\�����s�A@A2_o��Ft\����͂s<����{sv4��1��O ���� ��/À7��IW՜s��f���|�i^ޡ�͟k�H�C�"�,zf�����]��+Gm�0�JBI
�ˀ�U2��}��naݭ%����_�?V,��SD����
�m�`
�@�2��7����s�)w�7%%e��r�-�2"�!P�����L�����Oa�����?c����k���8�kg���O�1,�Q�F���41"����ǈ@�g��W2�I���\?�D�Ld��Vy�J]���|3>y��_��k�I]�O�N�VLbW���<��kkko):�<e�c�����h�]�0;���Y�JU�u8F\m7G�;�*�{e)�9e��9l�N2��;�;,�s@�Ԁ:Ԅ�����[+?�����9Wm���l��--�������Y��?��mV�G����W�})�".!�������H$}�D�'N�'�W���qO�X�7_�����}�`�h���В{����ߕG)�P�W4����7{��1�}�����̪[�h^с����o�&���O6�w�'PKJ��q�A����L�/ik��A�?�?����4���	 �^�������F��ˣ�>�\q���anPrk 7���	����s 	����K\5��B�?�r.�$�W@� .� �,(�ݦ8�b>�d�'{�TfёPrx-J��	�fƸ�3;�������\�����(�Cr,��Y`C�� ��|Emm��%���h,#,������
*+�$|�ff�*���m"~�}6ΟTO����(`� �7�'=��C���( ���PN��p}��e��{���x��,��Iٜ�����?�NcA2�|i��Q`�!��CB�3$艵��@�9c ނ|)��A�}��'�M�m(EdIVv�\��v�.���)��w.�_��x�����(h+�'S��d���Ʒ�ͮ[TwS�P��g��ם���5bQ��[���& ˆ<���m��
oد���dc 초����-��!(�!Ç��j��T;2������g�W|�8X�>A�6�_�	�����	Z�fX��z
w&�KcA�'���R�$�
���^
��"�f��W�&�C��^�_5��,�w7#&׶앩���Q�x��񳁿��w����*~W��(�ނ����S&�6�b�?�>�( ��<k,,�P�Kr	�6�r�*/I%�|h@��*<�N�Y4�8)u�M��1��M)\+�%��_�J������@�o	�}P͕��Z��1!�MX���?��r}֚���Ɂ�'�/y�Q�ɋ葇ӅK�c�C�4oi��#d�'�T�jŐK��ݲ�1n�I�t-�\��˂��*�E��mo�zO�[��?)��CO'qw��;�_�� �y��6���m�6�v���KdEʢ=��al����w��%ݓ� R���,.�
K���'e����w�%�{˟N<�B�?�?���rD$�Z6`���`i�    IDAT\j�'���@J������@ܢC��1��P.j{�ߩ ���s�1��d\1 ��y�.��<���������ɤx��D9�j�He��.R�ʣ���Ӥ��Naw��z"�-j���w�9��������:X�8�^X�p��9V/	�@��ķ�M��|�K/1���;����{��M/��\�2>�_U��L����](	��9�\h���� ���-rÒ�(K=d ���v��W^wwy�=ɔ���{s����3�.�e���R��t% ����yE:F$��y���/���x��������Yg���/�˳�7z�@^:�2���q�SEn�<�WM�,�'�|�ƕtɹ
����E�6��M�8hGɂ����ރ�Ҹ�]�]�y:�2��E�a���)Si�5��
�_@Z՗�'mjDux�(�Bȱ�iŠ�Mq��բ@-�y^ �9�?�n @W]lF5�S/��x�0��òǺc,�r+���/@�kh� �����k��w�A�(z������]EQ��/pI�d�駯yU]�LGb.s�*	? �,B㩫+S��52R
�x�z�W��ǖ&t[0p=�} i��B�P(�G� �T�r����}������9�w�F��Y�ъ�zRT�5j�o�(V�+<���0��������ŗ�?iꔇb����S�?̓��`�=A���b8u�+��T� -B(���-��O��=��-<?����<��s����K��d�;�?@��/}Ɏ�!��q�3�=\P��ML�7���;�$�K��d{�m�l3CRV?���~�^
@�� ��?�{���ώ�K�S�bs.P�okB�/T~r�F��5u���]d/�~��;�3�?��24ħ�� �mj��R.R&:�:�X{C�=�<��C:]L��n :��>�߿�GO=�D�w�<e��i�5�!��)��V:�
P#����\RH���XHV���Xx+V�H��U.����	����`s2ר���sp�ƹV�I�5���a�A?���h�"[�K��P��#&o;�KV��)���y��S#�<��؊����c�  (�����l�[)��v�gw����u+b}�I����#�ܐMƩy��� pU��|'ʜ@$4�:X� ��c� �(2��3BYI�!P=('��w����'�H�v,͚�{f���O8�������ŏ_?��S���5�Â��v-��@3�� K)�XH_��K��B��*vt�M��f`#�7���j�q�]�p �i)�����e~^�� Y]�8��a�Gi�P3:>�s��w[AwG��T�BQ���Z���P�� �m%�_�M���m1^x�U��T��ۄK�/V�w���a�J�����j�u��\�C����:~�Oz����O�|�^ �뮻μ����j��?��F���;ڲ��i�9�5�a�o�
���{�N�U����S���"�V9D�v���1"`|]��;����g^�0����|�]����O�')�vO��Y���*�d#�	A�{6  Ϧ@�-�ʝW{�̞��VIc.h"��s�Il:�uF0o���ҍ�Ld|6^p�9���`vu���#��5bx'��k�eA��I!�݄�/��T��\p�����r� P���S
�>�\|�V�*O9h� ����i���h g.�I�k�	�gm����?�Mx�4�|��Nu�d�-|��U�(/Q�Ɍb���.����j�����l=����x�s��a>�У�)B�r[cc�=�~XX�x(����mm����aWf�,���7��T<�VV�{������8�b���ӛU�� ���X��lB62uӗꇱ1F�1��6�!���(*p��#�1�?���R��ݼ��<��)N�˟��g�.���,D�e<sQ�r��$)�C�s���{�N�H .OS�G� �oϝG�U���2��N[)-Q4���߅|�{d\j�#ߜ ����I���]9�U.�x�u���u���o\��-���L�n��ƫ�T�OgJD�v#!�X�X�:��M�S>����tK7��0!��'���@�?�B}�y��C۸��5�Rg�jL��;����+} �j����Ac�Z�j�Z�|k8���-�K��6P1�?����0?�?��%�-M����8�Y2&o��e��d��1l|��	��t�WkKO(*�m�>�g�)��ؖ�Ke~rO�_^��+Y��TRyԒa�0�H���>���[����4�/N�k��������oO���'�3m~��!�m����K��4�":(�'V��$]�]s�VѲ�]�K�#��Apw�M��`���i� ��z��d��]#���Wq�֦n��.�W'11�dz�y��f,�yF2MHC$3��J|�Q�TO8��LJ�J�eZ�C�馛�x�����9Y��b1�7�с�2����x~h}WZv�er�g�X�(`e6�5�<gbܬ��;���^����w���a��3>,h�V�#{���O�~���z477x�7�y�O��7��Ͽ���^_������W���Now�Vs���Pv9V�<��5�  ��'A`0��O�P��݁��YY��=�!��( �� :�Qx(�8������K'�i��o(�e��pjn~
��W�=�%����g��y���`���yꮲ�>��������ᕒ�C\�s�Y���1�8Lf�ܹ�������J����&g��w�1�ͳ�<�[�w�ڢ��|�G|������l����=��]s�����ٰ�e���8d�����)k$},A>� �H��f\46Sa�t��`�ɂE�͘1���~hSr�� ]�E�qh�[Z2�0�^,h�rt=�B �����O�Q����k��?���y�I�ĲG��ƿ�� �W���Jnh��}d��k�i�X�6��mW�|D%�g�d˟uW�+��θ
����e7Ͻi�	�����9��˗G������۾� ��"���D覻;�+�(>�wQ�*+Y@'�7����lyv���H�� �A"*�`����)� ���;��������aEqo
��P��>H�$�"CF']1&�
�����߰�I���u�.�ÒgO�g.)�c�PH�A� J���w������$���o[o�އ�=�3c`Ȏ��x����.Yzaw���3��(��O�x����Y��P�]*�W��-vw�����С�d`(8���Im(�_�)$��͟6	��un��RN����c����= +�-���q= �L��Y�����KA�����Һ@ֿ{���f���8ԅ�o>�Y�FoZy�V�?��5'�S�H����'D�
�WZ�^$��?xg0g�l��T�2��ֶ�	��y��=[���5׌[��s�Ps�ҽ2b�Ӽk����_i�n_ײW���b�\|�S�gf]�gm<�,�Ϳ��J������a�Pm�p�B[��D�?ܿ2F\�E�|ƯϺq(� �5k�=xE�\�	TP,��]/��C� ߮'�{*� F��d�`TA��8���6̤%sp
��<M� 
��ۓ�}���7��Omʭd��.���rS�Y����7/�q�)�?㌕E�<��c�}��~S�J@���}������XG��4Qt�jS��|�3��<7cb������%�����8M�Hl,��*�����Z��w?�Z�����d4�����¤/�I��yEQ��"Њ�̳g�>n�:�Qv��?�?@��!������Vz+nB�k����ϧ� 뎼�P9���s�I���7��������@��ͦ�~e2�s��o�{�-�A�����ڴ����sX��R?p�z0ϻ����`��"q`!���Q
�R�5�LlO���SdD�/Y�
�a	`j��P�?�x�Ny������#e��w�ːB�'=� N]�tU~RYK���eZ�x����?�wPH�h���T�>�ޟ������/c�R�������<��axfd<�_�}��˵����q��յ�k��o�qyу]]ݨy��-����6 �pQa��%`^�޽�孱���&��f���t?F!�k�Me͕5!J�9���LOr������ٹs*��wS%L(�2Zb�����9p�pǀ����Q$V>Y.��
��J �'#��cUc�B��=�>3�a�ųJy���ݺ㡭6�N��3�����g�bW�G0n(�y�7Y���(�"�L�//]�9�O������~H��+
�2x�Iz~�p(l�xZV����]�.�P�����z����s���:l��t��m�1�c}Y+�*�tXŠhT�{dUQ�-���lsR����~�UH�b�T�j�\�ϧ�rʧE�L��i��[�z���x|�N��F�
���%m.ޚ�G>7�c[��[����'�! �r����>N�K�\��75nN��"�)�&�w7�����E_��<U�r����`�*A�� ����'U�X�|�@������J�T1���Bʏ;ܟ�S��HhO���<�h�J_Ei��g�� �')�/���y�駶i얹�p�s�J����!�#wj�)t7��w����m�������-P�ޙ����
��a_�l��+��<3
�y�M���O���ȅ��HH(�\tw/��XEvvvn3f��{��/Z��*ڇ�_�`�~,�;O?Myy�; ��E�v �F�:�r�7�Y��>xܸq铓�LP�tEU��˃E(�Q��m�UQ����L�|��L�cu,_�Zuڤrְq�f���yq���.��Kyq/�	J�MN����g�B�j�\/���t��m�V�*\h�p-v<z�C��l�%p銟0^�}��Ȋ<��s��3�ِE��SOn���sJ�?��/�0�̧*�W�[�gf�Y�&��-CF5̽���ho�b�ʬ� ����q �]�_�N�S+y��DQzmy?��dXN���k�O���O<����\~��ǿ��˿�ӧ�H{�meEZ�܉��s7C!�����r]^�,0�!��e�a�;6����Ea��Wm~��_Z^V�"�Ue~[]������TAO�M�>��yYm���㓲�d]���D҂?�̼(��!&`ѽ�,�^�	�wQI���O��z�(p͸�QQ�'��L)@�O�QAA�>���m�E�06�g���4ߋB�Y�lN�G�b�#c(��z����`�R�G"w�� \zO�\4�s_��%���}�q M���p����_��| �����U�<���^ߵG��Rm���rV�?��y���)h�����'�|mCC�%����9�J�]��K�4��D�ȍg��:�hk7��~�3fL�e�F�eVL������}��g-��� ��<w�)�9(gS��~7��sdZ��m9� ~�6(�Ϻs$��C�v@�����/����(%'�r�H
Yi�Fۙ�5'|ʊ�'2�zi���~P|tO�z�q+;H�,E!X�����/�} 8r�a3�%�Sͭ�S���_~W�T��p�G4��h+���kC���[�-m��ȋ�^d8�.�K+|ݏ�j��.�3k�Y}�n�<�ӯ_����_��#��ܓ�/:�gRx��!,��L&OE�宥�����=Y�\׈��e��a�6iA;��@����<����"j�,�_֢��I�ϊ?tw��y^�Τ�D{$y��M��pĔWT��]��d�+����w�G���a�1?�ݑ�v�$4�X�:V��x�_P�T�P��QO(��K�R>��9�oX�dĐ+O!�㓬��c�+ݏϋ�p��֓�c�/Y�����z��B!�G&�%=�C�א	��UUU՞�<���:
U$*�=�]�s!kY�e\娹Ҙdd�������s�(�C{j,'�A���sT4/��Mw�W �L�%��m�ng�J�gȶB����%���W]u�'N���^E	�����_?lٲe�&���P(�E�Z(�mƠ	-��|�����
�d��
���cҜp�rQv|7����wb���-mQ%����/@K��*+��s�Y�9bd,�G:;;�^�y�U�!Qc�6lذ���/ZB����,:ml�'�S�G@�^�������ŊP��6Q^����B���M�Pn4�#�5BqṸ���nZ�ƪ{�l+V�X���}�z��6TVVvvvv&����x�kkk�.qsss��7�<�����D"1�ϩ�R%N6�;ǢQXGY����E\/%�idz�?��}�dp���ʢ��mŕ	'�Tb���;]z����P�+���TC�ВiӦM?������E�L��W_}����vk8��#�b�Kg�t�����u��7+@R���h�vԑ㶩���=l e�P����Ӡi���.g�qh=C�����)P�(-��O���֯|�+����y���jmm}���	�*|r=9�f\�R:.5���)��,���<{�g]�s)և�9����Ҧ1�J�m��u��ׯ���c��3��,Y����n�<�L^TQQ1P��F@�m�P�R)))�LP����nR>�����^����I��C�6�#�S��{K���!X��V����>�Ogg��&M�����/;r��&j�̙_x��7~���|Ruuu9�� �+���L�uG&�7�u9J崓�uhS#c�y�\�6 ƺéM���V�����ZX�x�O��o��/�~�ĉ�͛�yPvwwvv� q�xpV�y�mv�����92
`� `}}��	&��\���5���/f���\�D�)���K�i��5k����WJ�QG�{b�����I�V�y���	<>eE�{��vw�()Ŷx^e7��ʮ�3%N#E�꥕����&L��ùs�Ο��H����Y�f�O�YUU%��!(�rPQ��Ke��=hs�|)v�J��pD'%���~6S���
���s�euf~�P��VvGJ�mPS�ȕ����1��a��{�wP"�x���k��/�uQ@o�fv����R�t�u�]���N8aNO���g���[n���h����d�E��Efܽ o*����\��mI5ֳ�AEe��� �:�*���������'��(9A�O*J՛H$:��˞�������:�����&��;o��§gE�E�0�:g��M 4�S���{�.gs(Sg�j�i�e���E�p�����M����8_�?���W�"�HcMM��ٳg_s��Gg��S���1���NS%(��L��<=N8�閿K��A�,׭[��c�=����|�w�q��yvuuUD��#cU��������i�lRY�/���˭�p���|�S�Ac���x�{|�ғrPFolll8p�G'k�܋/�8�>�5��;����O��������G�WS3`BWWW�F\�@�|a�I�m�P�����o.�W.�v  �O�}D�d)��H��~��UJ��Xuu����}͸q��s	��yh�%�+�1�(h+�_ ��"sn ���[���	A�$_��*풿�8��L�0�P(�p�'|����Λ7�Ɩ���*��?Q�W+N�o\HAle�Q���ԙk �2ʌ�� �έ�����O���gd�RJ!������C�wڕ�>sҨ�:�z	����n��sK�~�g�S*+*noo��!J$H��6o>��g�N����~�K�2H[�X��&+����t_��� p"[���i�a��[��kN:餜TOj\�c�<�+̯,~Q?���xBA��~o�_���;>7�@����q��{�8��C�P���:��˗W�r�-��dӧ�VTT�+�\oS
 �s��Bge	+�!��������A�G�ic�{����lR�*ڔկ،�&����k��j���5gΜ���^k�&{�=.���#V�Z������-+UQQQ#�I�-�Lv���l�&�|7�M�e�g8Qy6B��>�΂�$�������o��7��>�z���d2�`8>��� �G֒� ˾'߷'_�&��A/)�mݸq��cǎ�rG-�ǲe����_ߵ���*p��.�+��̜�H  �IDATy�C�T���>��/�V�	$v��Lr��^A�A�	��h9� ��ۦ��������:�����g!���=�͟��g���u���S�x_����D�	�BeA�Y��=����$�t56�/碌��L�l�dM�B����S>�+�r
��M&�=u�W���O��ӹظq�QMMM����k����,)
�h��+(�#�z{���9��3f�V9�1�S�zÆ�ǎ{��X�����ȧ�x<>����wSi��1�}�qf� �A�c.�WO&{-�4�S�D�o���}_�-?m�p�)2%����Æ/=dԨe�_}������%�߁�������y�o�f�ڣ=/1���r0��1������G[_���m�c������X��l-�d�+�F)���(�!zuvt�C�Y��b�!���dk�,GnL(�[�!i4e���I�?o���ow��ߞ����[��0&��x޿W��{�ҥKw(?��������YC��h�H��СC����&�Tjoo�ڰaC���2���E��]�,K�·��gw�}���9C�2g��i�������p+	�{�����[B��F��^nhhxvܸq�������˗W�����4}��}C�P�"��}�z���^YY�d!C���}��uo���߳�dS"��������(e���3{^��8����Ic�e��m7���D"������5;�Õ�}]���m��n���Vw�X���i�<�-�յ%�%�G��F�<��G���СC?�6mZS>k���R��Ʋǽ�dɒ����������6m����N$�
��D8��ɤ�,�3&	A�d�/[�掻�q�{���F��x���a��q@�1i<�Θ4.~2N���O~�߾��"a�ya/�¡d(i��ԘӲ��1&�������pg(jO$M�H���΍w�}�_�������w�jjjD�����Ӳ��pWWW����-�d�-5���ye�%�ɴ��L/0�LF��p��<����T�B!�3�L�<��o��S���z�k����9��K`�����RH3�]��u���d2�Qc�t��y�
��P�q'��L&�{�GH�1���J$�Ϝ�e4jMd��:��h[(�t����9s����px�>}jR�r�|��i��~�`���/o�{����>ӽ_����R�;]�lV�<�8�dKE}��P�}:��%�:]��ʪ_���TD������ͻ��]�0s�ѿ'.�{��k����m�lI�w��Qm���*/-��'X<��j��/�Lߗ�~N�Iw��~u����Q�G֩.�~NU�6t��Fc����q���K<"y���!��ˉ��g2ټ�OJLI[`��j���A����mP�C����X��9�?���cfAt��S�b�b��_)��%��i@k���1O=$���&,� ��~.�� PK   ��OX@��)  /   images/b4aefdef-6992-46c6-bd27-cdaf728c7c35.png�{eWM�5��I�� ��w�;�a��]�kpww'@���;�>0�溟?�~��յ�ԪSGj���Qj_�q�(�p�|�@@@"  �`��롭���w�t��熀����1��
W�,��sރ�ch�!��թb���A&��A怳�>���P1��c4�{?�ԗ̈́�p�i�7�o���q��'Tj��7��+ ��x�t��5��@�4ic����}���R�&�%��_�&D�]���]f3�d�Z��4�����H�Dc��K�j���]tЋ���2������o'*�k7}���������vF��*���g�u�ҴR��FR�(��y�J.���{���>u-y)��ȕ̚���7���/��L�B^��Yz�v���~rm�$�=ھx���%����$�p�(�ێ)�b�d����RW��#|t�#ge������&$5O�v}͎��l�<��էa```v:_��(�m�Xd��!�wgKG�}p�9��q��Z����*��Qp�!S��r0���t{�M�����/*��s�OV���1����3�eȃ0 C1�H�1��Z/[,V��c���~h�~��y�o���}��!V0oڦ���\�#�<��n�����E�v4̥]���<@ �!T���x�ف&dlJà�m������b���-�Ɨ��u�(#x��)���Ŗ��7|x�Z�j�S��(u�2hU����Y��W������ݦ���Ԁ@��Ga߾�X�Qm^�{0xy���pg����w�ל���/[��cu<َi+�u"��ʨ���۳��I�#�Uc�&�[������׉������ܱr����X�rAĈw!��/��6I�˻/Ty�O�R�0�,�8*ɽM*�}�վ���?�kV4ʷ�%�Û��1��[��/uzM�g�P��_a�'y�|�1���!�cQ/ے��恑�x���w��0y���#j^�gX��n�DT}ҨL�@�"9�=H�y_`�~/*�W%�L�kH�3DB�5,�W�@?{���<��������ѻ��껀��	��/b[;��W.�܍d~UI�o�/����R��6�P�wWа,����T�^Nw�A�֪�����%����t��'7��Iy�-�r�|��cC>�܁�������k�8TZh%嘙�k�,lV3�U��{��T��}@���旜�4ӏo��g�.��Bv���sfK=s��:����ʷ���L�1����]�j���1� ��6��uj�[~|�eĔE ���^���/�O~�бd��v�z�7s�2��L��xm�$dr~�t��������L��E4O���q�~�k�9�C$�@«��
0*�9�A-p����"���A�ݻ�ޜ��۟�6�[t�s~U��q��x���}Xń��y��m2ß���É���R����[�gb$Q3�AȆb���$l��TDl��4�m���NIͰ$��te��S	�)��>�9�'���B�Ѐ��k���vgCFt-*�P�ط?eg�Y�ny���N~�
�57{zz=���a�	�ãNݧq:.�"G���-D���e��'7u�\aww���jk㷎wuj,8˚3�"�/?*K��:�%�����v�v2�1�bf(1?���4.�I"ɍǬ��^��k�N���ɢ������"�ථ�T01�Ѝ=�ꊟ��:&2��f~��P�O�Lq�?���N���r��`l�e��ܫI8�������)�,����_��K����>J��r�9Ih~yC���)!���5�н}������[����T�'�-�>*0��ʏwLx�� ���8?�|��PK��O)�I/W.�v�x;�0p�R�l˘�)ո|��,���/��'��:,�d��T������u�b��
��%Br���w?���iI��Q_bu���qՑ\�#���#��(a�t��qeg�� z��"H����l�D���b���.�ө�n��\{[A����a	{Iq&��K�vGm��c��q�h9���
j�h]��<)Iw��q�U����դ�倛j��^ ���������\���D���->�ao��'e�讛���K#��L�FPJ�p���/�_"K0v��5���h�	�80�kw��t�y�V�����U���O�Gl��t4�ʱp�ll?%�!7,5:���n�(�6�,:��F�~��%��OVfJ�z����I��P!�����'�A��F�3���촗��p�(�?T�E݅аA�F��snA�
�ϥ�=�̴�#�b�gV�-�g8����;��'*.U{q��  4E�~���N�I'���P�x��A`�*p���C���Kښ�'��O��A�/6���ކ�5�-'_dD�ۦF����Ά�()��]�KLjQ�E�~NMq* @��5���C][���pQO^x�/�-�&y	��� ���e�lYfʷ�iߝ~�k����}�6z�{t����͞ �N�qC��:;1���ަ0��)�U���vi��C�s���W�C��e�C�t�4��zp�X�_��W�����|�C���Y�å��h,q�W>x����q�������Q���Q%|u� �� �!lg]���i:���x��0�2�p��Trchuy����^@�xiy�+�Aa�N��7���]@4F�&�e��Wl��ȶvu��4��J<�_�a�n���^����h�3� V�ɏ�0����f�N���;��iu�K;~���j�۱�
���	�p�9�����Ew�'11���>{�� ����Xi��n�^^���H��3�@� `���п�jYY(��A�tޠ�������S/�:c��a�l�z9�51��ǡ	���.�ɘ23��K��~�h����~<۹��c`��.-0�`�2B��Ť��M MH�c��2�동k=��y��4ع޻Q�S &&�0����f�~�Dp79y���b�2��L<~�/״���Wz\y�-VSYؓ p��y�5�m��(�uq���{��1��c�ɓ��Oԝ��CK� �4�q�j���Jt�ru��e��c�^�Ӗ��󅤋)�����iP�rp��������Ѱ��K��9��L�����l�J��,����@j�z؀�8��)�����:����P�@��Y��+�;���?��1�p�F_�ϟX����s������>s!;�K�.��?&F2[�i&%�,ߧ��AE�o��U���n'8���?.pr|��~��"�9������Be��t�0��Is��^-�����V�k��]�������~�2����ԗ�\���I�p��Ʋ���0�_g���)�t����N��SR��O�A�O���� �A�酵B)o�&	\��ᖨ�q���?CK)f �����}�Tz�������-wfm�J�ʯ��&T{Y3�E�\r����8[�O�����:L\�A��.�
2���N�;&�i�Ut�����s�e���K��C�
B	W����n���~��NM%�����Δ	[��]DG(9��(Hs0|��T��a>����{L�d���H�ю+�S���ʅ�'$X���P��k�ζ�iS6�huI9g�TݓKև�=�w��$�o����''� �;̽��������q������أ��}�GnȨ�D���Eϭ�z$�mv��C�C�e��a.���}�î�d�"��_:|�y�,4gZ�L�1ɺ�z7P,�eT�_��h�Y��;u=�A4u�U��A����8agF��!�@�� ~7[��k!߷Qg����÷�Da?)�%�UZ���=2X��=o�5�r�+�j3y����s�$Ʈ�}��������*9��2�p�[i����~m�(���n�g��Y��v����h�T�ɔibu�3�T=}�"�MZ�:-6m�_�>G����Ↄ1�C�����Wwt�I���i��f	F��P��8��7��!z�Q��Y䖫*K�_)��z�C�r�;j��v�-�%�%�XNi=�a�[����x��Dww�Ϛ�h����Jj���hQZ�;�|����ܭY��f�
=y�ne����ֽ���X&t������.���t�@ � ,�˂�s�}M8Y���!�� �2"��>���
]��b��@�16����iE���fO��Zz��61�Dg\F��,�N@� ��)舞J�����Mm�O}ɟ�C�`�}�!�7���5it �dC�lL�$�I�@0*`Z9��2��`�x���bM�=9��m��:��?���N�X��u����Q����;�#�ï[�~#Hqi�(�O��P�w���w�����"	���W8�@P�&�u�kg���J���;�z3����{'�&.�����zT^����l2�>M����!UG7>�o_�{��r�&w��/6Ey��~��<kB���׻�N�I�p���f
�&u������C�Ǧ�;����U�1�������iDJ$�w���v!sT;K�=Տ{r���Gj�{hN����q$���ͯ��X#)aG��Gy�^��	�4 �C�	�^�X�&1�O�֫����D)�Fg����S�L!G}���ϼ(nq9�2�tR�+��eF���#؉ey>�NR��g��?��tBy�L�}�Or�:\K��t&�,GY?M[q+1�R'S�Μ�4�G�oֶ`���3����|���d�H!E�BΛ	��.������W�ɪ���!}{q?ڃ{�fl�|�J΁���e�8�ސ��ìs}J_n��R��.���ι�7r/쮎}o���=���0��B4	�
κ��ez�Pބ�O+��MMf�һ����I��3��O6����L�?fn&�ٹ�I&�)�z����= �w;zm�)�'��'|�����\���~ݚ��������>�� �=����L�o��ę�r��{�#½�o�wm�?^���]�s-7��0�B�����$���\�D�O�c������&yG˓���43�6Fcq��dUK�:4����Z�X���(��A����wā���#H2��BLΔ� �u~� .N9w������o�^�u2i�x�5�5��w��<ay4�˳HI�/��y��X�׏�II�D,���Hė�>����S�����S�_䬺i_��'a�e׎3��f�֫G	�?Kо0l$�2�4��,���wItN��f��s]w�=ےqh����o��x�@�|Q2CX0��*o(��r_^Q��ֶ����2vf�=�6hu�B�M���U��;=���s���~	��z8�B��sJ��W��w�Db%�������{��2m�ݗK��w���R����&Q,����U�UL^|�Z�$�%���d�GҫwIC���.����~u=2jc-�e-�U"�mo���9����}?�Y5��8�K��~��b��(dk���#&؉�A2+��4�2��&�(p#�u���^b��}Vt=9�M�q;�u�����S4�9X���N�A�ӗ��(x,'�.��r�j���n�\��K�MI�T�W��2�����u��uP�l�����ّl	K���a҄X� Oc%%�Ж3���J�Sd����R��Yp0�0�tXF����0E�Z�T����� ���#-�B-F�܆�?�]�<�K����o�	�$-3</M�_�N�f̊��~�x��)�Q�En��k���?ĥ9�ZY����x����Ìi�{��d�W2O&E��_���'*�N�
6�+<�.R���S�^�G͊o&BT�7���3K�����ݍ�o�0~�0���Vd���48B�Df8����ƾ��Ѻ�ʑ|r~'�"Bm����wK�lN��b�-�37��:�������h:`h�t�2}���;��-�)
6}h5���LY�� ̓^Mj{����6}�:韬�sX��е���'�W�P�g
�l��LI��g"�P<A�9�a#�w�S|��1�H�8@_�����fP��qQB<��6��
��T��I�as��!S�����S#l��}�t������P�a�蔏���un�(-@��{XV�J�@="��u9�f��6]�8c�π�n�1mڒ����d]�^�h��c�M�֤�8�f y��} ��Q	���x�^�;۸���L��ܢ��:f�$/�駭��B��,��/!��g�cۓ7���:	�%~ �J�O?��������X�sG�</W��Š���f"�
�u�t�fC�s�������4�;tڇ	�c���;B�dF��3F��
s�U���o�KE}�|�	=��9�&�Hs��|�C)���	c��*�n^� �S�y6A��/$=�N�1&K��i0�h����ߩQ��L�\�%ޑ�I�u+'���U�U���/�A/3� :Z�AY#C�{��:M%�5�-�2���h`���B���fϩ,�f�K�� Dc���	W�@'B$7i���#�yDh��IoFb�&��_B�����4�� �#�\c�aA.�%��ھn޷��UjU	,C��^��=��EU�($bP��rq�℈�?���BT�Mm�)�Gj�d��z�㦨�OzG��|��U�}�т� �.����������wb���ٙC,ddD$�hQ���q#�� :�9�1=#�Ȑ�X��Ǵűo����B����v�X����S%S��!�g�VrLo9��/��:}s���~�<���j��h�`D=W�g�������|~\��<va���|?�=�ď��٬<
?�vJ���M�C�
%�� �T�h���>�7~�*�į����ȵ�H($�
�Zn���E��v��g[�?Ĥ:¥L{�Af�b%*�����3T������G�i
ߘ�jih���&��xY�O��fB�,	n*�×}��?��V��NeV̛ X�)�S�';*:�2<8B���:&5��їf+�N����=�V���2��/�)~Չo�u�&��N���v�y*�'����&����޽�\}��O��3�ןf]@��o�VA@�<P��]�:P��1W=���k
9�����5�o���~���b��J������qpW^�W����q3D��GX�a
���9����������d�o�S-|�>KU�@/�J�t���������x��
����shu��}�h���_�����|fv��o�M���I�>SD�K��/]�P|w��=�	7U�2��mv���٢�I�D~���z}��	����g̻�a�&zF�#u�F:��Ʀ�<CHJ�����m�{�|Э��Y�f10z��W+��C�]�Qz@R'a��]/	Q�O�����Gv�k�L~�x�Jn��ʻ�[��y���bI��H�lۗ�8)ώFnE�P�U�[cW��q�y�t��S��9�"�
|X��:[��J�������O�4���d�m�7�q\K�,"y�=�T��	C��'��c�J��ʕ$�&���į��#����1#X����p�E�.Mw].�K����1���	@���87�N�'Lw!6�ۀ�5���=�?D	��F�~�	ن�y���<9f[T�	1+�b+8�m�R�JO��Ũµ��Bgw��?�F*�.\��$�x_#���7��;Yn3�j'�����=]&϶��D��ID�x��>k�7�_c |af*PF!@7S�� @��o��]}i��f?�"x4�IwA7�{y���nwȆ�4�> �.Io�&�p���kަӢ�֌2VبXݘM����X qJ������Z��=1���q/g*0{YY����;��d<�/�����_R���*�[��Vݤ�*�ڜ�fS��O�ʲ1�)N�CɎ�'�������5�bc�s��ID�Ή	�N�u�\����7S�kM�"&\��2ԥ�^:�s��b�#�po"�V'-#������Xkz��^>������FR��Ν&��v� Ix7���^�Cf�� �H����|{�	�Ce2&�?��׵��l9�^"~��o7���C���/K��~O�w�&G/��qvm��(�&uv����7{��Y|3n<�#�Ɂ�Kl������v�X���(��{��!0�2qƪ��\�C��D	f�n��_4����Gx���^&���|"�V�-�N�����/1v}ŕ�����oӉk�]Z�4����_��t�}J&��MP�G�h�	�+��4O����Zy��m����[�^�RXi7kz9��\$v��V-�>�_������Λhp(��:;�{9q]sl��wy���x�	q}���EGA��+Sͫ͒D����A�Y��oG��G5T��E�]-��D�ep/CX�H�QY6��0�ة��hK$���J��N�Ã�C��k7���ON@���,2����l�r�����p-�'J�\���9�����a��e.
B5I���â�s����.*����=�K�?��4�f;�:�׀��B��B�aJ����1V�O�)��/�E��Fmcڟ��}��_��t�l�2��.����1��g������6R�������lN2,8�
�]�S�����S�}U�@X��Ɔ�Mve;��a�0
$��P)}��7#.�T��G\��lp]	>����%t.����V���΍%+[J� �D��h�li��z�X�� nw?�x@%�>JY�x��h�VP��l�Sw~Eji��u����|�M�6���j�^�n�JH�ؿ��dbMߋ�̬�����F��U�!�k\��O	˴�͌7T����r&�m10ͬ�:�j�����ז3fU��Ѳ��W����������E HRBt�U�(�}f!�JBN�,km΂L���HVӦxG 8t���h:�A� /ɒODO;���;�zo�;".�G�,W����%�D:�C1C�5Ŀ@������z)�Ɍ�#�2���OR*dҞ:����ıd�b����t�q���c�׏��q�s�{��RQ��+�ж�mi��s	�l!���UͿ�!�
���)�;�;��Y
c�)�PCp��N�G�_�E;Wh�̲e��	���̲f���56�eV%���e1�~숆�գ��[�+�������R��h��R'��F&��	�@��8�P�'H��E��KX��G"rr�[ZHK�G)�c6R2���=n:�HU�@6��{Q�f�aAb���<��װY�O�}Q6�w*���3��#�����I?I�f��>�%&>4��y� ���VrCｰZe�|x���'Wj��i�o8��e���V��2h}���=�)O�Qe�F2�!�45�L�4ՖuVj�a쫓ρ��j�+$���L�����BU�{�^���T�� :��vYI���
-str�gv�B{t,����kk3�hƃ/�I�'�_%߿��j�v�M 3�ѓOM��D�%�͸N�������z�MD��+���z�@�wL�5t2��_~�c�E�7��G>�w'*3\5�kImt��m���~Oq(^�˘��W¤�z��%7���C;�j����p���v��^N7	a�cz��u�o�j���'a�$��%�7����fQE	6c�c��|Π��|��&� LD\������Pu53asE���z�[_�&�W�@i��D�%���Q��kA�_�4m\��T E��3:���ÄGZ	�@E�YdF���-��>?s�Iz��b��m8�#C[�-�{�뢢!t��!���R����g�1�z��E\���Qly��1sF�;/
l2��g�(e����2`�����H�Bl/!� ��ޏ��ǘ����M�c,W�|��8d0+vP�]$B�v"��GO�����+E�a&$���ћ�P:�>K�P2kŖj��0ߘi������L��o��4�Y{y^t�<6:�V��\�{�}9I~@`��;5�W���o���j�9�ѩ�Q��t���]���k��ΐ�M�7�D�_8�<�C%�[<2��� q�J��ڂ'�B&܅1{�h�����pg�-�^�Z�����*bA�ʭ
#>���+��Bn��d�bksx��x�#}\֜q����|m~�:��'U���A�V-���8=�P*���]	��Є{��9p��Ɵ\�m�ی����o����|{x�[�h����k:�h�f6�>߂����j����<�'�(k�p4��V�I+�$���L��K�5ʿ	��J��l4���t:e��<�9�PU6D\�j��m?[nNp��)�7��.��쑙Q ��uA0��H�Lm��P�ݰ`�1�ixʧS���\a�Y� �~����i����.������|�ɜ��V� �tJvLv=rq�EZ�0+�R�b�nE�G��S+o�V��)-��жx'W~�>3�_[�x�����}�}�z~�ʃ�cQ�C¤��-	 �"$��"��5h���K����g�k�e�$Cjk*�XE}�>�~����וVBVk��'UR>�S����r6����8u3�p���FM}�ԟd���d�n�m?vR�ܼ;�?�~!�l�9�������Ti$�	�vp�}�����>�CөP`�^��,��]�&=5h~�O�{G�O����[�$�G�r������:7Rv�����IF^���9%�L�;���l���&�z�0,�Y��-S:�$���f�	9�)X����8_������O����9�O�k�塩\S�m���B�+X�9�ylI0k�����C�1{�^�� ���-4�8[��8�5N���I^J6sA����ʦ����j�QY������硖�k���M�(���_/uu$#]@�>�$�!�!����Ea��=����fw�>H3�94�Q�]!g3v6*݊4������ǥ)����t��T�_�P���6��~�a.���7",�U�K:�|/���βڶ��]�y�}*�?P��*�~_1�y�.�<���%�L=�-���X���>Ҷ��*M=9��P��od����ck%��x}�ȒMP�I�]	��1mS5�Ҧڝ5O�`L�@卬F�
�%�����7+Pۣk��I��,�G{4BI�0�1�֍�.�K��~��h0�4�E���;˺�~�{����,S�Ѵ��i��=���.%��o�˹�A 6��Z펩��Í�ݿ[�q���9�$M��<q侺ň�����+���������=ʐz~Ffu�X�|�?��}o��K�!p0���ur���8�lD��g�T�>�P7�����a�"3d�3{�
g�������J��%�����|�_#��N������f�j�TO��9=+qT�6�#�L��vf?Rk��|��g���qm������O{�֦<���K�ڝ�E������(u��տd�!�ӗ�A�vi�d݇����f���i7��тG��C���eCX0�h݀��A����'^X����'\�eP+�θz��J��A7�K� u����S~�Z4)��p�W6 �����$�+p�c����`&X��8Q�p��w����Ϸ䠊9�6���A�H�ӗ�u�pV���*}���F���x'�ssd�����1c���{�L�z��R"��o?E}pA����򩓲��Cʜ7���*G_���cv��U%[:٣����|��&��y�|����C�w��fv~]��__�F7H0���$��p<^$��E[BM8�NEG^&�ht.�C$�Q���l�uo�޺��`�4iM�w�q�j���cN9w�5u<ǹd'Y:��n�����.�m~�}S�֥���������x5S�-K��y�����5]G�_�R�-��x`P�8�v�(O�>�n�ݣ,T�XQ����w��������� yR"Y�#l5��`_��ݍغ�G!��f߅�jV��+�����ƴЅ�����
����=��޸ �*
Rj:m�z��>�XS���=:��uy��}F (@�ɽ �X}���p�&Ϩ-��a~'��J�'�:�\}NP�U�&ֽ�m6�n9B�����Z��+�V�[�=���:&���H����ʄ����wR--VX'����kT�g/S��*9 ��T�x�r�L�����J����#v�j15l��H��`����07��gQ-!���@}U��#ƽdL�6Ά��
Ȇ5��?�k�2C�r\`q՗]��b�w���t���yb�h�&`�!�+��k0x�í�ϛ���J�{[K�x�(u�J�Q���j�8q��j��@]"���z�8e�i!�#�Y�Y�1[C�u(��| WuFR��}�S�-�ƹ�0���Q���.�6wm[w$��Z��C7FMЙ���o���ZTnSfv�-a��i\7�φ��_�v��i�u,�eV�;�'ᶔ��B�	��s�a��5g����'|����%���2��\1v�Xk��_G��!��a��H�`����*�41`�~�u���cɈ��t<�	�b����a���0�$��e'1ί���e��c���
���fjg�*�c-z���m���ٚ�����a�fV��ߏ埞�7��-�cfN ���ˊ
��C�+��a��Ѧ��#���a:=i���ݦ]�W�ú�{K6����*�%��d���.�7�y3����-�ʸ����G*��N�Ѳ^�����}L�[��
H�9e���"#Z<��
�F9�6�T�B�ix��P�_�3�̪���W�f1[(��O�|�S����|=�$���b��X��٠�f���:{��J�p��j~��,��-ST�z
=C���+��}�?����X��-�H�k�~�}��XD:I��
�q�h��Dj9�+#D��Z83��På��{��K�?@݂�uq���Tȟ<���J9�!l��|�3#́T�T N_����"�4?���i������0���`����1�n�=�����r�(j�!H^�wp�e�<���\����haBxPXFiY%�Sgd�����f�*�ZH��ɩ2����tƩ�*�(RU+q�h��z��h��/�)ݳ�P�c�SPs�H6���i31�~42�x�Of��l\,���\���x}Y��>9=q�ґS��U�.����<jK�l���l1�#�������m̲�����X��u��Ē�)'�Y��G��}�e�����ū�b�3���n��o�\�G�wį�/m^��P0n�ө\��r�(/~�=4,��.�姚�LCn7AHB�٫~�#�y��cl�qt�*����ApCZS��.fe�s�6������{��BO�<ae:6텖S��:��N��.�Z:0�ͣ������o�(O�����'��f�y"��8���M��q�U�<X�^���>�!R��q��<������z�V�2"���s0�_�5E�HJ��ʿ���P�,5O�!��1��X��7Fq��̔$��j3��w� ���k��[
7��<�E�Ӣ��~��x�B
j�y�I�.yIl��}�-ɌNR�?�$�
�����&LC�DfP��R��J���݆�׈O���Ά��/���,[k�R�yEaQ����3[Ҕ�ڪ�B�l%n�k���@�K��fT�
��ٗ5G,H�ߴ�6r4�id�LB�O�[�j.��e>��f{ġ���@�Ñ$����'���䱳�yl�sZY5��s���5����k���7{� �c�Dqn�C'�q���Љ��S+)1�I&�4W����+u�8D���w�ʴ�s4�Dse���;tQω�{!H��$�����n��P\��n�y�m?���Z.�
5���%���+������/�"Q����K�K';�0+�O_���fpm�ֶ蚾C[%X�Fǳ�	��k��p��/ 5���Ge�K�;\�R�+��2)Ʌb�S��&�kS��R��%>Y�'�M������"��gֲ�����j,���<�K�p���Lz?���(�h���p��X���[zeON��B���J���qSZ%�;/SSr�A��RO�>�g%*V�9K!�����,�M���F�� �ね���ѱ০8��r��wa��'g'���km����G\�Z�Y3:��#�Mp��I��)V�f�֨���ˏ6�z�<#Y+�3�=Z U��Wں��-2⺃��>Ur��|֩^n��n'�Io��D%	Nvr���f2᪣�L�!JÞ���7����[����̖�����SL��tGy��i~�Et��TB6��O�Bz�-V*�A��o�Nb#W��J�,�W;�EZ�h�~-��:��
�H9��i|�
��󝾶Lw(a�x��ZG�(.��<� _�;dּ�5<�?C6���[�D~p��ep"P���4\a<�|�E4��CLT�Gz���P����6~)5�^R��4+�{Oc�m!��U@��s��~#���Ygw�Q:{ԄDA�Hǔj��`�l���m�z�T���^������(��y��yo9(^<iJؠ�X�D�H��~3{�Ze�hz�A/��ܬ&�L� �q�} �#j���U�ea����m�~c��J���l�
�R��3U{��a@ej������7��U����~kz�j���vi��&�h胃F��%=��o�ETYB��&F��l.<?�-I3�t�'aV�D�^�$�~ř����闧U�p�$�d}!q>ah�Ă��~t0�jn����#��)��Uqs���B�����	RH�	Z [��������U�;Lq�t#�*��9�#gCp�mX�B��bj�U4��ݏgY��,�}PZ+���OZ�YMh�l�dH���c1�]�tP-����
�jQ JAq8��|��Ҡzc�Gh#��p|����2�b���QI��H���;
W����	[�e���ALK-є��|�L8Aqrp��s岎z�B��5�Q��0�b·��5�X�H��w�~f� �i�p�Y�~�.ஊEH�4�/}�J�hu�[��1��k/o��|�ߊ�d�cf�AcpWq�M��oJJH���t~u(]�ݚ��F:VV����GL����4��f��'�������G(=Wa��?��)7���`{��P��s5b@ɠ�4	�03��+�߁�pߔWH��^�M%A$^9�>�L�o�NEt8A+�=�?1M�}a���V����ϥ���l�'@a�dI#����h!�H?�M�i��Y��Q�m�y��Sx�%պߙ�!�G��0m���ɓ(�B�n:#	ڹG��$γ q+�x�Ɋ[dO
�)�@y�>yS�-8.:�=�W4�k>�f&NWtO`�^�57H6f25E���vi��4���W��Th��� ���eۣ�ub��h��U�7V�7j��kc�{u��M^Ou����p��}�S�t��KSf�`+�5K�F0��G�-��ݴ%q����2�P��I�D�����-��?�i�j��"�lqln/aQr��[���]�d�XL�B�O�H�F��ڽ�ϣI~�<�H�8�q�9w����-pcRފo�5W�����6����y�_������yhiu/�pS�(WQ!�O��hn�@���r�|�U�Vfٛ��!�㵪�R�+_���6E�f"8�i�)bR�w�p��X�rҹ4�؋�t�vDU}����ΆCo��#���X:#9�.�%��7!��W�d�q�Y�5v[&!�/6�a���&�}Me���5��\�a�$�K3�=�Z��K�y|	�x)v��3h
I�k�8[���CY�9�"-��b��ʲ�8�!�[�ed�Ρ?[��m�gAX��Q_2!�2]+�*�^���_61��ΐ����F���c]׽�J0��;ad��n��|43X�����?g�/r��h�?I�tf���X�f��N7�i���:4�շ���T9�Tɝ�l	�%��5�J�@ա2Yg�t�<ԕL��KO��W��|І"Q��[97�b�;V��K��F�]���}9~��-�
E�AЅ8���e`���5�K�5T�-�J
�� ]��wE���d'�X��Y�{L�Ͻ�/��pd��Х7��ofM�$��n7�n��ƒ�P���z���6kjMx�>!�O��G����D�����do�� �����}v�zﺩᩋ	���=�05s�T8��x���T%`������f�P�F���1���i%�˥�9�`\�&�����Y�s����S�l���k�t�����|rZ����$7���"���C ��	�]ωs+5Nf����0�?t�k:�V�@j5��泥������hƄ��m�"ywc������N+�wa�,��6�9c�%��J�Q ��qx�e	�;x5��������HB�	���$��#*����v�յ�?9"M(��DV~��Z������N�^|�k�S�B���Ch�0�'�	����ŕn�dc|��`@����=���p�NkWm���F+ox�l���@����U=�}�Q�7�I<�`2��� ΑI�R�e���L�J���gA�^��-�ˆ4n��O)@Y.���߹�*���?nnl.���,?w{�e9xn�c�#�g2!�����ԇ�p����� ���֊g�n6jg�ݤ�D��w�k����<B�n�w��ۣb�=��K����O^X���+�.�L͗SOYf�j) �"(�����3��_����L>t��aݭ@����_��X��?�Vv��Y� �\r�B=��u��7+_a�\6�Z����oy�{߫��I�r�����{�<��	A^h�ha��,9Nλ�U��̳����m��fx�^].�`kq�{��y�{6��	���4�!��`��nيSe剧� ����|ꩧ�� ��yh����Zy��U�c2���7�?�,Y�D�z��������؈�E���}W�k��rQ�Ni�\���0����faiٿ�[3xӞm<W����v�1Md�̦$b��6Ԧ @������ܢ{d��sn��`�{3���fdS���s�|<�	�,���eB���mA�&)�x.6*aͨh�����Z���7�n	c
@םq��N*��e��?��I������#��r���m��B%��B���=�a^LJ�l �!����ݽ]
���B\�L�=���fM��j�a�[&˫/�B^{����PA��)�����G��C�ۨO��c��>�6���+L�I'��e���Ym���������a޹���y�0  pL&�(�ʠ0���c��]��ʕ��l�/Z�$�d���+�/��dD.�u{�r��%=��q�O��g�cNF���C悈�2��m���0.S�k�<��s+M�j���)`�`�N2V�"�9Y�Ƶ&Ș]0�7������6�8�E�(x�
�;��m��� �� �XS������/lIg��m���e}gW�(J-f�H�`�H�b��@�iZZ͝�/�5����>�Y�H�U�fLozӛ�G?����|\(8�:H��A�� 
a�1΁�q����{�9���uP�9|ͱ�&n3�!���VѶp,�t��Y|��CK�a����I���h#�YP+�y�+����ʍ���ovъ7�&Յp�={�Q�^�8�S
}�R�`q[�V[�y� �nb�?@��o���<�DW�[锉u��D+�� �mj�Ԩ)Ad�\ 2K�K!�j�Ԩ�ٓ�������S��B���jx>�R�pKoP����s][n����砐!S���r��D%��Z&ǘc;�)hf'�E%�S�;+0"���9���)Ӎ��Sk9�N)�ӎ[_c>3 �$��U�Vi�}��>4z0v|��|@���AK��xZ�ZV¬'Xp��M$��Z����Wf�c�!4�
���`�3�`��orB���I� C kD��=��D�Z]0�0AH�:��4%E��9��&S���q�>���Ae��4Z�ʲ����{��[�Fv��l62�X�ڪڭ��S��؅3�5�	�^1�`Xd�7k��[���1���9q���q�ݾ
��ϸ �}n�}U�c���?X}�|l`ι+�"�u�jSxP萑��\�����cxM*9n\�֔ƋB�D���*�V�}�>G���(u��.>$UyAY3߳f��x�L��@�(iM�V�y��k���Jv��M��.�}�z�ɚ�w/��:a�����^˶`�c}2>B%�c��H�A�������<hR�YK���Cca�F���# Ԣ�_e ��&:M^jVdH�	]F�����'�9�	�&7L=������L�Z�ٔ�4�8���2y��j,�}{wjuC<������c�\Ư��76��zfI�C�ɝ��(�x97�;6���q��Ժ����2p������$L�q��]?�мO��.�A���i�3��j�T�sq� 7��bl���3�q�C����z�TɨR0x��n@V�&ok����3g��!FѪX�3\: d�gRz���ף��F�fQ	����Ý��|Í�p쨔a����G`n�t���o� �7T.�4ak���ΑF��e5@�'��H0X,$�KޠT.EL<ה�����ӛYtA�ܰ*� � ��P�Z�|h2�Ajl�ri�R��Ak��1Q�@��}�?]#��
�4�kt��*8��s5�cw�i����� ������OF�Vo�68:��}��Q%V��;wFnBׂ��B�G�w�n �V�{b����.��2=� \�َ߃\��gD	�p=h�(3 !F��Z0xKbk� �lT�G�؏�DH2/�����*3�Y�ZdAֱ�����ڗ��S�k�PR%ݳRƒ���c�*@��芳�����z�5:�pc�0���G,�`����	�*�q�tsj6oh�R����M�h��z47DD��0Ml�FZ�į� D���8��R��@.�!���q=�H͎.�Lʞ��&C��v,۰)ߨ\�ճ�`��i��/2�t�X&<����oW�4炕S]�>��=�c7�t�n>7�]����;2N0�~UPD���
��Z�h�1F�}�_q����~��������8'��abS��x�-��d<\fH0��,@�0���	����������߯y�k���>C�_���� � 0@�l��Z/A��6��BU�޾^�_ 6
����V��,4�?~��(yYM��֏����
E9w��7ܠ�?ʺCQ���
~���댖�Zfx��s�X��`L`���q�����f��v����L��f
_A��R��B��G퐈�������Zh��k�>{����]��ɧVK�*}���Z�@�YlQ�ޫ�G�;�O"+-��.4-)��) Z�T@W��v�8�Mr�>��`=@��&eB	���q�\��K�.�x7(��+�g���!M����`�{隵�ۼy�BfP���KK��up,�{�'��\ (`�x�5e�b��!��KZT�:��"����F��{����u��S�į�_��g�2�W���rkn�"�g̷E���ݣgq������ *JVٲ�����B�yC)g�E8�T�xp��+�d�a׭��v��B��1*M �����#�礹Z�;q 2w�(�M��Z��+�B�ߥ~!��ν��COjUO�=��%��G�n]���f�$5Ϗ�:�7k�'�#�%������_Z�{��H����6͋[eQk����܋-��$޿�����w߭��:9������&����`ʌS0���Ƞ/��zX8�t� ��f�ƅ@n^������,�×���~���Gq,�����gsv��p<~ñ� �|�I٢�O3v��B��(@�U�u��SOJ�-Z�y��ǩ+4O�e�&��0 o�O����[��`�"7�H�����q�� ���`��S
�M�Av5|��r%u܅� #�@�Ƥ�ZRm��=��<���mL�Nm6�|����n��֐�^2�-���������� ���F�]�IYa��H.0B��B7m,%-�e6=��BW@b79j-6�4��z}�[%�;4�@�k~������� � ���C�	\�0?���� ���r���eP��Q?� 7�k�cG��!�tAo��袱L�U��k|�\U$��2o�+�j�{�N�/�F���	_���%t�Kk	h�����0��ZP�h�q�k�`b"������Bak��?��gRҹq!3�B���es��@n"�L��Ԉ�v�b��ohz����ק@�����\��B���6��w�N��]Q]=V`�B�n����_ށcC��9� ���h���
 �#H���g~�_����0��`&8�����Dt��."ąC2�ߏ�i�L}7�׍Q�� ��pqshE0Ǆ�D�ؖ��h}�0O�/QP�s��5�ǔn�1�u(��^`��5Np�:N��3Q �|}�b�� ǂ�(c@&<��ts<��606��/Aᅟ���TF9wno�C�	����΀�3qӻAN,.|�=>mdsp��:l���.�:V����W얖f�,GG��� �y
}eim�&۷�UV�Ug��:�4�7�X&b�� �(�_{0&OA@���,��l���Q�%��5]j�86;|��3�b��,>�8�b�q-�tuv�0b�<|��l:Zp���5>��I���q< ��d�8����?�=��83�)p4���\�ŭT�ZXcO������9{Y�v=���B9�bE]�%-����C�K_��&��Q����z�9@�C_|����q��P�y�_��7���+����omrq� 6}�4��F.$���k��(���M��f����Ѓ!U�[�R�5&j�4�=X2]ʅ�m�e���Z�X��*�Mii$��w!c���3�ʶ�.���w�[�����I.y�7F�}��`�6���\p��Ua�a��
��[�S&������`� O?1�y�d�T�������k}�k�q�x@�L���7D���Xo�jH� ��J�lI��1
$�V��gl �#Z�`�e,�*af}oݺMv��"�]����݃]M�R���e
J�) "���泮C?���T{���\��J�Pֿ���u��O�r����:��?����#C���T~�\<.' ���+������E�z(��ڵO�=��J��\�Y�[���
T�D�K��֠�. ]L��,uiycMsHd��w�� ���|�)2�?h���oFv	�
����;������#D�v�✘&�����*�87�F���:��lὕ����c�7�	��V!MW_}�Z@���q#c���z�*���O�T�&ċ�̃���@ny�������2�I������c��@c?[��{�V�\�x�\|�%�kj�b����Ui��|�H�P�����B?U�NGx���=��c*�+7��E�h���Z�J���*���\S-����~�'���#��-�j���6Lm�I\<�\��bc�*	Q��N^5��Æ-Is>-My�8У�/� �V�`���m���O���>�}AK��A�:܅ձ����/��PD;L���,Y�9���
,;�5`l4�/���'�|R��c�6���~����y�E�
w\��eR�V���$��K$O�m�����b��\Q��н�w�Cq�����d\L�" =�� �YXXn�9 ��3�0��k����.����|�[���Q������/̾��%G��_)�TE B�GU�T�E:���}�,Eb�=,��P{8�󬲩��la78�Y��M֢�2���������9V˼c�����C<(�^\�%f��N�+t(�2���ɠ���'/��n��C#hmn��^q��^li�k�n)4o�0P<�}�4����Ȏ۴�+�}%�fWC<��(��ۆ�]�2e_q^%b$�p���!�l�fq��$����+��@Ҿ�V�,i�(�b�����j�Ę��4��e�Wv#J�>�'Y� D_4QR`~``�`R[��8n�����׍��w6�p0OM�:��A��q5z� 6e.�U�,m����_�B	��Gg6�j6o�$�=�Z�Ο#���&2}�4Y�dQ�L?%��T��L�h j瀝~�{ߋ~�~�!��@/������#Z�T\p�w����)p\���I^6cW������^�sF;���(H���=��@Qjn�*�Y.��1�A����\�W��@AT ��c2�xr�)��+�kk�Ұ.1��vݻX3hԂns���u���e,�>���eR��C�\�Z]WPf�e3[m�\J�+��P�y�3���>ʲk�G��k��FN;����rQ��:tĚ>}�E\��`B_w�uZ��6�x �IiYpBt�d�1���k}�|��u1V�}�g2ZO�%b�� #�����;8��e��k��$�*d� l2�M��%�nj�����K�:JD��&r���w,Ǎ�!��H����(p�(�+������[*J�P��x�jts@ns<#��<�PD����V	�נ["���-�� ���};d�]j�s6�f	޳��y�	ZP�J���E(8� %��#d�z��}l)��ZO�ׁ9����#����R���׀򁜌׾�r��F��۩ �fË�v���5�'g�q��6�w���$�,��Ϳ.��g��d�Ye��^q��r���F[��"۷o���{��Ӻ�ʁv�9��Ur��ʹ|����>�#��b�]�9>Wl�!�/#ӧ��Ν�d���֔kֆ�U�Zj)ؚ'E���i2�Qb�fj�����H��"p\+����S�fi����X\+�����x��P
���j��j����V���g���XC
V5o֕"���	"���ȃ+}��``��`~Gȧk}��4�9V����B��92T�tQ�X�:��/L�4n乂����VY|�rm�R�x�W�\�I���S5��dI7K���h������_��_���B����&�ʤߞ�EZiHXl��񤣳W�|�qy�чuMa.Qtn���SVi>;���<���Rr�D�b��{�?���̀	[�p��y�*-�Ma��r�}��R� K�_�Z@�`�c`����m�������vO �#,5Lm�f=�7����yg�M2w�B�>m���K��κ��ul]r��À�ϩ�9�?�I�]�>lb�3w�2a$��Dl����1��A7���k-���R��V?��ƅ��!_C��HVz�pu\���� �u�� (�6N�r7�}���h�=��w�c=:�>6n�[9�*���g�]��D�j��=e��*֌��ڦʱ�N5V�d����J;kR�γ��E���S�yGa@X���1�p��1c��-�o�p1G�c��Ռ���J�7��=&;w�0����m�7���O?a��.9�3����SČ`Yt�t`�;���h[�dB��x�J�	�	�g�9�x꼱
:�&�+�}�fО1��+{�w�r�u��	?�St1���2W�[���Ѩ��|�fvw�����d��=�չG{���,r4}�ثha�r��c��m�c�	ƅ&:�h0����5p��D0����̰9Yր��A."��&�t3��Aӊ�@�B��tx0��	 ^�&�L
�=Ρn?Ϗ����ʡ�?�!f{��E�!KL@`�
�O�����H#h��$Jh(ˉ��D3
Z���Ǟ���}.��1��P֘@���f�L6L�j�)����K�h)���z��%��,�[�����1A�Cq<}�c�X���Y��D�pЧ7(w˾����m�Q�ɓ��W6��QZ2���+=����+.����Y�Dݍ��)�!.���'jIg뭫C�M�F�L: l�s�����)��z�̝�n&�7Z��P�����}���
�Ǥ��؄��N�5�&tr��sf1���H���0�L�f�I/V ��u� ��0=TJD�K�KA������e�����S2�K�/� ����7���������N8A��N���ʏ�# ������=�I�e�9I��C����o~3��Z|X�lr������k����w�|��%�i�����uP@Q,��}-�u���J�{�U� x=�����X�F(V+���f�K-�ַ�U_�������{J
�����Z���:�%e��������M4_~oo�TM���^������[.X,��:S�S((�z���@�Ρиg�A�HPH\�S�LW�	S)϶jKy%�:��h�6�J�5��.D�{dR�$ٵ��M���Z%69zw��t�x��~�^�E����NYֲ��im�I.m��r���E�R)!���o#��Z! �XOl6�Q�o�� >C\4�0@�.�G�+��:0Y h���+TS���������|�Ҙ6�]���2�pʤ�
�۷�h�}e�+�����w�B����5�gd)
�qpO`T \�)��������5F�s�O�	0B������
��A�J����j��]pġ���d�_��v�/�˥�2o�!�cm��P4?�s`�̜�D�F�+�i�T���s���SU�?.�7˖/���g�8m�Ƿ��-:�_��Wt�1Gl��?�vwȚ'�ŋ�Ȭ��e�_�4���^�3�=�roi��Ï<(�/]a�grdMn޼�Go�3͢��2P��ф3ƎZ��93�6��l�~�L�fi�e5��VnՒE�Ф#���7��C��\D�?�zܐk-mi���'�o�M�ךg(X �{��- �?c�\'1���h7!���nA5$>Aಅ#}���c������������$8�52W\��MX�((x#@��+��2�� 0Pi��#-���&����wn� �k��q����_/pK��ѳ�>��G�"�@�k%!��6r��D:�@J"�@a�u���%+��_���eS����e��Ge�	�$�d�~�(�j�%~�C!¼3~��}׮
���AX������K��	�פ�:��;�aƻ��ת������̄�
%��n6s>$
�:�q0~�q��=p��A�ɕ�If�E��[�[��,��#BX��Q}���m��_�����;�!g��)���m�ҴԴ�=#T����O�T4,�(�,��%}蔟Ua�����C��J��)*:�p(n������}6wN�4vb��2x���، ��]�	�bW��0��i��������<t���w��C����Ѳ�𾨀pL�}���;��#�{�6D.�����8�pq���RPQ���g�\7���<����p2T#�3�M�6���}u�jv���X�3��N�9k��q����[Rf���=���c�v��U]�{h��Gy$Z[ �0���]�7�e�+����	q,V�| N��b��?�y]������Z�{���}��0���o1������f5�b��S9�M[,9
Be��S�<����� �!͙��f�h�A�*�XHnh
�|.�Bɨܶm՘�״��V|iknU���#!�h��Y��|S����3���G�K%V�g�?d.�r|>��*�4�[4�-pr5f�,1=O&��{@.�хK�̏�w�%�(-���Hp��ܠ,����0��ɀ�c�2l�QQ�x�i�1�D.ѺaN��=����C#�K����@ �4N�ux2Z�1�^��a�a_@1*h�W6g��t^�����+�j6����X`�yͫ��y��A���,�����
���w��	�
����
�2u�qъ�eZ�Q���Y�ip9�I+��9s��!<�2�u�憛��?1��PD7 &�����6���=Ř�U��U4@5%��)��}$PuHW_��Ɛ��877]�(I�m5�!x-$
�ǲ�O|���1Y��t����b�5�͒�޽)�z�t#Д�2�`���M.�����9�x�.��ޣ�&q3MyW�e��������Em��Bf��� *�-��
>gv���;&�1a�P@���ǭ��<�D����/>���?W耈v"S#�g���
5�1�C94���*a�J���߾T��7J��Հn�Q�̝ky�����29mʲn��޿�Eo�EF!	�f�z���h�Y�e]��.C�M�k>���=�ܣ�/�ti	`<�Z'ˌYs/i��gsm��t�î����Im�F �x��3T �,��6�����z��?���v����}{�q�d�tvwȹ�](k_xFt���KS�h�d]f�m�$9jANҹ=2g^��d��ps�Իꪫ���D �����N����(&p<nb��&�M�����}��K�Lj��+����V/�@$bf����"�m�X�~4�u�nj�.4�ڸ���.��L.�P]+­�J���&�1^� �fܺ��5;W��o���� �����(���$өU7&�rqc�u9NC) |>�y\F��	��0Ǆ��Ұc^��B���R���9�|Æ��q`�с���d��^[�Y��ß� �$�L�9��0!�hˈ��4)�w�F�v�ؿ���kUY�AY�9>�' �~��� . ���K˖� [�m��[v(P��y��PpSk��O�5O����j��=,��>'�]���R��~0A�>���<����<��cr��UƼ�&}=�̝�H6o�&���/�*2�\�Yc�Z�ȢE��Y�\����{�N,��/~13�.��ԟl
bLH���vh@��~.:5+添d�ֵB�O�u�����tQ�j!�]MS���tv�� ���ʨ�[��M�'s��7�C�k���A.f�ǻ�DfF�h�E�Z_�8�v���d�|>���j����
@WP��Mܪ�'�I���q��߱E�`;�]��q�R�G�%�g�[!�E*���3{��s�z��^:s)�?��ޒ���<u�t	�e��
��ɀ��Lׅ�Ak,��)Dρ����>��ʧ>�)��~����H�s݊ p}�֚�|�lE�tv�ɶ[e���77	�VI{n4�Q���'���3t��ث(���r��R��_S�!.@�M�[o�뮽Fʥ@��Y �k!V�?��J\$U͘1K��XN9m�6�����[�zu���O�G`����Gsh	`��>�� ��!& �VS{��r�@�y���ӹ_U�\�G�v�����d�
4��2|�h�hM��ۀd0��.�k� 2
��e$W@���x\���s�)��!ƙ5\
W�P�PP��w@�_�}��u�D�w�X^�.)

�q�;D(�-�x�P�k��;}���U���:�@72�0g�8��W(<𗷷O�Y��j= �����E�Sr�+��+�`&�X3��в6Ϭ�q##w��._�ׯ�1�5�\�l߾�X�}�}��������z�{߫�$���]:�)|���_����2c�\��.Es�<����#΀�����rs_S���+*��*R�DP=���o�3���!�U=Sv�L
�&!C���.��~_xѥ�?{oe�Y��>{�]c�IwzHw愐�aPX��̹�8� 
.��\NG�\t)2xQ��W�H!!�$9@�H��t:���w՞��{����U{铳���*յ�7��3��ɮ|���A��� ��l� )����[�����1 �!���x��b��w��k<��M7ڵ�^�X �!�.��m=��-��up�+;�R8;&���%l��Ш�w�;x���-��m�52���aOeSfIZ
�Єc�^�ȩ�6ŋELD�DL�	��]�G�2AYeo��@�*u�T���!b�F���k��*Z�&5�Q(c��)s���i�e3�B*u����F��Ԥ��9�R��Ɲ2���'ռRf�k�~r-��2?�f������v�s.�|;c^Fs��9J���9i:�j��y^��C���G��7�ךA��מ�y%�s�yf���J��9��V��V�c繶�����x��h1oذ��M@�*A��_� ��mp�$�~�sx��\?�?kn\)U\�'������>�r���V�6�\u��$�YPD�	A�B���W9ae�4�O|�U��^�:_L�߳I�� K��ˎ��O�Uw�Z �� ���čMQ
l F�{[>��NMuY�)m����("�
����~"��k��Y���MoT-�)������W�kP�y�G��|�jhb\O��y��R�M~�7�c=T25Ʋod��
�@(�c(�bl<���I���¡�Oe`�!a� �&��0~1.�Ȼ� �^x��)�)�nP�}�	s���'1<1/�m�w+�5�)H4_�#�d
�;��(_�y!g��@���wx��pN�A�λ��]av�����	�2�hS��iw	x+���,�76�s�O�B��u��(M�g�p?4a!H�W\�_G��6m,۶�[�λ��3�mb���pѿ���v�|�8�,*��}���
��b��O�?����ߞv�Ev�3��o���i �$p#M�N>S�3bʂy����ӟ��8t�v���O��o��661ލ��s�p]\���z�T�{eh�U���n��׵��J��C����an1��.�A��.˒b=E�������!'B������pec���k^�':hD����P�5�%�=ER .��'�t!|��_��\�/|�δ�u�J =/{@8�t nDm8��Ĉ�׿�-�})���H��`116���B.?)�?��Ow�������b����"��\!"������'?��o}kW�L5+�M���LEH2�d^ٷ�SjӀ��¼0.��QB}���|����Ks�&��<�&�Q�{�~{��;7�fZQvdHs^g���N��K�p�g'�F)H�Յ�Y8#�S ��d����ǆ�ne��h�n �L��?�|�㡞�x�A0_���&��0¼G���ёh����u_�[o��g�$ʜt-�������������:D��<�h�>_Z������i�س�������wo���ZR�zh���V�~a�F��DȦ�T��ɒ��*t�<]h�v�i�>j{�;<;�\` ��o6�G��=�K��@t�Z��7�Ϋ^�*�w���*�A�%*VyOȑ�F�Ď�Di�H&���qe�� e��3�xS���D8D���!��nਬixaF)E�*ڗ{!���Y�� �C��<�@�#y����(�����B��W�W6\){?�a0A$<${"��#80؊~���=E�A�T?��O�{��^+^bh4�94	4��%�u����&�>�\�T��h�t\C�*����&AP&�ά�C�e>髊�@�`����s��΀�?5d����<}�ޙ[�瓋i�����?������v�3.�y��.4�hƌ���Z��f�_tG�۲�ϱw؇w�xR>��}�s͓���P�%�{�� �� ��D���N�CoP��Nx���uVe��$jB5�i^uhI�i����\��o~�C�!<"F��H�z���F�պ�a(�i���6?;e����>RN�P�s��	�-d?�������AܐH���7T#��T`	6>Ă�90�*ϒ������U$Z�	� ����1�)�"���4���B��Y9�"�����
Q�@s?��ϐ�d���B��{�~q�G?�Qυ�Drg��P�����{��!�H��)��!
��9��ClIj�X�]���ų��r�i�ar�9a�`�h*F������u��z��_�-	��2Ϭ�`42�0P�
q���_�����m�Ͽ��?��cR��kVwn"X�f��:�<�X�AVd��\J�� �V�y�~T���ce]�3�XWi�eQ�W='�j4f՛��꙱9���A��d�	O�����R��O\������K��n�9�HNJ6
B�懀�i{SW����������o8����ol
�8
�d8\��9x�"�mi�����7�CL!(%>��!=��#M�BAuVrۈ(wp/s1�:$q"D)�5�ZE�
��D��k<�k���@���* v܏���X_K���a�1	P�;c�Y8@�t�y/����ғ�E�Y5�-�*/2��nC�@�PY2�DK���Nt��%��w40�>c�Bg.y'��0�Y��~�E�+h|��4h^�	L����ݚ=�c i�B��ǟ9r��*�! a���:�C�AY�琺^�h1�s��w��?�A"~�7~�mx0`L��%�F�)�UB{\�����#f����M��'��N�6��I���I�"�r��>O��xD"/I���&U�������~[D�JQ�,�!�mE��J�ǉ|!@v�j���SL�u�!v"�����|�c�C���5%oh�$�8�X�9��Op,��1�*��sH�Ż ���x����,�i]Fb�R5�hD����^������@Ӑ�esк�/��E����|(�KP!��Ar�鏘&���i��^�W~Z�]9�i���
�VQxDI�k��\�c�b��aj�����p=�DJ��h�p%�;��jt��Ԗ��,��)���t"��V7�R��4Qf[*G!�!g�����<���c�a�s�s����5ߩ`#�I��ƽ���L����	O�����_�Q��æ����}`%?�^UL���>Tw�y��*؛^����R沴EO��/mz�p���ik�w\+��7iK����6�s!����Hlh2��2x'x4� |b��$m��8��Gʂ�+H�Z{f��:�`���,-�#y��� ��Wy�@�U�F�T9�0�a�r�4��B�=�R3�m��N0U�15*s/����+*M��҄�H�Q0ϡ��1m��	舾2F�B"%��&,�Q��#/zFz�41d���\l'$G+I]P%�����t�]�fUA`��|م1�O깕/�܈KQ�V�a�SGm<�{ͺӲ~������u�7��.ɽ���ޑ&�%��`��~�<	�Cc�ӂ>��M	�FZ�[�Q*,�?�'in������{��S�L�Üb��Z�Z�Y����\�����,I��z��m��Al�&g�!�gO��A=B�a��*C��(�=i��w|b�_ �0v�[��C��MQ��H�u!L�7��	B
T!�q��v �0R����4 ��3�:����-oY��h��5���g]B�W����p�.A��	��W�
�]�H� <����?�o��R!-b�3`���	�]f��[����L���O^6��Qqi�3��G�G�W��H?�%#��ɟ�I�����Ea_�y@;0,���3704�R�I�)�6k�=r�H�����^���ʠ�}W�����ϼ}�|�~L$K���=�ަɧ�v�yOw?�b88D�+�]f��	wj�s�6��g�䉖2�4��v�g_�m��i�^z���lP;y�}D��AF�?����L���I�-�0�I���I��,����{�����'�r!��C9�9\(���������S���6���0xB�t�E�$�*��?R5s�����+�} �G��!�Ҡ$#��H	�4���:4�s���Ic]�w�����>C����T�{�L��ES��N����n�U�A|r[Mm!*��� "#kߤ�f��@' 1�h�N{ы^�D��q��I��Aȶ³���=�D�1��Þ�d�D+�ko��-��&��{���	�j�����[��@`Ew���<����&�sS���]�ў}��8\p[Y{�,Ac���pX���h�Ae<���$�)�Ms/�w}���|�z�t&����N�2��Z�W&�7"��7������2���#�
j���1K*����q�/����>w�ҍ���f�o����򐧞&�9��呲5���a��ݞ�-�Qbu��d�4����aʁ���W�b+�'��0�Bd��!���NW�p�ͼc V&�:��Ƚ�T���+!�+	i2��M�7i6��& �5/{ُ{��/�K����9��D"f�䨨bދwRn����e<���K;����L���@��y�ޘc4i�t�w7�|��^S�"K�Y�xўpYe� ��V�P�n�&��Ǳ��C��N6��7�4�3� zu(��EQ�S�KEzt&5\�.��pv��m��aۅ1���^j�X"-ƥr�:W4i`��#���8�,� �A�R�u(!�xSc���_�i&E�=����OїZ���Ķ���V-,8,�CN+���?0�v���61J����*����r6[mXeh�#=Z0W��!�O����$:`y~�w�c+��%ɚ�a
@H��4���"�\)8x� �@���K��O���k�%sL ���X��r��; �MP��e��zJJG��i gA�!���`H�e�8;Fd�A�af�*��@3>�x�≫!^&bN41<s�ԯ�q�T�L�H�H�w��6�w@r0!k���f�5<�5��9Zo���-�
�G�O*��N��bVr�;��/ =@¿��!��5�U��Ԑ`���eƤoT͚<r��AraU�G���i�9?7��[�5�Z$���,��&�E6&�����71��Z��KsHQ1�Ԁ�w�N��\�4��Eӄ��Uׁ�MU���׏B��Y�$�b�z0@��B��b�i���F�-�t�fl�+y5k$�����m���?$��Mws�C��P�š�<����Y��Ɔ����Dh	U�H�X�6Ұ\;S��á�� �a�PA&��5�\�/��H�&pp�Va�;��&� =�@�C�\!Ykp��q��t	؂a �cc W�p���
��3n ps�*��H����0R/'EKRO��@����(݅��T:�9H�0 4$�|��(���YW���,�3<�����K��K]�����ye�06�S��-�CVnm���eײ����92� ��w�C�D@��`E�Z���4�V�Z�l4�*�B-V�Z{7��%�C���=)�]�iHJn(�Q���b� }���L{�@/�?��̘����B#]2�I�,$?lj����	��V�d
o�A`+5A� $�B�� �Ky��c���������I/a�h0B�ɓ��Q�j�l���p!��Ea੯�a4�t�Cͼ@�8�B�P1�H�|�DL��%�mAϒ7�pr��J���c�C���5���x�,$y�m��)���˚DF��cj���H�z ��a,<�Ƹa J�3n�@�8���������9t�'�PAY^���L����B���鏌��v!��k��3֒q�n�
?�Z�y��~��{�\�ϐא�ni����\���{�%�w��J%h;���fg�:׫n�o7��ɝ�';\�nS���$Vp�tzv�Ƃ����Z���H���9̛9��ʜ#����#��,F HL�Zڀ�f�����9�Ym0�r��'�+�<j" *l���o�SŽ9Dlt&�Ŕ���i������jZ��e��C��x�V~F>��}7�a���Lu5�yK|c��#H0�?1iw����34H��`��[��uO%��AG�aH��n8�*�1f�_�-e?_�P�KJ����I�$Bļ*���QZר�[,��3��He��3�+Y�=� �\AT�tǵ��+�>�LM{G��$P�lْ��!�K��Bc~�b�\��()]j�e~蟼E$}
����?0�UQ"�0�sn4.�$� �??����ĝۋ�Z�<����-��� �չ@��묭�,���I�d`rp�f݆��ꗿ2{j_� I�!`�8��k9��R4.Bb3ќ��d�Sռ�`���{f�G�ќ�a���[{��:��I��9�I�b�J�g��CF����F��<0��a���`�fa�	 {���������\�ؖ3և�Ƽ�h����?{�f�7H��M�XS�X�-7���D|�FX�E\�R%;l»M��tjD��|�N��N��4ikj�!M4i�b���I����jj��ׄN�����r��@�"�)!@Wq	�%���(��Ɯ�A��T�L=���IS4{R(?\#_��&�K�&C�[���	�2�,ͷ�M*!��6�[g��M�[�k[��0ng���:�����nrJ��sh8F�N!�=���oe��,�FsL��/�˺p���4ڏ�'R�'�'"��aR���h\��	D�'Xyuq+����˳D���W��Ը(i^�&��Y8�dAA��K���z�-h����>6���06�,��Fk�I��(mR�4Y�]<I�������֞�&	P�H�B�V1K_O�C?MN&)[D��P����B���AjH�O�����.��#@�Z�`�(I_k/��ԅ/��Dr"�i!�t�(�X�g���'iB��S��i��ԦEK������(���X��7�nh.��Rv1}���GK���k �Sg�]����:�ߞ�����/LZ����({-_�.�HZ��3����u�x �/�F|y&���H�hz|Ƴ��F�?��/�$ոE�?|MB��v�����9i�8jRW�I_����_���S�/�ik���[�x��a��3��2�B��B��$���.�"�"_�^WO=�	R�߮�g��`v�У�n�X.��P;�G0~�ż�f����Ŋ{3t�����7�I+��+C�6t��_�Մ��`��萪�ZJ�0��'�OR���Ii),�Fh�����Z ��/%������Hת����;D�b�2슩H��~�@�WذRM�=o�j�� &�k��X;�W z)Õ�"Mn���z�W�DsǵbLi��U�?��_���q9+�<�y��(N�K6>6n��l��yf$;�����ؖh���B���~���C��Ԙ�6H�b�i�.�#��g�g�|Ye�䩛}�Q�����~d��ضc�×##�~�/<�<7��ц�GiH�l;�?zj���	����\eC��9j�>b���ȑ�~�l��9g���=�<zȞ���|�6m�h�~֕��#�2	i�+Y)e��$ &�jË��0�"�b��9�d\��6�o>p{x���i}>�w�˹�<(� ���&K�6��8��_(/!N��K������P�T�m�<�f�K���a���n
��H5�� �.Hc�Y?-I�i��R�R�MR�$i��\wS5=u�L��Ik��9�qN��pa�?f#�9���I$<��w'�@Fa>���g��51�T�*¥yW_Rƥ>�{-Ո�YZ�MPRz����ƹ��J�.���K]>�V7�g�1K�;�-����5:uZeO��Yϵ�G�λ�2�Xw���C6;��e!�;^��
�B���L-�e�i�]�����3�58�����k����s\�����l�Ęu5[�9j߹�[v��~�֎#�7�ȁ��/�/�؞qųm�:k���b/��푽�����,��k�z�&��)��6W�q�.�;�l>�4��O���A;��>.��/���E
%/�p��\�����䬽����D�MN� �]�4G���#.g���(ˮ����x(8ԑ=l�tf�ds�{��o�|�0���f��E|�>Ҵ���#�b�"Rq��FUե6O�KR��G�<�h�B�4��u��_�/Ҕ\H$(��K��Yi)Ϡ����������R9+�Mڀ$s��&�$+�O�	6⹂I$aӔb��� ���������jIpW�N�R!���|�[����J����y���H̓a[���{ ��%���>i�cr<y��E۹�L��-�Çp}��8��`�4B]C�Ƙf�u���'Б'l$���h��q.0nn�a_��ce��_��b��3�+��qx!ur�l#˷��笿��s�*��>��O�5���o�T�u�u����!܁H	a�ڴ��i�z���s׹��<W8j�I��,�^�L�">��J��2�;���Zm��mނ�����unԍ�����OHvP��E��q��4�4�Ţ��;%)�9�fg�!w5<E��sK0^1=S^Tb<o+2l����;����Ѓ�
ߖd)"L���EA�~ˀ�7.�"����~� �ȷ|�!�#C�+�I�`=1 =���q�$6�+��1>b��3�m��o^��)����>o�L����5������	�AzG���uAӃ%K�h�i��3�3�^"���=��^O�G�A�/A�<Y��|�#]�N��-�N�f?���m��u�ٵ�Lв��/"���f�Uw�}����|N��p>�v����bXp_R�nX�6��V��x}�ݻ�m۟�tr�o
WG�=���5[Hw@ �ݜ1|�(	S�n��'�	~+sd/,Ե�|�E^.!}�=ca��0E}���u�~/�⣶������)��.�E#�	��I�٧��޷z=z��SY�p��ށ��@<�ʔ �CH�^�c=nsS,Y�А�R"���W� I�J�,���u#*�\?xa�Q
!�������1����<�f5�?aZ�/V2��� ��q�He�Nޖ�] i�g{��Q��w=9y�6�=y|�M����]�S@w\�O��د��hIr��@�8q%ozӛ|O����M���<�|i����q�w�=g�����졠���]�r�ssպ>r0��z���n\>s�9�o�#�|�=Y���'��N?�f��2�r���b����8a���I� X�����{��zo
�0(=�`.:v�d�=��!'`"n2���4�}"ps-�0�`�>�'�=��s��.�;$q|�\��绑�MWg!X4�#�+R�W!"���!�6�5sĿS<Y�3��P�]����w��`�0r��
��DF^?�����(jᤂ�dw�yH�Ja�A�O],ӄmJ�,����0��]��.�=�iH��M N�ϞZ��f�����r'eS2�e�9�	:_�e{��R5סCm|�~�Xs���(�C�I�x)�d�3Ns;�Ȱ��FAc��_��bm)��w�w]��z��9���g���Ja�y?ϣ#Ѱ\,��~᷂�d���*u�M�l&'<��bXu�
~hk8E���;��[�}�1�Ot�_����Q�[Bɯ$�B����`?s��h�	:IS</ۂ;��Ç�ك��t��@�5N�8!aa��!%����	���$���6��A�<Wf��8Q�[���-�Ik(��B�?��9��t�P����w�RE��P�,�ʮ�g�k�sY��V��!���Agh\��܋�QV��TZ��#��
��&�,6#��;�+�:��AG�ĖD0�]m���ޘ"�~i\u�J���hrm:m�6l���-��~܎�[Z�C���Zr.Xs��C?��:�m�v���\�p{b;�Y�Z�Y"�������:�>��KS�$�H@Nx�?��oL=�rcn�ȿv�v�8�-��f;H�%O�q�~ѓ��\�ŒQ��@-<��o��ou��J�KCB������!*¥�tzϲ-||�}�����+��E��|���/G/�����5E�Bx�f	6.��K�5��1�L��eRq���H�8��Ԡ)b+)�)H�g �@�!��I�yF*&���i�J�8�gTq$h���;c�u
xR�0�,���H{~Aw�;�Q�
B���֑����P�{i��5�N����6�.��'"?��/��~p����k����Ş����u�ξ�w<���۴%F���!������Ǻ@q�{o>h���{�j׭�����S�8����v�#!)���I����F��w����"J��+��:� ��D8�f��Co�Tq�=w��u�z�>���G�p�d�+��6�7����x�8:fa8~֯[k���7o���K�F�8V�z1�R �հ �� /��W�7>�r���� @`��$aJcL��]s��@1ȋԽkm��VµsΚ�fPU+8���2��-Rz�W(u7��`����FcG�A^;���.An�nƌZL���%Ė�����3]b+��&��|� �fL�l��́�3?s�����/^�,cQ�p
��{��Fڀ$��(\��U ���F7<+'�b������3`>Ur�4({��}��r�o�]NPx?������-��|�=���yO�V.U\3��)e�UlR��m!J���ƥ6Jҭ���3
sj��?��n}d�|~�W�ӳ UR�Qğ�E���i�mvg�����u�L�>:T.����mf�������W�ǟ��Uts	�|;�XȾl���0[A���^v�Ka���?�G����	�kQ�B�휟�)�oF�8j���~�E@U��<M d+�X�y�>ג�� H�l�~�n\�@4��~�Xx_���ᣨr����v�H�}���E�\�A�07u�٣�"0�b&�#�0>4��۶�w���a"S%������{đ��q�wv�k����`��,�0����������x�5�$E��������geQ�%�#��<ii���)��3`vc�+̃&�/5?�J� ��!M��������@a�	w�v�=D���`�����e�4�ǿ!H�!�[���"R�1�A�|�(v�2�p��}�=7*j/�-�	-���H��@���y�!���:���hI�'�e}��7��6�=�-���z�LO�ځ'{�#y��y��a	
��=��0��[�U��<B>4b+���B���x�A�ǎ�5Q�9g���89;r8�yb|�7.�g�{�My,���@_���F2Z���	۾�b����c��[��={
svȃ6{[��<i#|�U�� _�ڇ�Py�]��gن��mnv��ز�n?x�8=0���䙢��u�]yՋ|s�H,"��� j x0đM�	�x��?di1x�Æ������TPM�?}4�&�B=H9��7!D#��0�:!�kæ�c%�l�����@�k�l��aO$��Ę\-��9�Jf��a`���^Z�$ߴ@����:�%��7}�N ���b�� d;�w�G���CCX$� -�F^Z���y䅣��`�ߺ¯��n	����A+��F)�~C(0C@�
�/�q��ay.̅��YCT�O����uF��؉2YMa�J��ܰU��)b�zr-�C���E����>go�h<�a��/�@�U�����!�̟� ���P�<�g�NU�V׎]�b1��|5��#AZ�gsӁ ����
w�Q�+K��o�F�2B�Π;��+�)�N	A(c��p�Q�,F�<���)[�R�P_������oۺ+KwrȎNO�����OJ��9��߲y����/��Ns�$���vXj9��v��܀���5��l�����e��l��.xz؈�@?�X �U���۶�U�}�o�ѱxp�q�-`�&iR
�#i��?b�㏹��(V`p������!�'�?�CA�ǵ4l�|ۍH�Vؼ�J �@���ߍ, ��-w_��yA���ɼra�b����Z�x��H�lP�~`.儗�(�g��"� ����9$�)I�)���T��I�o�&8���AH���3���'��a�;�d�L��W-����@Z�����u�J&�� �E����7@��?��%Mr��~��k��� ��?����!���3�:0��"Θ ^0�MK�씌�uG�e�L�RV3/�a�d+e@U<wU����|�}����"G�ћ�^w�u��[�Rd���0ƶvݨ5֌�qT���[��� ���5�܂s�p>��͠C�3������y�u&��'��[�/����#�$�}���+���Mm�94g��k��=j��DOd�ư��watj8��h+���w��[Bɓm'<�Ԕ7}��	/�@�<O�����>������7�����U��x�Y�����-��@ H8<O�B��<3��g+��"�Lĵl$
�R:�Z���5ힻo�COl��Բf#fW���G����׾�]�<Z�T�20����Ԅq*~�"z�c	BB2�o�)/D7�Ad��H��F�5N��HT�$E��Y*j!��4Kg
�(��pPyh`���� /��#El*�k��͡
d�J����GՉ����>���9hE������"B$d� ��{�k ����_��B����a�XO�-��3�
�u0vy.)/3~��++�F�f��"L�70���Zs��G� 2����'�����=�;��,���y�� �ӷ˯x��>���֊R�ds�A����6;�̈V�W�U+�%y#{��d�>�����^��Z�����l;���W<�r+W
����gO��2���{l��=���;β��0�s66�ƾ��o���E���&�_��I[�:���Zu�֎G�M^�z�i_��F��Q鐺0����x��Ojz)l�@H<�Z�y���`S(=C��G��`q_n�]�u�ɥdU��k������ᾩ���Q�)�V5F4�[��3|�˓��≯�����UP�M�S�����T�����Vau�9)���)���q�D"T�C��	���i?��-��`R���ai��Ռ?����>�p�yS9l���i���^�g�p{�rL��F�V��)g�4D�[j[`�� %K+Ax���)�.Ps���N�����ξD�C���Ʌ�w ��H(������.���<��"s��!ӟ�Tu-���H�vl9h	��%Z�iI�?��ʖpO�3Ʒ��Q�Wݏ>��(�@8K�h�/�>�-�~#��I��<�e��W����0���w��{~���s��;�|�^b� �0g��@|��p>�v�eW��݀A��@?#���/}���_ז�P�����-�S�ֺ�폎�I���l^6�E]l�u��9;K Ҽcmn$�t\��$k>C��lⷿ����t����jc�[���o ���d�%��qVZ$�`�c65��L!+��-0���{0x��y2�h��-���k�Xz���p�qGc3C�f����Z��	���F�����!L���<@`�/�\�t_�B(���hi}U1gɨ�ajt_v�d>�V�z��`��Щ�������ijo�zB ���M�M\X3c��)����x��|x���<����%h�w �5�ɳ?��O!`���{�����+�3�:ׁ�C�!�h�q��ٻhPt��|�рphh�|�f���rb��>���_�^D�	��D�zZ�|����<p�9d��4�ݤ~���.�S�}C�!!��J���0��/p)��$���������|��a����_���-�ܵ��5�����2`Y�J|p�}#st )h5c�1���������h��:����7?_��x�v?��}�߿�v|d43�M��$��O]���N�����	���#	pPq9�GZ��_x���� y�J�ݖ���_�5,"y����A�}r�3�T6���_�MsU��[�!�܀- 	��i$�N��,��=�q8D^:H�H�ܧ���ڇ/djoJ,i�Xq��P�t�P5�����9������,����RJ����
�������b���]���d��F�	?��s�q/*���9���n�!���ј�Ӂ�	��0�o}�[�>��@�T���@$��e�<���<�Ϙ3�@��<%~|��0����m�>���o���<�,T�JB �g��Ә+�=�va\.�7��wF�^��=" բ<�A=H���Ʒ�F��uߧ}�Z��@P�]F�1v��_�_��~����(@�g�g�D}RT��cM����;�~Ͼ��[��`�w�3�y�B�A�~؞x��� ��'��rWЅ���C�?����QJb�:����&�`�>�s���\�&G�T�M��o��$d�H��ˠ�$��H�HLHe
�`��y(+d7�K�0�з�vچM6;w8�;���Tp[>���+�,y�k���^��(�'_~�����W�jw��N'���d�|���$?�Y�zQ��?�;�`��.UJJ�f���V�y?X5�1��H�iV��I+��@0ހ�0��� �!�z�_�NEf��yF��i Ҵ�r&�њ~\���\p7�̃�} n�� 8,NhG��U^�����}�<,���F̃
��{���T��Y�����_Q�i-
e>�[���
�×�I��{�5i�*��r�`�%A^*���%L]X�ny��9��zιچ����ѽ�������-�:.,�m�M�؍??�`�\���GJ�C�Ё!���M8�gl$�RΆ��8 ��R��F.�^�crk�0�'���}Z��s�V�\I��v⛷�!*`�<�l�NW"���A�'��z���| ³�9{�k_c?��{�U�q5�|!��L��Ar�4��ԋc8vQB�{�"�JC�q۸aKP'��X<&9���k�{)Q��د F�=�2��G�w�t8�O��?��/��s����{�<���v?�ֽ�E��?j\~�3��P�E?�B�^�Cب$0Ta0i���A��N{�e9)4�t�s��t�0�2�ʯ?��&��'���^{�΄xv���(+k~���p~������u׸0	��+Ulnf֦'��?�
������;��soz�y���/{�;��5���R�.����4׿`(E��9�ŰR��bR~����Zנ9CH#������,;m'�B�K]S)Y��|�����sA�:g��߸�=|:n(�sO퉖��6 GyF�0Tj�Ԣ(�Ja���c�q���ȜH{!y�sWo��`��sG:Y_�8��u�s�棞\�n#h�=+)�<�*|'<��*��R�ۖ�< ��7�������"�}�tM"@��#��
��:��Kv�X���Ar��q������"щͥ�h@jogѦ�7M!�R� B���1�~�����ʴ	�La�O����Z�]Z�\�
&�'D���P����*�U�&L����	J�z ��|8���Z�x"��5�,�f@���ۉ�	GNSU�,$z�w\f��q�N���;I�����g�����M� ~r7A>9;�{����TԆ�����B�Q��%,��[��'h��k���b��ҡ�\�RB�+t�#M�j�
ԔP�����۹��.�b��9U�}�������mQZY�EF4{���#������w��!�w`�$UEH䝣w,�:64��
�p���t�q������L���=�W�L�`؃>C� ���z`��4ߗ�+0�Ft,FDy�H2^v~���]�ΡZ+7��g�k"�\�;6����3��#��3������F��)"��n<�u�!aT��S6��
b�Y�<0"�C%gx9D^�00
�h>��3�A��Nޖ�ow��T�b�� �i5�iz"����l|�tX�u�+�=yȓK�&��z�U�.$)�Cl��[,��ڮ~�����+p>	i��5���c��=��l/q��V�'�	_`I�;�x�V��p���\}�cӶb�u��!�$�S��S��I��x$�
�Z���_�B����=�Vn2|��+����O��r0s�T��SЄl$�z��?(& R�ŝ�.>�&����&���G}�:�$L|�B�f������O��HS+MAƋ�ϻa x~!$ +��\|��/�4}�7Z� o��峂E<15C4 �ߵ���m���)%J��R1�0̑�#Vܷ�6���6b#k�ݘ�̗��A������Gr�T!�ԾM�4��*���qg���V|�O���\�rZ�4�*�*q������+xBը�3/�(�5MӪ�J�<�n�������=V��
.�P6[��s80(��
̢m�����ʃ��̻K'�+�B$�~M����J�P�Ӡ���ru��M��V�&�=-+)�1~�S�{h�N*wG(�N~i�"����Q�$d��]i!t���1�g�����!�4 ŀ�]� Oa��y���7�_���o�t���N�Ȗĉ���j��ٓ�r�������u�6�E^�q�}�8B[����p�����mG�J��jZ�+x�����m��I�5�-��޶ԋD��K���t>$]��<$$��`���\"�z�H�0Vmn��~�d'�y9:L�8E�0$r��<_I��X��c-��@�d������=���2p��VjE4��DL!�Z.�YZ��\W���ؽG�f����!u�@�U�K_W���Y�HN���i�g0FEz��k��%�IWM>LHbh��0ϐ�41e,=բg4�Z���px�N���x5k��o�38bs�i/��C	E?�H���`m�s�s�+Pp�m�A���~�	R[M;�u\M<q%�+�E�_���(:+O�]>�*�-���I�4a������?���\ j�	+H�5��0��b;��t�d/��uJ��!��k�@��-��iv	P��ޗ������.3M��p�r$"t҆�Ҽ8+51NͯR�^pt�,��ȴ&����LS�5a��GYYaH$$�xs��"%����"�a�J��E_�R�UeA��Q%2�gb'o�jQݞ���A�G$.,���P{?�z0<�H�{)����T�+0����ƂI "Ÿ�|��Śq}�d���=j�� �!w�=�1��l�_����?7�����vq�*cq8#l�\ڌT�M��$�*Ǐ2=�Z�4F`%�*� -ō�v�el�dÕ��$���F���6�U83ӳAI
?��Ē��V�9%]��%b�������@ɾ!C�r�H�#�m#WB�C��[IЋ<md3P�v�B�Xk&�Hާ<@b ����$�9�v�
`�$e��+6D����������j��N�&AFn��ߒh�Å?<b��~g �5'ؕ�׿.�x����]�/_tXO��D��|�U�����,Ы�A{���D����K���^e��TX�=y��'�9�_�è2*|;����(����cc1hfzzƯ��"
u4���`Iz��O	�
�N�`~f��w/���$��m�}��wY�Q'l�V݉?Iܦ��V��(�V��%��2�����?{|V����� �:�҂䛾��%>�)��Y�J�����vi��
^i��C��u_��O����`���=���Dwzf�/xL�.5"�܄uMZ'���=�Y�s�r%�ڹX�qdl�|U�ȉU4��n��,PP,�S���i6cpY������������Ҧݽ��w$/��^ӑD���y�7�Ʃ@�d�	O�;�)�^��C<U���g�s�:�FFǭ�P�#A�{�὞��۾��݅k��H��+zR��P4)yO�Y�������U¦��29{#��byh�3��N7챃�V]h�T�(��V�+���]iW�טSb�B9��k��Ȩz��jO��ǟ}��J7�,I<�j 6��Mw�P���oqfn��5�]��O��aÒg�`��H�7�C&c�����Od�cCn�y�[~���B�]8�k\�)��'�
���ύ����$���B��֬�Ds3s���cl20����ƀ=i���N�d-�2�	?�Ǘ�>
?;�>�xW��S�n�/��]~�v��A���K�/���4��
]����`�dt�_\�E���na�Hl�tNۢ��i[�U\�y�G�N���U����;<56���1�!5�۱�Ѡ����)��j+����S�O�w��%ҔN-O�'���Y�EϋB���Yg���m۶%�Ջ���!��9'�F'0�3�\:<kÕ	�K��+�3�,�w�K�/�}�C��L�#��!�I���{�� ��fi��3�lu�����);K��k�(4;�o���Z����j����)[����� �/��\��>�����]#l�:���h�T)Lz�"��ٺ��ڦ�6xpɸ���|%���7�t�둵��E��"�*�n�N3t���C�BP]�^l&o��ݲѱ���uWu�T�fe��"�?}ih��(<<M� ����+��jA[��O��o�|��%�L�����\��᜔����yخC�q�����G&�����\��0⮝Ĳ���l
�D��Q i�3M]�r�'�}�G�񩐓\}_��W�}dk-�"�E�!��l�zz`L[����rm$©O~�N|�?��@6D{��?a�#�dW��S;�������q�0p�g=�6>����Nد���{��'WA��{��^_�`7�s�N��_�e�5'E .}^�7�@HS���FU-@�Hi6h%*�%����s �'�-�������0���I�"���*F���T�[s����ک֧-c ���O�<V�˓�$\�-x����CONNۚ��6::�I�<-J�-����b��b������zh��>�������)�&�lg��L��5��}s8�s6��}{w{j��{���wv����3�+v�gۛ��3�����T��z����G+���2�F)}̉�m�= �nn�ff��;��O��������;�ܽ�v�=v��/�ˮx�5k��!���h�#�l�$�"������?��/�c`�t#K����]��g���v;p`�x|�MO�Y��iFEIڎ���A��p|i 2<���(�S�	JS��%���}��j����	�G�,d���o�6q��������z�*��@X�٥�=�ʕ1��j�A���Hު�Bb�����E�%����vw��l7�3?�3.����ܛ���%/y��:�L��$�i�����曾���,�p�n��[�v�z���v�}�:u���կy�}�3�q&4T����}�|;yO\���K.��Nߴ)l8q��s�MO��O�6O�7��2f����_��?8m��ɟv�<�iH�7�LyB��_�Wx`�?��?9�ă�҂TA��y�ۋPJ��߅Џ����n#;Ƭ�+[c�aL/<ݦ�o��Ҍg>̼Iq�����2�k-����ׯ_�M�G�ŵQ�g���?ӌ���_m5�S�T[�en�� ���'���ݠ�E[0'�F1�jں��v�E�:�Ǹ[,��-[�Q�
-e�(s]�`�5C,I	��N������&ug?F�׺g��/�T<+מ�C�=���vn����v�Y>�n�_��z�|�]��gYex��=w��w�9��[o?��;�ߖ�eY�� �w�9�������~sP�6�y�������q��yN�`�n���l���<����Co��%������~��=Ϸj��+H8���˗���rVϼ���#�i�U�]��:Y�x��+x7X��Wng���Ă��O���al�K��O����P����D�"����$#li�k=�T;Վ��׿��;��<���h�b.���7�5�ގiN��6��;�!Y��?����:��I����|�����{��p/��~�4�=��kҝ�|�@�����پ}{=�y�w���G\��ʗ�����}Ǩ?w׎3��;�<��;��?�C}� �E�۹ABŐK��G�c�6���[�G�]Dܻ���1�H��qr�?��+|s\p����o��B�F*öo�#�W��'�#��^|O���U2���}���X�QQgG�qQ����;X��X���y<��@L~�B���/��W���7n<� x#�g���t��RGS��ޜ�P�R��Ơ�S�Q�������)���U�:Ћ�NS���R�S��K�'_Fp�U�ߧe(�q=�+`KcS�ԗt܊9�8U4F��\i_���VAy	i���K���{�0�]1��$�-E�g�]o�]_���!M�R<���)�{����x�����FYG�N8�`���-Y��F��~���'7jYs��~ʮ��s����w<�~�g��fP����
��D֭Y�$�y��]�ن��lٲ&m�6_������7�j�-�����i���V�Pz�}c�\�R�tϯ���Ŀo�K0~��o��a��}��y��m[��������n;q!��������o��o��s�d���q�ڵ���N?ɿ��� -Tgڡ#���U2�p�dxdµ�4�9�L�D�Q�����PM�1���o�#��}���چ��tɪeL�)��C_S�_DB�S��X��mpe=��V��-ՙ[��{�oH@EXD��h]I�����ا�`s�*�w
��whR���+�9H�$���`9�+�\I�y�{�1��d��4��]j��zi�)Q!s Ƣ@4�W���[�S�I�и�GR�b�$��3�-%|-�豸�Z�1�l7ݦ�Y۰q��E���	`�;G��ƈ���6]�-����� �R���zd}���&����w�<��mXw�{��fBok.���M/�[ȕ�H�=w�m?��W{��*�Ɲ�w�b�y��v��N�d����XU�K�e�����AL�Ng)��г}�ͫ��!��0���P�|����M7�@�\��?�zB�c[t�l���=67�f��#G��<'���I7�E͉<�}�o�o~����ZǦ��m�HSɑ�BL(F�}�V{�������	�KlzpP��L*��L�k��"h�LQV��T�Y�.�g�E]��p�&���̝b,��k*ً���J��q�͈HZL��k|�Li&iD/M�O�h����x��� A�&02��5��B�T�Q��<VR/�TkH�N��1����7Xn� j@����h��5_Ms���'gё�Dl��}b�<R>SWg��᣶���m<:��5�Ǖ�
�7�%Y��esl,F��x�nإl#�?s����^�B�LL^9�8<S	���Ӏ�����`Lh8DB� p"dAspG'�"Li�R�r�'��e�(lT�c�ר7|qt�I��l��hZ,��TԴ�js�Te���{���[n����]WP���fQ�vO��g-��ZN����:��)T����(�ry��<L̉���� /$�|��y����H��d."N_qW}����Z�n��!���<� $�RB��M	�E8���ko*���I��N��4'��X�����ԝ&RK�r�W�%MC�!e
),���1�=�\��z�l�E�b�������� $'f��	��>����^�֐��]bip��A�RoTAEiiG�=e�;�:M�N~Xiv�V�]5�o���/�|�ݓR�M�W���B��ֽP{܏e���ZexT��4/���+?��#�#�c��9J���p~p�云�1��83�%�R#�Sw�6O1!M
B�u��9.��lxP��'��i�R�#�:b��G\Z����uu1HC�l�m$�[��Vk̅��݃�f�N�L ��}�s~ )��я~ԋt �����A��v�o*6�b��Z�0�9�	kRM)l�E�6O`R��3����,�v����Z���~�C�f!ց������)/�ą��`�}I׸Ѧi-B"����酂t����m��B4Io�1����N�s%�J*�4-b&��S%u����MꛘIJt�0oiM��_f�#�Ҷ`+����]�D�G�$~ER;�'�j 
*�I���<(��>�K学��Ms &�{5#����2�*�Ij[-��\��z\n�|��*�z�o3�?Vm���p���̡D���I�@/�������Jս�0���g��?�^���\;�0w����m:}K���@V����"i�7n8�?ɮ���c���K�4�{�C�	O����(�b�*�/�����a��g���a7���xҬ	� 'ok�֨�C�<b��[�T�3t�Dx��Xt<f��Q��~ac���\:TIWS��h��S��d±�y�c�
�]��6��Q�cY�T�f3��ii���`��}�K_r/ ��W��U����&�w�Pe����J�]�����T�?H��6R���C��ߒ��{H�ZYkŜ+�j�7ˈ*$�H嚛�r3����G�eҤz%��1N�2'1�h���~�.�`���UW]խ��/����uBJ�L�((�)�EED^k'����:i.S��bAz�$5�ߩ�Ͽy�~`��I���٠��-�l�t+�Dx��O�.E���ͯyJgR?��x�N;��	;p�q_?�w�w�%�������1�o}�[. ���o�׽�u��4^i���K/��|��#���5�"��g�T�u�6;�z�ӂ���iB�/��밖-ըV�Nx�?����k�,xp��]jc#�b�G��l�c�mzf���IĂ���Gm���v����!����&�j��w��~�w~� �R6��H[06� ))�F�֢�I�g�B;��KʡO������!��Q�����a�b�v���p����GV�č����
cÞ��s�׀�$127�Œ��\�P��Qaih|ǵ�G��Ԉ��#|]7���o�%�{!xz��J����E?d���r�|=�S�O�+���`v��u��������������g0~��7��>I���h(���d/�� �J|Ιgx�D���%H�h�A�i�,A]���>BK
ӉQ��@�觠4�*R�+���;�Rږ<���է�^�Do��p:��"G���O[����'�l8��k��f3��2�g��U�f\Pr�𑊯K�:���^W�o9�1����Z�?4 #����m����{�Vu�"��g:���6w���5�,�5���k��Bb'>��dtc"!ި��}�s,$��7o��[ny"0���P��DKk���?�.}Ƴl۶���1(P�߯l lr�5�4��<h���җ��Ŕ��2$��C��������=?d�F�8�p�5'���Ӟt�8�� �>�|�x"�M0n�'��D�&����F�ĀM�
��� �,�k9�h<HFƆ&�!๤��`2_�.���H��@8a��%!�-�l��!A���]|�Ů�+�"̞���w뭷v��@�!>0<�R�qE�h�It4�����A�!�`�3sG?��O/��wa8�^�>�����b#���@���x�'�42?ϔ��{��W�H柹�H�x L|Ƽ���\�#&s��A�b��ꓰ�ZJS�N�0w��&I?�S��A�EO��Ko�f���!.j�x��pK-��?g�N�jW\~i83hay�T�ߛ�eU2�ļ����3c2pb4�����e��A�0Rh�'���a��O��w��q�96_mط��M;x�q����Ex��v�%�k��,n�Z�;�;��^O�r<e^Nx�?����G������U��~����g_ye��Sv��ٶg�#{�ə�y��~#\x���áYX�S����1|��_����.���ȒhW6��5�yM�����Յ�-�����;ǼH�R!˴i��G�.�wo���^0�Xp:Q*,"� !�^�
c��"������5�saTC�s��0��I�A��������"9qX�~�p��< ��%X66`'y� ������Յhn�
qހ���?��3gR��ŕ��<�	.��ox�"am �H��ƚ2<��t\��[�������#���1?�@<��y6��y�X��w�ß�e�!в� �0�J+��z����H?���v���B�w�O�k�����ؙDj��Q�`r����=��nl0"����#�´��5�����9F�Zj�Z�	`�3`���;��EO;;G՘��J�8{��N��w�+~�5��.��מ�c&����?��.�ǚ�ߘOՕ�f�\��0`���c����]g�sٱ.���m:�p�+�a��kk�m�����H�n��˩
:��ۊg�N򖺖�0H]_���H
�2T�3w�gO��{�F٨�����t�MN(�"/!#��g>��@��90��]����)L��r�pl�E�ߴ�Pζ����*�@���ߎ�����+�(>$���VaqK��vߧ���o��*t�&O���
�8C��$^��A��;�⁔L�(BdyLAFK�ć�a <��z�R��?���l���BX����ε<��5��v��F��Y#�0DBȻ �Kpu8D���BZG��`\ya<���0��������\3��O�`2�����D��HPP�l*�Ë��H��^�җz?���Aq�����{�0�fO��y.�/���ó���jg^�/�m�� `�E����Fgh��"L��+���6�����Y�����A󥆯kP�6�`tl��ȯ7�\�/ʈ�%{��Tm�V�9?�N8t��Y�.�I^Br��������������~�;cK�N��g�3�v��}��b�]�%g���Z����O���1�+�aܴ�Ȑ=��>����j߻�6{ы^�O��G��9�g�a��c7�tC8��,I� ���w��UY�j��s?�sV��!�*�� ��QX�b�= A}��a�MR�uLK�(����V���A��s��˭��ѱ�OYA�ѹ�)o��֬�����F�5}R>s!� �8Iud����XUm�[Pb�D	�n��B�!��`y�C�3!�H�D'C����P"�qߣ���2�;#�N����!�2�)]8G:r���C��L߸��>�9�&3�0J�DzN��p�Xb���s��	�M�%�^�s�0�7�=�C������ɷ_�s�b�g<���	k�>��^<�x/ϓ��o�2��I�	�b�0��K��cXZA������vػ���;h�A�m Q�2b?���zw��w�c4�GZʾܰ!B{�G�7�}��Ky96�x��}�S��=�G^`�}�U~��:� ��e�Ұ�����/	�Ď19=h�Hē��q��A_��t0٬D����|SOL�q)��٨���Y��h2�	��|��ԧ>�Ź9���/����!X�WR�F[�7�����4f\M�b��P�e��@�[C/�\?Nl�O��6���B�|持��Ƈ�-�1C�������i�E�Q��q�H� �����ġ��sИ7��?�Y;�c�c.!�<�����!yq8a
4�H?�Fy'k!�O~+�C���x��$�2E`ƉF�{H�"��i�f �<�>\{��A���5h��E�1a'A��11�J���0*ր~ ��,	$"<�*#3sGc��H���a ����z a�AE0C��z�C�!�\#{�y&��z3_�����1�^�g���y�1��D�4��=���RD�S����΃�8;�By��]=��X7[� Ͻg?�*_'�L��g�9��=	�O�T���xff�v����n����Ӄ���Y��F�<��Y\�"��flx��t9�?��~߳�D󲯔��=;�+�y���^��9{$��#�_t�i%s�Ң
ד�&F9n���F�!��� �>�tH叾옺x}�vl??�3�67e<t�>�ߋ��ƭ�A>k�"����i-Vي��ϟ ,I���!��������!�G��F�c�:$Y5{��$�#�qCp�	`�=ćk!�ZS�!}�A�a�H��%D�y���_����� �a]Xs�v �:�4�OZ	?@9����!&̌�A�!�"���7Z��A�Ȣ%HC�9���� 0�����|���<m�Ly70�"M�^��k!��+���yd 8�Q%�A��}%+c��,����� ��|�o��~c,�V�j$�Ѱ�ܧ=���4�����4z/ۘe��y���u�].���gنM۬2<�I�b/#�gj��+:=2�| ��q��o��k{�A�!�1��)F�zMI��~�)�`����>�/0�=Q;�d���5������(�,Wm~n�\�s''��t�B��j1���/���
G��� wN��������Un_<��a�(�9_@9����u��D���kn��X��H2T��Ѣ�]�ɦ�v�7﹉���7<,�#�Qp���6z��J�Æ�@@88�D��o���Ɗ��R~��4\;-�.�7wfȔ߹����bǏ�R}����ɯ^��I��=H�rߤ��4�X;�ʡ�����s���> �L��&O��B�e`�/�[�ϣ�a�`��H��	s���p�>6�'����8`H�M��ɘ��O���y�x7��0�`5/�$�����\9�3Ew+e����@�����r>�qu��b���bzs~
���s�-�	����
�w=_�s�G;����ԟ
C��>���0/֗�����U��4'y��Cl�!ڂvkC�[���ͷ;�w;��ʼ�|v;���saP!X$r�,�c�Ĺ��&o�}���R	�$|�vb�W�h�4F�_��_�_��_w�3�� )�.�_wBɁH7��4���6:��B��!�p<���hƒ/e�7�"�|���4�q�����%��0u$�P!6V$b�{�l<gy���&�<宙F��^�S������C� ~��ȍPy��8$qy��7����lt��o���~����l<1�5�
L#�%	�@*��TiO��f>%,C"?�ٲ�X#��wA�h�B#A����G3�Y�xJK�z�4!}��ZZ�����$Qk�5W\�����8�vC[��J{��-�xK���.��ՊkQ.���z�������u2�	�ŹG�VW���cǝ�9C b_)c�������,h%��w�P���S'��-���\�K�nl��|;$�%�˝r����+��.^��|�qCG8�������A--�Ghg��)
Q��7�#p�x�B��</���p�W�Y�%Q��W��8D��`�N&DCɺn��B$0�}�E��d3(7��i~������o�I{�{�c��G����R�$u�ͽ��T���b�NAW���{�*`2��s�/��*	Sp^%�:�|�HV%HS����yz�,W;��
�V`��1�*xP�RF������� $��Rp}�s���� �Zl`�@�D��adozӛ���4��3�O����f��I{�A^\#�V�z¨�c:�2�k��'��	��0V���}���|ݫv5�5'�@����S��BA9�b�.@i�n3Ȝ�3cD�~P�.�!Q�����A]��ix
�ت7�}���2�6�n�DD*�?��So;	��V*��({����B�|'���R�ͥ�\њ5��� ����z�U8$�T�����ẇ�k���~w��˳GH���E6�.�K"�px�T�:b��W��'�nY�`�R�s���L۝�H�TAD��0p{��{�ԩ�5�D�%M��Hʥɏ;M�JҊh)���4�l*zF��&��RI�&��&`CW��O>��VD����oi�`�A��-f��c�g�)��h��]ஊt�D����ް��w�>1=��T�M��2"��U��[�-%���_o�~n��-�)�c[��3�/0�@�9����p����~��ֶ�y��M�f{�c6ng�n3˻&�7�F3��U���� cFg1O�W��񮶃���张̢0E��R��e��CY!�N���2�b!~��V��ϧ�+�\�&��Ri�Z�Z�v.&�r�' ���B&M�,Ҍ�:"N�p�5��:�{�����?l䃇��Ƀ67{ت�S���RD�$��v��5,�)d�I[K���?�%�J��Y`�TAT����q���H�H����C��xC�O�囘� �x�=���E�щܐ�	���&?�7ݣ흤�D��/4lt|��v��*hxl�S:S�	�A��k�-�BSFtN��i�i���\�f@�C����w��#��Q𿛭�f�t�
O�v�$5�jC�Q"m�W��w`�O�V��b��XʱPT*��E�)%y��3('�6-5�*�w9�Qj�l��8���x��c�Xo�@�|� �/dϴ���$��9��)#'������ϵ��q�?��=1�����sI������~���o��0��1�H�T���[;&v˵�-aM�%f�g�=�����5/�a�Uv�}�&�gl�m�7F���kڙF�g�`K5i3�UE���������vF��Eo�J	���\����^�|�[�J���d� $��m��A����S�q@�C�OE�e����� -2��S�JM�y��;���}���{S�}+��V��sso��9�����k���n�bwio�ji�I߽�_�w{��٢!(�8� ���=�y�8�Ѳiy6A�u~�l1���g������ ���o�׎?ꖂ@�y��`o��2"�ԭ�x.\y�%>c�����,b�CS�y���t(�"xMj!�C���� ��$E��ԷS���(9�QMk4�b��?�JX(��F�.��U�U�<���^z1w�d7�HǆJq�w2H�c%k4���)�.#F���2{_5�q�8/�Kl��٠�F�c.�[�,�1�[��[¿���{r��{��l��7��1�胱��-���/|ZU�jH(*-3m�F��m.mBY|��ִ�����1���w���ش���5t2W�mgƎ>�@�1����x9W��C���p�F(���K=�۟�7��(J���=J�
�5��}�m����(�!C���H��t�8��B�^o��C�l�S'-�rm��6��=�l߁63�g:�X��ke���BZMk���a�-�6�e�f .5�[/W0���؍��>�Ϊ�1KY\����l��_w��h�:��V ��*^� �8b���.*}�LF
��C0��'UX�s�=ç9㔰P:C�i6\�ѩ�C���J���{�z7kh��K�t�ދGB��&�W �e#^�R)2��Gy�i@��c����<��o?RlyY)=�S)������x��V��xtσ֜���Y��#�{�68�4
��c�`��h��9�i4�jQ�ˣO��c���֑bX� L�3zx�B.�(���p]O��f�GP�L���)�8��ӛ���pH�Y J�І���u��q�6z����\8��H���=���<?o�*�k���$ɷF�:ַ��M�ۻ�����gN�sAX�mf�4�jA1�4(1}l��u��l���^<i�A�GDe��l�m��Yrɹ��+��t�b���S��!�I+!AB_�~���X�ݳx84ۊEu#�a�U�ޖ��.x4b��ʵv�78�?¿X�� \�ctXO]�fpl�Zq����e@�H?�W�ݣC�v����ڵ��l	�DؿȔ}���:~���QF��l)�xQf�g���w�7;�9�(���[��thb����@��P/FF�o�s���դ)r��W�RC�9�R`J�y�K�q���_�u�Ycf2X'eg�t�C�+�q߾�v��;���	+v+1w8�~�3T0Js�(FEX�mW�
������� T{0;?��� d�H��9)��;;��-�'Y�m��Mv�5��=��a�y�aC�5�޼�;�o�s]O�hw��ʷ��O��Wz-P�����W��I��~R�N�_��_w&�^�9�?ˮ��*۲ꐚW ǽ�p���;wy<�{��.���ډ3�+v���x<��z�>e��,�x���꫟f/�����#�7�b��N?A�5:u�t�F��M�(`-$ �!%�L 	w^G�� �����5���^¿ ^9i���A.�?iǚs*!�m,�ȩ��SA���S�D ���}���g
R������?�`8C�sJ�¡��-���6�*�v-�5�d�<=���`��V�����1���E?�9�I�����2kU8_��ʏ����W��X%��9n�	�Xj��߲ҕ���	�ѽWE�O1(UO�ޫHOך>�����T��Y=c���2�^�:lB/�b9X�e
9�� h�M�c�a�XS�x�b"����V���&$=��/���e=c����y���ʯ��i�c��q{�w�]�4z.�����0�i/Ɯ����aՒ]v�v�,�`�o�����OkI�EO�%�Y/��/K��i5���`�o��K^�"p"�v{����o���M���~����.��R[�f�5�mgy�RH�*Q� �P<7}�o�[�3h���^+�����"^�q�	�L}&,Jf�y��۴����=웶������8
����t���Z6"H�� ��Vo�TA�f�k�8m�"�Q	c�$�T���u�W�Jx��ƙ/sRe�)ǉy�Ŝo�!���L\Li1��sD�s�񚠕4Q@<>\�^^�x~�)#Jկ���� .C�E��1�7�4����ž��(w��n�����7��Iqn4fmr�v�jC��-Y
mv;�,ve�k�f�s�&����f�n�F�4�������3�8�c�%;�԰��:���S'�ѕg
/���p���k�pf ք�si"��9j�zw(w�;lF�ú5k�&��z���Лv����W�h���u;~���DXl�w�];�ˮ�:�k79.�u�۱#G�?!�b�r
7^���|�+_��n}�m�h�������Nu,���!�=��]�a������lf�D�\:��6���OeHx���={���g��>�����݅�;�����pg���V���n�
ȕ�W�]��x*P�P`��<��g>�Y'�b�_��BO5U{C�!�̙�1�&('x:<g�X�����wZaxpD�FM�g��5r\|膁渖ok����"(�����4u1?Xo�������q쑱Q_�:?���D��A��uk�z�0�����gW@w���p�T�)�߅bֱ������ׂY�z�:[�bC�#I���Q	�:��kϟCDn��0��a�Řbm.J+�e�8��m���{���ҿ��;��!U�q�5��u7��T3�^z�S~�C��1�J)M 9��_잣�O/˟��Y*XU͸�ᡟ�:IbU�����^5j�.X�<:�z���C��׾����v���C��!��WJ��>��hr�0<(�U~�'^�^	���C_�<X)�ël��~��{�}v8,".��N�F���cq�g��i� Z�<6@���kEB��B�@���?��@3 m3��=z�K^����@�c5!�9��P(T,u���a� ��)�a�y9���պPMVd53W�)�!_�� �Ie�o���qm(+<<8͕ J��v���p��;�A^m���C`p?FǆGFI��������X�Pf����7����\8�ڱm�Si0w�k��͚R��<�_o)*��d�cࣣ+m3m��(�f���n,�,,��0$`�Ϭ���W�Q$cH-�'���>�g�� 2����e�U�ׯ%<�o�sή��
��w%�F���O}�� .��i��o{5��?���v���7����/�3X�q��:��YK��_����Um�u�o�� �&�R�88¦:v�MN�� k��M.��x����8�#*`�QYs����y
Xt�z)��u����EpO���-�u� XA?p��V0���52~���;|�#��H�r���2E��X�m'����~�y�#>���ѹO|���� ����[�l��,�Ga �x&��s%���h��q�5kW9$ǳ�y�]~�����\�q|^Ûcsc��9#����(����!���k�E����-QT\J��̱yM� mjR�|)�n��5ǽC�n���Y?NW�.��Șٱj��{	�V����q7��m��I�J��P ���{�)T9P��s^�a�7rl�F
=��]�z��q�����=��ɣ��r1��k�s�3M/���b�䄑X���������.��a��+��w�;�����/���gݶekx�-k�j�#��7^ikVӏv�ff��=�`eWmo��4� �og��+M==y�~���E�B~N�K��K�sW��)q�b.�^����j�����>�KG<b1/}��Kv1�VӨ)����'%KU�(�#�Dt&FL�����-�"����/ӿ��Ω"�p���J�yFT�JC4'������;Ne2BQ�Xxfs��~L�;׆���t���N�^���nܜ�&�0�3�=2=x�(
Un�lX�^tA @����}�QkD�+�{3J�/�>;���ZA` ,/<��銻}��6;q�S�[(D"8h���aO��ۥ#v�nŘ�O])��)���;��k�u�4g�A�¡ D��*>�z���Ԥ=��=�rŰ������#���v�G�R*ة'��ذ�B��}op^���z�g� �z�_��Rtv���XN��� �N�,����a�@fV�F.�"��v=h�a���dP#���Q�?��?�M�Pb! U ���Xo��|_��d!(K�x�Ҋ�Ƭ�*0�6�њ���ɰ ໯�p�.gt+,��l�B�yh������]X� e��������X�,�f�����P�\;K� �5&x*J�󲱸'p�K�=���~,0��g~�g\� ��g��fR������[�ͥ�s��=�v��
�d�_6=�k��g�ry���kF�?���v%����'̕��@�̵���kc.bC�U3z��2a]�X�W�s�p>�g��1pϸ/jCyn�QH	tm1�?)�<�X�_u�W ��=yb�V��|��6�L��I�pK=���l,�6/eee1�Y�@|�4s����«{��{l��Ƿ:�g�E�p����S���0�B,���W�<��̉���?�y��IY���(��̔oڑQ6����A*�U,Kl�)��iz�f#�T�u
f~����R��y�b{!��c���9;tp���}oX��66^��k���E��@YZX�۷�#C����+A܁�@F��E���k\/��DM̱���5���N"�k������:΋@�;Vp6��c']�#�Ԝ��،��^����.3s^�zE313�XPףt\^G�)~�@�o�r繂���|��Ԁ럘��������Vf���G�P&x��ȍ�qn�w��^
־�1��	؇�T�8��i�FA�5.͖w�b�;~Ć�ﱡ�UaM�[��{��k�#���S�����
��������a�������7����z`Ȩ��Ӛ���ke�(z�d��"��"�@��b,qxd��Z�"W,O�"���)��>7��l�]]Z'���Ց�)~=��K�r��[��7l��%�V��p[�l\�����?�������\y>wki^���e�?l�sAIET�3g	��E�(�"��ur�[͠h,X����u�0����H�s���j�
V��/pKA�2�
e���~b#x�pB8��`��^�ʯ�?~��杺���[�¬1W�k���.�q������#�jժ�֨ovܡAM�/Ͻ�9. 9��ب7�n4��ޭϸ�ߓ"`�dg���}��ܺ���+"$�7�.Jx��5���O~}ܓ���%�l|�F�m����k,���~�w�r|��Wlz�7���;��B���r�����(��[�9d�<Pd���/�y=�Y�v����� EI\��0/�~AJ[M���<U��0�RC��& Ȱ�qTӡX�֧��i���TťF�!���� �뾐d�p�[����xk{k�T�e��1[��v\r��׃< #���S1hɕ��q�Q�����[�?��'��\د����ۯ�����ҋ/� �����)��JT�%�@���Q�t#�X��t-�W�@3�ylx$�g�T�K���R�y���j�W�!K;���vX��9�k�{�iG�����w�k��9�U5�E����ի^�P�0ؼd!�����j+&�Q!m^64�D���>;z����e�*��$T�˖�B����Y�g(�
�m{��^
 �}bO���0	N ��և4����pN��9�Q�/֋Z�?�wP��,&yBx�2�a�s��fD�'�+X��u|�s����C9��zZ���1����J�L�5悧!aԣ4���f~��c)5��B������.�E2o5@W<F���Ҋ�MxWR�D�K��X��� ,]JR���v��z���PŸ���R�.='N�f@�3�^��sL\����(���8y�{�T��'�Z�S��k�(_������B��~Ϟ=�'�'��׼�[���-o�,Ω&���W=ﱆQԫ׭��bSӳN�7^̮ەV���ȕ�e���Q8ݵ�Ϡ�Wp��b�7��W<88����_���pݵޡ�۞���C�e0n���uހ�߰2<Ԫ�;p̨�A����K��y���wz0\�\v�BXW]s�o~`m�٬� kyfz������f��m��a;9=���iD��r\� y�r!�+�y��~C}dU��o>?���`�"�����`��]�U5C�H�_�zsU>#��&���yO�T`�X��6���P�����>|�M�5�y��F癨Z�g�޳�_躽7l�M�1���|�P��96�������ؐȫ�[V����^�PR�Zi�8	"Yв��B�@SN��	�*ӊg�ȩ��e��U�:w���ɭ~>j�����c����W�Y�4΁�H�H%& v
���DY�z���H�W�4��eu7s��\�X뭬��@'�?��'&��|���.�](؀��2��=i�&gmhxܠsvt!�Y���7���}�+�؁�/��灂�"Y\��H���"�L�.9�Ë}߽��ϼ���Y�x�6����AV��]87���[��E���s��n8>�?b�T{F�Ӽ��O+6�!��bx������+e�ґ�>�屑!۾m��_����:x�<�a����CA��=�U���BV�������.�!m��K/w�W����&vh&\#�3B�F�@{�	��`8/�
�C	�0�xE;Q����3�u)F�2�\�36PP0�	e�<H��~��x<���o|�=���Z�(pu��N �{� g(�����q��|�����/��9��F�=�<o�d�[�� 歴����=���=�뮻|=)�V7K�˛J!��}Rn����LxJI�8��RPEw
󤰍��������+�,a��+���-��!�+� �=X{����_�����a��iZ,�g�'�{�}�^����~�����R%�ͺ-�o���@x���<P��Y�����u�:�sb �Y�x��o��M�k��|l�~�k����4�A�tl�m�y�%���M604hS�s����B����g��_  �f��j���ȋ�O|���[���m�~�w�yd�^۵�A����+H���˞f�_y�]|�����qc�k��h��_�W��y�L��E/z���%
�C8h#�z�ڂ�ynz�>��OZs��!-��1����5@�<������`��]R��+��źP���z�k_���?����� <�������T4 
�J�K"P�%������Cyb�*�&�0L���tL�/�D����gȖa�!Xو(���o��m����i��{,8Rq�\?��?�0X.�h2}ڲ�Q"�x���.8���T�F�=YK(���7��9���7�1���^ )��e��%lH��f@�Eֵ�q�P��iuu<y6�w�
l�C�N���dm��.VZg2���{ �y-���?6e*���ݳ��{����A91��-/_�6+mbr�ceP����;mF�����'�vvO)Q�C��d�Gq���+5`X7�x}�C�֭�b���>��]-W|Τ��_�=�����z�&��a����g��q�q��~�
ݚ o?˹F�>��Ϻ۲��`��ƛnJ�{��~��`�+׬���.�e�"��E� ���ᘈ�������rx��a��Y�A!�$��<��wx�w�=_����`��:�!�(�u>zl6���rh!�Se/n��>�-/�1/��Qn=�M��MДkG���6���Kγ 12�E�	�b3pl�G�V$���*����̅{I�%n/
��3��=�H���B/�����;��fnT�FOf��/ރ�Ұ�����`����VQYH̓�^k�B����O��	b�S��Ҩ�F��'� ������[ǂ�u,>�='�h�S���1�*W	qF��W,@�[�B0����Q�<C�-o�����[���ӟc��1[�r؊����ʞ�I�;�=�5�6���yn��K�o�} yld��R*�'�w�?\�!��M�X^ׅ����FQ�$���Xx��֯�U�/��n��[w��?u��2��o��6m���0�w���ѻ?����+�Y/��ֻ�;�T1p��`�~d��ٟ��^��Av���k�k���HŬ�:��X�ln�VA$
�)��`RV�\������tK�E��������w(
B����Y�Oz��T�f.;,�/��S�V_�e1  ��IDAT�9�N[ذ�������
��=��3�&�
��,|\�T����@�\#�8��1Ҥl�(�
!���Ȇ�ް�8BOE���Gys��e�f�R�����h�3�g��E�rI1rY�\�,e:�����~l��!�Y#|��B��s=��ǣ��Ul�$DdK(J Kp��K(+� ����
�+���4{DB\i��e����|����$#�y�K橸�2�4o�)-EvU���n�Ev��WS�y��V���gf���[��+lj���1�|h�X��O*���tO=#�򛜎�is�>g�췗������~��z�Z^EVpr�{�����^��^�5<�<X�+l�E�mnfֳ�FG��.�+~�#=�ȁJ����9w�8v{��O����N�� C@��Y��@,�w������n��6�,V�ɐi�,��Y��>v�G\`i��0��@����q���Y��=�x�;��X��%J�%1#E5(�JǙ;K���
E�}
��_��]gb�D��oȃA�2#�	sF���#\�����pl�9� �V�ŀ�&�{bGDx��;���?`"e�7/�����: ��6B�\z} JE�[�����r~�q)���
��X��^��;�c.̕�t���qߠd�C�,��3PSp���|��ZB9W�U�Pe�p-|�����P�fjy���R8U��"0�#�B� ��#��*��uy|(��� ���y���k�xf\� ��?�A���c����8Ć���}�T����U�"��{h�f�Vۋ�ʵj�������E��@V�u(F���5�������]D�X�y�S�[����g]��-��]���62dM0̠�����=�v��G?l����3�ckiI����6��ހ0�&�ed�<�QK����}&XjP ಣP�G�G�Gz8,��f'���k�"E� ��q6�d� (X<��ۿ���i^�R4�u]YMMUm��	+���κ���wߧ��r�c}���c�C�{���@8^x�_��}�V�QH�D��9�"�6 �S6,��������TF�
������
G�1�!����B �>�dc"�`׽��r.�P%�|�7�e����>��7��
�p�@ �!�U�P�?�˵s������b`�PM0W��'k=%����d�=��FW�X�y��,U/�kn��V��ز ���Ǽ喙0�geYO���{)���=��e8ʑs��Pp
��.�4뽖Ѧ��R������_p��l����ɪ����2͍���)��[#��s��ǗŶ�@��Ś�B�}S0&/��J�X�������͠+ŮD�r��q�����,�L7���k����` pe�{�.?PQ�9�5 ^Љ�]j���
��?�!�{��͌�˩�x��	�]�ͷ4,��dq��45�ZeC�`�������/����O��
,�3�����Mn�⡽�>,�^�V+�>��.w���-.��5d5���E�@pE���:x�+_��닻�)k��]@����`T������T����l~��jV̣��:J���	kW�+c�%��W��7�r�����ͼ��:O5D�U�&�e{`щ���'�'�G��֑��T�(�+����\���&����J�w�f�Q���hrr�_S�XP�j�Ny�"!�'�|��"x]�(3k���W�*2���L��u�
��B��_R؉������kG	����5����J��u�&[�vC�C���F�f��2Z�ڡ����=�p�IH�0եp�����T�Ǌ��=���S�>�;*ume�Vx
"����no̿�]�'�]�5�e��Q24�7>ZT��B:5�� �X>���M�<��M�Wit���k��`�u�b�F�����Nc�n����pz:����H�Q�
T
���B~��2L�`����� ,��?P,@-Ef�Nf�7i����g�0r�<�ShcJ��hKA;s�ֲ�����"!��+y��z������*|�^H8����dR�^�J�F���q}�#c�-%����*^W� �3�,87�e��=��o{�E2�����`�c�
�K��p������\熍�eW\�ﱽ��t���=�����u�����f)�<�/$,��"�U��i��vs>�薧}�+
�#�?I���_z�Vw�����g�#>\��Aq�U��ǟW�]�٨��+k�_?���Ŝ��=�=8������xj���6gJ�Y/����q�t�eeҼ��n{�MۚO�K����nXWX���z˒����K�Y
��z&+����)g�B��Uv`��� )�>�8�AX0X&���gr\�,P M�N,<�U���lp,HÁ8��9��8J`#ă/���p��b�*$��=T�
�HlŋUJ��x��z���,�� ��9�I<�(���x�9�+׎@d���/!�g�G���cP2 �Rذ�|�����ٟn���z3��7� W�UB!�V��WU��2uXlz�9�Ph����
v#��\|����s.����꠆ף �<�����j�9ǥ�u%��5_���+��ݏů�n�#��9�ei�Sa�<��=�z�Iߠ{h4;q��b@5镲 ��t���)���?�'�5�<P*ts�گ��BLKu�"�X��sc������_�a�g�-�j>�E̕@K$K����<�����))��=<,R9��~�^���yF�K��#�û�M-gF�5�"��W���^2��,�Y�W�&��{�U׸ %�K�
��I�;���{�\���Gq�7	���0J�+��Pmx����;��L}�
����h��LP4�B���rl�N)�B��CJ�� ��9�
����5��X�j�5�f�w������,���

�`�ū̚�j5� ����x���� +J���2�!��0�W������7����1�N!�̑�@�F�P�iL(BYJ�-o.b�B�F%��'���y�*�z�b&��B���S
�̯����ql���(ԭ�l)�<���B���VF���4+�LZh���U���`�n�/�p��m��gPP����c�I9) �,��^@�s�e�� �2x�E�����F����������p.\�au<_�=���l�ѱ�3x�:E6E�S������M�/]kl�"��d��ĺEp��!���۵k����w |�4W�늴J,o�K�t	*	8��c����y+�4B����_A��H�D��u��7��F�� w�X�j��2R�s�-�5s�(3���ÛA90v*��!�D_�y�����+~e�(@�5�I��$P|�&�7����hE�Y*�|xA�?���\��E��d��� �h�����Y����\}��2���,.%υg�ץ���'��f��ĜQ�<_M
�i��"�no/6�]=����Bs�p�C��U[�:�̍���9O���Պ�n�� �<G}L����5������T�d���h:��E���0�b�9Z���?�������9��3Y8< ϭ.ƻ�ng<&����Sˀ�|`2D�'#b3w��  �c�%�=�J�;q���}Ȏ���
V!V6OS��-�O'��S�TQ*X �4�a����Z�H�!@����4]EFlz�� .}>�1�TʒM�<��s?e2�F�qQ8X�X� U_^��\�x�;�ax��L
#�J-�\��5�=�X�y`=��B��� �a>QAY�YLɬ vz�h�z�:Jc�+u%���c�O��&��5 'I!��<A�xR�>���m�>�_1Y�xO�o�פ�Vz��I�H��!�J=���N^���w~�b�b[�Jl{X�1��	*����.�r�_#�V#��Y+-��n�'U���Ih����x@�qnJՍ��R��]�օ�g":����3�.�g���������6`NY�-��}ou������W�7��).o_�5�$ L���m��p
k����c�lr☍��j�#�2�}��+͔�gyZ�!��<�����o�'m���%s�_�`�>��Kإ�����"l��:�G>x@-�!�!�KU���e��"�
���!��+���%��2��`05������ �X����=�n]*fJy��kd�xR^�zRПav����L��!��)K���K��Q��k(t�T����������ͣ�"�w���3n�նl�(�����~�a]�ךd.ɂ-'�l)*��g��]����������9���٨ (ҀX�N��)���nVx�S;Ik�">ǉ��{[��	߲��4��h�W$ռ�Q�h�~�w�x�2:a^�v�;�6�E��_7�s�ȫ7��r2��S4[u��|�U�q����NA�,�>���i��$�ѣlwb�03�T��5����A,���p^]y�l"��XlY}���V�v��c��J){Eo!,�f�b���=��٘�e���@�|A#�a�#���������6� �p=�{ѵ�]V
!&]τ�c}�#OP% FL= ��e ����Е)�Fձh��|�ǀ@�~S? U��ൠ����|AF���I� �@m�><M���L�Ac��&hG�>ץ�]�,�@x��s��f�(0�BF��f)\���0�fI	��N��Z�����ܴ�����~�ɩS.\f��5W*�zZ\�
p]k��n��sn���W��� H=)6�Ou�4%��$:����t�3���m;?W̕+�
��O���^~���-W�P%�ً��'B
u����=/�?35�ߋf���������-��{����F*��-pE�9wP&���t�)���9�X���x}��۹<
���k9�D������4#L.ndi�ܞ�8�F�"��z-���*���)>����^B?��+=u=a=zd"X�E��� h�5�A67\�z��Y(s��7�6�(��SgScR��,0	8��.X��M������0{捀U����P�g�����d���je� ���̊���s`�@7���~���>�<��96��<,w	@��T�)m����A�)�ϛ���R�����86�'�+�WZ�80��ԪR9�R�R��$,w\�.*�ytM�:��w���o�-�̇�������yC�c)���3�"D�\�=�}��
�����kIXCs����y�
r�6@���	�[z�L��,jf6x/��%��9/جt�г٘�}�w�Z����>׾��1sϫ���(dJv�R��f����7F�e�s��'O�c���#p���-,h��N	�c��Z�:�?����oΝ��;W����nӘ��3\���2F�%�.h��\�^5k�*?l�Us>t����e' א�'�[A1Ǣ�D��t�?�͖��x��a�
�xF�\*����U6[��M����d����[x��s��s!��p�4��5��'Rl�G*]/~�	�� �W.�R�<�e�I��}��bl�����	���X��A�my���,�f��EX����+�y�0�����S�B�_P����B']_��jϿ����#s/4[+��S�H�&��p&q��<#�%�;�����{�>	x���(���Δ���bAZ��պ��y;�W�$u��IኧI�N�������&[����{eͶ���q���M���N�\��{-(�L�1�b�i�펧���?<<j/{ɋ=A ��b^�������9J��^�g+�@c@"W)Ÿ��̔{Jp�7W� �9o�ĺ���q��Ɏ�_��������j�@�}����y�V�:d�@�w���BD
,|Y<
���O�X�T����,#B�-�������Q;z���;�E,�V3α)�FƖ�l�aC���A��#�U��֏Z��+g�4�X�??�@6�|^�b?�-A.�T�\�Y��LBL�.���\��#!�znj|�"2e�nR�+��\%����ϊHB_�A�H��o	���ы����(��*�!~bg�Nn�ׯ3:����J��/IC�&	e�-`.>����{)/����o�)����Z�B�����C«�d6q^���`z&�D�.�
G�NJM�a^��V�z�s���a��lnf�s����䐞��[6�Үw>���g�
8Oɔ��o�s��L��=�g؋^�b{�[���.�w���5���ZԞQЛ�B�əY?���k���$��Q��r�a�}�p��Y�7�Yz���P��*@���ew�U�r�j�`�\*n��_�����S�G��6��Y��cA�o	Yy(8����`�B�~�{�ч�e0����Y�B��g��{��y�a���K���w=#������x��k .Y^�Aۮs�p�'ON���H�јuET(�l�ju �{�s�*�X���l����`���BX,�
�!��Ț!HŻ�e0J����}�;((6��Ș����ȣG�g��M��S��>�h���e������ �v>����j�=�� �)z�(ޗ!�w9���k���0T`W0�`��������e M��DU8���9��;#��s��/���ۻ�ֆ�T��D�c�i�P�C��p��GF�TfAn����3J���V��@,�����n���Ea���Zv�����M�=�r������}ͮw�r��(��|o�˷9��1Q�P�P�� /�����(C��L�FO(���O:/��7���8
��# �Y�G���|���E1{	:���3��H�8G{�v�0$(����Lx#t�կr��a�V9��Lh�Ć��sa��'�&lU֭�>YK��L)�rs, �@�.)�i�2��j����@�.��V�;l��I���]1��`�ݒ�x��>+@�L���K.��5(���ov�"�2H�)��9�k+%S|/d�|�w=��X7��ʓ�(�����$%��$0xj��UK��%?�E�%@�(YJl.��$��&'<o�2!���,|^�:���%e �;�Y�E��?�"��^�qI]�>�*��<H�Խ��|��� �h,t�di�����}�(��	]�&�&����1��{��E�0_�����U����K+Wr1���mr_�kN3�� �'*ϰV�\�$�/������^h��2������9gqu�C���(���LLĊhkG�\����K�-˖۝/{�C��aR��c]��e[�f��ر�>����������A�]��ȓg���7�ǣ�x��٫^���za�fc�EK~ �~tt�Ɨ��-�0�*h)��1ɒa����E"�EJ0T<X�l`�}ua�9=.���W�,�bݩ��S,�4����\}*K�+�5C;�6��aS�ؘ󕅧�m��s��J[��2�2��AKZ%�A��M�~�(ā��E`Rp%:,Yb(A,"�K�'J!M@�cq.�T�у���TL�� �Q�(-�[j.�0`ŒWz(���Qr=	�r�Xn;�����,f��=�؍�B1�bD0���W�<�j�@��z�����
e�\"�	�4՘!�ε��P�j�.��X�֋��GZ4���j�Y����/��/�ڱ����x���;�d��������f��1���Pg��;'�,�P
JmOi6��4��i�}�I�+*��h�N۝�M5:��S�s}���� 2SN�Y�O�Ӏ��oϞ��>f�)���W����ړ�K�-�hX�ϸ�&�pi�hjjjL*/,c��j��9�U�8���)oϪ��Of���!�E�f�*�>Y�j�����{Ͻ���v�����Y	s%<��o����&o�c�E�1�"����&��g�gsܛ�A
".$.6��Rz�F��U���r��E]O#]�|u��5fO:��C>�*yJ�Sp׶P�Խ��W!��(�兒�|���UW�k���9#�j,N&V1����w�6%��M"J�h=E�%��EѢ8�.
��x��PЏ���pN	p6$B%�����h��$� ��s�������>���{'��MLsn��(R>U��w�f��1�dF�b�z?�M��:@��ޑ�z���2\R�����Q TEE��S�Y���KR�1��3KV�iv�Y�C�K��7J�NuY�:��KMg0�����H�����'ҘA�{�&&�����%S��$��
{�ہ�o���.'W�+|��J���
t�{�A��zXC����x���opo�����"��P��g�S�K���v��kS����#�/���o�kxN9Lz�u�������{1zX���G2���n��}��;ۇ����A�_v��v��O3x�[A�۳���_m��a۸�r�T���%���gϼ�v��W��@`�R8��J��(��Y lr�����l����-�4�s��-($kl��m�z�f��>n���¼���:O��w=��sY������a(���a�b�"���" �0X�@���{jW�k�@�3 -�{�E� ĺ>�7�e���`�J�?c�ca�T�~���Y���&eǨ��������� #��|�NA+\�j�9�h�sǺOy]t�P�<s ��84\B^V"
����?��� ���	�WN����ZZ���k�Z�>(k��9?���Ȩ��f1��S�ǳz��_�`���ՙN1
]�e/��4;Ią�����1�`���}���U[j��>Z���(���6ۚ���_a����C#nu:��V�I�����E��� ��w|��W�Ws
�=q��N[�ض��v�׾���
�t]�+"�i�БÏ����{�9w|��_����M7�b��~�ב`�T������/�����ٺ����M=����o�@�����8h�.wpjj�N��6�χ>�A�x�� A��sYQ�Q����	k���X�i%c�٢�z���b� ��Ҵ�e�e�k�7��2�x��0��sb���u��ӿ���֪Rf����Y����9?�!�U�L,{�9���_��s�4V5�� �ʔ��ō%����gs!D(�����a�X��<���]'X����y!��c�i����!��(&��uE�9�r�y�¶96�F��>����R��+HY7�(�aH�������7bJ��!�eaQ2�0Pe�}�e��:���a�k6����&\��;����2���dw���\�,y"��bAٙ�Ӫ�Փ^
���\;�|ݰ��s-��+�A��|{��[-��kT�chx�"kUƑ�Rd݋J�xz~$LM�8a�����o���p)��:�@��������W�x�����pҳ�%���i�w#�Y����T��˯��Ղ=���v�U��E�օM��Iϝ7?��u}:��e;����?�^���������\$d��ԉ��#�x�q�Aq�����¢��y�>z$w����}��[KV*EXyzZ1rxƍ���Ѕ3������rJGeQSEK�
x��d�ј�t��",��jD@#0�,BP]�Ԏ+�{�o6B��`�# �Q	�b)��S?�S���"WC!a�� Q��&���?ޘ�����X|�g̃2�k!��5���� ���>q� "`%�2c�\�ϱ��|��5A#d�p���)��Y��SS��+�eq�1�Tx:�JMv7/��%��En��o��1x�z�|�9I!�90g>#8�g�{|�S��g\����B���9e�Ⱥ��`<��G!YۋX=S�G���Z�زѱX���oY�V��`q#�wQ�ԝa���>��v������*������/��/�JC�!�x�x��`կ�fk¦�&���.yOP���<�^��o���*a��\����zљX���^����?4<�س;�s��:d�`={�CC1`Y���Z)z��MDe=��c�n8�?�s?�.?��B���~��XlJӫs:�?��n����O�KZ�d����U31y���3J�
�T%��$��9"�����H&����c(e���0 ���AEW|Ndp|����P 
�i��5`�r<��#�M-�2��=W�.�����w�����( )60J���#^�Uv�@H�(M�8�l�(�h="�Sȱz�S�[�4z�tXk�����=I�r/�)�9�p�0#J� �o��o��������yQ<�Ng��k����_��1GY�o{����\?�Hyf��{�r�5xq�K0���<	�`�s���y�y�]�(1=9�$
��cC�A@�O�G�@Φ�A9�xm@ ����܌�{NOO���
+Vm��q�dDF1#O�n+#v�gdU�&����1o���|��Wݐ�6�}�q�;d{v�
��B��jՠ���(�:k����{����r�3=^�^�:�}�b8Od����zc�1�]8��kqC� ��ix�O'X+v<ȄU_�2UySS'�����0p<��(����TH� p�����1�(-.�⧥�5�_D@O���ܢ'C���R�Y<cˣjV�> �P�i��;q���o橬���4�F�^}��2E8���%�l�3���6m�����íJQ-fq��`�����)}!��CmJa����b��+���ڎg�}q�W��ann&ǳ!��ξ[�J�;,L�x����q�V$�	]�=�ɿ�ï���9��������y�A���=�;�U�R�+k5-��9���y"��b�f�i�0w<�>���|�Z��
k��Z�
n�[����0��۰�yF#c'�@��ŋ뱩{��J 7�2���pY���`y _w�e����ed)u��g4X��@�4O�si��SB��g��r���}7<����~-v��n��
�X�[���!k7c~8<�Q`�S6��i�k�"��[��X�0KY�(�#p:0oa����h�BL@D��|���\�N��"���`���	�F��h6�R��4��[:��7�*V��)+9�#��kVPQx����̊"A
D�CA��V�Q�@�nZѫ�p\�V�'������[]��-*�Z̬�
`���ôЌ����֐�"�b)l^�󋋲Ty�Z~�P�������R�(�9?����MF��5�y��&���-�����P�����Z�x)�/J઒5-@C��$kIy���=�	����ow8�,1�jyF2���b(Z��w�M�ܵ���}�㠪�j�Ra��,8�?���G�v�X��Gl��N��iv3�:ˈ��N砤����l6x.@�p�?Yh��T��5�����+�jPp혵�=�v�Ѻ��1�Í��P��r�Ki�)�G/��y��!��y���d����A���j<�bL�D�V��)
5���c�P�	$�xpP
��	:;�!qq	b��>��M�⽲p�������c;�՜
�aN���i`�x;�zv���]xͲ&�=�(�S��`u;'��~	�Џ,e�H��yT ���:�\|5�Q��
�Dɠ@eJ��V�J���_/�%��*���)%�YB[��g�yu:?�PE����=�L�e��6���C�{!������ҌyaĚ�b�I����Q�T=�Y�7��ҕE�̓��	?��c����x�<��=R��A��ʘ�:ԁ}����K���"����}V��<�F�!�9� ��e��8Vu����X��O���m�v�� �n��w�\�Gcü���±�v���/5�W}�x��5���� ���(v+�2��ky�������v�8����������)���[zo�¿'m�,@��b��kæ>f�\|�ՃU276aa�jU�
�j��D����h�pW5��R�X,l򾱪�_���zVi�X��nq��M!���`��)=�}��F9�@m�f&OXi .��/D��Sh��螮�E��@#���|QG�k�*S�*�,��զ�q*�9����ɛ,e��m��;�D������"v���)��M+��{A*���'˞���NQ�oR����b���GE��x_�E�:X/BP�|GN�R'SG�S�'�R�j1NDy��!6J֯��xMp�FZI���EV����hR7�Eʇ���}5�)��ސ��Q
�7<%��p]��ĝ�_ۧ[���Y��X��	����7u��k)V���O>Go\�)�궜W+�Y���;_~��Q�"xU2��A�P��z����X�p�I�8yȦf��h<{otl�O�ѵ�[���=��9���h ���@����R���/��pn�G�n���%��+�28d;.}��~t��{�q�/�ff	tl,l�Ma��p�[�v�?��Nz[F���f�0�ʀß�?15i>������ٙ\�a�PQ.4��m"��o|�]WT�2�,�Y�p.Ulr�aA&��ȐMM#`��מ�b�i�}1�SV�E�()V'㪱{,,Zܩ[.8F�E��+�@l��(�=J3��L��������"}F�KiR�Bp�vJ��ІO��H	�t^��8H�C
�A�Y-R0e����|�@�E��\1�w�	
c�W�R���~��`������`�y���2�39硃G쑇w�.���*e{�?~�cSk���H�կD�Gw���"{��̯����mϣ��z���|�n?)��������>�1���
�5V������e�:�������O�/,:�w@>��OL7��)�mv�m��T-�{�1��I;r��a����t�^�5��K-���$7zPTp���C�R经��e�����=�����<[�9���m�}K_�re��d�uY�-7�Ɩ�&���m������&�����1[j�K9��˟�\$C�v�؃>ܫ�A��-��ԜW��߻/X���۾u�W���;qrʭ%pU Ua]���X�XTy�)���"J3:XLT�����qZi�܂�:2��`�dn}7X1mk461�p� ()�V\�7����J����к�BM��x�J�����R:x���/O3�FA��6+E(+���N{3��oY��W^�g_��)�df���*�:��C�Ǩb7e�1��
 ާr�c��CV��`-f<[ɕg�6�
�Յ���k��u?~�F�3�{ ���Η���V��}�/�ۺ�B�Fl��v�ȉȔ�U�
B\�v���b�����dT�Ѷz�ӥ�LƐ|����>�����F�e��I����^���UNi;kW<�Z_fG�ǵ�v���~�F���9�m�sX4XV�?�a����A��X_4W%��q�I{##hn&�2�����߽�A�������
��@���:	�em,�����^�:aِ���??��C^��7�´]tA��k�� �`�S�@l	�
�C��7��qA���H���(�B�ě���<(�{��R��|d8(� ؏��a���SRb>Jc�����?��n��\8�(�J�U,E����<�y�.���LA�³�÷�>���r*���&�0��۶^l/���Ju�9���q!��Zf#m�?�On�(���`�K�*V��T����v�R�g|��mlt�6l����똚8�{��ͷ\���ꫮ���"�C�'���͹3b�\j��¿k}�8*�&����{��?������k~��ʾ�m��w\7`��G����#I�t�����
���l��A,86A$gY,-|DiZ.k�J��yN�<<6��I���U���������d=kA	�J��XP�Ƿn��XZ�J��uKД�F ��k��De�G, /��18<�4&R��_�k��)�f1l��L 7͒b�Aq�7���]r��8��ķ����e�(��Q�U��K�}%�Pu 1!Ȩ�`�/:<K/��m[!^�f$�9d�ʒ�1��_���;�3]��& �Eߨ��}�?�Ǐ����g��Ipu)��`OWka�+3G�nt��k��=����l�5�7��-+�ݬ{.�<>OL��ۯ�{������Ïtء����=g;y������I�G�9�!;v�����ĭ(.鞠/��%C�u�����ұJ6��4��[�5�UF*x+/X�,�i��a(ȉ%��R
�-����*2�_�5kW�f&X)��
��9�aSԃ��n�*�����Tc7�蚗=��������4&� �A�PP��5(jkՙ`m�D��&댵�\�X�.��F��J�e}��N�=�¿�c���0K$�TZ#�t�K�{Zl��S\p^uv����d�n5�Q�r�@��g�'K�Y�1̼�pMk���.��r�`���Vm�ӵe�c����50�}�@'=/�����S��?�u.1>��G��j��P�4sQ��I��f� >���ڱ#��Ѓ��[c��68�6"�Yg������{����X���=����Y/��^��0{��ĉS���7�Nǃٺu�kjR�H�"O��*�͡^���ȌtNh�y��M#r~�|Xboy�[���H�� �U��1���
k��M�)<�x|��a�u��bFbN I��,�X�|~|���.@�X���0������ e@!$ș'��
�2߅v +{.��9>� ���M9\T_����W�@V�����C���J�5-�c@l((�c�߷϶���^�ĩ���^��AI�'�
H12*��^ĐY�V�����=�����͆�K�[τx=x�����F�!�c�p�����s��/X�6OTP]C��J�#����z��:�@���l٘�L����p�=�e���C�r�������l'�~E^1x��ȐkV�W�?��a�~���9�m�k9g?��MF&@ڶN�����]'+@�N,!�m���)�,k��+ћ8�ųe�6�eu(��G���7i����N�5�_*���`�Ȳmx����J/L�۰�y~�|e�Ɉm�u�Ќ�M��^N��6��5mө5�{� A^�q�7�<^���C�����\����<&�@��7�f� ��@)��0g�S�
���O�U��b���=�sq�*�3{�{1���"ݼ���k�>lr[��0s�T����g�Ůt1[�*�B�p�{�3���&v"��稩�~p���磔g�~�����>�E�r0�����h�2yj��aϊ|p`8��`?�8<��
�sS���Mr�dYɺa�@[1�փ���j���E�r�������1��Qx��%� iǔ�*��HpG�l��6���w�c{}�S0�cp�K�c;�J&L:9���4����k��a��!V�z�:�8���EN�ų�b��HM��5�����Kҁ��-9�T���lԱ����w��e�h�^_�җz���80�x�"���5��]�g
Ͳ�T�+Д���u�*�4�3����C���H�lWk��y�[�nS��P��b�K��xz�Vu��<n���*�p��u���T:��xN�� �r�ʼ�T���^�y�{�{�.�(��^�w�N�)^)|�Yz ���P'��[���%#�F�sb&-�/fe�N�fy�_�b(o�EΆ�J�5p~�a��}U*8'�PV���uc.|�+5��+�A[�b�M�<n3��
�����T��F����ٯ���K�D8 �`�KR����T ȿE�&����`����վ��3��,��CL@5(	������{�;�5���u�`�°��\`�:7�Tf�F��\�I�~+�o��H��b�9{�A�_�i��[���!�2�T�����#�S/GM
�R�c���m�2h'��AM�u�����}�7�tP��*�3��ꭺ����n�"M&sJɤ���(�L�������}V�>ޅ��� o��B�4�Rʷ��B�"��&�%�M��w�����:�H���q&&��Z
Mͳ�x���݂c��^��ѷ3�g�V�^^�Ƿr�/Y���
_�W�g��r��_�,�aQD �U�+�Y���`}i
�x�u���f�ȏ��.<Y2�87q+���y>G�&s��L�}Z����������x-�̤>~�K�8���ڧ��e���]�:Ԥ�R(+A��	�P
���v�N�H!�L��lN�c�O��{:7= D�!�������E�O���7��_8�D����WK6O��0����yZ}��7��]b8S��X@,l�XNlB�(cH�/�>�g�8�ڝ�X���d��˙k�ͨ4��Ջ�Ƿ|�x1��@(L��Z-�9.�X΂!����W��pf	
�S,��ǎ�m����>���ń��k�����W�5}z�}�Mp��H��~��6^A ��@U��b�]�X��&p>C!��Q'/)��A,�Ua�|�T�(/��N%bX7p;�X��r�t��WD*Z�V��ͨ�ݓ�#6T�g�gڍ�^,+R�g�z��ݷ�H���߽UZּ%�P����t�z�_xB����|"i�����v��t*	_̕�,
����S�8��#v�P,D#�'6���I2O<�y
�,��<��m=�U#��ֿX31��h� B@�����x"|�|��e�� %��Y�+_��(��k�@���Y�{<a��+6!��6�|��VsQ@$�b�s.���!
׈��us}�n�����Ҍs��-K;3��GOZ������И՛���NKy�q_f��ќ��p$U���PBJWr�C��!�o��}��3K|���z�U\Z����Xe����HcbStr��f@���g����]�}�6[�SCT�5��>u�U1����6�)n�~�Db=G�f����0����!�	��u�]��?��?��yV[f��8�)�|:r���g�������:��Fŋ�,9��S`]#�	�-N@��MQbc哵�<$������ �`�������z!c;B�Nk{���hp�?�����;.��1}����=�R�
̺1�윘f��+���b�ǐ�#��Wa1͢��su��q?g����ȫi{č�ajh�*�Gd`��Pڨ�r^�q�[/\3X�O�ɩ��lLY�B5�y&C'�T�f�K����dXv���v�����������3��e�,TQ!���:R� �bS*R���pLΑz��-b7Q���[�kJ{�w�J��G����`G��Ҥŭ��BOEe =~�u��.�0�V'B�@si6;�6u����e60X�L��R����S��~�=��RA�������k�57bY�w�l�'����	�?װ���,��h����قֆ]�*%��!KFCʡ�i�����ڀ9�s�C�Ϯ/^���<�Y]7?f�0�Ώo�L	Q`���N����4ax|�C#ܜ����E�	^��#G���NT��GP7�L9.1+�C1CF|_�\���W���wߝ[�@TdqM�3S9�������A�F�+H=Uj��STM�E��t%��Ub_��`FE^�j^��ʱ~Wῢ_o�K������HcnE'Xd.�ã63W咳��ߙ�H�j��ɫ����N>�؇� Lɍ�?U��-��ۨp��[��0SL^V:̅w��OG��H����O�)O�,����}Ѻk�x� �
�B���Y�D�um�`�5\Ѵ��ULS��� �v���S��Vp$�oz�0���9�$2|=�,�_���9�r*X�_�S����y��A>�&�K �}@�Z�~�&c���d��yۮGq�PO`�� HU%��'q��a���"�H��b��z� �S:���ؗ�={zF2rZ�R?|���޵?Ҡt#����%��2`'NM؇>�1�[+q�r)ҳ��xj70�HNq���8�����kg2�S�]�W�-�ʧOg�*F�`۳^�zV���ز����L�X���l�b�\�X��Y�~]�y&n��CG\H�2m�~�r�����Gg��I�+���f+V(f����>� �o�^8ǅ��Ӷ�SǬ7PX0��N=��<}�X-x�j^㪻���ȩr{�4�$��M�et]�0�|��G�A������w<'�Y��H���� 8��n�B�N˶|�����/��҃8�T��� hUg�⫵���	��ˮ
U�9E^E���[n����҅#��������Kw,踆��ګ���^��<�)pn?CŇ��87^FJO�2>�q�t#́��S�/�#|�68j�����ÐPQ��������V'�g�M��Zu`>�P�j+8w��}�R/8�\��G%�u�!���2��G<@�j�1[Y<�kE)׃bf���E6��l�+J��7��g��/�������lm�-8�7�!�O��v�~}�T(	��8(���]Ps��AҎR�"�Ry�ί�"�Bvn��e���v�ѱ����63q�]ڊpڠ�����v��1�7Z��o!.��OC�~��2t}*����L�I$����jCҴ]�wޙ	^X��)e�T�3p����%Av��AoX���sX�@5�a�"`��w�ݟ�����?T��^���G��H��X�R��<� U ��Dv��Ӵh-�����xq����+����Z9�^.e��ю�9/�(��p��XYO��� F�������U�G��������>+���Ӿ@�(�;�V���W\��Ä�����{<��޻��yH�����Ԟ��:��'�Q�S�*�p�c��\�dd�^������	њ��K����6�zԖ���۷�'?���O�J�E�+���,���jv&�h�������~�� F��ќsvy�x���#v|�DX(4np��J����-"aQ�pN8��eC�Ñ�/���,n�w~<�!.~�������� G=��D�),�!/(��5��Y���<DV���])"Y�b��wxM���f��*૶�i���֑��hX�Bܣ[�;y�n-�:�Pj�~�]s�e��m�;
�v���ܲek�˷#)�"B1#���6��R��ѭr�s��
��`+3Ii���]��ee�n��Y�������;^���	�j4Ȣ[�n�]{�u��ؾ��/�}��i���a�I���^�{D��۞�^�^Y\���ӮZ�?3;ִ=t؎�<�^��Uk���>P# �����0H��{���ܕ�7X��>��O{���:�&���`��Z��ێa,��R��������U�"�x'+Z���w� �W��I.�b"K-��z�<e�S���^N�x^��d�H����~��7k�կ~�c�<?�J��@a�b�s^�5�)PSz֥:�!�H�T�#�X ����Z���Utυ,.E@�F���9׀' ,�aD��9�3V��?�)�Mk�i�,CZ�Qw�(f����Ms���l�����٘v��z��s��@�o�{,��(OJ��w-S������x�N瀋��	o�>�Т�
^��V�U\�ƾ��_��_��m0����U�7sYr���z����.��U�9v�O�S'�z���������}�P 2<4jW^y��t�-62�<�Ղ=�Y��Ŋ++���@Ѝ�����@�
�Op�~}���h�z�С����o�ӥz�A�"��l�s��^���^@7���\�;��3�"DbKq?��lY{jB�TF��.E����xr��M��`�eRk{��g�D	M��q8���{�oe舁�2(�3����Ӆ;B
c��Y�<w�8�a�C���j_P�b�NF� �C���"@�F
�O<asF��c��I����7�r�l�!Q�_��p��o���N���Vl��Q+6P�ᆗU�
h��Uʶ�.{�*k�>�2��̝���E����a�L��=�;�p�a�^{������g�|����m;l����-ۂ2\m������c�֌�ٛg����Ӈ��z�_����ş?��˯�ʞq�Mv��^���G�O���/�q�gT�6�d'�����^��9��%�@)da��*'X�����������{(ɮ�\x�[�s����F3#�r@�H��g�c��f9��᷍��l�1^^��<�m9'EF9k�&O��t��|���s�ۧk���i�3u��=]U7�{Ύ��6�<����je���Mo���IY�Rs�̝�d͊3L�U��et�������?�	xu1Sis Kt����o���`�ca�} 3ȹBW�
�=?�%�aB_�(���H�Q�.J���C"B�j@��ר0� A�
���8����y��F
! ��~���8g2?���*��_+}q]8<R�EeP0`�1��4X�^�O�Z ��������Bޜ\���n��f�sޠB�O-�N#tC���4��L�RN8�@�2U7b8�f!N8-�\G�n�e���O�s�(;�C�w0�Z{ը&O=��<��C�k�.��^�z@
ټK#r�����]���x�,Y�'���Q�������cn<Щ/��z�����JcґO�����X���e|b�P4�5K�Y�bqT���?��O��x���C��&�Nc��R��8L��$�Fֱk��X��C�����=%�܀���C��<��~�;9�6�ɪ%G�`4�^,�-@lѕ�H�
g
v'�5���k������=7�	�P1���;`�d!a���I��*]��� ���� � X��
�TL��H����9�]<�&X�P$x���964�EL����E�Dx��H 7���Nd,�b�sa����f��`դ�W�y�j�G����Xo{:�^'}�+͍���l\�Z�5V����`�5,6�D5�>�A�HO�ׅ(����6��R�A��1��wE��j�T+#�����HWg�Tj�תқM�T�.G����?�o򋷾NV�� �V�4E�o߷�Y�/£�4������4�X2`M���әH|�ټI'z�2ٻ���.�0g� d�'&�TQDr�h�/49�%,X���〛qO,v4u�{���bs���l� �U�������\WW��s]R�M��A�KJ�c�D8�U�E
n��K�5
8�t� ���%*��%� �c��AE�nPldN`C7��P�q~���a�@���j@b�x6pg��W<8'�)�>1�sM�"�����H$*$|��̑����)�	�m�b�i�G^S��Ϫ�*�CU��Ra�,{x��}Kep`��������S*X��Bz#n����Z+Y̽\.�1\�=z�GO ����U��ɸn|�P�z�>���^�v�^GE&ը�zGw��G��d�X�cE�_��l���39s�F��{���q-�)/�-�6��BQ+�V�IOW�.��F��$��QT+n�Z����,��`��,-kzՄ!����P:q�:��Z�܍ՔH����w�i�6�&Zp�4'�[J�$"��jm*!��u����ez�hm�|,a��.X��Wb����,m5�^ ������sI�8�/x��$�&�V3>%�����B4�����}�vZ�Q�!��i���W,�����J�|�FXc^ ����������a(�C�^=6��v|� �C�^j��](��ߧ7�VZ��Ĥ|�d�����T��	|��޺�e+�������·�#�x1w0���IÍgxp�n��s�:�3���ۗx�&9
������y�]�s���M�����c�V�ϼ��Z�S_��3�< &���C����
�:�L6�`�@b�V�,Zj�<>�)��vx����}���l������©N[s��UX�P�\-
�x�FT�D0
x:���E��~*0�7��ix�e��!Y,~��7(YI�CқL�m�ϳ;��v p��b!+�ɷ��h,�:E��!Zm��S��}�����>R�gx\��a ���&�}( �����8��7�zQ��(�ώv��U%1X��~�a{���G 
��f�}	�j��`�խ�5�=��-�S�խiz�܂��
����rV��� k^@���?�cy�[�j�-6�G.�=(?��֮6��e8�
:�!
J.�1T!
��+�*Γ���Ge��{�
��x)����@��#)W���V���|.)�w�>��^�x`���QmG��.'����Q�X9ࡀ��ݿ�8���˧��8>��J"[�#��ȡ]r����EK��j��Er
��"RQ��"�T�z��p�� ��A����	D�A��ˎ�c���T���2�7x>��b<|�B����]�Uxn�,~"�$�'����r�}?Nx����Yx�n�v�f  �K����
}	��N!\#'z�8P>���:������nB����?C��D�W*��K��uOEe��2���C��t�%|����6�~$�VUϿZ	�=��S��;�}�{���pohbO����"e�'=8���f;���T���CϛM �$��>�1'�*�(F�FOθ�f1���9�S^��4s��ɴn�j��X��8��o&r\aUh��x�u]p��@�,����x��K�\p@䰘QJ�67-Y=����=\5i�8�o�^ߤdԺ��"g��8H�X}GӖ�v�K`���0g1�5v\�\�>�*?XC��;=dȇ������=IZ�P\|nx�a�@��eX��C�/��&(4d�� � ���%+������u�p�����Q�Qt�B�v֔�|w�}��
��q���ճ���o��8��)����Uu	t�E"jm�z_wv�˹[/�J��*�T���O��_�.)���@٤Ru?���½c�c[%naZ~���?�01o].�V��~	5��ať*R*oV�[#Se��Z/����i��~�m�w�AV7+~���~�*[�H���'�L�w�v�Ly)tvYy�Χ��2v��i�+҈��G������w�y���w��][����f� !� �a��tv�?2�o�BKf�4�Ua��EO��?��B\x8����Z����`����2QeT�~�C>�>�n��,ߘr�J�g���b�����Ig@4
�:�g�BKPX�;P�q����hL��a�T�����60M�F�9i�wS��EE �z&e�8�9���U'`1���H�m=2�����,�G  ȥ ��#���!�t�2Y�j��Ke5�ft�ܪ��7�vmM���5�\��A�H��}�z !^.��������X��v���-MUd��{e�sd|�\x����'d|�l�7����V������(H\��7�� ����E ��<������q`M����z�굌��ş�2z��1�4T�hp]�J.Hjűw�q�.o6\u�<|�zX�،p����I\��'6:��yv����ρ
�O��sD��B���0D����������v[�x�X,#�^*��|����W��(8*&�휺�p����w��@���>�)�V(BDØ�g�ٱږl��
���˩�V��=�#vC�����C���0%z(#B��q���l+a��6{`I�Ž!���G>��%�5p�}�c�R��m�](���P�ꀾ� �Ī�e�Y��[&�;�-�$j	�=���
��?�8����s���A6�K�bz?�C���iY�f����*��2tx���&&F�d,�.Hhn�z��u��$<?b�L�b��� ��͞������&]w, +��?�����~N]��y�.�$��8Ir��K�\i�yZCjX�ӷ1/�5�����p�c�(6g5j;����$.��a�ǯ�3���%a>O˟�B�,c�8�6"餱|��iE`�g
��(?���{���!A���Y?�����-�F/�`���U}�X=�%r�Tn�}p�O�Tq����L�#\w�QC�� �_��_J��0ҡ�$l֧� 4��u���Kj��a��AȝBΘ�׆36�5��h�ò����C�䓻��-���Fr�q���uq��>�e3/�FY��? _����u��U�rM]���iG<p׮r��ak�GͰ^��Ns)�q�C��p<��|�3�7�Ɋd �#�V�+^�
��W�l^+�i]�ӗO�v|R'��dCv=�CjU��֝��@>+�5���E-�T:�����Xp+�%��'(F�W�p�P���'��yQ��µ6����0"�Ճ9gXe����e2lCd�X��7C/[�Z�:��q|&*B;1��҇g�d-�E ���Bx#�okk�81i��By��l��R@�*Ž�F�#m\�į �݃Ec#�q���ڄd<�1�E:e׳~
4϶XQ��������A��0�BD(��Ї>��ϸ�gp�DZ]�{�!�6�����J]��d��@�����<8j�����l�v�z,��� %�m�}�d��5�i(x�q��V#p�bb�(����N)td�%/y��k9Ier�eW�Y��&IN6��*�U�����1w�?�c8tP����ֹ���k���H�R�����k������X��Q���]ۤ�_j�Ѓw�#�X*�:�gƅ��J@%�d�.�?�.�@�a�<����r���ܡ��pNl �5躓��վ�L����7��S����?���~׬Z]S�@y& Q�=6z̅�j�%䦳7ʅl3c�;`�j(�񊅐�� &�>rԎ�Y�0�rd�����{l=�
7(�8��EBki��a����V����P 𤡸 ��}�8�����Xƫ�Є�f��ի��[��FR>�����è��F�[^�R�3%5�r�K�������ռ�`<��/���y9�c�~�<����84��+��I.[-����\�(�~��!�c`rtJ>����C�<x\�x�(l���s�J���}�0�x0�L���p��T&�~��񉒹��t`�@�����pb�@� ɋ��x<,�~c��*!��.#,�|v&_���6���ŴI7hd! @��
S
�C���,,*�zc���D�c���  �ň\Y+`�!,�{D����m�/n�ه�an���<��>{H�;M�	�i�3��:,rҋ�w�e��_�m�ug�  q���7|���Hр�`]�<�'�>�{"�k�9(!��\ӣ���v`|8+W,�m�oAה��!�`�aF&U�wu�[���j7xwu0���$���ɸ�g쇛~��O~��	����J���M@�Q �	��,�[�J���$U,tv�cO<n��@A��!_0׋Aӝ��?��e؇}E��"��K�я~Ԅ?�
؜�dY��H� Ə���b3zǬ>,�?��?�ςW�f�|�4��bq�����gB��⛵:�B�T�'Tk	-��h�`Ψ�Q��m��CH���j���.�s/ ,0Z��� H�`�ạ�|b7Ɗ�����i|ZgZ�0&��� 7���7�O饢0	��[�����ǏkA��A��w�wm���_��	i6H��>��4��:X5�A�c���뿶�!��ϡ�PQ;T���&[�c���9���i�5b�sd^���p*�^�Z������\���s��z�"�^�|Y�|�]���S���j�Q����|����8��q����D����d��/����b��)/��d#$d.2�Ҙ`,>L>�U0�c��7,J��ȊȒo�ƳM#�}>�O��C�~��`�����;?��D]E��=$��b�r�@#�nD�"����C��Q5��mm9���h%B�����_h����{��d
d��j���XD^��/��`g)���>�|����h���a�\ ��{�]���a,����`������8'�C�<�������ll�C>�=7�R�,�FՅ�@��ϲ�{�T�޾���⹌�=��F	��� �R�*ܔz���?���9E�0����������=<G(W��^ �'�7�1�02�9������:��|�5~r��˰i�4�7��eec���Y���������0��I��k0�E�&�	�釞����EuH�<��s��0���Ca�L���U��2��m�ԋ��&|��ZG�o������m����Hos�~��o�+��aeb�A�����p,��/�.,�w��]	���!�������c���#$�Bˇz�ӦWɦG����i���<����M���Y=�U�@���7��ֿg���۴Y���K��[R���*�S���64�JK-UK���~��Y�HH�sG�������C���O����-���bIVi3�@�EzrW ��S^��7�Z�/Fg��������d�9��O���,6,�>�$P��d �Gr�%����o��L��:J�;��뒎�ZS�qݼ�p�k�}#���:�7��!��	��[�J ���Φ����>.��8�AC�\�X#C2n����7���a"EaϺV���%��3Ɍc5�c��B�'`�1@t�F�*����A�ǳR����'���w�Q��f?3�Dm�r��V�4�����m�:�+ӎ�>�0}d���������w[��Ph��½HXã�L���C��DC
���3f(��c���c��b�i/�1�L\{̰�9>���
�Ho��\�x�X�
��P ���U���[� V5?ϟ�l��l}���oTC)N�%�B��KnNʕI��fBG�4R�ؑ�ſӨ��F����n��D-�b!j��LaDWߧh�����rV���X}�(r�P �*��q\*,����J���P��	M�@������@1�G\��J��%��ҟ�]7Ce� <�??�R肇�ew��fA��y�汦,\j�9�_��P��q��=�1�"(?�opݸ�}�c���7�5��"�3�O���lY$��>�~=A+l�?N_��<��R�\Z�\d~۷Z���9c�<-��H�!��W.x,j|�)3�˦|�87,�Z�YS�	� ��e�?��q�wa'�L�l���j(�0� �AT!�,F�i9?l��>e,�n?&;�:k��(��!�?��}( h�0�DCk�	��6\��!b�T4P��nR�!1��3�l��ռG�Q��8��CD>�r����Hv�V���!��c�L�d��P8a���֫�7���q�?�9~��=����?��$J���L`ؓρ�<�$������<��fΆ������Nߘ�|�_�>'6�o��	�kCDxDJPX�'j  �a ���[@̵i�$�oq̮�&�՛����~�)�nE
9wO�c��6E��[D���,��FvōG+�����s��%�[t�3n���R{,l�����/���6��/0(�0����g���}�LBC�x��|H?��?�Z�~�����ѐ	F�/s]��ܵ.\�а��Z��n�\V�"0@�{F�����2�t�q�)��2K��h�^)ǐ�ؓͪ�E�\<Yw]4����	��g��)�i(����7&������':N{����;���VN�oՐۃ
�V�����	��l��e�p� I?"�=�S��Q� ��PO���ftb�^�D�T���F����9c���;�q2G�e��o�QPxFC̅w�1��\���;(MT�T��F���#�?$�HoϠ�^�A�U5�O(N��%��f��	z�T�����"bh�ъ��|N�"�@Z�E���IfB&9�,�ހ��i��!Z/P���s����T*�w�voeA7����r��n]��DTܗ���V��Cf�l����� �Q7��@7�Q6��+Z~�M{<W��kQ-q���ټL�F����K��ua�Fv���9cI^�74tHB$��h�3�O�"�3iT��4ʡ�-�8��a蘈?�C3ĕ��Ӝ�8��|��ӧn�`�#Q+��LK����f��|r�3yǇ��{<�}����ύ�$�,����T&[z�r�H9��(t��
c��b@Ӏ|�]}�cm��8�cv#��]����n���o88rW�Z:���V�e]]0ҜYŔ�4 %p�l���}�*x��"F߈�	^�b�:��̣�8i���"=�٨���4����  ޘ-.��Td8�w�h��°-v��|<.CA�|~a?��\�KK�_�R�ԪGb\+Y �b��Ѐ�Ti��LUʒ�,>ZE�_��u� �'���Ӷ���6f�I��v�t���)[S&4a�u>U�X�s���|Q[H��ܴ�vh��˷�����'8� �a�Ic�0�I �oȠtj�{��TP �L�_?Q�[��<O'2Ny�?''r<U���3���	.�����Xt�(�}aތv���Wr0���#�J�xD��k�f\%��
�TC,�+99U�kba������7Bc\�f��Ԙl&������h��5Z�HrhX�rprj�5H䆇G��Iވ���d�*Z.�^�W\_$v��'KR����d&�l͠��p�&�g�f�0����~Q��_X���F���?�8��f��%N�D
pChd�3�A�؊�������a�M<N
O�]��Dt��&u����bh)���D[��{��T,�F(�uߨ98_�~�]����I4��26Q�#G'��k��ϿVV�X�\/��M��'{�Ʊ1�T��w:�����ό�J��zcK]��K�O�I�Z3�P+�Z�
��:T�ҥY�'P�����U2Ĝ+:K��x���]�`}�^����V�Npq�fU��F�m˿����� T��1�6�\�p��er��73X��&�7M����y��կqpb��)Q�ҝcl��u�`Xv�6�Å!:ؔ��y����ʰD�8��1��;��T2k��U��C����%/�ŘH��5��7�~'�W�q<܁Mb���dE��>�d!�	��A�h��Ȯ��Lޗ��I1P�g�t�������6湟�;��u����毙�ol�56wMM�y�Ӵ���<���6&*����<�Y�ef/^����Le�4,z��Ҥ|���_��~/e��W�6?�/��[�o�Z1A福u?�@��1�f(�����8P��`�.�#�����d�gZ!�o�:����ϒ+.�\���oX%1��(�:����x�Є�iZ] ������U����'�z����1{9�r �=}�d`�Y��=�׼V�{�L	�(+��u�Ԫ�U���#�
�Ը�FG��L�wMi�Fdx��f#2%e���;W�V��b���d�X��K�����G��^3���
�f:���2��%�Gk@@4*��<���(x;���T��3�!�V�7{���ǧ�f3�ڨV�,�0��,��V�..�!"q>���n�.m>%g^Ohg�3FH�7�����$��$�%J�e�&��I��H�V^q򨤲*X¼Y��;0��E�S.H�����y�����y�E�P�J�)r�/Z���@��@?�D=Bz@�`/�3�Z�l\n&�c�PF?�FG9mI}�&�׆�J@�����u��<Fz��?�����"_E�������Ƌ��c J�JY3p��L��z,E��V�?,GF�4b��.3�4�'��(X����Z���L[��D������7��g2Xc�$��|�͇tC	ԬaRl��=i^X3���X�˰k!�]������(��aPV6tx�>�d�R��R��Ȧ�Ζ�k�[�� ��ߡ1�N�E��E^QԂ��r�
\;����*��ꄏZ��O���k�����I���/�X�ٲU��XeM���j�`e� �h�fO,�׽�u��YD���ˇM��D��d�"����0b�ȬE�o�,��}��45i:������czh>��kL�h�!�'%&TL(�@d�d:�_u�?2��@������4Bm���7��u��b�/�G7r���w�h/��y����HP��JkB�}&��#'\U���&�èG@��g2ܚm4 �.���\�}P3u`-��}���~?��*��ç�-���	BrhP
�j�|̏��X�7l��Q�h��dVn΄P�2���Ϫ������ร�_��-�E�Е+_M�=�x��GT���8~E�F�u0.�鄷	^���GS�h�X�O+Q*��8�c��T��p����}g�/���(�}�1t�1�U����T'z0'&N����ȇE�?�}��(䬝㱣#*�'�|\�������q�9r�ŗ��3j����?޾=!������u:7po阡�I� [��u�\�|��pJr�H���%w��=����K�汪�h�����^����L}@Xl7�|�qsӊ�5 �>r�B�;���<����_�z����[,c�� oj�+����Mق���"I�b¬h4��E����&������|�=��A��t#����ZY��U�(̙�`a3��1��V]qI�zL��n8P��YG��7h՗a�=4�?	��x�e���sq3�,��~���5,����F�	�Oڊ�,~��±��	Ⱖ�جi"OƦ/tmQ���҈��A6gE;
�nK����������R��G�� U�j���5m�tʅ$Cԩ��~=����P�t��$���g�W�<AJ�����v���,O^#�a���$�3��E�Y�<f��;N83��0%Qz����Y�C���k�5FS�����@oP���������߃�����7!{�<!�|ر�I+P��p�9,O��>����] ��Ke͚U�8��'w<������I�)/�[�}�[M��<O7�9��f�c�%���[�˭��"F8:<l�����_Z���{�g�a���2��6l��.���P�o����Qs�����o���a���d%8O���>� ��:�ıZ`Q�*�'�N�B�gI�,�����QF�$�Z��W��I��.����P�V���<��*��n�JY��B��9"ׂ̡�G+�!�{� �Z��j2�|H�S�:�[��j}DJ�q��(�5e���;oT��Vc�!��]X�8_Ը�(;u�"�%�!�jჷV�U��KO�R����E�*m��N��`mG�0�9*�ָ�U^�q�:�*@Gꗊ��Gus#�l�r΀���V%�����U3�d�ff
�|>Ãa��-�Vፐ_:t�j�ٺ9NVV��6���
��e�u��ީVc~��ǯWFr-�����Y��>��"��L�����`���"��_��������@��=����j܌���!��I]�����3��(�՛�*���-�7��笁;d���0W��
~�S^�����q�s&��͛�ڄ���ʷ��e�ֳ�uk����	�6fdl|B����	�y�u�]g� x�Gy$�h�F̎�V�h,�p��2f�����2�(�}S*�U�,D"�j�J�B4�=I�f�E+{���M��5 �j:���F�4�.<�r���g�/��Jy��+׮P!1�B<vC�p^�:@���ty�*���q����խ���C~�
��� E{��321Z6�epi���,Q-���+��v=.���p�K�8�B;+K���a�H��UUL��0p���T,)it˝j�g����#�^�#�s�'���/�;������REcޢ�wthJ���άtvAY�1<�I��g6�#E}��[��u�ͥ��)�� ϰ&��f&k��,��nTu9z����O�9<t����N��~,������cR���r>��I{,�1`U}cF�k_l����8b.�Ǽ�����n�[ �B���z�{�k�;�������=�\�T����񈮑��Y�D��)kh?Uv��K��������;�'+V���/���m�'���>�ih�e�<兿��� ���U�;�Q�������q:\(&�l-�p��B�S-�1k�v�-��%�Nm�����	�^ U��݋�/��/��@7%߭$wG3�ۉ�f:�f��E��I�m�ΕMg�։�������*�.�_7�V��@U��C�F�;������b�'��R#�.�ۈ�#uRy+V{��G��w���뮽J��ҮQ7�5��Z�D�#�������wn����u�Y�e�:U&�di����*��>V�o�^��(ʍ�]%}��t�۰�W#���kBqa�'Z&Ǝɒ%r��W�v^ ���\�>�HY�ꍤ��Bjt����#�ߴ������*.T���W���[=� �8�s5>V�o|�G��^p��?�i�/��!��IC�c�׳����m�,W^u���Y�9���	�F��R1���}Xʓr��[d��:?u����[�}ʱ��7��GF�^���K����<��E�����0���V��O2|�B�������~�+v.th����Д �������#r9C�航���xTe�r�?��q:R��2/}�K���蓣:Gw��r�%W�~h�ʕ�������f$���k1Ny�ߒ�'r�-Xh��Uj�8p�ڿ�P��֩��::T"n��*�qO
ZZ"����H%
��;�y�?��/ؿ	�d���\�6�
�|/c�O3���#maX)(�)�&�,*��zք�6>Si | lr����VQ��ch��k��"��Q�o���@Za������MB�%��e�S1���ʢ�	ز*�@/���`��-��p�f�︡�
�M)XE����q��B!{p���Y�5w��]C e@��oOA����Gz�s"��a�,C�j��u�A��~�
���B��Tծ6�BөF$��6�8!�Qu�"2�IxO�������Kh�fG��(���e3h2��zQY��	bNcsGx����p�0����@	�z���Hf��q��b�q3RH���kD������F$�eMJ6������L( �u���
�9��!t!C�^�7 �@����/����jҮbxl|D��R}�i[��a��	�$��󙔮�kk�DgGo���:�q����o;�����Y��h��8D���ߑ�!>��x8��@1��o�����P2l���|/����Ic4[K��ɒd�ŵk�yF9�؂��'"5WSV6m(���+"6mEh%�w ��<F�v�C@�@�{�X]��Z��[,��>+��Q$�1��	,$N+�)��ͨ�"1�#�آ�N@:�G�a��į��\�ؘ�rQ�6*��UХ$��}�*$�E*v�Z�b�]U,���M�EU�����nT$V 4K����ҁU7!�S��͍����`���K��T�~�
�|���ME�Y�Q�nM|`������*�lƞc��C��)�C�-}h�':ȕJS�iK�?_���3H�\�F�"�i�0��.Yh{*c���ײ�D�I�;K�B'��b�'
}�A`�{�{����ޒ��?��^�*���lﳾ�͎X=��Z2��^!��kA-i�$���&��,��`^\�:��n�2��3P�Tͪ&�R)���>�.�	F��	���v+�5	:eCnQb��+-g%=<�^z������7-.�������/}�K���`˾���}�9Z:���9�9Z)��,�kp/q�˨��E��*��:W�Ѕ�`� �Ě���3b��#��Аad �g"V["^\6��x,���5�Q�)�@b��0F��s�H��0��$���g�TW��6��nө72U���В�����d�D���x��A�ϪL��.�	(�sʚ�l?D筼���E�(��'	q�!Y=^�����2錛�c*劕j��	{�~Y�5m	_�S�u��z�����\C)�)���=8�qEP�_#w�$�[�<s-�~�O��a�Cj��:m�P�r�����Fw�>!�Hp߰�Br�gfM��c�Ν������oΫ����q���8�RdH�l��F�*U5�
�NWcr``�<f����=.'�E?����?�@U`GgA�����Kz�j���V�[�{���Y#���L��DE��V����6����^ ,�������K��+���|�#����\@$��U�ܠz�6}͌��۳5��������B�)uOIU���`�Y*X�CG�&�!���F"��F�j9v���\�g �[�`�a�NQ֡�fE̽��N����D�����>��g��ʆH*������g����1�u�������]����%a������5�Vv���W��UG��r�p��BcYU�cG�z�D/�`�����16Z���^��;t�����|%e-���hk�3��8����
Wmj�Gz�X��$�#g)�JU+�����̑#Cv{� B38�SQ������U��l~�z-׀�9S^z�\u�T&&;,��/��B������wK?��Sjh��W�hG�L�2#'��ǖ�+����q��gn=�Ċ�0�^��D w��;��p��� ��?k�~���uk7ȡ�g���V�����n���~����I)�|��[^���zpL'ͫX�8�$�%aN��54я�s�v��7�+�-W_�y��{���.��]�K,|�u�u�M[Wv�aX�F�W낯�ӟ����P7�t���o���0�~s�"7�$�o��o���E鉺-� p���b���˖���:Y�|�)��v>)�?-S��%E��EY+r��`�2Y�~��%�?�^FT��ԣ���c,�L�
�^������;e��5�v��1cC>�o�ZS%#��d:,�X�5 �*��'�fQ-[�Tϻ֊���{Z���%�)�\R9C� {_l7��8,��@��߰BV�Z/�� ���'ǆ����,T�kjD����������2A�D歹�T �-Y�v>*��~R�"ٲ%�%U�L>�)� B�%�ӻB֯9[ϻN��1����U>�T����K>�ڂ�)���\��Ⱥ���Ы����?�C�ј���p���R4�����}:��e�ʵ����d����Ԩ	�P�	sVL('t��Pa?�B�]+T���9����^��\6{MHDW��؈��4k�DӍ��j�}�8��1�.��ϱc�~��_��_���E�@����Rٹ�aٷ��Շt��V+��;��e��~y��'u�����,�F��@~ͼQim�EQx��}��#
m��bR�㮻�˥_&�j�#q�~�9rdhL���'�ʭ�1n�p�W˦�ےb�{��\>Ұ����`�����|�k_��Sf��1��s5��q�-�GN|D�C=!6�I�Z�Thde�곥�g�
�N�9��aCڬ��#G��sm�����L�����9c�f�����W�궚
c��Cf����X��D��2��@ϹV֮ۨ�YH�3Ղ�{߯
V��%��q�����w��sW��X-����JU��U9��rŹ�, ��^��N���M�.TA![P�Vz�d�؈^g�u���oZYU+W�wْ�r��3�"�ϓ�*��� @�*F��Qv�O*g�w����z7���*A���;/��R�Z������Wb�@1V��~�w�Z�)Y��G�?'?�~�
"�ʺ�v�zC׬�?��/���v�U��4 1ͫE�~c�����x<nq��-8�A� }Fh�۷\�:{�z =�,;{d�*���wD�1m��P�5Pn4�T��I����ǯ�hQ+Xf���]�z�z���~�����Χ���5�y�����}�3 ��[���!� $���սT���(���W	dr��Tv��~�U��s�7�h�Ȱ
�$\dJ��1:s�Q�Mҭ��#�������E/ԍ���^)W\q�Z~=�l���[�����.6K�/~�f���H�7��|�r�ԧ>eP:|�w~�w���a[��,�&�n!h.6���.���A�U�ꆯ��4fbq�n������.��YQV�ZŹ��~��4\��b��,��IIO�r�n�ֈɺ ��(O��c!�jC�Z�pܜ�TEܻ_��B-�^�2��M�b�UƻU��ˤ����T������Wk+��2���:u�;:���c&�sªY��l�*1�x����kM�@L��V]�� ����4mJ�����0�TC�W��֯�"#c���ڛD�4��F̀M���):O%��"�*�^�R\����H�`���z�=�dD�j�58�ӈg;Σ�s��J��Y��jYv�K�=�d�>��S%QO�1�U�T�w}E.o��z���Md�h�=�R�3�@�!��3:��~���X�L�
�Azy��y��F��Ac���%�F��<�P"�x��<�b�WR��q��Ss�2,tp}϶��ׂ�IՀC�����?���z��PBr�礝��<~Ȋ׼���[��,]��y���}�?�Ò����r�5�ɖsϓ��X���>�_�)����e�����?j%�<��U�� G�O"����)/��Fc�V���kn0aE�Sk'�ﰅ`t�z� �	d�X�@�� �9T��;��~�#y���-+W��!@iU,􁲦�O�2>Y_��X��<��,�zF^���e_'�ͤU�Bh�^��
��7�u����׾c������j��q�*���U2e�6�I�KRQ����m��yz�nٳg�\r�r����E��`�U`���{���&J�Id�����˱�1y�^��?_�EQ�mJ��
�@�W��MDQά�~���^��]�����ea�[o�U�٣Ϸd��(*������yq��n9g�6����S;���[/���&Y�r�Z��l��.[c��)��`�U��7�\6o�P��|�;ߖ��k����s6� �2B2��&�`EYl��h�֨�c�paC��?���ۥ�җ�D��id�t�B����*r5j��]{�z]c��#����9�\ 7��")輢�"�Ϲϫ�����R]��.ٲ�K�~�K_�b��oy�іXD�i��_��z��]��D�r	�^Bk�C?�ӞY��î}&@�R ,�\�
}�pѡ�:��S����ȵE��>X`����@fpO���� Q���A��k��P���s�̳Αo�9�������iN��d�$w�u��w�vɫq�~�1��g�o��=MNy�H+Ӡ�����y)����|�2Zg�;� �����N��z��g�����.��� ��g�/$w�	�C�ŀ�x�Ï>��lC�a,Z�-��8��%��	�@����Y#֟c��� �DW�j9��F������r>2<)˗ʹ[/�u�W� ,��ZX�g���Q��t�jA����19phH��v�
��,TS�ؽ
�2b��4�,H��D5�9����e�X��.�B�ظV��}��rV��87��0��eЩ2��Uo�wTWJ�l��X��b �ƘP:��0|Y��2}�y��'Գ�+�ܢ�|�����Vv=�A�!��"Jg����S�6WeAP6��@t��X�X(-g�EC(�]w�t� -�>�J����BY��K�QŠ�H2#4�0�Td��U�۷B��T{r���?d��\v��5�B���<G�0���e��Y�"/G����[^�U6��Y�*�.�Y�8�"��!��ݳD�Z�z+Crtx��vδyH�a�#w���q�.V�������9�p�ؓd�D�Ίeˍ��!_|�W0 �
�0��rYX���W\j�H��;�����s��##���ʑo盦T��;t�M�1WP˜^��K�<�pp������Mem~��ߕG}��;V�Yia��jo�;'���wВ�۷ߗ^r{�!0v��8>��Z%0*{�0�)|�S�4�Pr瓆�ս�	o��<���j���f�	*#n�r	N��']B�^u�!�9���㐁�$2N]-�RmqC�����@,�6�Ej�Ud�h+��JĪw+�X!mU�)K�A0cn�F;²�LNLY���c��ڋ�W����jgü�[��l�f��A�r��>���9���}��҃Ŗ
�"oČ��Ɋ	U��1cNZ�8�\6o���*5�r&x�:�]�H#�� �',i��@11��h��C�P!]��˲���c�5㺪��X>��Ƚ�T� }�g4:6ay�FX����n(��Q���x��F07C��y��F�,�B��R��ks�deGGg�9|�L~(R��=:iV�Ɛ�(YL������>"�"�P��8�~�Ϳjt ���� �9�����Y�c�+�
|�+_��M�e��.Dɶ�!Tv�ܽ��ͷ�q��ۿ�h��ET*1P�1�ZgA�����.�
���"&��V t��
�q��׿f�<�:� �U����x����ZR�0��i�� Uox������k֭�߻ݒ>��� �/��/m��B�G�����E<F��b�%����͊�@�WtE7i��8��u��L�"���$q²��nk�ё�!�mxR;G�GIP���0�՚��;��B](	�x�{n}"ǜ�U�?.	Cᙕ�QRp���¸f�Op^��
N��������g�{�.�7N�ȑU�K7�y+�r��(�M�TP�������I�0ra���Ūa]���)?\c*��Z��t�
�i�hV��P˭jJ7g�s�X�*�1Q��-����F��rE]��F��%��I$K5tךN�cZr��A �2����m�y_4��i����Z��>L�r?��e@=�?~ߟ�
X7d�>�Ʒ�������>A`㻀h�3�l��`�=�z]�o4��5BX00-�{�-	�#g\�l�m�>�[��X��c�R?RO,k��uu��B��[�(�B��׿�����`0"��'4>ڴ�9��2��2�4����a���&�1�npΨ� 4��̊h#$R��>.�g2nz��������n.X_��������/����!��^ ��@k�����2I�)�K$�`(���>��D">����2τ���["�P�g�OX��ݜ�*DQҎtnn)Zˁ	m�1 �,����"b6�~^㣅���ʙ�U�m��3�<S>������ߟ�� ���>�9�� ���D�^Ƴd�ܽ#�����T8'�|8h���s��6��aʹˎ!�3��Ȋ���ݴX	�B> E]�Ї�w����躄M'pY��\W���~�17]�t�O{ܪ�Y84�No|&:_���{Z��k��5$>����54�H�s��b�3���b�}2�{籉�'j�J���G�h���量>�-��AZp&�G�b�mmb�B�`O=�>��>�k����}�'��Z�v�F�욟04��W's�s�<�,��:�+rv�x ��>�,9�0|zOT4Xg8����|��8�k>�|�M��40��P���zh�aa�+`����O��L�=Sc�{&i-S�(Y��s�P8aP���rS(���>-5�"�{���M���~��;�w)l}�#T���y|AO��S���Ӓ'j������ p��2!Tدi~�|^�5�3�p[H�p<�ab��B��ÿ���.�G>������yoD�  b���-/ �
^��,����Ƃ� ��c����hNFs,�����ɤ7�'�m�i�yc�Vڇ?�a����}�����͍�>������7�s���P��L!�6�/�}�I���'��Mkʷ�\«��"6Z��5҂Ǳ���hnxc��y_�ӛ�s$�Wz$ �W����d(�a)���򇉀�����2���sH͖�o����}�~Z$H�4?,⯋VU긎�DyF~�g���-'k�f��u�w��N^��#��yDU?��y��ו�W�>���4p���q����O�
�h�%��Z9=c��
[�M<<�������>p�xA�#�e�^ ��6|Z�'{���!����+Z0��Z}��D�-�wz�x�gU�|�<���r��js�z|���|___b�3�G�L�B��p���A9Vw����������\�����4�3ŵ���yzE�Z����q�B�
�G����g���O:8�4p0'�(j��Q���ż�Y��+Þ�������9�=��Z�4<V��6�ۉ@�hٙ���Xsq/��/f��_d�6`% �	�I<
��M�\�}ف*e
!*1ߺa��0U4� �.9|d(&�j�X�͞�h���	�5�����c�3���5�y����=2|Ԅ�/����A�{�@b_���{�6L76�o��:g���Ő_�`}߁�"�s�u�b뉰�ߙ��@@�Ч���5%Z����>�(]�������-,��c226*ݽ=��:p�����87���8�x�~���:������>�~�]Ιڢ�c��:��,����Q"�S��[��g�dz���a��k��c��h�y��j��Kn$n�<^�uIRaa�c0AI4r���'�]��� �}�In��7�Ip�����l$b����L�����hY�@K���b��ap�O~�3�r4�f�Oa���.U�B��U���3ă�
!��.`�Y�CagB ���x0����܎�s��)�}t�����ߏ�7���00�Al߾݊S�5@1c#oT��n�5����2����s�d3��*w>_*zz����yP���<=��Ѝ�Ȍ��}���h�Od������ډ��L�Ml��+�u˗��Ń��H��p6)�
y�)q^�8�no��	&?]|�~8p�\�/?�����8�މz&�p�΃��_&�y���jm��9?��G��������ix��G�c���Ƿ���l(��0�
��6p�L��a���OC�
��Nǟ+*Z�;<��;���i�%Iq�A�`��V�)�4�4jq_+6#Qb�"�/�3hm>�� h�Rc��e�_�ͮ��<%]=�I�̚�x�]Za�d`�b�۱�ߌ~���Lt"j��h��76b�� 
����Ď,��~T*�d���;�8���<zܒMq��k1��s�a�#���?b��0����%T�I &�zg耉A?�K���R�;3|�����{)��x�����G��|�|��W�6س� �ņ�Oy�?Ο�/^̔_p�lݺU�����gYSr��!������S;-�%��'>���F�{��x��]���+
�V{��s{�'�g��3�G�{m !g�
D��oȽ�w�}VD�y�o���>Aˬ�ʳٔL��I�?/<���u����љ�Ze������p�g�s�>tD���;��"y���70�1�D�0��dCD����G{�������ʬ{1���g�^�k�J��_h�a�Zy���#i�a`":1��׹�|����i���J!!iֿ8��/|�M8NWwG�Ks! s����@ׯ_/o}�[�c��ii�~���Cdh��t�~���¥����h��h=f#h$z��믗[n���	�@0�g��-[�X��Aw�u�) �*,��Ny�ߘ��
`jr�������w�g�nk��{�N�x�K�ʦ�g�E�\f��(�B�6@�|�I+��
������_~����G�h_}�7�Bb�l��h��6RG4ú적~�K^�dFz{�L^ �������ADa��A��W��UV=��������F���
9�A����W_)��21>"#��r�]w�~U H����DL�<!�<|�zc�o��Tڈ�n��K����J�/}�|�ߴn^����jU�h�N���NȘ��o��h���O�3��W�C���GOW����ܿG����㏘G��R(�#����\x��&Pdx���lE��n�8b���Qs����s�\t�����)�V�etx�H�\����4���l-�j�>����ɫo�o���E\(w�q�'&�T���_ϻ�
��G��*��l;�<y�������޹K����h
 Z��H kBҎ��Vc���^'g�`�͓B}�g��^�23�ц!�B7t���o�Ċ��Rq�%�ʚU��V-�qZ�����cCOKg�*ݝ���RW����DE���w��񆛭��ٛ6�k�<��&�|���*�����o5l�!̢�}��_�ݲ՚z䳁<p�vY��G�ذR���ɤ�Z�i�6���P�~\?[S�������ꪫl1��G��6$�B^�}�{���7�2'�3���e�k��h�>�0靣;���Y�- r0������mo3��=��h�CV`�W+E��أ*+�j .�]�G%�	\߈L��O��ب�i����++V�1�Б����,>�:=Q�S^���a1�C���ի�J�^5�s�S�f������J��Svr������ݵk��t�M�;�Z��v[R��&ޯx�+l� ��\>(P=ca���( j��o��x��3�>��C�7�7I#R����W~�W����}��=],����<��òn�2�~���J:$�=-wv����49w�6k�y�g��e+�����/����-�g�
_8K��T0�)�I�VD[ɻ�O�oe�֤�!�0m�ᒱ*Z�����xa1@�Ӫ���+��������ϟ�V�!IZ{�G{���
\둃��;o������9~�������x����qR�<�{X����+�FJDVƋS�C�\iX��{�Tt�=?�W���Vk�T�K�Z��c!!�S^�A넯�42�M���{�|�;�J�h۵�C[?�'����/ ����/[|n����>=�y�<�$vj'|O�A�.l�9��G���>��gL��;�A�S�oذ��;�������-~~X�4�l�֟�0D���dJ��L8ցj��EǏ���	�5�Ԩ���,j�'lT+K��2����ٙ��֟4���0N�0H'�Ux��ĉ=8Y�����q�Xxn"�?2��]w��C�����0��h��;��Qx���ַ�%��ޝ���T�-oy�y�0����]�ش�'��P�̎�!'��Xod�4ʖOѤ�#�$�I�����r#�N�"�(j͞��4Y���ʥK,�a��R�Eƪ�J�%�q�1�ή��d�>�B�%~H�X����������\>򑏘�G�7�����Ѭ�����sj��>�0�[����~������G�O������˭��j{�`ޛ6m�O}�S�؊�M�H���/�5�֫LI����AQ��v�9I�p�(t��XY�_�m۶%b<f�"?�0[×V�/�a���
�y"�Zk׬R/��}�<�G��0�U��/.�JoO��-H�|P?7 �]v��e�>7
���`����"����=��K��?�qz��m��>(H��=컀����{v�o���MX�$y�������ꔳ��,�G��ɤ�,��υf�����6m��v�BG���	
F�X�q��iKu��R���]x�
�,[�R�ղ<��ӪaG�qG��!眳M.�����I\.6r��~`߁���|�8����wZ���ɇ��}�p�c�N�ʎ��q���W�'���ty��"��$V~GRg�d�YB�0�o�1[���,77)����8?�/�ɉ�K�������y�1�_�2�JƻX�J��5*  ��P�����Hދ����-$}��o �?&79�lbC�z2T2��gHzs�}!�
��_��s0��k�:�iP�����y�@��-��y�_����~��,��<4�1j�������?o�j�$+d�X��{:dO'��U���Y��(%K���_n�Q�����]O���s�}��������XИp<������=G^�����1Y�t�\z�UF�p���Y��T���˖�%����bIg���m�<t1$k':>������ :,AI����ÇfsQ�Q��h�gjpsb�#?q�����E�M�E��^@;�/k�B+�\�>ԕ��A�4�����m�=(x�~c�R}�/R��^�7=�`ǿ��կ���ߟ��=_1P]s�5r�7&�W���3���]���j�H��e/7K���&,2�DA��%�B�G�߉ޢ^7�F"�}#ȓ�o�9i��+<���$i$�U�A�1^�\_��WY���0#�a��?���������{����<�B��������0���<�ɟ���gC �y���׿���{��{6Ǆ{�a"$���"S�c�y��j�wȗ�����K�AC�=��/|�K���_�x��s�]�?\,��2��Φ��*��k}�s��z�^t�ҥ���yW��e�^���JZ5m���9�Q���6&������-��A�nX��n m�o��o�{����I�+���bwl�Mr7�W����!�[C52�%����䴾[?e�9���6L�h8f�7+}�
A:��Z���(�sB/D?\}�����/]�tV�����ph�ؘ���&�9ر> ��}�I���JdO?l7�kn��|A�>�LY�r��3O�^j��W�=��q?I]26���
E%9�u���S��ӛx"~��38z�b�	;�[�͈���k��<P��MG���,������gϊ�J?,��`�����C�����dQ���k��mF���d��+L�A��=��a�!��q�Fy׻ޕFrmq� �eq����TM���׾��\W�<e�RД��)�G~L����q�d��F�q�� ZP�<ɚ���7�pú��߿�v��B]f͆�=�Ѓ��s�w���L���zF�����#�=jud�%���~�*&
'Z|X���o!�b���UNE ���R�c����p�v�s-~��
����ϰJ���ߧ�dώ!!�W�ӨI�~��' �q8�^�{���`������8Y�ʕ��?/�m������}�[��l����=��a/���'�}eϵOO�k�ϖ덞�=Syvqs���uB@c�RI`��'�y*1�}0�_��,��y�fS~��{;�{ts�X)[A����g��/�����i�珌o������RR���f\!&Ъ��/+V�2W�O,���a�����zUd������M��0�?�iq�9n�W������l's����xa��%c�rȑ��^�|���� ^�������}sh�֧��I5X�xQ�Q��q�p��S�u����a�ؼ����xp����1i_����5���=�䥳Ё��f��rQXO�+9j9�T*�sCh3:o���뇑�^D�P�B���g�Y*.��(� �<BZ���%�^�'~�i�|�s��yŋ���/s�}��)=ey���>ԓ��~����7��]?>��}$b��Pq5+J�#��a�֭r�X请�[�T�ܷ�LV��l��~y����D��Z�I6?�C�NS���rv�:��\�!~%� ���?����d`�	',V$��.C01���OǌX���f��}�!x�,xp����7[�>� ��O@���͍͌P�� �i����`��%�������7==)��5��7�,T
LB#���~7���$)^V^��ot|,��)@1�D#1�!6�zBPњ�9���0mV���9iı��1{:{���B�����Iٹ{�k�L�/|*&��=P�C��8��g�|�)��1��c68'�p��s�����g���3`�����b`?`��0�9�,{V��y=I���مD�yqo����tp���կ�#����~�~G����)-?�Ž�^޵F�x��\j �B�^1�a�����G��R�Щ�:���N��F����?h�v4n�u�k.�6`E�Ʉ.�ѝ�j����|GN��,X�VD�`#�DՇ?�����w��xӛ����̈́�/�N�`;J�#64��f�Xf��惫⸰��=P��l����D���a�;=\6�e2ˍ�����I,��}D��+�(�yh�IbZ��Vz/��1�ZR�^�C�E��XQ��h>��r��C��,P��J��*(N�p�<��,p*�f��?Wț�ea�8yJ�M����� �`��s�;��|��dqds��� ��1���i��� ���F>�=L�����[z>Jέ��TPիr���A�,�$k0N�Cr�5����ú�0/b����"	,�=91e�	���U���I���p�$q�t�I4�ߍ���X�e�2 ��dŊ���Й78ق���k?��w1|8'��ߩ�����r|�()X��_h�j�Э���q+�D���q|��6�����0�ޜ�W����(`}��l��Ij^+Xb-Y7�0�C\�)���{�� �,H��_=���{�Ռ�3gB��������[�:����\�0�G|v\���p�?>>C�|���S�g7/��J��珠��:#E�%�ߢՇ�b-�o �d2j,�l����&��8�,e�dB��ϲ���{b#h��u��ۨ���?V	�^d}1�0m�� �;Xh�]�X�hcc="��x�ܳ��f�=��C�@�x�Y� a�pQ�R���̑l~q/��(nf��Ru�h?��j�q�)���KH��Й�}V���%��;@ZY�R7��������˾��i��L濓�ϴ9tJ&�vt a������)<�P�<5�����o?gp`�#Wt��Xx�� �\g&��D0֜����3	�3p�����Hl�ÿ*?�M���8����l:cs��17��ʦ�4�e
�,��!�Ű�M|���,�<�߮/�p�=��a�{°�	�<�.����u��3���	�`��&��ǉ\�9|�;�� TuA�Z]zR���w��m�W�@�$��� 7��o�/}�K�w�ð���c0��_���>��ǥ�ǩ=�}�C��
a[`�ִ�o�qӷ��~��k4b���t�7�ik×ʹ�?�8兿�C�0s2�sq������`��ۿ�[��9����p��C�dl�H��!������g{L�F�
lME���j�z�=~�G��>L�'w�3LO���A�������� �+fr�
�f����9�F��D�I�8����6��)0��1<?��G��虑	����d����(L�g}�b�q���sz;�<��6�����Cs���������W���y��<������V$�O�q�8�HY�|O�3 Ny��A}<�`6������b?�O4F3���P���ΰ6B�D�l5���������`��,n��(\�h�}�͖}̤S��1�n�3n<s^�1��;!���Oo��'�s{�c��ii`�u����`}m��Ux'#r�ۢ�+��)�g.|���'�����M�4��h	�0�w��k�w�l��~� 
��
^
@=�io��s`���"�t��|@{�,��Ѭ����_���?}���Ж�-�F�	|�ٺjSP�{|�%ףUT(�ݻ�����B�R=�P����B|�,��9}�d��s�܍ފO[܌��B��z����MFG�J'��Dn�|�x^=(V�2\f?��̦������|�����x�,��I�XC�b~�c6�?9JGR�T+�����������r����>�oQ��lI�l�7\�1L��I~ ���Jȟ�E YR+!�$� �)�1`\0`\�1��]�,ٖUn�w���g��9����;�;��+m��\͜9�-��gW5�?���U+���bZfO�*`A�Ey����.1�l����[)��a�;�l�5�GaY���H(���cQ��p<�-���k��7����Y��{�ޅǰ�����"�{��P�4�y{^[�w�1~�����W� Vڣ�#�}c�+m���?��UuN�W��ZE*e�|Qq�^�-�w��m
c̊;l �����+�u'j����2y��؊S��Y�ąN�*�����8
��Mt?!c��D*d%�ez`�<m��1X� e��8�}[������0Xm��%K�m�p�Z���,��D�sT�����sl�$���.F�<�
���3�56Z��(bKgRzL�Z� ���#�(1p����JX�F�A!Bs��.P�Z�� � ����Fh�ز�N�b�(qL�R�1�B���9f%lR�v����G��9�t�b,��7���x�	���8�}.��sj���ϙ3[Fǆ��zp���A�]~��q��ߢ|�VK��!�дg�A�WD۱�0Y���}�\v��N���Z.)�b	Mݻ
�Ig����uN  �1 @�l��
^�fc!��Z��GX�YL��Iu�����&��N�Q4�U`0��Lm��u,d��dT 2A�q`�)Y�KfNm�V���"��Mgb�:��Η��,��d��r�S��N�	��1��2��Z"���ñ}�5�Ԃ9~�'��ٓ�<�!S�q*
y
��5Pج¦���R����� ����պyO[0�}��h�A�ь� pOj��5HAa�/�OXw���7�Y�
>��,=�9�u.���Y��sf͒׾�5���\���^a���S~6��4I�Ƅ`�g��`yL֟z���Ȭ�3�f������=�ec1\��c����9�Md�6ky���._���b$E��� �a���B�Z�&��D�$�؁��K����d5C
4ݘn��Y'c�8�#0�!5yj�d�8?z�W)Y�O��M�sw��59���ٳba���иy��[�%
�;�.BQg�g��92�����b�3\PL ��X`�cQ� r� b�>�bT���xˠ^-�������G�f"K�L������L�������a��D���&������cl�P"�Nz_�����t����]�O�tQ9!��U���_�����%�8��ݷ�٧䷿�[��t캻���h�)9��c��7��u��k~$/�� �@z��ml�i��C	�z�8y̓/<_�͟-��N����~%[�>+%'�!e+���9&O<&3,ǝx�t��ҎPhG�~lR�?��]�SN9E���_�m�K퉌����$���"2C0	t.BĶ\�ϟ�-�;p΁e4ٽS_�j�\v�eu�t&��Ʉ�&��ǀ fs�A-���.���Q�̟Z�O~z�jRV3�1�
�L�-'ў�`iDs%�0 ��o�a��Dc�p�b}��K���.���C(�X4����C��U���M
e��s�9G�=(ȒZ?^�=p��z��x���S�Źѥ�!a�R8[��>>��kY��f�{B;�3�<ӯ�Tz�rD`3��%q�/c�A��ޤq.4�w���O��|`\<Hm ~���uD�� @;̕+�;!^t��O6��<������(� �z��k�rB����M���;������B��`��� ��YS�  �A�-���\9�%R���}���e��s�;����-�����'w�u�l~�Ey�;߫Z��@�>9�(�t�^{��7����_�z�h�� ��_�<�7�abc�'�	'�0�1�Uc5i=4<S�����8���<�+
�]n�yO��غ	B�q�ʬ���jo��0�?���4��P�h�y�\U�����f�02+�0&`Rt���E{>�#�9s��r��hL���)v�^�����}�m��*��i|=���cM���E;�ItS]�c>)�gŊq۴�������Bj7#��&�׮�S�y��C��82ִ�]?6 ͽO��Z����ZQ{��1f����G�޾��o�J	��P��k�S �,�?z�<��S��9�;��~��<������ʍwEN[�T���=�|y���Um�|L{�6���is���渍}�G�s��;n�#W-��;�ir�ed�_��7�G�B�� �<ޠR��6���>L:�p`� &�@7h�hm���7�u ��6֯����t�n�6H���b�H�9��[_2!0o��Q���vM�ic�Wۀ4�),,tv�����b_./]td�60=Q6�2dtn��|]O���0%�źk+_p>WPE��@ 
��1j���0F��gLJ��͞�-3�5�y�:����S+�A�ҹ���x�Y2ѵ�?�k�
,�Mco�8�vp�úB������WW0�� ���|򓟔[n�E;�q��~a=�=��?%�g��Z(7=	�(�+ȩ�Y����W;
._v�
�#�X#����[;�)W�N{��,ϟ�L��×����twed�K/ʑ+�Ȍޜ̘�U(]��LAd�Z��c�ve��21��܅	�f4�|���Lr��.��b5��XsP+AýMt=�O�m8������l���7HR�M4�z
�����Z��q]��O����y-�O�I��P�4ux�
f��x2Qjy4�q��lf��d��k``� ��x-��6�)�`��ٜf8"�}#�$÷)�d�xv4Ɂ&��r���B�)����^���Q�̙׎!���ϛ�}p�����Mg���|�l�5쫽�?x~�g� pK�.U��������Ö���B�p(��7��`�6�>"�g�d���2w�wÏ�X�hA�����-ȝ��[/\!�3g����e�aK���Ti�3�f�����F��;G%l��-۶=�-HA;F�v�;I���[yL�|�8�S�`�Ϛ�AƑꈺ
�����_�1����Њ��翐����̙77�Y??Lln��I4��t�������y�|��Ǖ�=&���s�E���q`�b����:'s�)�d��]�
�����X��6��f3ڋᩧ���$�;�L��ܺZ@����70(���������3 ��
w�r���)�C!±��êD��fy��6&���঺t�z���?�-/k�P3��q��d����a�ARY�.*úRk���M�m��b>���*��C��MoR�/�� ı  ��s���^{񅗜U��?�(�g���NȎ��q�"�q�Y��ky����.�M�����_|�y�Vp����h�3�Qbb�v�ʦs��Ckԁ��lJ��ɡ��c�5�ӒqǏ�n���Q�ƄM�F�^2w6��d��M�l�9��=a�a<�,��5*���V����O�qܬ`�}um:� �^��8��Ա���}c������cj���6va��Y"w,	0�fy�,X��F�<��gצe����%ƿ'"��®++���I����"�f�q��ʰnЫ�3���|�󟏳�p����ަ�~�/��8]'N��#w!Z6VkN�G6W&���J��`�qp��)�t2���5�6':b<��O��B
d�8�ȫ^v�
��g^�Їv��wҵK���ag��iSK��;�ͬ�X��p饗j�j��@0��{�y�7d�gf�X_��$n4�dL����J܂�%6�f7>c��L���[�i}��\N �1�c5P�l=)sh���8�3�+��
U��-�i�67����%%�k����c��4c�v�9�|>S2Pm����#�wؾ���xnd���_��j��v���������g?��c|i�0#��B����3*�rF{���ު��yi�Q�@]�iY��-�Ҡ����S"kHR�0Г������x���	�_��	�/=��=g�̞��i�nӧ
jrժ6 ��K���\�Grd�5�ό�{�G}��}�k��;�6rva~�+_����7�f�Y�n�6���Zs���u�-cO.�F�d5�fZ0�ϑ<�-@%���Lx�d�Q+4��B�g5|^�~�8s�h�Xo2��˞�ײ��^׎�i(�~3�k����K�}����J���L�eb���e@7yO��ܛ�k��`V���뿎�'�� Ա�Y���cb�
�×.��b5-�l |"B5��I�`����󥧷�E�>�E�B��[+��q���?&o��5_������3ϐ�;v9F}���}��9)�#�fuG�+9YԻ��Ԟ�.+V���-$9Z5R+����P� r�!>����>�1�җ��ھ�ٸ� h�l�7�'%�o�_��%��̈́�ua�sY��M��Y��t3q��2jF�1w���|�y�6Va��V�?��y�ɿ��������
�f�׎5��H��9��[?=�����co�CA`c1��j���]�E��MaGK ��9���{����p�����@	��dՑ�ep�%���B�L�vVB��U�Y9��3���k6�G�@�>�X���$޳�0L��P�����\Z�{��.7��{�L5ǰ��966$4fϤ��v��r��r9�����0�M�6�@N�h,��.�*`��?���p̒a�������,m'�!��Z�e ����2U�:HZ�>�L�j��Ѫ�Ԉ�l�E���&�߼n+���&yV��3
C+x,��cb�Jj�,���P�ot�V,��{.�Z�1Ѽ�m���B���(vC��;3߬0~�ޠAw�&p,���:J��,;���T�Y�R)�M�1�h2�ͻs�e�;�s�tǮRK ���[�QQ�k��:o�WUZ��r��r�mw�+/8_F�Z�d���"�������c
]r�I���^"s�-t����wOp���_���wj��~�� @̶m�����l}���bd���w�/�9��i�$����ؤ�8Y�����h�[ �%��O���ǤO�5b����`�2+k�7Ҿ[y������3��cac��ڠ�T�2�F�9?�ț�[]TlƘe�������v-���������KZ�M�EV,y$s�uI%�{��塇�SO^'��,9��N����]���������b�r�y���k��r1����]�=*]��b�Dn����?�?I~� �'��?��P��c�s_����\�������ŭn�f���9��8�U��� ����=�,���0�9|���*�׮Q낛�n �q�O"^�D���Í�{�I�}���=�s翭��U��H�p�m�)���p{��>R��粩�I����
~N렙�k�u[��<&7�s�T�Ɉ�g�xr�W���Z���fa �?��?W�>g��f�� H��;{��\�J
�9��3�UGɖ�7��� %��L֬^�, �SR9�%��#���?�ŝ5.��s��V��=�oF~��9L��\u��w�Z��	��9G�Ξ[߬nB�ق���u�}/�������?��?>G�=��ƍ��͛b�.d���.Y읤o�L���`l�2�F ɸ,�� �����>P#�ОR��Z�7I�����ͮm�C��7���jF��1�&��~��o����a�k�m��k� �}?p�Dw�2��ـ�����A��
O�������7�M?��gH�[����I'�.���xP�]#x�P��n����:+�?��� ���S|�����^�.`g#0s�q�)�6�}L$.��6l�GyL�=�0���l,�w��ݺP�@��8��?��'�.�={v�;5�v��� �8#i�X�8��QV�>D��`%�ka��}ٲe��|�f=��E]$?���!�ҽ����{?��b;�q��b�
�'2��/bk
(N���=���Nhx��g*�B�z�N@���u�W� S�7C�vI��}� ���u� (��[�@ ��>@j 4���|�Wj��Ƣ @�> �z�ߨ��XP� Y'���
�/Ns���Q0j �vb�:�S�a�#U�C��Z�@�E��x�`�Ŷ��a�Ê��������C? �;aR�g�2�*j�V��R�r�_����ө��N�N���G0�Aq�"Xa���&
�
�Dj*�7Z�����& x!ЋB.��~�a�馛tB�����f! �:�����Ad�eQH�F������Ƈ��Ob�������ܢf�+����˿T�
�u���� �l����3}'����ξ�}o��4SWÈ��aӞ�7���<`pA, �xV2ٌ]@�����t2Ku@+[}���h�$����=����;��&�M[#=��"3�=D��`%��2�M��1����������` ,	��{M�E+�?���� �֮�����[��gS�q�FA:OL�g��|�8�!���Zq���.��-�3+�S6�[ڝe�������XT>@�"�EĎJ6ۢĸ�f��%����{��E~���v��!���p�0����}�s d3�\�f��dVF*^ڗ��BOlex�>�k����PZٞm�g3�OGn'���R� oZ{�z�|��K�4���E��v���_�O�ӊ� ��XLHE��׾��* �o���ЮۅZ?�6����l6������=n�OX��`05||��O�~��/����f��|�+V|L�1`��
�y�@N�{��LZ����'���D�i�	���g�M�����]��N@*=��"�Whְ�̜Z�L>�����҂�}���"J���4PJ�$FK�f~�h��)��ŋ��� �������E�<���5�O�8hNcކ��ֻ�Ѻk��`������ҩП����/�l���m	2��=��f�Y�E�3�#�^����7[�kB�q��>��<]�A��{K=B��/��h�	�+�@�J=��~�z*�׺�ƶRZ�D�02��@<V��oP� 0bҷ�ܡ�$ѯ�ģ�3���(��^s��=C�;�X��e�M|*���y�X���cŇ���@d�X��Np�=�j��e�,�T}+?x>�r����z�����β��J���촞,Vp0E��^)'L��3��� ���ZM��N� �k�]�ijn��1����� ���[�)����U�xR���@�琡ں�d�� (�$Pf�AV�K֊���bƎu��,�m��?����[z��]��]�"~�N��sLg�S�����L��aJ�����[�!�hzІES�g	�,w��ò� N��G�x�z�"��Mz�p��DGc�^K��s�0��շ�yj�48'�o�vl�
ٜf̔��fh�K�k��cJ�RHd��E�ð���;GB'�*��ҹ,L7񚿿�={G+Č�`�Kѽ�:�e�J9�-��0�}G�����/�K�_���71H��t+�Aºd&W���@!�%P���s����O�Ly<{e`�����R3EN[�"#d�5~>�,j�_���ղ��T�h%���󟴁�����5�)*W�:I�5`/GЭ�jݯO���:�m��V�"s�����M�DR����A����YRp�*�����O#�F�;����>;%i����;�̌��B�t���<t�8�T�u�A�,��|���쳲t�ar�y��9�,����NP k
̿
�B�1�ZQ��[u���-U�W���H:�J_��|Ӎ
ّΠ�O&������q½w�*�8>��F�,5��}E�_0[Z�!�M��(`�x�����T�|�[8��dd-�F�t+�L ���5x�*nQ�O�[�,�EJh���i��C	�b$@���ה�����3#n��H��V5���v�I?i^'K��6ɓ�k~x�Ө�ҋ����n0f��i/�]�E�Z��eo�_J��ݲ`�|��;�i@�R-"���4�XK2�Ǚ��;�4�Tg������E(�� ~��3�����	*���䶕���fc�nӹ�̘�#��,�o��Kp;���@�FF��B��2P$0~:P\=�p���&�L L�%���SH4�R?�J�e���GX�z���zu�R�F��z�(�<nw�Z��k�!Ϳ!�}zٰ�1�rMq�1��C�n�u�.����(���}n���wO]���mTQLַc�{Β�YrQ�?�}�i��%g�h�Ϩti�W�� ��,�h��~{�/��Iw���Ԫ���^ɧ�B�He~xǂk���!��.�9&0�"NVkS����g�?W-�� ��T:$�ZY��9uE�
y	�Z��Q�����"�XM�ʽ8U���Gx�LCf=�Ex%fՁ^����
�6k���Z]�&C�X��w�8X�*��4Ѱ��������5p��A�=4|,("+
����n��w�1�Ë��M�����	[���b2�}���G�9F̐l�G��Uefź�5W��xn��3��*B�^Vj�蕙s�h���`���%�<:be�7���9���gܳ�z�%ǐSmdD��i���ԱgYcN<S�FS���	�J�397�9't2��S�b���|�ΠӚc��D���0�FOk���`�׶4���E~�Sr�'�1��؈,�?_+���fb\��B�W����6�ӰKQK�\1�������>�h��[�MY�l(�)��ŗ�RN?�tQ=0J���>�9�u���jr{ٮD�dU��Pۣ���Į5.�ae����$К��������1�*�����o4����vz���hmX�8m>���T��y��s�Nh�Kge�1�.�}%�I&�չ��v	�4CrZߝ���
��sK�{�.'�rRvB�\)�X��!˖.�MO?�kb;4I�4����9�:P�%d�̘�#�'.�Ŝ�3ئ�:5�3β>��3��sϓ�n]A1�
�`~u��ZIL�������}M{���3hJ�ޞ�����sΕ׿�5Z�U.�jZ$�%�"r!k� Z��|��_��6m�tO[���i�j���+9F��c����qV����U  �"�;E��ct%�}���p#�qi�PkN�h��H���tI՜�VH���G�2V��ʘT���v�;�0�B��˘ȔR=5[��-Q�eU�⳺$����L*�Wh�1��~֢� 1,�c�����u2 69gS�|�Q��ýv �Dֿ�72Yy��ީ�������ݏ������w) ��UGʯ�k��m��|��.���D_L{���(f��)��"W��M�Q:��M�T�n���"}�}�`��Ys��Xy��dg�q����ۿ�[\-�I�$����?��?��~���'�&�ැ�>L՛����3L�Q����n仫pH��X�� ���{ѣM�8�B������$,�J�����R�8�;�>K�J-3&Eg%Hۚ��}G_�'�jydB��H�+�Vk("s>@�T�9�WM��+O�������5P��n�U{y�`2c��݊{���P�t��u��l�e�{��J{'��I��� ��Ś�~���mJ�e K�{�ʕ-��P�9�����K��a�ڬ?޳���1�������6Y�z� ]�/tV�}�<�ݼ0.,�#�X��u؍UY���Μ��f�k�<2�n�3��ɾ��x��*K�,��^y�t�s2sV�lټQ~�>y����o��Du��'�g��Qǜ �ן����e�]����s�9��կ�a�� ~�t��o�]���oi�7��Y"֠��h�M�{J��:t�F�J��8���0�i��U�V�-�·��L@�&�]x���>�.�2��Z �4�`Yw���G�1��%���R��ߖi��Z����tYw�M��.ٚ3�L�%�J>�M�`�<S-z&]BG��Y+�b�St"���H�<@� �
{�9�����p��_�=�0 �/��r9�5Z̈ڢMO>��Z��9�:�v�nY�r��~�ٲ�5�,��;Y1�  l��Tb�Ӟ�7#g89�c�`h����Ҷg���[��#����h��Ӣ�����V����}�yH=��3�_ߩ�`,
hӐ�-^"7�|�B�b°@������=��3yV�/j+,m�7�Oj&)��\��(�pZc>�6t5#���K���s�������ˏW&���VI;��7橥*�ʨ� ����^��� ��J�$�6��d۞��m�62(��j{�&�M�&���70��ɸ�M���?�LP��ReS[=K8�N=C������rꩧꞇ���/��b�����=�ZE�ݬ8��ի���O�տ�rܼ�Qyⱇ����+�?,�-c�J�������ΖSן�	
�7>����r��^'t!�)��g�M*|�Y��*U��a��淿��yY�l������^ �<�B�ᑊ�x��r�jY�x�Jx4kA��>K,��[��Yg����������?_@<�І����tM��{*�aG�Qq��|v�P���@Z�5rbld؍u��AT�&��K�?��?A2�j�pM�R�Z��u��b����1�q�5W��ـ!u��+�Ȃ'2���2:��0%�{��G�s[�oߩ�C�c�ȯ�JH�H���%3��;:�&�e1ЦA����*~��R;�1J�C|�d��?^>��O��c���Au����~m����^}�,�x�*�]��2&�f܊*h��wUah���䦛n��K����T�@�`~[p���nA�?'���eK5�6�Ч�yR֟r��.[�̲�8������;�\�J���>���;��|�n:�k�qD��"��w���՗�n��F] X�X�����$�)n{N�l"��tE0�6N �̘׿�m��RM�-��*�28�]
��#�$��|4�ew*]S=� R1��B�3��0��V��!H��ޅ�S=}͇w�x! �P�RtLi�c#���ޤ$���j�I'��4A���?'�4�� �P����:��q~��~}>�ʗu[��x����b�Y1�2|@r���2]tP����	���к�u�E�{� ����/|�ʨ�	H���ʕ��yxý�d�Y�h�����;.М�+����s,�����j�W_�Z=Ǌ+���v��V�m�3�fD�����ӧ����s2:��&bT*U=e�\q&fyX���� }+����I��,6Ӯ]�T@@; ��{��^��0�&:����l�@�|e�@�t&u��$Ԕk1��~���'^>�rԴQN�<&)7���ՃYb��`��s�"��? ���PqO�ӵH��"�Зz`�0���T �� i�C��F.�0�Ɉ��9�8K4ɉ����,�KNͺZ?��.i��F)d� �8X�\�{ҵ���<7����ۥd�&�O���x(rK�.�7���կ~5{Z`���Ν?~�ȥ��m��='�4�n��lA^�a@�c:�1}��}�=���/����W;�0,���k�Z Ӟ�������g�%cVq�3jv��	(9T�l�riDjUg�� �3�j-@*��ɬ��^��T쟋��O�S�����MDs��K����[9t}�"���BA�cHtu��m"�����h���͂^
�ﯦ�W��UV<� 5����%��DA�v����Dh��T�sBp�v�g�����^@���MnR[	�,��-n<�%�y��$��[�&�̶K�G�;��y߼w
�����a,��If�gc}���+�}�ϡн�oTW.��ڵk����C'�w�Ճs ����~��R��}NX��Kh�@JQu5�ᾃ5��R��c��S��i���5sa.1����TN�xs���������� �����G�)Mgh�0����oD���h��Hjm�ק/�M�1�8��h?��f��>7_ǄC���Hۍr�c5���5��w�g.�CuL����!��(����
����gS#��S�o���#_��Pg)�4�S��8rt�(�ã
+h�M�L-�W�g���p5�����M��mj��NQ����Z6+Ǧ�RC��kƽ�p��a�C�>�ǴK6k�����L���%��O��
=���NS����}M� ��e�ݧf���W�������og+I�si�	�2:6,3zg9!��1Z��JM� O{�N���4��]2:R��+��KfΆy��4�R)#]��NW4ҷ��Ȁ/RM��/���1�!��W�*2!R:i���X�h�UW�}�&�d�%�.�OM�����2���̛�)դ�������	c�"恳��+ձ��s"�240���,p� ��F-�� �vL����W��uB�-���5�SH`��J��[T�@� X.元fi�����r26<�n������QAd���t��y�Mx0Ƥ4VԂ!
u��y���� ����|���V��H �:�<���$�BbO	���^�����تZ���x+��o�E�������[������;]W�����E�:�(�\a�޿��䆛n��R�6��4Ȏ];=�������e��Ŏo8K��B�L�o�ҘS��&�/�X�ם�>��%�Ok��j>{B��BӞ����cOl��O<N�֟z����K��]n8!���M�O�����)�y�n9��T���7���>�nL2���ju��
>Z�數Mls�4��B0��dұ�b��N�F�r�i,��1~�؛׮�;7�_�j3��+��(4m�<���������x�1�Z��,��9�|V�n�T��L!�'��Ouų(J(�Jj�D�%��1�����J��r���u�:DQi�Ϟ>|*rxG �>�|��?u���آ��B7���;S�=�x)�������~�2k�B�(��E�9�,��v�ˮ�a9��ӥ��[�d[�<-�7=%��yiFmߠi�bM��0�P�q������Wʖ�7��%-ꁦ72:��9�[4K�=cr����J\,��^zI6m��4�L���ze���C�c �yx�[���e��D�����[<���F͛+����is�7	�-��)t�E널�H�<���x���b���{��k��KP� �Xq�1Y'ra�Z�g'�Tݴ �\r��C.���X4FS��f,�mړw`Uſ����ܠL��-tfKe|��������b
^
�hjd��<�%Ō=ya@!���lJC��'?����}�,=l�<�н���!w��S��d��T�Ȃ�K�R�ʪU���/W�cht@�{�Y����'�i���������=�������'+^�����A��'?���~�+SJer�x���կ�E��Љ�tG�|�4�p�򗿬���1����?�o8G3��

ݲn�:y�Wz�(���3����w�� ��K;w�=�/�n�VՔ���)�zqc��-�1�7`�1e��%U ���6�H�1��z���l�dr�,��F�v�m�]�WoF{�jm�"z[�YhX5�a�k�E���;����d���3&�̝׿��qj7>g2�7��͚��{�Bb�ƍHϟ��.9��u�םr�-�r
�f�UK�\�]
/���s�=�Y�0Y3���Ɇh�QOWs�"���_�d���85nH��{�1NS^�����i�ٴy�j�k�>F�S�1{�cZN#t��-��"w�u�8�%,x��(?\<G}��@�lذA#�H�1V1��%����u�a�d8Y63�L��E����X^1���%$������w&�3�Vא
M=�ˠV���/�Ɯ��%��,��ze�PU������vR)�j�=R^�=�ŷ���yki���K p�iphX7�:��(7]�t&j���U�}�L?��u�?2�Ps��B���ه�d��{�ys溭�-��~��Y}�<�Ѓ�e���e4&�~�z'4f��pEQ�~�Q���~���.�ixƔ�M�;5i�D��	#��������G����n�3w�6MX�t��x���#%�Q��M7��Y���?��?V�����r饗*x2���
�Bї�a����k��ry>�b�����#��p�t��h���6�{ob%��묍�'}�04l�!��2&��(/>����%ya��̎T�U�3�xr���'��3�>�<';�������0S��rJJ��t���������MU*v/�C�&Y�$f ����Q�����5�X �:R������D�R��P�|���hm��×鱳fg�.��pX[8N��s�	���Oʏ�cy��-*l�u�����R=	�06R��z�t}�Qg;M��x≲b�2͂A:&�VKI�1�ǞxLn��V7)��0Y���DÒx�k^����|��؝��я~����.�H���!@��Ru���j�2�L./�<��|��߈����,��b)����3d=�:X5"NۥޞY280"w��^M�����ל�)���$�	��������f����K*�U��x
�?��<�V���w� + Up�A��|Je:�#a��Y6�-�h��m.c���R�h� w��m��;��"�}�yp��0�];�� �p���9��p���(bo�xޝ�~��/�����V�i�3�s���B��]�9�����a�͘5S-X(���v3�]��eǎ��s�7��n�219�D�Ϣ�|`��|,X��H�p�$�7p=Y�f��C�=��(\��	��)bQD��!M�+��^�i�t̠���z6ױ`����Yݕ�\
n����K*'�3��҇�/�dj2�/�
|�.oqQw�s�V�*�=�1�uTS
5S*Pl��gZ-y����>�O~��'��Q�뭷j���ɟ�7����"o�;�Lxf�32tː
�U�V�+�T�`�=�͛6�s��
��JeU��+|a_s~�������QGZ�x�	>$F�ˣ����;�駟�A=)����Ro���(s{Y�?�����%D�V���3�tG�ԑ�j:b����ݡ��s���q4{:=��u*�����4+Q�^��, �U!��u�⎫��X�`�)�RZ���L{��)���x�P-B_��Zw\{a�{\CP$�V�����i�v2-��
�\��tF`3n�v�&.�)�դ[ (��<?�W,�u�r�9x1�����~��T�����;��P�
�7�7
���}H���'u�m�7!]����e�6 ;�v(N���(�5֨�)�u��Ti�R�
��ct���2�[��3|b�KVPE���.0,>�>�я*C�������MM?�zDqd�"��Ͷ��m�����	���)��5�`�&�mj����}��
��_�����>���e�M@���C1W��+��̰V����;0+2D
������(�m�ʒhU�ձ�x�,f����$i2&N�TiV��Q����;�
|�����a��YP������K����BRp�"	�Z�/x��ʑ���u���ǫZ���p�=�oV����2e���#�1�1'��X���7n� �,lD,@��p��#$�+H�0գ��(��[�����ׯ��E0��[�'�֩E�X~c� Ўc�k��{*J�4g���Ƨ��Z�lJV�-?��#d��B������g��WŦ��*�����ݽ*[�`tP|��`��[�S3�ռ���4{@TX�v�=5��A�'�GsX���D� �{��+��)�Uů皏B�.���f#�i���u��g�惻�o<%M�o~���S߱���ޠ��WH�[|�����ˊT����R��~���?92a�����7��.�`7��CVӷ���$Qx�+ΕE��-*�?RG�"��K��G,j͚5��!��$ԠS�:g�&���I'�$K�,��<�ξ]z�]���F�3�=n��A������(�!g����y����{$v����kt�ӕf�(���\�!�P�nӑ���h؉�9�s2���qI~�1d�5TZ)�̮`�O�'h��8���K�����e�Ų�[c��/S&���b��[^����Jf��9\���1�w��}}����x���'1��Jd��] M����?�~Z����&�?iER��4U� ��?��UK%�&�'R}� �糀�����8���?1q��j9��3�x��`m�r����JVp�E�s" ���~V <|��u?P�������O����_��3И��5�-�	9��g���.����C��lAl���0�B,\ &���R��o�y��q�Zf�� ������1ל|��˞�:$���#�v�
���h��&/���od�=���2�aЗ!�HZ�E� ��v�*כ�[�xOt�C�h-
4SɁ��"d��פ�<Y���q�����cQG��e���n�p�?;��x�y�6���.� S�����/L�s&�SS�i�������:9�c�o���8��͟�b !(f���\b}pS��	;aj7�ĭ#Y�x���,�i#��=�8k���� f<@�bQ'��*���@{�>�V��z������RKK��o�
١�B����z\�`��7x4�kLW�:�dĠT��ֱ��!�ݟ|�ɒ&c��;��,$4�k�'
��-Ȅr���wr�;����O� �j�������>�A��7�U2��2a��%5������.K� QK�o!�9�,*�ֱ{O�ERs��x#�_�f��e��߇l��g�}���ek�a܆i�w�駱�t�A�̔?x3  ��IDAT�^b��YٴL2
�yR�d�N:;��e��K�Rq�!2ie��t��h;tY�	�;����e��{A��B�;��ĽMal����g�F��_��EAPW�gQ�2�%��w��V|��hL{�?��'��(%w���b��	Q.U�HWf�T��er��q���S�b���Q۲B�fh�o��-)�*���2��)u�XF=�9��ŜC1�=dD��itD�*�cΧ5O	�^����5�r
!�J���w-ܝ�m����):^�Y��Vp6Ef�6��rkѻ$�Sѻ��lΤ��9�c�y�f���oM*(��1?2,e2)_���	+�5��;\3͘';e1œ~ ���uL���je|FQ��3
N��P-���F�* ����;����K����ɂ�L���+�?,]C��	���e�<V���A)� ��|�7�r|A*���3~�<�fn���$b~���Iiyu�7�@g��bE+q��2����hS�#�[m��G�Ķ����ٱ�������?������}t��� 
�f,)�fY�(�R��|j�A�B�C
̠�3kQF�z.�&��B���|�)�L��g�5{����m=L&?66o\\{FO�2�z���H�g��}���̦Y@6�+LE�ء�Z�z��`�z�S�����l�;d�螱��{�8��Ne��:���;�7v��9IE-3٨[w</P6�b���B9T�#V�/m[.M�ާ=�o��s���DE�:��A#�#��/>L����64]wf]��m?�mMlLl�v&�mۙ�v&�m��}�u��9g��]�]]���[g�֨ ���p�Z�+(i���Tߖȥ G�M�qdM��2�0'��^:x7-��R�af$eS�[���"*D_٢U����	�&uj9ad-Gv%N(BJ�J����
�ǎ��B�wh[��zZ'.u	3��c$��6:qd�l��&�%�#^��V�z��˚93�ٷ���g��Sq|ܥ	���ʦ�&�8Iz-/@<2��TG���<�߬[��X�j�jZ��U�������q~y�J4C��h��"]�j����R{rU�R��4ǣ����T��9��w�Ļ��<q�;�F^���.������LT�"� =����<4ƙ��+�����"�+1�>��T��$-�*��y�D5Vr�{�l�:�r�Ԋ±�Ey&�����1��d� u���b>�ѐ�N/�7AaU��R��o�tY1�7㻇X���pNcf�Ov>6��þ�p��wH�\��lI�`��I4�+�=�J��!p���s��ɰ�F��X8E�8�SԞ0o3Ĳ;(�w$�J�0�'�%v���
������ 9�:Lf�Wew���c)����p�"Ϟ�Ê����Xag�5&A�H�� !O=,��{�s�Лπ��.�ga#6�J�	���������-�%qH>Z���ϗ0_rP���R��٣�!��H�֛�P�E���7>�ic�����v��:w�:�I$W�kj�o�*w�[vq{��ͼDM(��ʗy(�S�}.�AO�?�p�����i2 X��MB`<���P9:�1o�}0h����6wp �4�\t]Q��@
&uUS:F��f�fD�*��y��Q�y�kSnq_�W$p�^�����Q��R����^�_�<q_�e�}�B	���N�o[3��!#b��V��.�e���	�Ȋ����~��e.�a$�j�\k�����l:�a�K�8���d�X��y��e���s���	$X��D����Y��S���p�?��B�i�)��F���Y�*
P`:RQh���e>��!�mN8�Ev��q��B6�~#����3�-F��������2�������ҟ� �R��U^��~�+�^?p�������濑B�����ݗ��o˂Y�Ws.a�J�b�Q�hT��'�]��M36�U��4C�'G���{wj��r��F���!`u����y��)U���>�a;����f#���UԚ�H6�뎛*S%�;ڼ<��3�Y<K�6��������C򬷟���d�=w͌�c����b��e��q�(_��1'@'>+�>�]�@���m2�ΜY���c*�x�z��T�S嘎���Me���Od��3ǔ���˭:h�l��1O�k%��S�:��쬧��SZ�ݾ�]?����S�ܽ�E�/�	�\4�M1��6_y���d�j���Ue1���ѐ��Z���,�j+b�4W��d�aɞ���D�����qAL\K��_@�q���s��Zn02��k�4�\�k��<6̵���[+&�$� �>���k�������� wf�:�V��>\�e���x�����*�;�M����F��g��K��;Lyk�����Fe+� 5iQ��.����4�������/1����Yj�4n*�����u*�֐��P�ɿ����w{�����ϒiF�7?=�h��.�bW:��Z��.�� ��U���ˬ1�x����Y���Ԣ
�W�ߤzB=Y�B�^_{��9|vڤ���%LuyU�e �-r��Jڷ���n����(�8��rk6��q�Aec�\�L���o�*��DP�m&O{y۹�o����8�3���Bi�H�~��P9�������/�*����3�%�#nR��ViӞ^0g�>D��,e�T�}�:�9�i,&y2��^�8x�d���4U�pQ�0��8a}�K��``������F[�2c�K�QW�n?���9�>�~?��nkw��-��������}_��}�8>�i���J�� +��L�=c
�+�X �kdw�4-�
ʘ��9I�b?F&�s��ל��本�">�IoL检�*Q�[|�ɖ����c����8�&,G��d�}wJ5
	;�#���q��t�� ��{�P��w�-a澜U�� ��@	���?z�˸KN�|�}���͜VK_�Q���?����ZE��~��}�6[���f�f��ߟ��U��0Wv���c��Ev��Q�	�YH�"�W&�W�B�xc�����RkV5�-��x���������z͊9[w�<����e�|Pi���R�<��q*�,p��*6�n������&��R��q�
�v�s�z�q��=�Uv��u��\�'�������i�H@7���I����ӱR�V�֋���q�$�+�Sw98H�t"�y���ݳ�|�@�ٴ�p�+Ŗ���P���u�m������Xzl���Jp�� ��B�m���=%����:��"������&k,4�}c��I KW���Y1�dx�O�ϓ��zM�>�zUn�Hv��/x�6�XE��S9�	O,�����PP"��i���(BZH�]l�n�"�Pnr0�i���b�o��$�Ѡ�j�Q���T��.��Ѵm�~�1>E��浱se�2^��$��w1��P�h2�Dt�oh6y��:ltL�3}P��<2����t�	�/��N�(��#x�bL�����Q��?0RI~U��?&[g�3A�� �M_F�I}7F���}a�A[m�/���ؠ�p��o�qD6-"'�_��t�_O�ze��sT�妅�t[ބ���؂v��~`��Pq�)�)��&�鄲�~�2-5ڐ�# ߫�D[��QH0�P��e~�Vy�I��C-�L��Lnk�6�a��s�7��}օX3o���b>UY�3}ف�u��ߟ�V� ްU{���@w���C�t��t^��w�*�gH���Y{iǑ0�\��~X��6�:��!�_6[�Օ3<'lߌ��>���'X�&Yy�4xOʕ�5�M�iDc���`���k�`�0qA	�7 ����I0@��w@@���'3��: �D��q6Ap��uX��R,�7qş� �N�����9{	#v$)�8���Z*��s� �������=�[�9�[yK/]���ZI����.D�܂K6�M3��,��r��G�X@lv]��.˹]f�S��T��,E�pQxོ͕K�m�'o�;7��\�1!2z_w�lN��������� ��&����v[�a����Ƀ��
�d��-J�����,�vUP�?�Av'���/-S0d�����l�2K�A�ړ���u�N�咕���N(����j]���O+"٧6�<�O�7��$ޝ���L���,^!=60��E�9��}���agM��%�O�4���b�ˁ�^b�H�{
P눻�#����v>iX3��#W�^3�_I��r���I�6�lc�����p��n�2��v�����4(i�n�d�N�ˢ�3ރ��+���Ӏ��řp.p���c3�]�b��]�5\'0���ۦ3�C.CS�k�[Ҋ(>{O�&1t�/��ȹ��f�{5'���Ϛ&h&���o�^[,.g�t4���?�cbm�P�%����X��'��ۧ�)z��
��7^��?�{�S?w�)LК�;Q:�3�z:,�13،J�toI�J���{7&1Y?���=�����%1�ޡ���V�p��Vè��M@����8��_����A�V�F)�ĸ�ު^�WՑ���*�.ܙ��h��c��|���DlJ�S}Π��ӊ����?m��,���T�&�%����������{�N�m���#_@Gc�ΙA%x�����6ɸ2���
�e�;���,��u�2庫���������~a�/x�IMyHvVb9�6�^��̨(\��O|�*���t'�l��U���=Y��?��P8g����^i?�o�Xy��3�"aZƟ;XGT-Z}����wy�f�o�侓-��Mq��lL0�R6d	�_�V��1$���i�c�OB�0a��� @b���2 ���i~*1���/�/I�M{�����O��_�y<?�xJ-DP�����qrb�G�ǂ�������:0��D6�:($�#���%X=�il	q��%���}U=�MG*/�~?�.�WQ���^w=��,��$*(?���.�����!Dq�*��NI�<��]�ǥ�T�8�7,F�i�����\�W��x^���+7{&����<�`��;@#��Ϯ�,h�/�s���K@��e���I�6U]E-�pj��a�58^$[-�3��.��e�$�������!ѫ�l�hO��91[=պ���\l�&@�u�2� %?�DX�s���bYow�����H��i��l�">V����B
�+0�[�GAKI8	�m�[�@�Q�̈́�X:Z�X#�O|B�@X�^���xwh��!M���E�q�QAsJo�e/гInv�{�������a�(Wi�5�>ig����}M:��=��b���W>�����Є�De����+TǇ�	t>;6�y��l9�F��v�6�������W$J^7K�W���`!r�Q}��%��ƶA�� �q[���� �A���M)�]�j�v���C�ڂ����ې�oS���bg7���C��|�خJ��}�h�=u?�.�E����Sr��T�ݸ*{�ݿ�%<:j�ܹ�o1i�y~5�Uq�d�D��kf���_�rAc�����śᅟT���I�}�a&|0e����?�6WN�t_Flr����1�y���?��(��f6�����7�[l�Gr#
��I+7� �Vk2~����L)��z�EG���x��W�Ӡ�~l ?�-ؕ(����Η����2"�2���ԩ��a�������(�Q�ffe�A1,�f��yj�a���5F�j=���^�ŃS�_����{|��ҎOj/ ���=�p�6�4ͫ�B�+ͬ�`��[q�MR�Z���S��gt}u�|X��2šT�W���#>� I�C�v�-�r��l'O��__q6V���N����Gw��1��x�����y���pP�Ӝ�鞐��ogiVģ�A`ZڻJ7�8��z^���H`�L74|������6E�P���GJ>DJ/\~6�]M|]`2P���q8T���lF}>�g�����6ZlFe��M�2�´�뿁�g��c�����Tڽ�z^�������s,�����|2��/
 >0�����mp��D��V���#4������ G��4�	�iC��Ԓ��tR�L������P�"�
S���ڷ�ڕ�&��<'�����{�c���t��ð.���Y2C��+r%̇�f�<�0/c����k����և���� E/-F&Pɫ�{:G�ifm�T]/����$_#��s�lBi�[��^���R�Eb$ZiF�(�#�TD�4x��F*�$�����p}��R��k�X���n��E�Gs�w҆�<���=��͚��;����e}Z���#̾�!4���)���	p<�v�0K&��\�M"G]Z���gf��?����%���7`h��.�P����m�ҵ�}v~���B�4�����Wg5���g��|6<�f_�=�i�;Ё�t`W8`}�� ����Y�۝���^f xsL�=��Y:��W�/�2햌nr�r�w���R�A�[���T�b6N�m�X>�6�.}|q�Εf��MPl�O�+�Y���R�oQ�l�U�.�H�����!8�'Fͼ"�EC����)@K֓��lY���q��H���;�^�r?+��/<տ	>Oěb ���i`�n @����`�!X�~�AFepB�04<7H���Fh�ܼ�iC���$�o��0*B`��oScU�<�K�*��8�B��Gi��'{�"��ί�+&B���V�`�j�����& Ͻi��*+�|���4e9��4a|�����������93D��;s�*-9Uܳ���$P�O�����*ίv���!��?V-:Dq�y�0�O�G�<@_>�nyo�X��D`;\L�9����xQۂ}�;T~��V@�(��4�ܰk�>��T)��1��?8kMi��Z8?A����y�D�!8�M푕�4����s�2��29�3L{>��q��3}z����8�-��L�Y=��@>�d�Eq=�BZA\\�s�;2�Zqbc�\�N�^ՃC�.�r�X��&\��ό��Q��@Eg�����DW���+!$1��P�O��9��ʟ���	����q7yi�u"���53Сz�����bs��U�:�sb,���˘\��W����!�{?5��c���Sc��y�:[>��4��Jg)�l��
�M�r���(�����&��b�@2�33�͠Q�Y���!��U����e/�\3@z[�5��4�+��MUnw/>��J�\IY�׃��z6E9<�F}ŭ���2K
��?
_��������#�lfE� #�k�^�7�&u�-�A�{5�{�ߞ�**��rI�$;=;�V�,��Z� F��/Pd@��<��6T����w��p� ���=���)�h�����'�3ٴNr�d��8=}�����Ue����?����k��t������G~�@�`;}a��){พ2ki.�R|[-,z�0�V���ex��/�2{��.D`�6��t�G�.��?ו����&$$�(2���M��l���O��2%<y~�,�s�I�i��;:d쫮C���[(�O9��KW����@�Ԛ�ݫy3nd\`��@�!V��>�XT~p�uá}sam���!*��F�� �B��2.���l��,��ȋ ��§[�7�~�YD���yj��Xn��Q��Z��ct
U׈��.�^S�g?/E����}%�	F��z������z�:���8�A7�Wg��2ݗ�E������d1z���T��(e4�#���\��a��쬧�<�~�Rٞ0e;6>�cO�8	����f ��:�y5X�R9��[ۜ?�%P�}�/�ҋ�	�Ve��]�t��!Xգ�[c�����k���!�th��c\m��	�EE�f��v��2G�R���5�1�π�vR
KJV�&2115K�T]Ϭ#I�������O��PRel1�&�On��N@c�ZcI�)���J�6��e���)��l��"�H�T�Q�V6�`ɼ&����A#��e6�!���<����Q�&;g��X��X�P*�+��˳"FOX�+��b�!L���Րd����(������p�G�.3�Uƌ�0T#f�/v�9�թ��0��|�����^+
���ud�]�,�)z�BOG���^��%y�=��'����i��u߅�*�:���1�i�ŝ�J�Tń����6 D���@�Y����&����+��(������� ����3�������L��DO�%+�½d�W�}R3;c�=2V�|��[���
�c�.�yf�B�BK-�X�А�s��s�+����MF��P����!NK�B������x�T�aӠ�Zbsݞ��:��e�%�;4�p_�v�0��ÍH�X�U���{�pa�jbi#_��	RԩybN����N�H�߼�y���"2��V���ui_�����k�X�]j8��w������F��~j{і����5��Ԅylze�S�{�P�P�9q��x�ۦ��Ɉ��ᶉ�ځhP����8\���j3g�K�c.G��h3�*W�a-W�&˦��/a-�Ȃqm~��CBZ��f�k�⦩E�5�A��10��h��&��!S��q|���t:5Lh�<8���P!�vxӻ��U]{�y�7����ЩyI��k+�&u��o�f݀��,���41�����;U����˴)9�q�1g���?��R��8a1C]����^?a�˶�� 6����WMDA؂�֟Ɲ�-�E"�W������������Ǿ�8�:��=���i�o���������|ʩ��'��,�vz�`s�(�J|lG)��џ�|u\�S��2����l������r���#.[�m9�<��%&(f���]�"#<R��o��X��1�ϥ8}�_'Mf�7��G�M�ƌ��j����*s�PR"3��	r��S��m���X����7��+���3SbV�	{ ��+
�fN��v���/�����/ΐ��Wl����SOP��_��|�)�ف���+t ��'m;�W����Ԕ'[Z���ο��h������)g�,Or�}}����~�]D?��+�fu�'���R������t���lን���< P��k"��i����jND�����$8oњ��ǐ��a��{r���r=�r�!��N���� ��Z��=�'�	��7À�x��vs&u,�Ѓ@��w����VʀS���N�)���V�h��d�C"�ĭ���m����y�7�@�N;��G����(�P�*Ćh�L��6�������;$����ʢ$�;�K�2g~�D�\�qUu�p|�*Q�]�5��8�	D����o�Yf?=gD_S�o�	΋ꮇؘ���O3&2Vi(��:+u$3��&�ځi������h���"vA'�}~,���sݏ�3�!��0����l���Eٌ����]&�9Xq�$f�]���h9`rM3�1��l6Ĉ� Pʔy����(PW[ n����u���m:6;f�q���7�0 ���B���F#�e_L#-����414.�sZ���0֙�`������VWd����kc��N�vӜ�x���
���z{Ðn�R�ya�qE%��r��q�}�,���L�j�"W<(�U��~�]�giդ4*�Wo<k�~��E+NР�g�>b�f,O������c� <�X���� į[�ѭ���1#~	ڞC��x&����{�M��	
&�d�|%�@'���^̞���"�!�|5 �	����V��y�z<�(kN�jj��p��>��`\ g�r��%�A ���y+nM�F���|.���{�I�L�-S�l�%z2a�d�f<��ǋ�<�QxY�	�%�'dn�K�-�P����֏j3�q�g�2ܿ��Y���1ط�Ƈ����#��ʻ���C:f�+ڶ�5+��C�H�ge��������}Vai���j�@ݤ�|Aw�q��K��Ҝ54&�ɣ�����)N5������{����4m�g��(`X�~r�H�H�\�����S��+P�4��ЉhM@��N�*&��o`��L�YB�����b���M5���"��׶�Ҝ��":�� u�'��[U`�_^��>_f�U���\�,V��������}Yu[
�g����a[?7��n������n�r#������F��ϣٮ[D-�O4�'j����9�^�E�O���:mwHeKB:�J�']#��e�	-yGK���I���yg�dm�9z�K'�x�����,<�t����1G�؆OE����2�:�Tj"99bDE�w������m�f��m˳���_m��1�1��Z���G<�@{kK�
.Ԩ�Eۼw�d�ctɾ��%pƃ�b�~Y�WTk��-c��
ED󰘆ou�2��]צ#*�QVK0����b-��*I1Ê	�r�+�i��1M�
9rU�hL8;�;٫�����c�^��ȴ��������a���(�}�FEiAE��h�3k�����faF���M7��Y����|�,B���)>�^�E�sU0�1_�	qrݴC�!�o��Z�2�%GRs]5/�X�]F�&>�����AX�M���g��P����[��:?3YLt���:vH{��R �C�b=%VQ��sa�^X�<U!��a�o�c������9��3��6w8v�"�Q(�\�B*�V6�\y:�ߗ�#M�o��4�>���ګ> �څf��� �����k��^����MW���p�N߸��n����A��Z#����8���ԨbFFn��mR�y�W�ǵGA� �}`���N�q�R*���L'5U,�ċW�L�ZiM��wծ#N�|���f��*�j8���ru���g�����ɚ��T>n�\��;u����q	��Ǆ[���_0FZm0��K���	���:EH�Y�G@�O����]=_���T���m�r2Z(zz�(E����>��ִ�o쨈�U�*���B ��[�lk��r4�-?��t��8�o��+'z�C_<�3�� ~@t����eveP��Ui؊#�;��B몀�^�-��Y7�:~<_G�E�*+�j4�G������s�~}r5�A� sq��z�������[��I�c�!�vhJ�����R�B�4��@G�c"�f.l�����jUbA��ݱM�����hz��ǧz�t�E��醧�N8p�!���ud��s4*�}"��b�Y<�6�S��`�����$C�(�JV�#�QD��e�TG=���W}P��tڼ�����&q���u��>�&��ڞ��dY+�|�)����&�D�_�4�L�Ԇ��9{��k��'D�	+ۼ��4����0�~��hd�u���g�{����xD�w���`j���0�(��~�޴y�Cˡ�ތ�#�w8B��!q�>X,ލ�Vz��������O�V�P���v����5�x�ٔo�rY ��&%d��X�qm/4#�PԤ[�����������K�~�V���a ��%��f��f�l�y���g��Σ��TR�gE�.�m��-�)���M�u�w��Ix�+�*��l�+�iSD>{=f�X�
/f���V����#���Ql�>���6��j0��5h��E�~��a�����z�W�����M�f{ݪ�JL�tqp+wK��]��觰�:m����2p�H1�q!s�3!9�����u�y�k�/��XZ,s_���|��Jʋ�k]5!�8�`�e�Ì����b:��~'��Nu����ʍ�ڻ�(D�
�8�x��܏�G����U��J�Fa	4j�i�`����1�L�f�P�Z�YOxĘ�B'�?���,��S�D2HR-�_���0�����a�F����jn;�r��~ʊ�Y?�Pފ��#�J�&����pe�� I8oo4MkRp�;�4��,��S���ͪ���l�����Ѭ\ ���Tc�H̦9+�R'շ7�����8���Ź��A����A�2(���F�\�;��!�4��ܯ�܋q�O�%VR�i&��!1D���~+��z�9���i���j9��_����V��0K�<�3[�9[����� L0���q�r(ڷ�m<t�φ5�=�!P��(gN�^*F����d�GN6ĺ演�Q����w˧�ޏ�j�Ӷ�Q���4�ph�L ��	��w��1����ݝ��"��.Y���$UL�R����O6߸@�=����X�˖F��@���R�!u��v�+� ��x2���(���g�͸ �qZ��P��8�	ru���-�#���~�#>��3�jC&2�@ӟGv�C��lV�w>����5UM,��+�4�M�`�h��R���4���..�I0f�?�,nT�ϖ�>4�[�<x?��}G�%U���0�D��0=馒����Y�4��t�lF������ ��k2R�Ԥ�^����GV�~���O�'�Ŗȁ{`������?=4�RzخAI����\ZCEj�ϔKϡ���_�sUX�$=�]�>;nfQoP���({��܀�l�H��՛�w���o�&��_�Aq�[�н�Iݟ��kxG����wi����F�B��KIh�o�S�Fo�����q�7xz[r�{k�˻N���@wN˂�+{q���Oui&��*ٸt#�LpŬ/���L�5���W��xبN;�W�n�'��*̗���֞�����1�*�ZnUt�h�ZӰ/ǳ
��/R� ������P$Ɋ���d�f��,K��Hj��Ll�rQp��:69������gi�c/̷�Z��K4*S�uוp	�땮qY�}kϛ���:���dD	l@g���#��E�fq��Tύq�s����KU'(���Q$��t�zws�"oh׉��F(V�MC��x��j����+Ȗ���5�j����?s����hu�,�0���=��\}=��d�
�c)>�&�����d�칤�]mҐxc^��V/tE��}t���aT�gn��~���kͪ��`����X����h��|��QGb�{9����E���cE�Z=�U�����Ø�C�C�e���K���k�0"6�d�}hʱ�}��5u��TǕ��G��\��A��K]��=��h�]�l�E�[_1+��Re�Z�ݢ�]ã�m=�]�,���
��]|l�coyiJl��	ǖ�1�VN+E����;�7$��٣#�&��`J�!bh�^���`�����IlW�0���W�3�ƺ/��q�b햢��ũ:<�MS�I��os���L����qFv��~���aDmlp:�Sۊ�pU�0���U���W�NC�d�t>I,�ě�����j��usi�O3a�1�j��gc�Z�Y�y�9c�U��mh�!�7 R�e��v��W*��<���滻J��\FrR���b/U�����*d]g��M�B(�K���L������s��'�(�A��&��=�����G��_ys���S��rW5�]+���e�J>��vI��.��MJ͒JM���F*R���[���f��+d,|Qee�B/��=kx�]���`Ѫ���9��uCX߅��k1���-y~�%k}�=�@�x�!p9�g��=��́���!��`�����'瓮�_�x^�o��@��'ұ;�u�D�oxS�rY�k�0%�g�^��>�h��=�#.U��_ay4�}��R��F?�J���}��rq�D3�BN�:���[��$���o�E�����&��d ���s�z.�7,"��������Ie�9��J2�fqLR��ņ�&�:�E��{���3ב�*���ĭJC/]��fd;��,J���\���
�5����{O�H�%>�O5���ҁA+�m�mB�8$�4�e�*}�j+�)����{��s����g�y���7��r=�z�S���pl�rϭy�z�#�׻F���[/�/f���R��m9[s-&�1��/R�%��l9�D���%
h��e۰#�u�kB��t�reM}[x5)q� '���sGӵo��R�n�|��"��)�{��;$Ӷq�m�c�Y_A���F������k��v���O�nxLg�m����"�3�*1�Z a:���I{�L��Y���kX�5���-�b	�	܃44�R�<R�׻�4؞�G_������#��͉�a�;̘���l4�ݩs$��kͮɾ�o\��� KR����v��3T8D�m꫏�Akc��TE�n�u�}�@Y?��}�� y��Z�4��c�)MG�ї:���=\�c��J��eV�� Q�	r�뢞��UʥOs��꿼���.Еo���z����t&���9/G!GJE���$�cfb�t㻗��b�(���Nɧ{�L�²��$ط2\{��	X���<�8��C��1 ����J Q�L7u�_�n�3 d���C���ݻ6�:��:���0����<�K�x9��7����w�jZTn��&�9踰a��0����ǋ�T1�����@|���8ːy�[M�Y����g:V8ݿ�f��F��[��r[�G���p��軨�y��˷����QP�ˆ���mu�3&Bf���o��d���0\A�΄V�@Ƨ�����Ӓ̋>Hg(h���Xg2�ix���}DO�4m�x%�̌H�����]-�?�Idր:NPTP�\����5�l��ѠC�YC�?:����~ޠ����u��y�y�8�$�;�+D�8����c�a�(I�h�c�;��r(Gcs@�ĵ]�+���%�`�'�>�#��4ٮ��G=��h�W��Ψ���~�~kW$	�q��x��.��� �m
Q;�V4}��,Ű�;��j�*�*��K�I�����������?�X<s��(�v����ʻ�sBA|���1��oY��}�'m۷2��f�V7�43��X�m������R��y�{�tbh>�CG/DvP�C�M#��O�at��dy�N<�ȋ� "}���L}�0�)f�� ),��0:��6C�Ҵ�N�!i����Q���d-�ؒ��x&~..]R-��/��e.����b�[�E&+�{;۾s?	I7���#P�ߡp��'�{��;�~,`x������6&Vpg�F�����\Ы|f��3W��؀��n�il��Aư��b� �j���f��k��92F��.v���ya�#I�g��m��_�*�����P�ߕ��a�^<�89"�A~*��J_��bf�Qҧ)[�i�V�+3*�z��*O���2�r��y��m�i�<,��%�྿7�Po�`�1(��O-S/�X��v{�M�]sC�zw5���Yt+7*Hb�㾤2�À�O~ZЃ����m�>%/�ZyZTw)k������K������j6��~�~>��b�@'��35��hGAB���ß�r�k� ����N�h_D�~m�g�"�$\��\�/�A�I=���\Da+���������Z�W��%�ʕ^:�I9����ȷ3eE��6�lRҹH�@16�L$�P��Gn�?�W���kh2A�^�g��$x^7!�&�������� B�LjA<��"R{^y�<��<N�U2�z�Ê����ɚ[���V�~:+��}|w�1���_ݻlߜ�XY�B�#A�,�1���'?�I4�S֝��3#���}�ヶ��k��ֹ�E! �T��?Th�'�/b�]�����R�*Vx��T��uXB0o~ ¦q�"5M�ɫ��os������%�(�Y����FU�����/��y�r��DѢ�J~ �t�{=�^��$�	��#�_�� ��E�ơ7����ҽ��#�EFn�ɸ	z:RU�oxx��X�?�06�oZ,4p��XY��~���	
�Ӈy9�%HkĄϑk�O���79� ������eK	��!Reo��a�'[l�]"��%��$�(�)A:�%����9qRl�{l^,��<r�-_v%�R3�J��2�╌'U�Oבb[�G���8�
���7+�fء68�ɅĠ#)�B��2L�6e�R��}�>Q��"�V��g1G�3I0f߶�qݱ�Cς�c�7VOS���ŬM����cy��Y����!B���ɀ�1�1�����v�����ro�Tۧ�����\�4�Ut���֣�g?��?�����\#�>�9� {���K?����s�A�����`�r��u��� h8U���)n�Y�N����R�]h�*��*�L�+�m}5���+�_��%��*u���E��9F���y��a����L.z�Yu|2fͮ�A��&D4�Z#�)�<"��䌦����'�&�A��xX����oӑ���I�FB���������5��|��0zw	t��7�N�m�{�仐Z0Z���h_����;��w��`�G��T8�O��������rZ����c"i!X�����Du~�he|�T��d�E�3\������eۏ�K⫻i�g_���ޅ|�c���mqY���Ѵ�>�*8�qX�ȠZ�f�|*Ԁ����O1��Э��O&��qᅬ!�^f8 �b���]����00�xՈz&S�HmXkU��~���w0>%qP�U8Q�.��[�*<ބN�v�Y0���xdg�����4��#L�kh��.�4����#^=Q��6�
9 ��o��L,�ߙ	k[ͳ�Z���l�CIK��]��=�zN�V3L��<# �6����/}!�(�QN�R�Gj�4ǟ��n@��w2��
�,cջM� �cRxB�ݫ�,R#)��W�m�����}bu��s��(V���?	r̴%�=�1�n�&6K�_��ˆ�=�6��Q� ��0�����%XĒ`0!W�b����[��G�Ə��=�5=&��
���pL��}��a/���!�b���H���/(�('�,d<��hϏ8�0�b�2�ڶ&dݧޛ�s@T�H+�$,t��2K��G�X�^EMcFv��d&2ۂ�eYM�8ZI7=In�D���7,�'\KXŐ��qa�6�^���V���.s�Z���t˜S}�����@��#�b ߖ���it?�ca�cp�_�D��"Q0�Ӏ�*�DE˴���qA g��@��a��Z��Jd`�d�X
����bP�W�4�����2�!H������c(��hS��+Z3q�U����� w@��n����\OY�LADٔ[��fQ �L�Q���OU�2->�ӅvvW����4�T�X�Ey�۵�F�  �Z�v��V^���Y{����Wsº�����
��xd~CP����_��o��%�y�J��E���s��t�Iv�'z͍���f7����,A,��/���Dd(�AA��Z߂~�<&�D�%5��<��|&a�����`��]۠�2޲�y�t~j<�9~��G�?��!�9�Aa����@(�L	�~���g��:7L�/�����u
<
R���
$x3���y��Vt22���KVy}j���-[��p�p�1�Ⱥ�{X��֮;2��<�kj�nU��=�=ϩ]�O�m`�f[�n�]#��Eg��������wXc*�����!������#E���	���z�B�&�C`-!gT<R1 ��5��>���;�$�9x�+^a�������L�=�8�ą�llv���\�M��#�o��j]�!2�r��R�����G�M��N�`3#��f��M���|��ށ怍MYo}�rJ(�E� �α��T3L8��K_�R�`�6�5���aY�z���\*[<o5ptʔ�n8,�V<�%���_�<��4��7�:�vf����>�-�3r� �+{��m��͙�O���3[�G�-�G��jj���P���d{hƼ�E�r�adF8�9�}���۷��-74y_���}�Z�t{_Z�u�Mo�2	��]`�Lf���X��h�Vv�5��cc��z��|�� Z���B�O1AM��!�������P��[�/n��-�#��=�	N�t��!�ʱXt�1���!!�b�ϳ��*��k-Oc�m@$��!$��eW �to���ޏv��ɺs��/��pZoI�4�lr|4}w�W����񬍏��/����DBXR��{3�\����,��莴Ӈ�w�Y}")��	� ���Ζ'��{��~�j�P'��C��/��,Yk|���kr���it$��);�3=�り��[�¿��7��u:N��{���`/������$O��g�����=��cNGcA���:�l��5���Kq��|��ڱ���Vڐ�)�zc��}��!��s
�}AG��-��`�}�L���y>b��#.�����0"�0B.������9��KC��]��{P��W�rn?�!��7�e�gX'S�j�6h͵����*�{+c�����~���dm*��]����G��~��Ie̜Y���=z\���G��O"�/��iC1�\��U�����{p�~Z�>zZ�s戮�?fc�۝�99Ѱ�;��W������^ ���[y�,S�L�{���66���$ͫ��t/ɣL
��(�t\#��N^��K�FQ��=���	.���l'	��K;(6����l�F�;�jW�ȚfRV�&�~����g0�>�\;㌳|--_���~�/�Z��[=�����z�pݢ���Kie������<+=��/�'�x��=i�֘�x��~���i�G���k��u{�K/�3�8�'��LJ0^%6q�#�8>�h��y��z �\&kQ��9F���0�s�(x/�|��f�tfs�����+�'E�8�<		љD�0d��#�,�ى���Dƙ���	2}�����"h.�c]����'�*g�9����SXO\O�qRP�!�JO��ݺ�lw$���k֬����:A�48ɡL�v�u_K�`�v��Q+�j�Z�CIy�%,�q�fV�U�
��u�s��DY!���R�>b~���M�/��j�aOm|����$�������Z��{vϝ��ӛ��W��5�`�,�+���6=����;�\�4�^�[�'ּ"�g�y��Y��v��e�n�d�c�����Aa��Z���i�sɲ۽{�v<7f�z�o��N;ͅ<�:mv�8)��đ�O�=c��G}����SP��^h��bzc��a(��"E6&�D�+:^��oi^��
�J(K��<���{��X4�!�ň��D4}�<���P�U����,&������,�邔�o��	�$^5���=��g���V�В�[�K�,K�g��O�ã�+	҉�,ڪ������d�����7����[*��wK�Sʼ�bm{�(��L#sK�Z#����#���_�`4�~ޒ����lI�'á���NL5l|l�x����/��b�y�a�=>əg���9`�����F=��Sltt��4��v;��c�ϱIP?bc��aU|a�	�vW���^���y�l�&y�{��]�轉r �o��o�k�q%��_~���D)�S�_����z�������S �K�ySB�	�L�
D^�ޏ�:#�^�}��)&��K�Y��)DhH�9����~
$G��5�ZP����5�,}��r����j(�e�A���-]���E�7�9� `hi��p�+4iY�4���\�w��6>9���@s�.���|{����o[���M�Y�E�N�sK'.�c�ȹ^}�7/c��/��7��G{ ]�|�z{����y1��Fmْ��s�6Wp?���SN����8RJ���;��x��"��^��zp	E��&�k����㫛6=n'��Q�  Iԝ?6e��
o��+��	�V� ��!������+^��g�@�cA��Dt��3ͭd��1��s��`},IA�����;���nd53g��&�R�c<� :�,���{#<����^S���XF� ��^��cnH���J�f�zbI���z����FV§�,ٵI�Z�ɾ2'Tp�����xF�M{?aɲ�~��oM�=̓�H��MP4��BL��t�������[�P\�Z����˿��EO)O��}��=��ԭ�uĞ���C���ڱǮ��kץgٲ�RSHG��/������?��O�|9�c�Gy��]s�=����L{K�]�¿Y��I��o��>�����b=�١���1�oƴq�&���O�p�|�^m^�
����GP\w�u�pp�	��A��c�wdg7�e���)��i�,Y�9FPJ����`+�+�N�U�Gʇ��U%�c^�6wL ����v�9��>�����=|c��{��v�c>�l���";e�J���,�Z���w��$�̂�N.�'y%����+��!��'��K���=�c�-s��R�J�����h�t\XK�����+�}��;�<��_�U���߁��xd�>�{�;����Xc�'Ň	�Ï�pX:��k}�<���#�<˕����ֻ��kiM4m��U��bMD�g�߳k�E/�{�RK��N�/��/fN�&βɫU��M��L<15Tw#�*���~�!*7��]�C?��ُ������U�)������o~�uW6�V|x	��M�yC�K(F�����G e�g�}U��0�!�!(F8�KxpN>ˉs����j� ��x&h15��"ry-}R|�+X�E]P��-���پ!�)}���\��,K�VYe`iV��<@\*W���=͖F��e{���k���L^t0��̋�5�I���l`pvڵM��Gg<%2�.��b�l��̅�#HX��G�I[X�R�j�����x.�:�H�7�CN�����d-M�-}O�^�ٞeH�B�]�¿ԍ��*����X�: ����g7�p'����崨�_ZN�C�)�Sw�Kբ��Ұ�y�L=�gV��63������{��`�j�� ��m���C�6�K6Y���ñ��?��O��uϐU-Z]�dp�^�7��ω�zXj��y�!�����*՟s�z,�qy��g	l��ܛ�N�.���k�\�"8�S2��jȒ�a�wZ}����R^A���t:o١���cɫ~����d�[�:hO<��Tyi�HR,��Z�]���\�YO$܋�U��F�9w{�x���퓶eێ,�ײd��h�;7Hs)��%�!N<�g�<���c����ەQ���	JY���+�{/�rqT�Ȓe��z��}�6[�r�mٱ����X��?MvO�<�Mأ�<��Q�O�Y}hZ��41#Vo���I�Q�vȊ[�{ܶl��欳�*�Rzy*�Y,,=6���h�(h�U��%�����C�YA�K/����R�S~A�?C�y��emɲV�%����0�����<G)��ȸ��T4N�:k
1���m�g!l����E0Od�Ha�}����׾6S@�v{S���ط��9$3U���-��cTbw����{�/�R��ozf��6����$,���t/O��q��$�К�q����K�+��4�7���j'�u*���i%H�^�mS3�k_��~����!��!�0(š����S	���^����d��x\�5�j������������gmbr�ο�,[vH2PmԞ���m����M�:)�4�?����W�>�,b��|�N8~��%����`��w�m~v�'bd1�J	����$�e�~�!�iXlR�{UeѼ���׼�5E/-"ea�qם�����w�/���b���nk�^�\�1cFA�Nn~dIȃY�A�J��>:���]*��f�!Ų!�.�Z�*8'�qxZS|E �q~��
���.���u��攋��4#�gF�TBV�ٰFS �j*F�ߔ���>�{d���`�Y�9��\��_~V�� u�/��H��V 1�+��d�`(�����v�/���7���������=H&�u�]^:f�-v���m�s������� O�֬]jûFl鲕����;�زQ{�)'y�J�����{�"ٞ�w�V�|`
���/�������ڹ��V�X�A��?�v�x��ȳ��5�竖���O{�����t����n!)���f�����G�f�����ۋE<:8vHX��M�9<2���Z�I��Z����I�߼�< ,��2�ʊ%H1��t}X���Y7���i���~,�s�<M���m
�CP�9�
�P6 K���R!���� �(2V�q��hgҔ؞`��d�QnA0L��GP6��J���������B��[@!R:3ɽr� �m\ż�H���Y��{��
 ���y��fB��Տ��Gp�q��e�t�HoH�߿�6=�ɦ&F��Y5�Om�dK�bkWeW\v^:~m�%{��-�u�D��c��V���0�)�΃�~�;��;���68�o�#%;��b��m�=�̟&�1�S;����/��ի�M07�ζ�~���{��%�\�A ��x�^np�7���H��3�����CPV0�1�X*���rW�f;�uZ���`I#�# �sqNA>���'��Pք���
^T^�M�`
�F�c|�-�׃����HB�\^zd�]�Cu��$�"b4��HT5U��,����e��T:�j�2ku�Y�	b��
���\��_��@��h͕ 17����+#����}
멼6�!�Q̳�#5d�w��;~�*k��ǜh��%v����Ș=��öb�!�b�Jמ�^t�u�zOv���w�{]R��ҵ``�|X��?���ߦ�\���j؏�3_�o|��m�в���^}�v�k^�Y�XC�w+gk�0, ������X�:��l@(�#��f0-66�~i�}pt�hl`6�\|��W�R�� ���H��Њx�b%|q.� C���C�V�`����Q�]���cbd��^QQ1B���׃�y{H1Q�2��}��z�R�S
��5������x��&-�
�ߖ��
�>]h7m�׳�Sn��f��?�{�
Q��r� �4�����9�������x�}~��󁒅�)
hdW)��*����y���=j+Vn������7$I']���G���F���/����v�=^�F��}�.~��*���MF�ʕ�=SʉA�����ܶ���.��O~I�*��<0�ԅ���pM�5��޻��	"�N�j2�l(�?�я��� Y���{.��U�����V7�F��o}�L��_�Ln�R0@��ɳֹ�{�O��;b���� ,tq��W�0G(`�5BT� %֮����`ۇ�r�b&�cP\��(^��W�ҹ�%%a�V?�60���<R�5@���D����Kmf0�C@y=�v\K���;�tx)�������f}�|�H�-r �=���Tn�09<(]�9�F~^$L);/�9^��o;���]l�Y�k�C������u#6�d��عծ��Z��G7gl�ь-V��3�X�¿�h:elddgf���&�s��o?��v{��G�\
�أ�v�N�e$�fvo��6{���{,�F�SD�����?�C��h������KH0x������_��p�YXjxp,�P�U��SO=5#t����'�E#�폘?CBRyZ��Ǆ)�}h�cP] �t>����G���,�I�F�JHIgA������>Q,JTV��;:��l�{�<���e ;���ؙ?�Y��Z���]�ᡒ��l��{��b|y�f?.|N�X�>�6bM$����I�p>���"���gV�����x��<w��7��	���o�=���u��?~��vc�ݲ�5��!�n����o۾��ȕ(��G���4�����7�X�¿U�N�ECg���W+W������2͎����h��@ڠ�b�U�z@ic0�X]*��q��;������)AE`"(������2 8�`a������M&�Q���+P+H�y��3��$P	�ך`�F0 x���q|��W0v�S+�22��Jb�7V������J̍TO�Ž3��4�P�PD=�{�k��_�F���t�l<��P*,��&� �C� g��A��R#h9{�����,���m�pD~�1��1xy��{���+	�������A����	ni�3��k_��?+�Eo՘nb��ݶcǮ�HH߅g�{x��T�̳Ƣ��GZ�Su���H��#ɵ���0=�:����i4������d�Q.��=���ܥF��D��44�����C��O��Ii0�0��#���M��N�'V��KL@��|�`�`�tB[X�k�軕���=�ǜ	A&*��?����x\k�vQ/���:��(�I�3ޟ(��B&+�*�C,��;dH �r�:����J9w
�%�Z>
�b����l���P�]�>?��`l���<���i6
%��(XS�\�6��9y/���l�|9+�9W2W��Ox6q9�}��H�s�4ʘ+Z"��K1���z`�(N
7�����=�����q��栘�A���G����"T��0XC��Qʆ�c+}e9S=�S��J��l�����d�Q|�+��E���z��ڸ����"b��lŅ"�7�\��K�D���E����BK�Pcq2Q�|sV�s:�>�wxE
^
�%h�������l��#��m(kz	d+�h���E�b09���e�k>�<�%)��ȥ㣱 ����ܷ�T�,�u�NA���	���me4�y_��tEPˍ�z1z���3V#.�>/�@7�̸�*<s*�:-�ޚv]{;b�yUڧĀ����@�����1��`��=�{�̣R����{��E/�{|go=���:Ӛ��6��?�y���aU��� �������>p�c[m4-�H-�9��mp�Z��d��ǾЖ�(��k�z�k#d�=�Ȣ�A���	�U�G-9x�U�E�by���Cשu��v�ɳ�x�X-�	%Pe���B��!ڦbU�������*��"�\D�z2��s9�`�}�&���aȋ�E�m�Iq�kjgHO�=���sYM����ڰg)�c�՜^uS�o��ٵ�bn�*Y���y���g3��s���]3g�*F�gV���_��{4g��sE�\Q��C@������r6�,G~�{�.J^l�.�@�p�v��mp>��N(`(��B`b�r���c"�Y�);ݫ��7�����b��u������0�O|�^�G���m.���:�_��`4����r�3zF������3|�*��8A8�Y�4AN�֕
�EA$�&!��w�N~9,�}ҋ�O<+hܫ��")
	J�U�b�n�2%1��IyZ���htXx����{�}�D͌*]��_aD�b��wQ?�)�U`����^������(�p�	�qi�,��YQ��ͭ@��T6%���*�Å`.�bC��Ҩ'X����õ��׮T�,��χ�/Z�P���8��hY*Q}%��g(�B0	�/���S���΋*M�0�CL��9kPP�2�uY������Py�����0�C�`�x�:��T`�)I{gEC��P�Vre�r$�cs)<�K���>JvblԿ��#��ƾ�[�x��5��PW�\�}�'�۾랻3je���3��"�.���yD�;����l��!o�y���G/�f�8��6�bD���m�շSC�J�Q�`�K	6Zp��TS�H6�m����h������X��}uǠ����Z����9����{#���|
�	�ݟ�{�C�A@$zqR"�^),	�s�~�o5fU�k@h��#HBВbGz�N��ۇ���w_	y1�$�4���nCumtm�l��~V�.�1R#���l�[]���%̹�Q���L+y�*q+�F2���^�c����X�¿���L?�g�5�.�Y��̔�� WPM�{��e9�/�_~Yb����f=��n�%��X�,/p�a�~-��u���L��r�|׎�UU�.s��9O�%Bϟ �,8��g�u�c�	�^��ye5*CT8�����$o	+��V6��:�X&b�ț��8ߍU�^��"�7]�O�S�A��P�N���X�VJ���,"�:���n�R�i/��k428�k5g�Y�	���3�� �C����V��a|1�C���ǿ�س��L	�1��o�/{�m[3=���L��5���Fĕf�`�j�ֺ,5Yڰlq�%P}��zo�XbX�.��r�^
v�M�0�F�L���k�cD�������� Ās'�R����}|��T�-*{�C�,oi#{GX3��n��_�ñ�,)�5)%� Vf0�ٯ��
Q��x��̫n�W�)�:8/�'�*,~h��>�=�r�6���a���O#�Ә��i�hOkϪ+\�w]�n�gX��sؓs�\ا��nf��T(ɐM�H�|�g`��|�X��h�S��j�K�F�/��P.qt�5�����V[xE����,#]�R� ��\ӔM��H@ĎO�4v��=]C'��=Yt�0�|C|�j�p����eD;��g��֊���1�1� n�Ź8V5���9��5[��,~,v?�FLYE ��T�?*w5v���X�3i���"���nR�P �:c�X������in����U��e�4��_�1�O�gQ.�Oĩ��L��֥�2
}]���u龳}���~n�Cy>�d���6�!��"_ �����@E�^���}(�P�fV�X����f�)�x�q'dV�Ĥ�G�mٚg�V����%�!+�����Z�F
c''��-vX�q�j�+`k�hQw~N���3a�^�NX�ҧ�PbP�G���GB!2g����PB�y��+K�90����a%_͵ܶ�έ��3W醨�Y#@�
��<�	U�Gx2��O��ד>��se�F>�=q�W\qEf�4��`�S������z) )�+�9w�~�扌d 73A��׭�ViZޅ�����K���~R�=8_�z���'��1���^�-҃Y'�p�y��g��@V�i��K�����
`��V�'C�4��7N5	��1�:'/y�K���3���)�:�&��d�y���'K^�	.&.��O>�j��~{��fcSD
!�[����`Y1�Ŭͤ���)dU����GL#Y��F���QK�G&	#*3)C	����!O#&��߅V 
�I�<"�F�Ne�
��^P"�G�\
E]��1>7�^BZ��V�̺&���:G������JT��!��2�״6���:�����9���z
ȫ%�Kq�n�[�Qݓ�Kk�כ-���u�s��j�+�"3$�5�2���G��^��N8�=ϥK�����n_?��Ńv������lyY�9�t>p3|���U�gVOQOG����|�7\��H�HL��f��V��&k��u�i��op��L:�~��~�7��_���\i\{���]Dlu&�Lc�4{�N7d�kX��%������Ɋ��YC����Z�Ŏ����N��ڬ�.��(����u-<�d������,AS���z��u%���6��/(2zCR���o��0^BK]���u�μ�V�iD���T�UDl����Dh'Z�b��we�f���lC��O����~ �uZ��W��(���!&���d`R���3�p�oȕv53��9�l����䦧�_�G7 �U"�P	t_Ǣ�y	�YI!�Ed�j|/��"��񤝫e\�qۼ#�j�e98X�ɴAN9�$[�f�O�����ª�P��K�����|�7ۿ��������^�Sة�	Pa�sI�P	C_MA�� ���1K! ^��C�G�j)���'�
�ٯ�r�3v��,x���_��(���Θ��/
�s�]�ys�L��zI ꘨e`Ȼ�=d#D�s�L*Qu�����y]�	����n/?�ZPRН���Q�1`�ƺ֩F����Y�KAc=��&
\x5Z����4��a��⾋Ɣ<���Ø@���կ����J¨lN��(�8͂$���ڵӖ,�����>�[�/|�Kɀ�ϖ-Yj��#��q_Ǣ������˽�����^��+��9�H���n���Y�W�\�=8O?�,��<X)Z+^�	D)<��#>���_����|�#^��f,���� ?�5��׆CyQ%/C�v(�'�9��~�(9~t/j΢���5����lV,,e��������Q�Œ��$ "�����qi.��z�h�Ȑ0��=�/Z�<�JR�1�'��R*�������R��bs�H�t��Z�E%�EZ�s��'[U+E�YJ^�+���q�6"�罠���@m�7%�̟����c�~�^ӱm<\0��z��ב��нy	���0������R���7�>	~��~��6nz�n�����;}n���=�<[��P'�,Y:h�~���_����^��A��v[�¿Ճ�59Q�`��]#v�1G����d}�U�?�arٶ�q��Yv
��/�ݞ|�q;�e�Y��RW_|�G5jg!bI���p!I����ۇ?�a{����3ZGmj�|�6��(l�}"@X�����k\�h�	o]�g��9Z�q=>��X�jT@�8�\	&Q��[B^TG0N~7z�Xx��6*�X/E����xu�*1���u�־p`�S�]T�A�-���y=Blj���C�3&�˜0W�a���=�X�ū 2ǣ�E!U��FC�q�Z�_/��@�+��(
���e�����'wq-Y���;�1��3'W"(��<m۶=�s�C�����h��=�y�k�A%��g��w���2I {n�3v˭?���m鐕�%{��_�5�����^w���V��UW������vNI��Ƣ����dc��\ȍ��N��m|�Qk�ǒ��O�t�UrL��o�޴�׶l��w��}�ݑ D�M(�#��F�W4<�dY�
|F7�׈L�N�!��M��T�b�Y���М�sa��@8F��x��
�,S�	�X$���*!#Ꟛ���D�I�="^�Z�RFX��	<:���l7�' K[ޒ���.��_�3w�F���������q��3��U0a���jq]��՝{���7�!�-4�5�>��Ϻ��� �8���q��<��Ig������ܙ�+�?�
�zQE�������o�o�q���\��1��?�>�[�y=��Rԭ�1{v�S�s�6[���zkmbr��Z��}�����ˮx��AA�u�v��?rJ�/�K�3&��Y�kIz��^nL$��u߽ގ>v��o8̞����L�?ɽ��)�oO�J��Э?�Ņ��ظ��8{j㦢 ����)�.���B�_����n�tz	8Q��^GFE�5�G�g)XJ��\��,>5���*����BB%$T�����e&�@4Eᘂn�#��`�ApR�k��vX��/4癝3ǡ����i�iw&�u+w���Y�\�փ:o���v*�^�J=(ʔ�����&R�������|�yWp;��el(�4>9QԧaD�c�F��@�ր��+Z���״�bn���]�J��v:xql�O!�F�<CFRr����oذ�~�#u���o*�;��Uo}�-Zb_��W=��o
k�b�z�+���+�mz�qk��؉돰'7>��~��F&_���-�����V;�S�_���Jo��hvx��@�������;��;�V�\�&��I_���u�G���6�`�)X�� [��1�,(K���kXO?���@*��𖷼�q>�,����?m?���E@/�ᴐz�N�Yt�8{W���B� ��,�����o˞��>�@R���^�Ғ��+!
S�uH�I���|�>�];-���k�gAO,�p�^Z�zL�L�Z�+��|�[���gd�Ǻ2���	B�������&6̹+�r�5��	2�ٹƤf*lV.5�&�������A��KVt	k_�����s�X�b)
����?���Z+���~��N㦮����<�����{ϝ��C�@J@�S@E�����T� ƭ�2h��� qd�	':DM< ��g6�A��+Ib��v�����R�d�?��S��-�m�&3�Y�T�R���L��h7�@X
Fbc��	�b�}�;�q� |�w�w��?�)��Ul ыJ7pd��������H�0J���	�$�)��<�J����ıD#J���P��I��@4��D.��1"�U�
���+���������;Q���>fbGVH�̙�ye�:� �ǅ�G9K�k��(
�v>g����g�W+X'*9-�W���fce־_���ݳ�{+�L�]O��:��ÿć~x��n��!��e�ā~YGxyt��|k�����m���y�!i�ҟ���N��O�s��=���o��VK�x]�\Ǣ��L_���0D��rˊ��Ov�����I�*-��!��X�C8��t�y�{�:��ƥ�'-ߨ�N]{�L��@Y�)��ׁ���
03x��4���V=�$P�(�)I	+}w��kr���B�\��b�;RW�rHiʒ�	Uz��+��>���6��ˡ5֔<��{���k� �
d���?� /�Y�����%����,�)gP� a�
���Q.�z9Nީ�J�=�L[6� �`���c��BI,��3�bє�u�O>n�F,@�%�� �D���-PE��O�S��4��i}Y����<:�ÿ������OL+s�)�ۈ����i�>����l��z�ȏ9f��t#�+K"�L���db}9������H�Q�H���l �"�;�3N����Z�!��|���ǚ�lv�HmhY�F��1�����Y��7R�$@�����R�n�SѱN��G^�8�ԘG!J�1����������6S�������P�q�ְU���yMA^�Q�C8��"��d2�R�z�/(���oֺ�ː�I�����?��X�)L)��-TF�c���$���O�q���-�׫^~�S�K��p��ۿ�A�w���M��w�y������>�o�!���[Cs��_s!�m՛S6���Z��rr �ג���2���Ĩ�5�!f��9�E/�ͺ�wgg3`~�a�j�a�;�OѶZ�VV����Ln��'m�ݾ!�p�$&M�*�t~YbJ�<� �"ZR���lC�����`���q 1��6	l,D-N����q�����=���c�^��V]A��y��"�^����%mJ1pH���+Ȅ��f������^�g.�_�M=7��
ݕ��uQ2���Aq��0ψ��=A2~e�j]�X��o8Ya{�F#�k����xĠ�����i�=͵�Ѿ�Rkv�L���mHc��{�s���W�ʧ���8X~�m���<;�XO��������X�3C�������,����lt��ɦ�|��>gcim�Tdh�
�&E2�\�¿٣����l���^y�����s^�lOۮ��l�����F�(��Z�R[����a[w�R��#I�[�8�2�#�KO,�E1(
�ن,���`U�W�_�;���}T���X���r��bPL�t�$KV�
���A��C�Kx�*����v�������n�M*�D�LP������υ�h��f=��1��
��2�A�1j )���`p>QL���QS�L�Ab�b���s����]��cnj��r�v�ry�z��0�-�=�N�n1�00�{���!}�!;�%��3���۞�F�φ��:��4�v�I�أ�lLϻ�pF_2F�3��w�O�&����;��9�i��g.8��$�WZ�@5�W#���:�t�?�g�Ɇsp)�v��.*0m&���l0�?��?م^XP�b���G{���ͯ`�\��%p�0�YE���>��f�9����H��s(���C�0F֢��V\��͓!�\�AyX/�>�5<��"��h���6?���$%X��P�e�� �,ƙ���A����H!w
"�Oтǻ�F��Z;����C���ľ�,��̚��o��33��o�s��&�^�9��3��潔@l���-oՍ��z�a)~�'��7���>��[�;e0�&Ӽ�\u��ܽ+}~�m����J�犲�f�d�Ye�^v�{�z�<{�F�����/�Z����'�BIf�;��~�n��&��5�Nx��:f�/͝���'7�3<n�rՎ8�(;��uv�y'���MǺb�p��^z�M7��"�gS1�K��B8W���Eb)0���lB9&����|�7C��K��{D����uQ�-o"R�Ua�XH1��x��l�wO O-��cEHE�L	��6��Y�M���3R��m	r��P�;��g�a�8����D&�����W1�"~��dp>�����`�2�*�9���i���b^�_s=)�Z����z^ܭ4͢oN���\���zT��*ʹ���
쿈�NRӿ�����\�h�����/
�ꫯ����ﴖ�<;��+��,	�I[��4۹}�y�i72��ɲ">s\20/����~�	�������n�G~�ȍ�t�N���*�¿�G�Y0Z��ot,���K�y�?�X{��׻u����/�ڵ�rNu�l�L�S����X�r�� ���o���_��c�4��;X߸���o��"�3\�cb�	A+,D0bY��,�IٿwW����/���<#a؂��6�%Z$�*�~�И����?
��Y�<�'��7T3ch�ƫ��x��3mB�<X���_u��.R�,e�
�g�x�j��8֥�-1+���3��^�?�x�.�����Ox�bŚFsabE���B��B�%��J���L�dk[sR}�ݾG�K��BŖF+�q�Y){���m���Sݽ�^^����~eE�&`�}�_�ߏS�eyƬk%H*7C�c�Ĺ�/�ܾ��>�ev�y/�����)o��x����������lȊ�ױ�/�>�wı��Ѧ��g>�Y����� �v�����8*���6:Fᬺm߾���o�օ��ZL�����x���������.� ѧ>�)_���]��ψPL��Ŧ������ fHH��8� A�(PX��s��糲U�AHΏb�R���
���:�%���M���D�,T�AX�|��2�D%�
�1)�z��_��_�k/%ſ*PƘ�k-v��Ǫu�kS��
�	$�.a�3D)�9X�Ϫ�C�T�����JaP���_��`!�i��>A�F�!���"��`��H��9�%T�NtL�@5��`�:�t�&.������d��Y�ֱ��ã��̳ٺ�r���2�;STޑ�zŹx�=O����\��x�rX �7q�o��^%��K.��Q�s�)g�`�LN��̵>�����{F��j�k��V��_Gg@�QY����W�CP_p�Ey�⩂~���?�1woQ�E4K9Y0X����Q�෾�-�.��B/�@�@��
D�E��3,y0,BY�
؉��*E	E�D�Q�/����|��F��.=��r�=�C�"����@
�r��'b�,4��7j̑� L@����ΪT�EtI��Z�ipN�s�)���2�J��9�[��*!+[qU�d�c+P��c��cL`�!E�ʶܻ����c���x/�"&҈�(�]p~��'ltx�=���6�kGz�n�[��R�"@#W�<�,�Q돷#�8�cqO'��^zzs�-͗,�93�=�,�'��X����Po��@�-�l1��s�v�w��x��_�m���a�g񙆓���k�X��sN��?�Yͥ��q��/u���d��M�\饎�e�Ъm|j�mݶݾ���x���k4�%0>�Sݙ�����
�J(�E#�x��21�*( b��JP0*-�6�'˓E�LD%)H(]TQ����'�������#��Y"A�� )$��n���V(�eM�_�X�!���w�k�Ϝ��{|���3a�#`e�G�q���C�Q"�N����wz%��x��ށ��4Шp����5�Dzyg�\u}�A�ɱQ+7�WI�F_��+�Y�MU�-�D���X�]J
#c�4�mE��h�s)�/+�s~��l��r�AG�^�L���y��
2�JwH���o�F�G���xR����p���y*s��N�j#���x����e��RT�^�+YU$`d�{˃+�mg�wʭd�!�x��;�g�UC�e�C�^u�U�(O;�4�H���T���&�5r���| )��X�vK�ɢs#���d��'���|*=��Q�?�ѹ7�AX��? �]V��V�zY��k�J�Z�~��`���)� L^������)oa��TyS��UDN�[q<[�?XW*/�h�9��b�sC(���'��@&�kdl���wHA�
*l���E���~4�C�.���%i�٤��[�}W�fΓ���̠R��M���ʜ���{ �v����6��=���J@g>�|�W�*&�{docpѷ� �bzzf�ڱ?y��2�3Y�6=�%�S�!����݋�S{h�sT���g.̸R�t`Z��m�ˈuWD�t�%�_�k�� ���`���`�F<�k`�I������E���'?�Iߔ�A�p��?~-W,�����W�v&�)���,PY���c��|4�N� ת�c���`�^\R�����p�E�YpLE�8�0Q#m�K s�Yo�f��|.�iމw���L#�de%�u��iK��ol�+v�0�N\~=o�yQ�D�7oRק����T�X��x����p�u�0o��$�T�GU,X�s�%�e��X7F��l ��{s[�)7�j�	�d�I�yyh��@溪bB�AmdD�����y}��_�}N�7���������̟�nȐf��J_�&��V�Oϴ�ɣ��~�ûlp(y����ʔ 6��F�$���&K���6Z�"�~�E���f��d��m�z���K�1���R&,����� e! (���O���-n�IH�d��h�h}Ja��#��%oɲT0W�Q�'z�+�:f�"�x�AB���E� �K����0R�N�
��F0�@�R�Q)1
Aל�ZKi)�b&���<������H�a0�7��%�5=	 ֔�y�����l#�1⻕�a�r���I!���g#�-r���X\�ۂ�Ӝ�f�Y�i�%%�%~a�;%t2p}U��t~�Ԫ��!*�8�W^��ɑ<!ŋX׼Ϗg�潒�HX@`��dՍ��'m`{��J�V�Z���I(Zg2L���Қ�� ��}5�x���du��Cm�ܵ,{i��H��Rő4��0�O����[9_p�^��w�>������M�{d�S�c�,�����˳keMŠ��T HG�B��x��rs�Yd[%�D�dh�r܇(�x*׀`'\�d�q�QF��D��7�hΫz4�.bYDG*cy��[FgPS��C}�f�u3�ۿ��΍����s����<+�*q� ����ׯ/�S�]�j��bs
&� �G��<)��R"XΚq6K~OJ��[�E\ks�,b,"Χ��2�ߨ߇ ���N�C�VL��<MQm�3�۩�1���<��|��6F��~��Y�H}���+�$x�PQ��<��QfK���0�־A��\��G^�d��3{�g���y������_,�i*��^|��2�a����^_0L',"�}ڵ�r������z,��c�,LYw�?`���>���x�*� �BP����[��#�&��,J���Hu�`�}�m�y�G�x�l��1"J�P̭�%�n���@���8V����͛zK��,TxO��I�L��Qָ�4t����Cl.�A�~���$�8�g*�=�f#)����ߏP�{E�¸)&#o&��ϕ���܇��R�ϲ���D�p~]��}���o~ӫ���?�q��C?���eĐ��׬C�劯!�F�}��1z����ح�0�j@��EL9��큪�k���/��/�ܲC��h���;d9��Դ���zt�&�F<9v������mL�(j�oh��Q�H���΋�#.f�
��&P�Y׫�$�#g_�X�F�'���{���s&�G���*X-���P�^��+Y[H��!K�&^��Y�xK(�X�ZZ��-?x(O�q*)A^S�G,I0SPV����-Ԑ��<f�S4�͖�"���ͽ���*�`����-'k�Y�y��5���%zp{��kDa��%(��vT�Z�>�`1����6<�*��Zӕ���j�i,k��f2�H���HY��}/�r`F��e){������Y<\�@PDw�!�u^4%ܦg��R�����9GW<ZȲ��Q��b���$���~���K(�]�ML:k��_���;��$�:�[c�}_�sӼ�p��7�SA���@y�E���yw>/A"��WF�^cJTQi���s�j:�֞����4�߹���ӳ�wLcy%�G�n=�z#=���*"��6K�P�-*W�,�w�`�����<:��)���Bs~���x��PL��D�P��zS��s�[ƙ���dzɍ�"�n�1�:iN��|��¿���5���6y�	(հ�ZY<�'�]�/��z����fV�g�D	�J�m1���[�i"�:V,�SP�S��'���}ˊτW5�κ?1o�㗒yH�JTN��,��Y�m����ڟ�=�OV���b���)�d1���O|��1�S<��D�%�y���He��;��G'$ة����^�������b�u�T��'w`b�&Y��$k�{�f]�X_{&y1��z#�1�ǲ� � ��ڂ�<�k��;h>y�R��baC`��@�xn������9�Cc/0�����F/2����,��=���X�¿�m�6��$,�k?:U��m¶թ��6Fw�7c\0b�t
�ο�ń�4�C����F^�������5�f�ĲuQ�IE���_�F+��F�ә{=�,�Ҷ�ע��:b#��<���&�'���a�#�FU�-�!VL�W��(/NTP�(����� ����wu
���9у/L� d��Ne;�!ť� \1��S6����,߱d=[s2��	�	/�W�Z�!�\[�j�-]�̃��t<����.�O��ؒ�����Plѧ�*%�h�id�Ǖ8D��g0t��)���d�������`�9`���E�pl������/{���DV�m鲥>�Ln?cc�6�d���Es���
�B6�Ц-0�N�W>.Ta�L	�t���(�'�vۣIVP�s�⎐N���Y�A�N��Xݓ����+u!GTz��Fe�n��4���M"B�����.��~XX�w8�o�D��9����w���{^ÇzD�b�������\���y]kGA�R��	r�	�ס:R
x�� 
 S���p����jVճ����o��=�P�m�>b�G��i�
��*�G������|Kqʛ�BVv;����$����iLi������u�o$'��%�<1��o��\����y��'-+����ױ�k�n���vZ��	(}�}�km��徙֮]�Ʀ���f��[�~��<-	�G6&�@�տqkK�D���f�p����v�
���`m���i���xq(����"�9"]0ޓ���y�qn�:���v��y�}����O�J�"�M�﨣��F��w�^��~�Cr��,?������sX��\s��7��M��W����_��_�b@���}��zPԮ!�Tɂ�����*�G������5RD��5�C�9+�	��O@�G]޴v��p��,�JF��9y�q���=mKl�r[Z���J��)����$���MO�j=�G=��b?�'Avj�Ɉ,��
�F�q�Y���>���m��?X��%Mf�_�'�hc��?Psh��j7��ױ�?��f7�VGI���s��n^��Wم���d�(�sءk�g��)�'�z�]w�u�%�41��o����o61�෽�mnݱX���/yIg5[S@uY�>_��~�~7!*7�xV��18�4|-v�K���������{ /�	9�����VR�o,�D�����:2	d����C� k-��ɉiMTp�D�Ku�ԴE��=^\$ŦGy�8< 	Ш���5����E����iT��?���(�����n�����.U2�%�Ջ��:5s��U���k�:L�\y�u���-�\��ǾZ��w�@~����,bE|�w��C=���_b�]�^�EJ�ܛo�E��=���v]�����l��n[~��=�ȝ�>�~ g�v��=`䙝Y��$�)u�[�f�x�Ŷ|�R�ԎO��&=�ӯ[Ln��I8�����#�����޸%R����]�S���?���`_��ל��~�Wx!1<	Tc1<R+ƓO>�/�>�����3���ҏ
����	��Q����+�O�����;����R��I ���תe���Tc6���j,��CQ����Vj/����}vֲ���l���:)q<��K(&��}}.*o)J�n���uia=�n��s��݉-��-�J:n~l�^_�)k�WD��9�6�VS���8i����������#��j����'�3��ח��d8��H���E��e�'�,Kط<�E/�K=`�r��V�q71:n�sn�'}�L=�ܳ������m��<kU:yy��zꙶ����C׮�+��F�=��;��IF���>�9��N��3N;���^{��Ǽ\0�T�+����\d*�L��)���,J��~�}��fk6�Q)���
�"I��Ijg�3Z��<�x�#6.n~6�m4Y�p�I�X,�o|cZ���
.��`��Nq�9)g%�}�"svr<���z�Q�����VI����}���I�ޣ3���l\��{t,�4~?�WJ�)�K�)��g�3������͘k�ǈ��ێ��Ȭs�w��y�������q��z������V��hbZ�d�o�fO<�m۲�1�ի��I'��%����)��d���a���g��c�G@{��V���\�d�Vl��ەW��IcjĞM����~b?�$ؓ�54�'|��m����9�BW e,e5ؖŀ�Ǌ�aA�z�E ��&j��I��5im�[^�="_XV�g�Q��6�P;:�Pu2p4�	ୈ�a��4��HG���y�+/A�wI��r(Ы2\ץ��=<)���p_L��1�O�ڪ���;h�e��[bj����b��mt���^�!Gk�!��������M�~��ݓ���^
ts�>^�k^�;��#lb|��Fw�/��~�������l	r&I����y�A;����QGW���w������.��|��>ϑκ�c�+u����Sq���g����u62�ê��my��$䟱�]f}G��� ��:"�w�����9�W��J������g�E��br�>��F����{�x���}���*���;�Y����k�+�$'a��6T�+6c���덂Q���*9��-��_��L�+����P�G���"��9aD�"���1^2�2���|�
�1��n���(���X]���2�w�����GM}�za�0x�r���w��&���3s���gG)q�?�"Y�q._����*▍���g�d)_�k�8��f N�y�+_�kO_y����?�coV�o�Ϳ�?��?񹈙����?:6l����Ϟ��H��#���Y�i�9�A�뮿�N=�,;�����Î�N8�6w��	!���;ow�!����j'�t����X5�?��F[�jȎ?�����4�c��J�W�1۾c��%�Ɗ�k�a"�ُ% ������C�1���C#0\�ˢo�34]��t�c�AZm']��Ϊ����<*���������Z�^fA�H����6��"]K�������X�y	��>/ap����e0ڨ�
}�=�s�;���E��k@��;�����;�)ԧ e��4's����#C�f�3	o�S�����\�����^c��#���:�,�����!u�t�MN � 6��u~�9�V�f?l�=ro�)[�n��?��F�G}O��Q����ϭ6<2a?���X�'�֭q"
��=�Yi�y�^��X��d��v�y��iR[^5���n�7��r[��{k���"ob�N�ɢ�8E�Jε���<xKa-�9����*ңW�EQ,7���p8a�ެ��Xp���ٽ�����}s�M0:��3����R@ΌH���Y݆�U��N�������)�/�P���ΊMlP�*��y��*�8��ň���ǡ��ӈ5�E��#�TВ�'�C��b{	�={�uf
 �N9[ڿ�S$�u�?�;�:����)��X�|'xM`�[�pσܗd�2[�z�M���FQ�u/�����a�Q�u�s���`��w�{lx���v���E�����w!\��g�ޘ��ݝ}�����NZ���`j4�=Ѣ\��-O=h#o��/��{׻��X�� Y X}�����z�j�k�GKMp��ǋ�'��%�c�_���V6�h�6#ŲS�+�+�!�XL���*�|����U�}a����0��RL���k�+Ll�Q�C
4�q%�s!.
���	�+r�9��I	h�u����B�뭲[�e{aÜ�q��}W_}�{��f���|�����ݣړ!�9�{��s�l������MM&�0>�{a��¬zg9���z��f��
�x¿xT{�����{��ղK�V��*�_�����¤���P�ȳ--���
�����eu���{�m_�e��K� "mADE�b�h���-&Q�����"��b�-�`��BD�FT�" ҋtv�������|��~�9��{������ܳ\�ַ>�yN���]�AY�x��%/	��������,���k��qՒQ�>N-��U.���f��Y�x-C�(N��9>�#_%��lk���bm�m��R�f}e=�l��g]D�)t��8�����|�]���g��X���/�:�|�Qh))JUH���<ήJz�ĸ�X��u v�׫�<某��c`YW��؅�[#��i�9~:xp�VdG�.}� �>�>ѧh>*l�e�;4`sk��q8�}����Ͻ�֮���2d���� ���zu)^���oV�':0X�n�`X�|��$�H1�É- �r����� �F-6��A�bn�\~�_X��$6�`}��Q֐�?Gǘ�^i�öYub[�2�═��Aơ8h 9.�Hʿ��|�X� (�FP�V��H|��{�j"��~А~���x���V����7|ܾ�8tͲB.tL�`g<LQ5�L��;5�,���h#[�<�s��ʿ���a��Yk�=eH���\�(��?�nr�c�Q�hw��.ŕyvg�5�7l�Du�n$���Y�/�"�����X��<�Jޑ�nl���۲�J�2�eO��)���wo���w�)ny6]�W�8�)���1�0��+R�ʩ�|�{ʽ)�#���I��O���]�7{�����E�Ѣ^5R7�L2X��e�s��$�|�IV���Qԋ�o�L{�4��e�����ްt�n�)8���kV?֬Ò�W�9�^����%�Cm�3<��6������������@ ^�e�h�Ǡ���/FȂV�2mi�T�b�J���bT�H@_!�H�Gh��RӾ&J|XM�Q�y�b�",�u���.�-PW�����`R����V=�Hx�I���Q9/���JX�t����[n�3t��y�Q�T��r�%��:�[�떱��X�^�[���7|���8&�tW�.�v�����~�oX*ЬZ��/n����Ï�vTN����7��Ƴ8w�q9}��3Xy�ќ�MqKK�e	ζ�egY��|$P���լ<��I��S��OsǗ�����>'*��������|�0��.�̌=��>��]tQd�6�o��݌qu���¦�=Hݑ��m Ϙ����;<�ȣ����]����"�2�z�O�4 |7��J�և��7G��~�3�mrg��w���M�{�N��`�5{n8ꨧ���=.,^�gN?@?OY���s����Y��E�j����7�y��=�4)ShK[���p����(#�Q�=��l�Դ--,�5����WD�8�a����m�<(�����%��P;$��u�3CT/a�=��fox������j�8��#�	+��:�ظ�u����?����R��"��dfZ��&an
��/*�+���85�}��ap�?�ߡa���	kW�
�7�7��yX򥳣'�^Eϓ*K�����0��2@��Q�*���}p{P�L�|M��a��2��4�k�TO��C�7����a�\���e3�o�6jz��Z���`�	ƭ�>V?�"���+W�Pm>�⇹_���I"�s�!����懧���s@��Ca�ڧ,��v�,�=�[�(���Y�B�7�䧡�ws�M�Im�����vا(��	�	��VC�˾���j�S��SN��˼��¬��aϐ��VK�x��|�;V��V���e��x��h�nv�@�ɏ~�c��a��Z�CP(�n��۲������M-��q}�-ʈ�K�N{�*�s�����{J��n��p�Yg����}�d��#�/E_@��
B'�+�/�z
�^t�������9+,�u�%�}�'�,�������_�첼��r$�-���E^�&���/̒QI5m���L����ζm蝑Z-�6eE_�r�e�a�k�+,_��W��>��O�M��T+�_��B��@��mT+����g>q�rN����ծ[���%�r���4�<��wɋhDR+	kO�,KO	6_il�`����%?��U�V@�?0ʒ�_.�x�ڟ���U��:0����y�v���(9��Q��Ch����E����?/��� ~��*DЧ0�{(���;�x���g��Hݠ}P��_�����|.�J�'�]ͳnf �:�R9>~�!�ED�o�`�P��}����eM��R��c}�N��4���~�㟲���^�|O��Ю���#��!%)k��MB��e,K��O�h\�"b��7�#̂��0�ꈕ�+6=d+
�}��TV�k�b-�����yN�f��G��U����
A���3���n+�&������O����?G_d�Ϫ�):��/���i2E�U��v�IR����i���f� �{O-"cf"�r�?�A]�=B�_��W�k����eFY�E�<?��,3\{�V�s��#?��T����f,�_�Ѷ����0��=���n��PTG���R��&��o��P7�6����yG��޻�W��+��s��i�Q��C�AT�°H	8 7S��$�E� ��J���ۙ%�dmx�6��-B@=�M~OG��X4"
�RĈ&����j�,OO�e�����h'���.ޞ"[���5LjI�GA����������&MGƃ����i���2N��E�k3kV�Q�Jɐ+i�r�r����W��($�y��mA96%w5�՜E0l��/�B�&�\��%�7���1�ph��~sK�H�:���>k�H>Č��j3�ᶞ��?U��9�����P����z:�j)q[�,�tp*$ �k�z�ue�{��&Fb�t��(�d7���<�y ��+�q�WGY�ry}�F��� =7�?��s��t��X��u�v�U#j
�� F�LDj���m�r����H,
o(t�SnO���UDcK�Y�'B҈:z2E���;�1����KII���@eT�o�q$�~�9�OCh5Q�0�<�@��H��QJ�s�/H�[� ���/�c�h/U�(s����z���������>���)���
���>M8;\Q�&WR�,��lT϶�,�� �b���k!�|�;��c-fċ��ѷ����',E��1���[�Z�|!J���X�s.B�t=4h�Y�:&Ÿ5���h��=T�������Gu�X�;���Sr���)���=S�xD�!�U�Y�IcE`_M>٢1�á$;���б+��ΈC��ԒQ�D��'��W�u�Um��)<�n~1��8 y�˅�Ȱ5��f�%BX%#�K�~���=X�J
�n��M��Dj��V�K�����?KWm�MT6��ь��U]����\��)�	�w�+m͗)�Q4ΙE^�p˾� �$at�W�}*iE�h{���qkI=e"��m&
/�2%�\��EMqT�Y+�;�[�PQ�Mݴ��L�z(sQR+�9ޘ��-诮k�/�m1f+�w���dS6{oᘸ�,TB� >�篙Oו,�&o��y�	�Q(��s��)�Сs�O�_����2gNOn�#D4��Bm7k#y4XN�Q�/��C�1�a�V�6h��e_�J=�7��Zr1�0)%P+��>?���)�jV�7W7��7V�Z�u����4T���|����{�M��=��1��n6�=)"OC�WT�Ÿ���0��l-�E*/�,�re�v�0٬ �os��$����>,�d<��Aw����U�E/�!�@��C��X ���/}I�m��ro��]}��Vs���dJ=��Ʈ���/�xw�dd�"R� �'bl���$2BX��x��DSH/��-�7.�o{z�,�P�s�m�W�(�]�R��!:�d�y%M�p�J�J0d��\�aK�A�����~�s��y=���<�տ�Y����@۰c��3���Ot	B<Ǹ$�c��p��Q����b�����n��-��1�T4��șlM�k�B8�evi�x|�+��T��RMR�w���B�#d��q�$�uHť�b}�"�h���Ȫ'�@� cJ�ʾA���d��>~��*̼�9����5�8���d+���IG�*�5�&���Ƣ΅��k1�$�ܟGQ|��������x�5؂8,�Kc0����馪[ �a�m
LʉU�1G;;���\(��P�\�|LZ���u�!�ƿ���Q)���l
AC��\JW쁡T)��;�)r�W.���(&��A��H�=�C���{p4����h������g<>��̍�&��8Z� P��j��eU�I�s
x9��;��H���9)t)r>�&�硲*���#
=�O���X�"ߏ���T�E&[��ĸ�CD��*��h�Z��
z��-T�̪/%#�Gڽ� 3J5����ǩ=V	��~��&��[����\�W�Q�y������5)Z��������aJ�T����E8��Uμkiv���~���7�@�����J��9�ƴ;�o+2��x�::+Yf�ìl� pߌ�;k� 7Tqq���F��7B?�Z#񿑞�ږb�����|%<^��5�h �M*���B�c�R��������H��EM��\�{�"�7����;�;O���;�֌R:;���x�o��!����iҎ����g�C���Pv�Vݛ��g���c��E�wnM�y0�chA�}�g&�����3W�N���ם����`�ީea+Bf�yXI5A}}t��2�s<a�i�����z�IM�3���L)[��m�H�T�)e0�5��"@
E�SL�m�_�BXF%�)�k�c��L��SD~x��d'���O�z�a���m"��V�7c�X�_罴����}K��z'��|��exoK�TA��[�mlb�ް��'=J�x�޷���ֽ�tY�=5��\�3�֊�(?'u���|�ӣ������ȡ�S��Q��T�F������Z�q�CU�$��y�Y3iy�!����o��Ψ����)nx޼���a�:KΤ��(aҹ����M��h�7JVB,������ ��/Z�>f_T�� ��%哽�8�9mmry[$O��J9W�G��U�x��=�x��<9-�x
1�Z��S�L�xX�{=�Z��S��)q�v��&)�V�I����"Aj�a���[�$)%�v��a���c�h1U�I�� 2\��&��h�VO�q�Q����PV璵��r��y����s-,M(��`s�V����:`�A�����,�ߕ�����p�QG��sS8]�\J�}~}˯��<��Us"J@M�y��3��{��lq Aʊ��_n0Pߔ��58<���@�b_֢�W96S`�|����~���� te�q}szYt�WŅu��3���
!�d���������d���־��V�1�R��� �c?��f�7���crkI��b���?����j�	��� �[��ih�/������B�Y/*����ہh��K)�)��;��}�1F�ĢE�æMBGg�l�y����52+J�X�K��a��/^b<�rw�m�d�v�a�����y�T�9�~��������o;��W�J��q���w���ۢ�"��|ޚ�R����)Z��f��Dy���yL�"�u�$W�����.Y��&�S<~"��H�z�/U���@D?,�e����{P��M��D����8/�4�y`��+�YN�o-��A��-��Uua7�l���x}QS�1T�e���3�����~�Zu+�
�y���c�1Ѐ�)��y�q����~��[r��$U/'�iXq�I3��Be�%K��A� ���AR��eɀ%{W�^c݆@[tvw�=�\�X�$�_0�������������{��^'�/pMn��_�j���Q"�R���/���(���b���=yWq���B�ޢ-�#��믿>�
����B0���U���+o#���xg��Gl�	��ҡb\�;�L��E��Uա��>g�y�s��1�W���>�_g�>���=��¶���q��?�����=蛡t J�����'>�<Q�y�E(���;#r���[��H�QI�D�澰ے]ü�¢Ż�����ʹw���R��k��^������J�ț^��4gx�s�-�y�TNK�~�âӢ��O{z�k�ea���V���f��C�A��.}<�ce��DV���6@��XZE_T~>\����mg�Z����?�c�¾Ta-*
�;-@=	r�P���*>?��#I4&fb��6�B�\���?F=lUU�f[%��,a τ���%����w-(|?��s�T�2?-����u��`h�m?~_%�Ѝ�������*��g?ks�¿׾���P�P?|򓟴�#T�ƴy<���#?�@'��=em��֭��"�i���Jٶɼ��l�΄�ǳ�O{��L�ɝ�g\�l�p�����&�|�/¯o��ݐY�������=�����p��Ǆ�p��X �|�t�bWEA�k���lٲ|" �JV�౎���'��mU�H�6����,l!���F��b�ɡ��呕�a��}�"=��������~-�o��|��0ط9��prȰ��Hj!-yL!��rHߏvr�c���g�����և/~����LY11��ΒmC���ů;���SO��:8���^���/��b[���7m;�9A�������@�>��G�7�����'���=��~����"�(�:!�C����|{z�V�a3^�w���`�شV���n��e(*�êU����-���a��e��]�f]�ߟ�8�\�.�}�����'[G/�w`аYYY����c� c(yؖ�+R��OwԶ�jR�*#�oB��;�p��z*�4�)������p%+�V�U#�z)q��0̖����]��C��ې0�1E8������'yY\~�������ֳ#�0.ޠ8���z�E
LCu0��ۻ�=��*�a�����Ɯ���S�ׇ˿�p�	��7d�'�n���p�]wY$b[��i���&E^p�E݃��|�����/¼��a߽w���#a��}��b��֮[���p�?	���ߔ; �fbrr� u#�+ĀO�]A�����}�(i+�)-�e���"�C�������~7S�s�N�<GOs`CV��5� �~��hd%��Y��?I�Y�U[J�Bt�kr/��HG;�C�����cm���߹"�wιa����&Z�ᔓ�̛֬~*=�x�4*UxҊ������Q�$�a��Y��:�?@+�p��>�W?�fU�я�.�=��2�p���L{�J�#~��K��i�{`s_�;�ۚ*<�όx~ظ�'fq�rW6[l���u�6G��Gm�?�\A|��Y�SLX�
��'b5!�|�H[��-�l��hY�SY��y� ��X�a�0�ը���8��Ba%��b)U�fϙ�'�ߓ~/.���^EV�x�V@�/�
�^w�u����N���뫮���,���^>���Q � @��#�S.U��o�i�c�°�^KB��ު1 ���\w��`X�p~����-w�{����@B�ΪUOm�M{�_
�M��;��sٞH�C�#��0��qY�������\�a[X�<'	,�/��~�����;��=��!1��f1`��җ�d��3�I�D�ôe��p�J��h��^1׎DB5�bHJJ9�laӭtf�
��BZJ-yC1Z�n� �؜ΰ��Ѝ�T��I� ã�?���B<��Wq!�hFZ���O��-���7�l�n�Wy�w2�V�ZV=�xX�����t��l������T�2n�Zm�E@����L/�0����c�3Ꙕ��p�7K����ņu�CgY��MiqqʤV�6��$q�2B����� |F#x��|�.����t5e����
�Lm�W}�#CuYM�=�C<��"�r�`dl4./�åa�XH͈ޔ�5\F\ �� �M
?QØ�@�P�ƅa|��;�y^�2��z����s�����/��'�c��) Taz�CwO�u�d΍%�nI�4�
�Sփv�k�L���o&)?�4������Z���S���:-�M���v�OWGw�<0��ss�ӀQӖ����4/ݼ�+�s�9���~`�_����芧��֖����K�no�<�4�b����Q��r<�h�1��D�G?6[�5*�ٶ��u;O2�>)e��Z�	`��::��M�_砤����@;���Ë��E���/�x��q$��k���4�+c �Q��e �}�O<�.�E�ڊ�Aӿ�=��Pn�R����`G+{����ʺ6̟7� Vs,�?��tǬ8@;�������M�;��I� �"�Í�"O��$�2 (���#�?���?��?�/|����W��/(���-����S��{�.���6<)Z�C����V��k�eo��������'�������2ۢ�j��;j/(+%��E��*tQ�y���z.�����WCw>#�G���X?ߡ0�a�
ݺ��tu϶�J�fx�����5{j����ua�^;�6�gI���%�R���C女p���+��nV)u�q�psX�vSXs�TI����6�n��=b7�?�b�<n��ִR����t���Ȩ�;�n�.��_�o�}�C��N+\$���e�cnˎ�ɄZ'�TQ���(i��0	�t'�P����ڐ%q��*Y��?�i��xF���O	��`t!�d@���.� Ý$Y�_=Ҝ��-�fT�:�֦�����a}X�~]� \�g����x��C��Y��N4 ���MF�F����	�6�
�V�����{-�#���;�7���W�5�����Īա��k���ƀ�����B[�]K�i��s��VD���p�aO��zsX�a��*����[騄����~����ͻ��s�N$ox�����jx �@l����g�"�EEBB���Ԗ����5/یs�_u���������uM��RW��U�P5mi���j�����\��_���Z�v���-�V�%�<1�j�ق�!v�����I�U��9�<]�O�����{�Wx�oSX�iM6�g���U�[I�ݬ�粽�I���Z>�߰1�u�=F):���d�S�eȚ>몃�?�C³�����Ǎ��'J����3kd8����Z��QO;&�Ǟ����k�F����mA�g=�n����j� H�PZ~���t����-h�Xpmi˶�o���� ��w������y}���z���ʯ���Q;{�_�|��&(o�=*��>�ݴ�8��_g��W(��ܠR��\H��/|���^�2��R�c]�$1��0�|�~��������t���/<����xU2~��v[N{�s��
s�.�c�����]w�6�t��;c��5���T��!�w�WZL~Y\�I�{���|�>�Ʀ��G2g��ea>���ub ��e�p�~���VOa��
�ָ}(�W���:5ߞ�(�����J_O�M7�d�1ա����(��� ���O�H� Ҿ���U��J�����i��R�导� ��9�=�г�q�f�!`���A�0���9>u���W_}u�m�Ea�ys��y���f͞V�z2��m�r���|�5����7��^{ì�9���U���o&iB'����������a�����a��9T�����oF��~�j��FTra@��+v��;��U�<h-�do[vv���
w�[U���o����r����zܨ��0~r�?U��ߛ]�z3�f����z�*�J[7��,���
�b���׿��]�O����(~y@ZL��^~��-�=k^\ ������@�ي�2cq���QGt�u��{��U+-<T�3��m���q���Zޘ�%��/~�?����7�����q��W��6���ׄ��+�巈���������fx���;�>������28���w;�Iy[ڲ�ģ{<���jCi�ݼӮ����m�$���y��6��gaTY\
`Ͱ��l;�W!��"�c~����I'�d�Y��	�b�Q�N��������O<eq'|�;��:t�;(b�i����On��y����S��*�^�7+�R���m��fϝg�W^n�����u���LY6i��?��n�:(-'��!]$�����>����f�q �/\`!{�ψ~�c3,0a _�5=`۲}e���L(��̘������@�u�E��8\�`��vBj�S�UΊW;�ݲc2�Y��r�c�D2t-~��`��>I���_���l���MA'9�o|�F��^Q徘z�B����|�*�n8萃��˖[�?�G'<��#�E`4��\�6ܗ�3�B 0s;y5asey�jg�ǒ������X7��?�x6,2���B�=����W�j�\F�O����
�����G\�mi��*��0��ϕ���	[�V����%�����{.F���O�f��Y�[��A�VT��OA�5x.�³4jBA���O�~�к�{�F� �
���Y���Z����O�G{4k��:+{h�����z���xB�X��}��]�5�`-tf�a�q�ש�Q�d
��J�!i�!�Ց���^X��/�� $9������e��V��(`[L�V�}�X�FZ��w~K�@�������	g!�<��/�	���5�暩�����:�*�B*���{�"X`% ���~};P��HH�}�mn{J����3�Z�V���Xv���ζR��Ŏ�ي%tS��
QV�(�T�b�'�ݡLq��ϊ���H�ߏ�C�{�Ï~�#�ü'����J~r�$����c�CF]�і��7��V�e��vU�F_�P��J�⌝�ʟ�݄m�TMNu�g�k�E�Ɓj^,}�9��L>�z�<H� ���FZ����7�).&c	�X�WyAS]�#XQ"Ucb�
y�y����C��Ct���#�+.�;)�c�>����[�o�_�}*Y�R�o���']F���X�ԓRP� ��^��͏J�¼s�k&�jod �����_�����Ð�}��`��<PO~+䞌�����1�כ�(���?.���Qyc��^ײ�6�^:9�܅b�@�(�z�[�j. �[�����e kLx`�f���N-uo(k/5nbK-�$�G�=��A�K��N�Q��{:�f�Ų�EQߓ�>
j½p�[XB��Z�@-�gX���u����MI���/�B��g����D�@��(} �]�V��9
�3���[���;��1���p4t�J6�E��E#��5��(es"d��>q�_#��j_�̜a�R���w�{T�W�͇?�a3�t}8jd���Y]-;���%���]u��M���p��W�(� ��|��A�í�x}(��hpȂm������0�({�Ϛ*�r�?�V�T/2S�FEp(D�b��𚸈��=^�Π��E��<(zAh�e�6F)�d|�����I����ڱ�A�����D�_�GJʟ��$eP��@%>(�8I��WD��͵���ͱO��fVO��V�Ŗ�R�fd�o�3�<7]SY����~�%�Y#�Zy`<��m��fc�^��k�u� MhgFf��yK��rke�+�Z��/^�r�/p��`<��ۥp�&D�%$&?�#�`��R@^���5�e�*l#��lb���>�*�U�Vc��-�֥ב��B�d��R<\JQ������^�F~�����Pl&/y##0�P��țsF�)l%Ũb*?~�@d���K�Y�v���&��l��ª����Q�@�t�t�b��+Ua������Gख़��gˀVV��f4��6���暊��z���sm��3����tq��W����V�~������R����uq6?��=��?�IG�&-����($��m6)E'%���>�z�>�.Z1�k��&G&�X�:�֑Gi
��@��>���}�/�]�\�ue1s��7�Z>���H����
e"�N�FU���0$����jH�Q��������1L��������<\�7m���I+��c�!/Y��pH�o���?��&a;o4H�3��a~�9�;ƒ�����FyzJ��#-*�Qa��s�O2q�~��W�IǺ�z/r~c�(H�,�}�))�)��G!yإ�<gx+�_�c�X0��؄��,�~eD��M�䔬���I�s\�dI�O�gAn��Ip>'�A�)�t=��gk������,�f��ZȔpTX��%�s���t�:�9'�!#�EC��z�#�����M�K?#�~�;JF�2589�]���,5lJY���Y�w���04�.�T��0����tTlQiz�uBz���jg�j���9���t�VR�Q��ku��ʴW���8�}�Qc}�V�����z)g%"�KO�UB���C�DV"x��+7����?
DI-����1��krj�q�b3-R��z�rC��5cA=K�ԑ͔��x:&ŏ9V�[H$��PD
1�D6��;j(�筧�{�~GAWh��=��A#��b]K���Q��(�;�<�&���`S�V�J�S�HcEH1�-���܄�Ac��W3=�~kԱ��fe�Q{���к�J3�߬·R�j8�a��ڪZ�IȔ��:-'O-B�db�zG�k�'��/�������ڷ��5����J $q$pa3��w��h��0)�=��::Owg���j�����5l�^i������2���#-*����^�h�q_�&���r�0���=e�g�CǪ�i���PЊ�9��E��YH�63^�o�;
����N��!;ϸpu���?d�,�t)�Q����@H�{�+]'��3؊95��0VA&Ǖ�sOZxձ/�0�E�;�.�nʍCc
�:�s�OǤ�u4�Oc��i���a�&�c��]w5*VU�z��Q�d78M�=Q�����h&��w���o�a��e��
ӣo�(�&�b�<� դUa����)�YY8R�,��$��ީ�gx,�����'/O�s&�
�
!�R&��QQ�����ߔ���(�z����^�+��<�Ƃ��p��<U�1�h|)�%e��������RE�'#�X��?�C���?olճ�uZ���e�]L���	՟�Z�9�:�����PP�'�Y{�4��	a�Y�������?�䨄>Jm�:ʝ��m7?���OJ��P�E���_V�x�]`�KC(�j۷y �}Κ+� �u)b �� �_~y>0&�:�.�&.�L���g6Pe�kA�v���,]���j�l����W������=TL�
�M�ܟJ�'�T�7�wW3"��b�0c�q�x� Y�Eԙ�c�#)�E~"D	LY���9yT�Dqr���sնx�׻���TG)�V��/��\�Ej�:�K.&x՛�!5M<G
�)�$���+�cW��y�ᤓV�=��==�J�7�m��Px�Ǭ����z�Ø�[XX�ɴW����]mC��3�8I����n����M�q5N3�==i,��U�BϬ��Y0���B~<�I�l 3�T ��&���Am1L\���Kp�f	[m_1��!��������O����b�^� �$��$/�Rca*����(�K�$����Q���E�(�F���R�0�S߂r�a(D! ~ON��2d���z�������﫝sJ�Y��XT���t����W�e1���{x�P��T���q���q$I��!r%[�jIX�d���z�<��p��ׇ+���NW7׫�<i���6��M���I$��N%��o�J]�d
��|����c��@�%�l�ޡo0~?��B�pË��v����D�&�?� Y%*�A��'� ��K���	ca���<|t��欣����u��ӻ�
oy�xkE@�[T� �(j��7����t|��b"EJU�A��X���D�U9	��(��Έ3�3�󂹧0k��TU,�w�qǍ���ʯ+4+��T��74&tnԃ��cn��؇�FOPV�+����ܳ�	'�8!�KI�˥Z��;�d|��q� �6�<�0�<��ʧV�cc[e(�ZCӗ��l	��>��/�ma��w�yG���_��}40�
;����V���?�~'R'7����&�,f�;�!�� 4lrtt�A�i�X"�e�w�.U�
��f�2�����lU�����
1�z
��(>�������M��SY�:&�z�F��>Wa+�����1I�,��_���S&�x!�B�SS�õ������4��&�����3��R��������[��ݏ?.|>��`���o��d�bU��v�iv�4����(s�'�|bڏ ����3���w�֬[�ſ|��ê'�O{�3�ҥ�����-^�]���Ӱnh��e�Z�%cc[�|�֝^�����љ��
+W=���DK�?t�l�bQG�7�p����Uk�QO?6��*�R����N-�<
Y�~Mz�bXF`�{sT���#耱EO�J�AU����G;,|�<����ĳ��8��"R��{x��d�VP�����E���d��ZBQk��W��ZBaފU�x�V�.��'�=m��&�E�|\��Y�F��ys�KKR/�m�������4W��|������}O���Ҽ	����V\��`Q�oi�R����/�{��a]T��w���9,�M}����~���p֙���S�@����([�ʴW��	@1���Ι3;U{�o��M��H�Kw�����?�)~��.�����}���?��!y��7c���z�^hȋO�y6YXF>��cͶ���#4�X4X��,⛅��
p�F�E*O�;ؤ�*\�7��d�Bl���a��yy��M+�UQ�D���J�
�H����"b!-g̞�{�y�Ɵ �����֬��p�C�5��r�~<�Z>^}������o��C�f_��O��p��[N�s�?�lI����
룞Y����_�bx�E�	wYl��#;2<�Уa<-�g���	tW��K���m
s�v�[n�U8���򽉟�5k��;	����as���zVX�nc�����z4�<� m!�x�	<4yx�^`�#{�'�MdYy���������O����C 5Ƚ2���h�d����^���tN�!:��]�"_Q1Vު�ڑ�$�����mC�WJ�U�L3�7�"2�\|ިH���0��[woC�	��d[9~�ܥ�{�dk���И���?�"�EO��^t���1�c98�F�0�U�m֪᷿�9��	a���>4d���ӈ���V�z<>�V>��z�r곭Q�A~�ӛ��F��Z�.ȴW�I#��RͲ�W���3<�أ)�H�ue-�Y��G��ąN�E �o����`g�y���TSx�'���/�5�җ�4��_�e���'ێ�j)�V�r�-,N��aq��M=�d[�SY|�{�e��D��?��Qdx����˛$L���ӱN� y���i�B����~���r�O<�8��
�%��@�+W��{�p��ˣ�9/.��3�� J�[�TaRl�J��<��,���.��#�?��p+���W���PO�B�ء,�����!+��������>��+Z!�ërχ|'�/I,P
,x~G�׿��f	(^���b���M�����+c���V8g\e�QԬF��9��'ק��L�թ��D�PR
��o�C���y
)��~����/.J��0�"O�WI+<Hn���%��+����}���Q�j�ĸ�GT��
�R�3�W:�EtpB�8�fu�����A�E���<�#�^����jQV�j�u��7����՟X�]�ܙ%]C�����qM�:�8�,wA=>a���ĘZ���7B�8U*�jB�4�!w+�˒Ŝ#�gC6�ERS=��E
��'baf,���~�|�m��62
�Qb#�0��&Y���IǦ� ���檼`<\B?��Q���+�'�=x-�a����\\l���e���`^w�Q���OL�uk���W��ು�ƥ����[ݳ���`�YJ%�!�^*u�M*UR^n"�{!atS�^���O��2�L�>�{���y��U�F�8�BGE�f�E���L�\�ĥ3�K^���O~Ұ� '�˼=e�A߶�GDʟP�^O���Cё����~fFA��B񵒱�C@�`
���G�&��	'�`s[ʜE�ӷ�������T�������ƅ�V6�r�_�V`��j�~{��.:�3�#
�&���L�z&}�tRp�kf�ww͊�¡��Fk}m�Y��h�f�QBgX�;�Ǯ�W���?�'}�Ї>d�>&(�?x j�۫ց�(�y*%�&+b4T!�K�[U�;j�E�����F��-*��)  �G90U$���J�W�J�z��b�Ó��]:v��!� ����Kx�0F�(:'e����9�ȧ���k��5���:u�9���u����-�bŊlA������UO�L3���	�j��O��]ʉ�3���{Pxr�C��G�aH��*�P����[������ ���Zgq�f�q��)��(8٧>��N)@�>	5��2��l'%(�O�xK��
�R[;�0QhB2�^�>�-��4��c,����\�\�o��2�h�񊮗�E4J���Q�V�}��P��u��4�p��>���'<��á .��]�E	�gO���ݢ�K�,��E��v0b^H��<M9"�T�_ٴW����#��}�s^�={��5�+,�.�~���~���Ҙyq�8���1ǝ:����V�V���
_��YU	"ڽa񫠊���<jH��2A�Of�_��2�t�bX�8����w�(�;��d�c�|��4变r���ɂ��fAP������@�I�&���������������}����k3 i;��cC�^{Z���ݖ��_���0ؿٸ�6m���ts�qǞ�v�3��p��	�@J��3*�g.�O�2��:+�B��������0{ޢ��!G�E��m�;V\n�.w5���h�@�I%7���d ��ӟ��n�����  ~� Ą(E�KJ����SF䕨���b�0����D������־�4�CV�����lq��
������A�|�q��L���D�w���	>=���¼{e��KϷ@�v���s��>Av��n
#z�~���1��%���·{ "��>!���Q�0>��������]w�i�Ϳ��?��N�,�T�` 1�1��$�İ/`�%M���G��M�
!�k�C�3�f|݊���wb��Sqt�d��zvO�O�����X��w��k�i�j�A%��aNT��.�?�x��E�=w���:��|�!)d��6n�W�ϕ�_c��]��{+3��O����K�f4��=[��Z3����h�����E�ȨU5��j�0�:���M�!\pAx��^��o�&\q��k_��YLLmW1Q�&k�S�>b�����K�"��k&n9^xb�hdbiۂ��կ!��j���I�ce��NQ��s£)�*�@�d#��+�b��c���$�}G�yOD��"+��'���WwM�P�B��E�+��B�B/�h��_�<�����@B8��������E�r�,
R�x�į/�����;�1�c����)��H�D�9�1����s���crO�f��o��`*����d�׊sa?P��M����4��/_ȋQ�󊗽܎o�Ż�9s���?$<s�)mC��>�9�P� І�%���)4�zjB)#�O�z֩,J�:_է�7��$(�!_@�]Y)bGT�NJ�6��`�Il����@r���>` ��\��p�r����0Y�-�˕U�;߃�.J��	Cų��H������{r�RZ:�S�B�Hd=QX��/R�οނQ�.�G�����ENVe=���}�zh��q0V�@*���+�}��Z�@,[�0�}�7�*c���£�������LfOx�P|��zECq�T�KIm�k�����~��_<�@;g#|G�~�Be��wA{H���CW�f�q.ox��E�C,<���/�\�1(P� ��K�~��~z8ꨣ�;Jx~)^3���/䞆�Ȍ%v�����WX��z�M7�
#i<ł��Z!��TYV�D����o?+�Fi��]v�e�\�w���h'E�+\�5�Ӕ2�I�q�9�+_��m˔t�:�!0�Aqބ��;����;L���t0�\�Rǣ�g�{˓�c����(���̹�]����X���z0Cmϓ�),e�C2��T u���gE��!U\ �u(�(�;�qSj-����3�Q��\s���/Xؾ�	�
�"�f������?�+Xy8@�Qp֭���	�O���Y �sl?ߕ{�x�o����g���O�$�'bM�}��,,X�Z��6�	p��싱��x���x򋱮�t��w,:��X���g�5C�Z��`�q=�y��F��Ɍ�zZ�Dq�
kEn�o�"�M��h���{��)��b|>
�N�@�L�`Q��m-��@�M���w�-&���x�O~�܂`���/�{�7V>��$

YҜ��d�� N��eeyŞW �}Ja).�܃����X����+9=�2Tx̋�ڢR��)T��o��d�_�t>~�-��Ň�t>�影Qצ�IP¬�Q��΢ �C]W�	{0�x-CB�E�Oޯ���<y}�7�a#o��Ʊ�m��x��[����2�ѥ������m�$�6ʱ��x ��?����{��^{�:�	�1�(��A�����9�ЖI����3~�G��c�'���C�EI=]\YA
mx������c4W	J���X�X*��b�a��O֤� S[;3�G�_)|3�'��%��%7ٷ{�y��XM����x��5X��GǨ��rqY[���4pM��G�z���U�P�6R�XO�c��ݓ+(�O��ׄ�qY�+�~�H<��,:)1�g���|2��̞~z,eQ�#��Z�-�~z����w��[�K
VcH��C�}���3�SCH��@ʠ�exCL9,>c�1t�����Ka�H}��G�t���9/�/0w��_��WٱC�v����X5�}N�/�X�bDe[\C�O��P�)%��6�><���ذO�q���|#����nAt�"�|q�@#%��.��P��J�MF�Y�?ɋ�d�MB���)��OhY%rk-ќQ:�[ ��z�%�BԾ��P-Z]�da!����?�SM���J����$X9f�l�� ���D0� ��x+�uU��{����Qܗ����a����l�+FΟI�dS�h��'Q�,��(/ΗEoO�J�EPJSR/���ל}���kxl��d趾��ay�׍k�}��5��uQ�����cD6�[J����!$��'�M
�Ѥh�țf�a5��߶��·	������K1yY�7�ٟ���;�7\3§�w>������w�Q��uև�Y�Q�Ωt�s�y7{�\�� �cp6�z��a�&��\`o�!B�ԋ��X�B<�#�G��� D���`>~�d�,���QP�E
PP7<�I>a+/AJD������}�Rg�qFn��!��J�Q���cb`��!�K����-������^JL��(Y�LL��e>���d��Zם�1�u�@��mOׁk&��~�m���|�3��/6����d
�Ca��C�0Iz^{@?�|���X
�#�|e�)<H�k�H8��
s� ���J����'��SO=�ƙ��
E�K��s���k���4�4�=�*���xd�(SZ�8O�����d�)��v�NT��%ijOpj��a�>8G��]�앰ւ�ךk���n@縵R��8�������U6�����2R�>��x���b� �()[M\�A9�*B2%KE�X�P���ؒU?9�ө���R*��� U3���ۿ5�Id�*�^�W���T��hC	̕���Q����(��4[�t<��|�+��ҹj��9�""h2E��#�J�^0J��9�z�ߏMY��������gD^'���'>a'��v�(k�G��vAa�X\r�%f�{�[�iy��7���"��BCR��X�}D<�Ya%b�,:��\�����{!EM��d29��H$�-��_�a'?������Y����Lsр&~��镧���y<dybrJ��5p������Ʊ�� ���#���N����{�]w�n�_ F�m�]n�$��R��`��*(~Vᕼ�}�3dぞ�J�+�Ȃ�� ��N*�=�n���9:�f��q~��"�?�S�I���V:V-��/�5�����%��-�j^���,s�÷��"� ��R�4%�j[v�裏��|��W�DM�g'�t���p�KɃ� D �������*�$i+�F2�y%wQt,v����{����o�KȊW�/��bJ� ϕx4��%����Dj#�6��^"�<���#EĘ�e�����'j��v)��\�;�5�\����CM�Da�Md��Z݊댧���
eP��"IG|]�p��y�"l�U)�c[�7ҙ�������X�BQ���R	b[�����A
�)�%�4��fA:6���Ci�UO��	��|�BB�7�Rj�����
�u�%n694h}�M�6�+��F������*�qP�O�KK�3�U-�_�1S�L��>mIe[c�8v�R%����ڗ{�g(
�~*[A�YӢJy���C@��e��Q6�3l,��k��������ߓ��WS��Nŏ$�����Ҵ7�(V-1H�C��U�XWL\�4)���~�����b�m����ZX�@�����(�w��?�m�Qm��(Y�L���,��s�U�3�����a@���E��1���Çu�:>�x�0�_,����\xα���y����D=T�T�i���{�_� T�3������^n�{_4�s�Ө}���Ry0�<N;�ܪ�ّE���J㷼�-�}�z�8�[��m�6Q�{"�` ����+_�J��!�O|߃�(���/�+����R����B-�����q��m`xlM/�F�P�^��TV�ȴW��=�o�!g�D�z�*��!FK�"b����CDV��T2�Α�,�?������\�h<��x-cS[ƖV8{Z:�H�׼�5�ȧ��<�*h՗ZL�(�������s��/��3Qt��G�ÃT�f�*�Y��yHo#)r yU������/	Q��2�?@'�����d�Ax�5��0�ô�s	���	5�:���B{��G!(�6؟&ߨ������6�,��a���>=����d�����o_�p͵�U�O�tWg�q������MZr ����+?&D�i��&؃���[[W�R����B��b4<h|M~������X2�Ǌ_(���
K�"����`�\��j[������(�ָ}Cx�����k�r�=N��y b�_08Ny�~�C'|~�G��A�!Z T9��=��XX�,>$�	E��R����G���������Sjܔ��Tf��/%;�寄����!zx%!b��Jx�b?ȥT��e���-�&�`z��9���"���B�!o����G����.E1���6a�f���bbX���)���R��<Q��W%F��4O��b&���������o��
ay"E_��{,���C*�!���������X����u�[��Vر�xE�%�N+�B�o�<�?F`؉E�@�T��^
����ʁ+�䘚ë+������9dWPȂb����rDC��[c�f��I��}c�q�>o��V;z��H�n7�0��m$�ے���3x. H��o�h�IE�+���}�E�����ٶZ�"���V�%�g�D���E��_�%j\� 
���k^͇<���rQ����+�s�8�����M\vV�ǟ���ʿh��l7Ӈh'[!,!^snX_|���'�{<N�X���˲?��g���|vu�\G�F�o�zƭSA�=�xA6Fs��E���7��DSma�;�!h&r�Ց�S;p}��s�?�g[R�u��1(G�X��ͮ� �,�,�(Y�� �4��<+�((*�����18 ��,�Z %�C~�Lh��&d�3���2ɇ)?��T���(�ڷ���ۙ%���TM{��lugV���n�s)��9_Q�X'
Z�Lաk�I
���iʚm͝=ǬtQ8�j:=�����r�-��ũ�dR<ZU���X�g�u�uR"�� ~x��!�Z�#+�,Ă*ب�rK�E`��/Xo�Ḋ���U�3ް�?��O�7�����_��_�؅�����YX�4Ua|���4�-�U^$h1�Gq4)���2��1I:�!��7F�ƫX8U�"�-Q��z�m≰�����_)猻;��k�TJ����������Q|��^���M_��}�K�o\V\]�$s�`�z��>���d��
b)
��@Lo��f��O,�F�����!V��a7�/y[=g�IQ�y=�>��R�x��IֻN��#Dm�X��(.:tѪ%���7�$���XM�W�1n̂��@�?1��lC�Xǀ�[�2�+'����u��	H&���DH�?IGwG��ŴW�q�k��������I%����'��-Z�>���dՖ��N%ٔ�U��1}�6D��Ќ�5�W��U�Țc1�dl$�0<��9�Q��W�V�~݄�����L�o$j��ppO�N�?��8��҇�9�I��C��#���F�TM�Xt�z̿��=�� lKy.O�k�&C�J�<Ť�3��.�b�?�fo�K�B.�X�r�5i4@}`O���C���)���7�֢��M����ĵ���\CV�g�(�3AU��X�R^����D�阽���,E˾���S�Һb2k��ux�8�h���W�D�"P�9�43 CUOy �k�Lݷ<�ƷBA2<|����YO���VD��+#�-wf�T��==s���ٴW��Ty�[�^	*�3�E3$#�gE.M�9����D�)�llk�%!�����xeQ��E֥�s��e�Y~!Cl���6��˛%�&�/
�
����+<!k��J����\C*TI(*	�1#��S��s~?���י�&	UOR���:��"f�b=�>�\�:O�_a��G��O+���U;Ey�y&zD����n ���$��Z��K#�?U��E4n��"���_{?G4�$;��/gƛBV�����{.YR� �ښod�����7͟?��M�Ԓdf��+��H�Q���׾6\t�E�$D��r~��sP <�LEbp���z��$�'��T����b"���7��h9u@Sӟ��!�g�#��8F���Y��9%�E�,�&�4�t}�U�:MT��<:mp�����\�׽�u6>�؅n^���ã�?6�8i�։<o�5����ق�n�=������O��{�d�ƍ��w�&�T���D�&%���Lpoa1�9a���Ț���@�(!rI��	���g��_�z����R)ԉTVń�Be`�9,y.$79~�!�bƱ�:Y!���3Q�L�+��W��ն/q�����h� ����7j���˾�e�m�ehK#Q"]p�Y�O~��+��v�+���-��Z�7^�C�"k˶��1`���y�ؼ����b��C��v)U�i17�p���k� CNm�JHM,A'�'�^��c�'�������
˱ `q�|W��^��(�a����J"��K/5���������}�5�� ��7����>6�����!�EcY9�ٳf�{��'�-Ӟ�����O��v�i���\��5ض�'f[FD�F5�'!t��=R�R������ʿ��  �IDATK|<_}x��Ǫ�E����C$F[BO�ࡒ%EZc�&�΢0�^Z�|�J�m�d	��ZQ��9��0|��9F��.��2k���9v ���+̪�C߄�[{N�.�gK�-���u�p��ϸ�W}��o���GN?���]u��/]�p��(+� �k˶��v�!t���A��4)N�EL��_Oi��P%�s�,F*�����{,dB�����o�=��_,�B�������*����.�U���eL	j) <�n\S��e�b�E��G޺�0��x[K���CG<�w���������W+N:��xa�V����.�BJ8*$E]J�����x$�^���#Z8>
�(tCD1�r����%�&%E̽M%��P�6���
�����VHj,%:Q��J|q�GSi��?���jKt���el�H7�`�{/[��?��?�g����~��߽�_?;��T�����˷'[�dbЩ��j�	��LLe�'��)&�z�h�Dr��5�����)�9L�xxa���'^W��ؿ�f��F�Χ�5�����ب�=��S�s�i��q�����ZX5�5DiKs��F�E���U�|�W�n�(�s^�������>��p��܍��L�3�҇z���r���1�})
D� ̻�cҲ�FB#F���g�T�����"��p���#<�J�[����2�$�
u���CY�r�J�������dm�߱@;}���>8g!l��6������p.)�^�~_�s@	�j����}{�"�Aq�~#�c��)�(rA0��]�a}8��s�Yg��~[.��,�_����}g	ܡ�P��W�@��ZĔ+R�]�FW�.uƶƱ�PZ���:-ORM��S�ҟ�\������ ����贿��~�zvϬ[�;�[�v�(���E�\x�_������y!����3n���������Y)�XNr�Q�ziԓC���'V>�+ioU�m�(�,w~���z֞��K!�G0V�/v��C\K���?��k���J��x�a��^���:�!X���ndyRؾ�I!�祰�/L���J��gG������Gы�Mֺ�N�C��Їrg%�=lјѽd~�}������^DcQ�V
�=�P�M��>����<~�,�>G��Fk�#�2e�{ Bu��2��5����.�����6� 9�S���{^o�y�Oc��^��d��j5�h��"��ui��a`���:�+�f��"~�_�x /�1���+W�H1�>Q�)7�S�� �}ݚ����Ś���G�Ņ�,��x��\��r�0-
Z@����/�rjF�_�=�_�I��2�����A�؁x-z_:N]#]��H����s?���=#&"h,�џA���C��gh|	��חmiAW1"�)�HV�Կރ��G��M7ݔ�85o���}��;�h�^1��8���/~�w>��4�݌R�тz��o~�7�x�aq@h�0=��Y1�~D�O�q���R��)��&�,:Y>�z�]�c*���v�R�2(�B2J&2�e]�-��yJB��Q�C�аV=V˵�-�~~�P���Y�=�s`�{�+^a�y0�:�΅B4�g�������0��̈́��,jfy��q�������*�H�PD4��Aޙ@��}���c�,7VaZh�D�x�Ɍ�Y���&|}�T塘�5���C��3�<���og��G.���?��ˢ����'Ƈo�T�鞙����Wq�vu��1֎�&U��\<�rɬ�v��L�<=l��ΏG��~���&�b�b5�����6����{�"�_�I�&��5���-=����
���h��G<��o�鷃�Z������J$��B4�Z0u���4v���Tϓ.BZ=��b�ڎ?�/�k�,�d���l�"_F�����4ߢ�A{�0٩*Zp�O�Hظ�{|����[��S�q���?�㣟�������%Qyv�϶�?O� �#7��S��DO���\T�|�Ᏺ��p��h��Q���G��w�����xp��U�+�h�vw��C��Z-�,�Ks�RZ�aÆ���^��D��v*�k%���TW0^��r�|}��DI���¥~(~y���=%c=ݶ����B.�7n���v�/Nd%�Y���Z.��̍����0v ��xF_��+dO��Yq�Iy�B4iq��i�>�����@Ź,c�'�=/�S]��ո@��q���.�<��ȌS���_���~������V�`�EG�B��ʯ��OZjB�
�sd��z���'�����)��p���|�q�-#):�����̙��W��e�~����c��c)'=IG)�UX����k�w*)���&�Ox*<!�89!!W`�$�O')�<�W�zo�����!�c�9��9�~�Y�
�(ɫs�sy ���/��/_~�G?��w�m���<^��ZT��4 ���X��.��ҷ$õ?�;{�"����:�dF�g-zr�XK}�L�^cYqx�'�����1���Nr�_����h�X1�1�O,�����/|w��[��T���_�����߿��7\s��M�o�T��RXr�YU��M$}֊����2�a�714�O<?�(������q=��������o�г���Uc���]PH�k��{�`m�+$,W�IAR�bŊ�ɷ��,h%=�7�=ďC�p������V�C笐�^�|��7��y�I'���&��骫�z�%�\�!n�q���1d^h�����},_�(�䓻S�D����g��[^��x����/�QP`-�B�y0����P�ђ|���{sl�og��G����7��w�m��6�n:;��]
�zqmo����+�O) ?�䎓��i�mb,��b�԰�jõQ
�Oબ�q��5�dg�GY�x�_�����G�R��0~/#������>��Ǉzd�J���RH�ڄ��zƆ���?��?�Qu�x��Op���;��7\{������x^�c���șI�
e�=���O����ւVTƾ���-��Iw�������]-J��9}�y{���j���6Z��L�D�B���*����y�����[�����~�����-oy�O��M��^T��R����
�Qp�V���sl�뮻.�p��H{����I��W��"���o�#��څ�כ����x�O4���81���>�+���L��^#����Tq��vi��9�3�_y啗���kg<����4+U��\A�+��зU<�����pǈ�{�ޒ�I�W3Δ��h�f�;�!��� FyGq����֊�W\������n˾g��G�K�ȥ��M���OƋ��Ύ��!�Rф:T���PK�\&Kd�kr0@�!x���p�
	��Ysf��j��;n��N�O�&Չ�+tuu�[�[���w�p�	<�y��{��8P�[a�}��YR��r���a���	����7��E[s,�{���/������*q��׻��X�2�a�l�h;��*�v����z��oG����9.���줮'��kL����d��'-��������u�kf �)m�ɛ_��W\q�;���/���G~�O��d~��#'d)7��<���x|AS�2�
u�}&.5��"��Xg���)/�XY'��/���:�c�)~N��؞����}r\q�f��tW�^+�-Z��YO|wQj�$�?��u�\s�����q^����W�σ�+���(K��m(�������#$R����d��z��>
�f������M�q�^�]y�Ag���l+'�w�����y�{����\saT!�tw/����Cx�f�{{����ng�q�s�����y��Y�U1�r#�6�Y4;�fʩ�ҁ%�v�����+_�J�c���8;�.��{�0fY��9�����<�Fֲ���!ت��n�������:{������+�,����#������^�|���H!-e$��x�\&���*e�|R�I����h�<�`���8a�G��w����}n��n+�:��������ݯy�k�sϽ��q(ύ7�8��;Z�'���|��P��^\����M����m�������ۗ/����u�Y���ٽ��.�&�&s��=��me��]<��O?�l�n���mrmN?��M�������O��O�|����&"i�p���P:R���h㦈������1�&������=��1������ӎ���ۿ���+���}�����?+ޭ�{�����7���#������{��7g�x�:';��	�T��	���|�é%�QU�B�H�5I��3�C#�+_��׿+Z�+C��z��Z�kD����+��s)�����a!FY�8�c��ړa,�����>���;����x��ZI��"���7�a��o=����-�&W4�8&<�x�6Ɨ���g�]��O������{����	�w[�� o{���>���~��{�%��y�Q����dxy\v���0]���WI$CV~R*���L.8����YSa��JI�aҷysR��`F��,,g�rV
S.�=���R*ل��;R�YRuk�4�`pB��RP��;E%b�����y�m���@���x�?�;g�G�F�#��wߓO<��/�.]J�w��Y�f͉(�6'������q(��bի�#Wz���z��Fp�Xyka��%�F����x��h�sSk���^o�F�go����9ȧz�Wuu^�ˮq��R�G�X;���@�}��J�8G������m'ʽUʕ�;*b���Qf����8�x惵�����rg�(���R�RI�zŗꎇ�}����'�\J[ܛ�{T����j_<��{�������C:�8����7��(m�������W]uUwTB��гf͚Yq0΍�DԡS8�y\��%j%dcJ�n��f+��w������7�3N�2Ǥ��5Ǥ��/����&�4��1��uR��'������~v,���qL|���K�������x�~W�Egէ>���ƒ�x≏���?�hT������R��n^�#�e�m��3>*<w�7�d��g�W��H���Low<^����.���,����w	r]�d�Prz�K��^Jo���&��4����@��@�����uB3�;�Z�T��{���;z�I��ܶ�1�W�XfPƱ�~�u����gOs�1�V.��~z�;����y��ٳg/�ے���.u-;^�A5~n��{:���������k6��㸩e�|>_�h��yvM�l��`���K�=*�����54��M�D�%��&��9r<�cw .��K�,�׭wٲek�9���7�%m�?9�l˶�
m��r�i�Q�{O�d�&�(o*������k��Z�%�z׻n�nm٩����ҖqH�M�J�������[�Җ��@i+����-m���V�miK[�2����Җ��eJ[���-mi����oK[�Җ(m�ߖ���-3P�ʿ-miK[f����^��2�R    IEND�B`�PK   ��OX�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   ��OXʪ��;  6  /   images/d8ecb972-58b1-42b9-bd6b-2e1505532ecc.png6��PNG

   IHDR   d   �   5��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��pW�	!$�RB���4���H��dG���P���m*�V�tZA������c�H�D�8�V�TfJ�"��B�_����ޣ����{o��ݻ���Nr{{����������Q�5j]�p!����g�g�}={�J�H�Pv)��]�|M����~�}�}�}��&� ��ىToz��)
S��ȑ#/�/� ��5�O�'��ag(_�t{�Z�y��i�?�{�;ٻ؇(	���sɀx��G8���3ط�od���@$�']�~����+{3{#{7��B��u i@\Ǿ�=��A
W%�%�Mv3{-{�_b'�=�&k@Ҁ��~�}��uSҀ��]On��(�`�$�	�`�F�:�$̳�?�'��%P )@�W��~����@��Y��o���و��������4{��٘O.�%��AFK @$W�W��Snj4�g������7	 �fWP�����V�o`CP|�`|��I!叐E�Ʈc��~��`���姐x��(�yl�����Rh7�~AO��6�Ք��!ȕ��&P��H0j�m3�zk5����.�6��ʯ\U���-�8�]���@��X�KV��rG��@'JL"�N��d՟�`�Dn:_YJ@<с�����ı�	�%�r7��S+5�An�{��t�<FV�z��⩮0��I������'U�-�AⰘ�t�3'�z��u�L!+SM���`��Cde�I�;����+��TDc��ߎ�@�謌�Luy���8���[�� R<��RZ�,�@V~��\��cF���H$��X���O�6�ZeY >� ���/�L8n������$�*K@��.����Q:~J�^%VfU)Y�L8v �z��sY޶�J]��tNh���':�gEh̵��"�[�/���'��"%�ҍ�"$���V,��F�[u�N֮�.��A�a���Y`�ý��0LOV�� ����IV�I�;L���ĉ��J
�dذaN�a*ߗ�Y��7;zV��Ȫ�,�����,�����,�����B2t�P***R�`���Ң��2d4H�}Z[[�ܹs�B2o�<���t�*B:����8��>�f͢��j��+`8�֬YC;w*_��B�����L��e�uM�����尪�%��'�W��\*U��U/b�F��
;d�����b�d�@� ho�M�F'N�ո�>y�$mݺ�rA��ƶ���O�n*��HJUe!rr�*��|�1�<�D���s��Ç�y2��b{ 8�cƌ��K��|��85��a\�D%䍆8^��@�T������ �"$b�4Щ�E��S.(6@�po۶��?�kF+����iʔܸ�]l� 2v��E����S�Nu�O�|�wl�@���mϕ��
H>���r�X&�m��� �N�>�g;@<8V	Ɯ r��є�E�M�Ν�\��8%'� ���ё�]K�@2� f]�7Y Sh@0�F�GeE��֚T?��ŊvUa_�U�A)4 [�l�ݻw+��		�����8r���:t��Rh@���.���ݻ�q\�
$��hK��I7�J$G���[^z�~MJ���_�@�+3n*֦����O�����D�e�U�Qȿ�1~=���
u�����]+}�R�Q�M���de�ߪ�d�?��b����*#���u�����$�5�<��~�۹uk6~-�9��d$LU�t^�����=��T�<�-$EU���SmAO�g���U&e/�?�f�9sF�E&#o�B��^IV��5r�oZR"E��ٵ�;�&��������Jc.�!^(���s;::v�_�HX&B|,�())Y(]������ﰺ��g�0F�=���UUUO2$�r��kپ}����v$�2M�u��������sw�cǎ5�ٳ��Lӆ=#F�(���~���Pyz����mǎ�[[[[������k�ٳg�0j"m "J���p]�~���q�&M�D+V��j߾}5�mݴiӲq��ubf/��O�N3g�� '�|^>0�oذ��7oN�τ	��������q�NV[cc�����Ç;��x �nt@F"�8qoB�9s�Psss�Aq�t����-J����˝�E���g��ŵ���	H]]q�����೗͟?��'&�	�['֟��F�d�DL� U
�g���8�\!��f݋x
��}��o �耞���z�N<�(�D���}�A1����o�+���9�4_7���~�B1"�@
�4�u�WddYX��9�a�E�k��~��`��^G�p�@�"��7x���_�o'w����A���B�MH�cF�d@(����_��`��
���w��&P���p	��U�o�p;۹�}D�h��o4|=� ���F�sܐJY�d�RJ@�*
�|�R��/^La	gq�;�a����←�ȋa�۹$B5Z�"���?&7:���-=��}/�큩����*���P����L�|��?�x�ׯ<Q�g�z�
��~�=���l�/��%-	����M�_X#|)�uIo�`o"��g|����SrD�	J�7�`L$w=�5�_Xz�^L�������u��ȭZ�
��½��+�P� �`Ԑ�[b�"�)��F�!J0�$(��m�@�8��h�w�RA�D�����d6r��� �ubCaIP�����P���vd����E �*
F;����bC�aIP�c���	e��W�r�&��q���R$6xt�mF0����!6���m	�]�`�Y4z^h
>�v.-P�6^!��=�M����CH���VrS,�}���dy��ERt �a�/D�lJ҇�CH��<է�����B9(s*�{x#�,�ɿ^fב��8���������Z�E#ł��ic��wɿ����wC.����=Ay�{|�BqAT� �${T ����!	
�~t��|�G���� t%� :$��!	
�(u�v��Q��U �	�+|��˯z7�2!	
�+��K�˰H��n�>>�G�����11�;�G��@&���%?���o��`a/RD���o��!�ko{?X�J��)`̃�2(�@L���3���@�.	��)5���N�<�� V�<P�����@����>��O{ȝ��� �I�FG
y��� ) {���^�1Y �1���B\Ez�Y�U`ڨ�w/n}�P|t��~xI�B�    IEND�B`�PK   ��OX:����  �     jsons/user_defined.json�XkO9�+�|XQ	G~�ͷm`YTJ��E+�Pe{<0R2�Σ�B��z� UZ>���k��s<�1i�/mr�t���d6/J�%��7[7EU�p��=i:�m����?�Ԣ�{6�<"b4��r#�j�]Uw#�\���&��qRdn|Nd�d* D�J2�
0m��PI�Z,�Җ��6|��s來;��٩mL],�uڻ���q�e��i��P�4�@X�S.�����坛W��\O�T��m
�Rb@��@g8&Sy��Ia�Iug/+��5���;�b�����(/ʼJN��[��r��O�����1�q7l��s�п�x�!�tb��]Y|�ܪʋl�օCw1�US���y�#6�Hb~L�;A�H�P4�澪����͕����)L���ǡ��?W�f yH�E�#��! ���a(>��?���`!�4v�#��"6>��OC�e�	s/� ��zd�"���Ŗ�9~��T �V �"�(V.ίN�A�@т�������b%��U9�bI}��E���������"�m��PEɍ���7��;�ڻ����|�/ ����h�!�!�w �����	I���hX���;�hz�5آ!�w �&�wi<$� �D��D��?!D�(�_p���&��>MBd��P�/Ubs��)����v)��h='�j%!BG����"t�{Φ~�����,�������JuH��������'����P�����=�����b�w��S�o=L��^wm뾹��k���^�`���B�,�$"����/|dS@`����ZJ�Dv����Er"\(5Њj`�1<�HQ�o�V S�<�	 c��j&�ƐC�-ÝJ���G#2:��������8���s@�^]�4:*J?��z�Z�$���M�f��;�u5/�}S�nU��3N��A�G���+�~�)����S9���l�J�)�B����~�V9����*�\���m�S�?>�&�>\�2������UY&4���JɁLmXJ-T�+��6�f 
7݆Zqyvz2�~�F�q��ֺ��|ݪԩ%�`S@'FHҜK3��V�P�O]��=��8��K�lX��rr�g��DB��� 4����^Es<i_��m�y� B�X�W�­���lP%�P<��n�?�,T�*���C(O
+C��FX7�]T�T_�o$�ߗ��0���}_W*sl��\f�[�M�:5@I�sPB�)ks�~#W��W��Z�MѴU=::{?y��g�U�9<�y��ր�\f�9rD#Pf["�,�ux��$"����;�J�PZ�Ż�3�-TEt,�2Ȏ� �KE��vQ��+�_e��I	�"��� o2/��U�|8�P��R��M�T�5��|���蹐Q
�tc�H��F�&4k	tƝZ� c[c�L�ۧPK   ��OXϚ�  T�             ��    cirkitFile.jsonPK   ��OX��8��9 z /           ���  images/11b938df-2630-4b82-9eb5-abaaeee165cf.pngPK   ��OX��g  n  /           ���E images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.pngPK   ��OXhT���� ċ /           ���^ images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.pngPK   ��OX�1.:�  )  /           ��[ images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK   ��OXǐ]zd� K� /           ��z* images/972a987d-5ae9-491b-9c1c-35ff468aee03.pngPK   ��OX@��)  /           ��+� images/b4aefdef-6992-46c6-bd27-cdaf728c7c35.pngPK   ��OX�GDU7� �� /           ����
 images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK   ��OXʪ��;  6  /           ��%� images/d8ecb972-58b1-42b9-bd6b-2e1505532ecc.pngPK   ��OX:����  �             ���� jsons/user_defined.jsonPK    
 
 j  ��   