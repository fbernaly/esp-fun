PK   (}OX����  Ӑ     cirkitFile.json�]]oۼ�+�^`W��/�T.�mX�v���H���F�cg���]��>R��c�>��n�Ek��9��~���櫝��imG_m=����&�����7��[2���ɨ������!������'��ǧ��N�Q��L�I�E�c!r�6%q��3�s��DW�����SW��0��BZE�<!6Df�����J��*�erDI�P�p�s����\���q�J���<�)�cN�R"�P���х�f\sa43��>��4��a4��Q�N0#Q�b\��IF)Y\�����t��Rę�2g<c��ޞqո���T���h�>��4Bs@���m�;n��\�W\�+\q�+��S三	K���2������~~�=�1��^ 1ĨF�o�����?��|:����A�i�P� �D
�R
AHYvK�r���@���BuQ�)�_����<9�M�T	��"� ���.�M�B52�W
���o#(_ۏ(����Pu��@:@�a� �U )*�DJD
=ܑ�dfl ��� ���C�	�7��T��ސ�Yc�%;oj3F�	�D
?$L&�R�L&�R��E���&x)�L&�R��r/`2��r/`2��"�HQA�� R�0��0�a�K����0�`��9������b]bTߣ+��oUmg����m1rdcZ���n;WqRci�U���BSg��p#�2w�w���b���Z��:�h,�Dĩ`$N��Y*DZ��_8�T��i�~|��F՚�D5�8����S���@6��5�s�>�@�P��Tcv��ӭ9���s\�F5E�F�,E�ўy;,�Tc`�<z��ҽ(��ս(C�[@�ѧ:.[Fb�ĸ0�Z���i%a9-�P��P@�{��Wg/��ɽ}j�#��w�Q��I� Sp~��^L5r��E�)������,|�28+i޵�'+Pgnq�pP'�ZC��[=�Ax/Ʃ��[
���M�/	�����P��Q3Lc_n�����4ձ�����|m�_m12��k���y���{��@'I{8��}kBx�Е�iA�D���	( `71�H��e��,[��P��v�c�g���k�9�;�`w=�`7?�`�@�`�B�A�#�� �1�7 �?�� �Mr"z �h��Y�k�[p�m<��7{Pp���e���B� �a� �OUh�/_�C�	�*�m۳LT/��/3o� x���� @y�d�F����
��A�,���	2v�e�ɦ��-�~<�G��}f	{�d�u�����Н��-�@�%�h�}�R��;E(�Fz�4gP��۷�n?�������0̥A,��K&�L
xO̅����@��k��~��P�?D�=Ⱦ�r�f �	O�|8>Sq���%�"�e���`��Xh��(���g��Igs~x����</<6흢�c�9N�b}f�r�"<C�̕ �g["�By ����	g��S��\���y5Y�I�~���a��ͫ{]�5t\E��BC��w����K�`��^�Bfa���Y+�g�B�|����M	�)�W��Ѳ�	J�u�h0��ס�����σoDÔO��%��B����)�<}E__{����P숌��M;B#�6cL���D��U�鉓8��2z��=p|c{���C�݂��3��=B���� jܯq�H�ë?��w�کy{������U;[m�o�����/��/|6��w�hqM�N�B�r ���!R�����ݮ�{+�����N�2��5}�T��F�1�� �oaw	�5B������W��榛@��k.�&�c�vU�7ۼ�]��Il7�/��nR�LJv��2I�&�e��M��$�.3��ښ"��y�����Ѹ�5� ܟ�v�쏦�#я���z�d릲����4��y�;����&_�=��}� �j�s����c��}>����}�=L�}��s���Ҍg�%�l���U�خ����Um�誩��U��L�ɛym�}&<϶��m=5��N S���Yմ/w��L�LU�j
1TY��_q�\o�{'!*3e9�܁31q�y�:��*nEAh���֍�y�r�A�Hc&�B��i]9)fam4�:�e#�r�����z?��"��m�V�M3/��ڐ���#�۾Id2$)�z I2�Z'J$[�H�XNc�9q�Ӑ8�Y�<��4*3Yr�[�tF]}yhv�����z,>K"�i�|tua|��G�=�ųG���Y+�H��P��yovI"��j����nU%��E\abA�$N��3[dF���1�`L�֏���N]��ee�s�p�p��ɉN�J&�h�ޑ��+�kn���[�˙˕Z�JR��4U)�ʥ���׹�3EH�����C�z!� a���J�;��X���⹎u�HӡHE��P_��t��`T�l��\��TmecC�%�|� �:��+��tK8&�~ZnL�)q�$\뵬�jw�d�j������m�����WX��I�Γ�;y���&��Q��U����o�Hn>$$fo>�������oޭ���c��"��P�p��ؖ�����-�n ��1s�]̱*�če�-�4�����e�)��&=��L�Am����Ɓ��b��!y�4�O�:���GF��vyhlK�|��!�.2D�"��y����(��l;޸�Z��L۲�_�}K�_�0��-ޮY�um���ϕ��ً��?�������n�"��hp��d�溚�/ڤ��˭4;)�ʂM�[Q��v�6'�O��{�V���4��www��ɟ�k�p��љ�������Gہ�g�r98)�W�Z�mr)�W�\B��\��ˇ�\-�ٗ���]���Y�*�E�
�.
ؖ�nLzL.	�,��@[���a�P��^_4'�lΗ���������5݋��0�4�!�ѷs�EHO_�&0dO�{:��i؞Ώj��с��$�e3�|��N;ruCc�Ր�c�AܴPL�(`l�֌�-�=�K�N�ۮ½:W���,���!������	KTٱ��j�nB(���Wq;s�}�zxF���<#0�ӌ��8�e��+�����|1���#�8*��98�����G����ǥ�m�h�q�ek�z��h�ab���r�ij������Fql�o6F�{#���l�KjȊ0W���[�\����j<�T~4��+3�EWy�����->��܌�N�7�q�s�3��PK   (}OX��g  n  /   images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.png�xUP�u��{�;�)�AZ����C�I)�-����8��P��+�{���tw��Μ93�pfv�,B��*�  ԠJ��&��q��un���j�	 0�����z�Hj/�w^z��^�V6 ___>GOk+7>W��S) ��AMI^�/�$���Ġu����������1�6�b���w ����(:��9�A�B`hz/�抉���T�K����%U�0�2!54����+|������#�lI�)���ŶE��V�c����m+�h�@.�����9UF�*o�@��Qt&��t�t�DA:2�L��K�H�e0�j8"0��h�����A�a��/�b�V�D�o��휞�H���l	}� }L�~���>��t����|f?�Y�����0)�){��`��o5����1�䩩��-��&�{�6�P��54v�J*c�?Ν/�yޣ���;_�����WF��� �z����ܻ���1)�?�n��9[��j��U�Ҫ|[;9�K:�D"�m�R����7 쟟[�ެ�68��<Sic�"�lM��ljn6b:m�&L��}�pj�������\����ֶJ�U5�tޢL���n�l�)�ox;nx�TY �J��y�I�@��y?E�ʯ���zZ�Ҍ�w�;��T)�?'Q�63�������W��:�@��e���4�R�I`��V��ʿ׋[��^��FS��'kc��������k����$C��7HY�T���H�"n���v+k)6���2�& �gg���;�>=�y������SAJP��f,����ׯZ�:஀[�?�q���Ǚ�UGtY
~s��^�F)O�\��Ý.�`{��3��b�$�[��H�:/7(���D��Y4�zV����;�r�w�Jtw��t��iYuI��>~ɺ��%�^4%����o}�͊��!b���k����PP�N�˺���y^�i���	?	�<��횇
���<疗9ϺN�s���Y�S�nF��r4J[���松>���]!faU����3�:ːG�q_�
���?�君���g��fٮ��v*�	���P�������)��Wic1�&��
�*�QB�#}�,���Jt��Ut6�c�Y�RY����m7�dgF����w�9f`z~���������4�)�n2~��m������遡`W���g'�x���!���+�y��Dx���/ǚ솎q��0�ط��S�<�+�/@� J��,jnn6�FB�YW�1�z���0i��,[����zUiQ;�D���ϽL���HN[��|o�����\m���UU����@�Q�������g�3Y@�/���Xޏ�w;�s�n�%߷�WtMfI�0�c�IUr�{��K�����a�u:S�a�n|�IY��ARĈՈ�:� ����;4�JMP�64���g �6\]a~��u��E��5M�e)����N;�Y���@̬�{V��ɫd}<,�� rp��!wL]ה��V��`�|��L&�E��LJSKy� ��V�;/�w#����(�.��o�L*��P�,���L��f���n*��/f����k�M��C�I��V�{��f�9��e��x�Wڜ{A���S�z�}������:L��3�DR���5s���l��x9�o!�b��9�!��9�����ӖJ#v�2w48SݷwӤ�Y��VL�kR��NX�I��w�L��/�����}��ͧ���^��hx��x��|Ԗ�+�鳵�	��H|:Cu��*Z��j?|8c�{�|N�1)���.LCCSu����L���(���(]�:��@-�/!�7�?�X��M�-�p�.Jjߺ$�s/ls͂��Eg��L�8�:�?���{t	)�|��V�~ܟ�����n��Lu	�gAOB�����Դ��>
�g���xԂ屙�WȖ ��#�!��{�8ğ]�7�F�G}^���8�xڎV+/��f�}�X��}�,�<cj{h,j���~f��gi��Z�陟�`�c@�3��8���`̂܇�7�7+R)wQ6����"z���:�*��F��7�|l���nI�o;u	%�_�ۛ�?>܃�Ѩ&~�	 ��:#K��6
n�F���4epftg��(���Қe��M�o�#�a��%�:$�O(���SH\'dn��DN�O�)�Y��"<����?c�Ǫ���	Y��;���ª;�lH(�)x[t"�"G��<��㬖�r®�k0�&�`��C.�"0��<e���a��@�^�c��",N<�s�9q x���f�\WOL�F����j�&l�f� �����0����=�����	�@L�6Y�Ed��Cy]���N��5?'?_���Y�q|N!u�ʜ�s��u�N`}���$~��g��^�z�qr	J^b�e�T���ouVT6 R �zynZ�e���ۅ(�0���ȗ�<Y�/�hm�K6`ϓ'�L4a4��{�щO����������"�M��8�;>������m+2/�O������2xS_:x���S���P��A$�޳�l�ϞY�(���5��l���M�'ק*������w�}�����Zq(㪯��ϣ�,�݄1��-����E�w�>�k�O��$ܗC�@x�j�]��O��'N�TY���"\���Q��K�iJ�y��1��欎|��q��b�ӽ�#W��T�Q��ݪ�6�E�#g}v�\|)&�Π��!��S�y���k��i�$��f�*����˫"T]P2 Ȧ��$-t8�j�QG �7��XV��#�{��L�v�&g|�|�;I�Q+>T�f�b�+��s.�	�]t�ۃ�cm]N�û8��z���׈0=XX���8l����=�]��x9��^$9�m��r��/���Ɗ(Nwn��X���Ea��z/�ejǫy&�G�A�1��u^�U���e�Rv��	A���L$��t���k󴊧b`�x�`�`m�c�[m|�q����%�`���tl&i��{CwC�W���v��3zB��/�0
�}���j�FχY�e��QeUNh/�e�违:����y��',�[`�Є���l�#�w�-ܳ�ע�yRx�DE�����.B��l<զ�	�b(Ι�O���5i�K��Վ���R�'C�2��Ut��v���R-�U���H��Sh��W�\h�a3Kf"!N�PyMlOB��	��ɦ��T~��p����&��.��`�|S�����YP�H9B��7���'67���!�2RT��l�K>P�����F۞)/���� y�I���I� ݺ�
혷7������v���4��YH��V~8�(�y�E�l#� ߄ϲ�̲�'7@�eV�M �:P�����D���U9&��*(h���p��`�V������Z��ڎ@����Wu���T�xhT� � �ɣ����w|��n�X����7��`���PI�l�� ���}�wd��.�Dj�z�P�1�sB���E�!w���Q�(�����z�Y���H��-S+����D�Gb1N;h	���4A���	��73o��Z/	[)*�PV�"6ӱ1S�$RϠV�+��_��A�>��2;DU�l��
r'F����m��;d�7V�+�YW�H����4��5K�/���z:©��/ؐ�O��n�w���f�eD��<}�?�Ҽ��_)��dz����"��Y(v�+cZ%,�`�UH��(4���ٯ�P�e�+�靑A*&�4Xf�%�#��#�(�C Tq�j�YSu*r.������K�<>5W179>G��gf^~�Xݹ��������.+Ը�.��� �	Y&Ic0mu�]��;LlV���ֆ]2a.�|�K�FE[o=�a4�X85�=�%�P����V/AK�Ndb$���
���(2�R��t�b������ޜ��R�~�kbs�ۦ�]�{��&S��Rk\B\c��#��o��x��cK�\ۖ�1̥܊ou��p�rZȠ�xu	焝��9ȟާ�F��|nG|Wo�bhp�Y��`��sb+����IK�h�=�6{Ǚ:_���������ߍ����B�"@sMGK:�`P�Q��Ls��A,p|��{'�ڤW�/D?EWp�c��؊�o9M��
��M�'�c�{y�z��e�#�F�l<�B��]O��%۰O%��<r�e5C�f_��!>�ν���g��_��/gL��f�#�EgN()-#\$�\�Y���DB>'d�f��d?���@4�7h�
ǉ9���x�5�������:V19q���WxQ $���%��56��	�2��ea$�E����Ғ	�tlRh��`	d-f�Ԓu���:&�h�S�3��я.˨��v�ٜ���j$cT��	�$7~U4��Βy���&��=���Y��!1b({�o��rz3Pǌ�:֦�<G4�R<E�e�̼螪oJ�e�=��{�ތG���#��Mx}I�����G���1[g���X��p��ѥ,ߋu�e�&N��<.Y�WNH�k�|c?��M�
�t>�,�s|�2#b��-j)�������o?�ǘ�}�U�ˉ�V.f^��q�`x�9��K�!m'�������7�-�QMs�E�`λ�_Nz3
?�;�e�͊��~�]T$r�Ɗ/U��
}B^���c�k���~���7�jF�.l�g��^pr�3��+q#��)������{�{�H��C���c�L鈈�B��\�c���ġ��q���jh���@d^�Ѯii{���;p��e}w9��l�����YT�'_!ߚ;���¥HfH�+�2k�5�ASF�j�ʙ·P:{���s��	��d	��pT��!i����x~p󂭡�RS�R\o�"V�XLq/	@�U`,0�������""����*܍u�P�xC�|A7K�e#,�b�m��:��*�8�NB�������X��[���J汁w?���h��09qװ��~�g�(�5�׭�F�J���_�J���b��5Ƹr����z:P^��kϹI��\��7��������%��|�SB�/�[Q��"��ƚrK��T��(�R��T#����-K3uwUi�4_I®g����x��t�S$/�������v�"'V��c���)ʮl�R�Fp�I�xrQ'f$��[������X�%Z)	��t7^�RƄ��g��:_�ޘ�K��������.���*�|�!���K��s�?��Rl9g����fr��F���f��J�CrVZ��_�S���!�Q�̛��D'~�A����W�E�pP!.QC~:�/�y��$�c��3��4��֋��ULM��W0Q�v#�C/�B�9��q�=�݄	 S���E���}�AX��a��*� WMa��ə�qOu���EDO��k�ء��NF"|V1r�>�R�ʨ+1�T��@	'��x-x��ˏ�g�ea�{&z��6=O5���p1c���X+���cQ9bǆ�����dj���[���d-*b|Hvցޫ��i�zeG	{i�*.�P�a*`��!���]}߷NM:V�hR��~�
�v$|�RP����(����'�c{!��8�[z��!p`�����B��۟�֚�-T7!��0 ���A�Ԑ��@�$�9	��#��AV��ZO�TL�����N���V��@�2�x�M`�w����@T�'��B|�T��)��J��o��))��9)ӢD��s�a�!8t��le�%?'B��p���?�F씿��������_6_=UbkN��Mj��Y�d�_|�{1D99k6��Z8AM��ƪ�����rF�Aq�� MWZ��m'FM����;-��<|��t�mN��a��O߰�O����O�',���;_�h��u���sm��$W�S�HĊ��ԅsv�wث
�� ��2E��4���a��y��ܖ���䒺���x���X�>/�X������w;Q��kG��J�ի�q �6ǰ=��I�u��F$���س]8���3�F�j��)�/!ݲr��Ք��4��l��hgf����c�&�IK��6�!�Q0���x=��]=���,��d� ������0;����=��i�@w����sk).�sOvA�y��W��oh��6#��Mbۍ	Fm�����F�F�2��PK   (}OXhT���� ċ /   images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.png�|y\����Td�D�+!*ZD˴qk�J*E�B(�F��-��"d�V�j�s�!5hE�(��}�]gD��<�>�_�^��m���s��z_��u�3~�5�7od߈�`6��(��`60ƪ���/�싿��8����������7ت�s�`v�F��)�����vCQ�������/a��Z[:�_��$dcoE�a�`x0�
�u��}�R�8��w��`��&���`>�kq���x�i����-�S���q�A�rg1#u�]�u�\��ʖqѽ��D���A��뗬M�N�Wj��S�1N�0�����^a0-ⷥ�^2�;R���@�z����f����n��=S�u��x^����:v�5��+�5����;����w������;����w������< �M����R�̼��CwR_y��ح�|2��t���S���]o�[��}��C&-�Y�5�	Y|�F/	}<W�|i^u��b�ud�MK�e��W1�F�]����F�I�G������&Zꅽ��c������7����Ϳo�}����������lY���и�vKr������?���dfE-���aƪǛX�nd��z��"��&�99����]�ʎ>��4��u�8�O �d�%���	g�}��&U���x]a��{+�;;�٧xՏ������ZB�����A�ca投�B��䠏����d�������l�i
^�QHȤ�����[W����9�9�nj賍q����#I�_��Y�6l���xrR��Ӯݙ���\�/_�Ħ�:�|lB¾���FB�q%%r��~ۄ5�*����i;�)B���q`�~�*���;gF��:+�l<�'�%o�9�I�?�w$�+j)��˫�,ѺU;�_�vRU8������Z̕�~�!rMG bf(��ْen7�����^ &F��}��l���^
�ŚU����M����{���M�yWVRPPP2�9A-�s�[���4<��ʕ[����!ܚ�v�������lb��ˊ������x��e���fii�����C�{����ޘ�׷�u}xv�n��Z�iĔS���߄{ƣ��yL�Q�'L�9���\-q|���M�99G'�~�)��璛����Y6%-y�c0+� 6&C��uO��\v�zK�W��a���[k�L_���g����sRv��Ǒ<St�fF��d[h�J�l߯}Jv�OP^+5+KԺh�J�`{�����ʬh�}{��٤]&��oү[gnjʣ#�w�f(A�N��ŕe��>298##\Q�jtS}���$Q���7�|���	N�f���k�:9===���h<��uA"������o�aDј��\Y�v�
�U]�*�SSSsbb�≔C�An�U���vRڑ��k^�7ݺ�3���k:�H�WllB�ڔ�>8xnۏ?�{W���o߯Q1?\�=\<m�6���˽������^ϫݧf�^�L��@vp�4��p1���5�u%�m�B���뿼��/-�K۽����I1��$�]��WX�֐�J@���Z�;hTp+-�M\կ��r��Ü������~]�!I��0?��f���󱣃;��ACC,��������l��Us}ͳ	Q�J��`�mk�������\gF!�?77��au��[�I���%6��76oN�.?��֢e������b-��3��&'�sJ��{��p��;v�����R!ս����r�#̓㐣sRY!«
Φd����hur�����|r1�;�l���M�Qd:*��D"���rdY6g �&���^C6dQԪ�U0�h�i/�^
��]Anb�.��������?y�ĉ��Ϧ��Q��[��;^��\�Ӟ�,��_;:ǉ�w���>>"!Q�.B�+ڕ엘�H=қ�w6�t�,/X�	�}s����6Zǌw�ڔ/,--=OM�c���-����A���I�'z֐x�;�\&�KܜQ@R�.FL�Fʝ'�͇ۋ����b:R��Mi�;��)��L�� k���;'�MB��m������[@~�	FٽV�S1��Y��,�3���-	�'��j�Gf��ή��Q����RT`	l	�^�4�$i�]e@j/��~^��QQ�)�vLJFFF|I��.y~W�Ǹ��{�e��i�������335�M$J���6:]�,�4YZ�H���¿�n�E��SR���eV����T.f�}v�0�ݺ:C6��G!�Ĵn��p���Q%���uuuN��������/�Mca5�=}��o�G��~+!d7$��#��H��n��F(W��8l�d��G�V�8���.���˺֘�4����ݺZk:������Հ�q!r�,�"0����l����D����|�9MG�A_i���Q3Z�ɄP��������y=���7��[����㲑� ����Ӆ���c����m�/]�v��{�.��hW!H�g������O��:�8C�jr[a�XwM���=Z��;�vG�ef
���h�! F��-�a�� ���d5��0�!�sww�Y��ʺZ�x ��T�|-��KJJ[j/�.��h#��N8��JTfm�y�?��s�OԌ�%x6�Q�jn�'.[�TI�	�]o������ͩ'x/rߏA�-��6O�=�&�z�x��8_p����C;�ߣ��E�/���Us9V�ºH�o'��ЭoM}C��2�
m1Qd�c�b }��~�ª �	��'���-+>�����d#C[�j5)b�ޅ���e���G���V�E����mQ���7l狧v
��g�v?2b/�Ĺ�G&k�l�ׯݔ��dIOv(2!��jf����
�Ľ��h G_J��?��@ �h�Y�?�m��I�^[�{`|]�I1�ʻ��1�N^^Z���|���@E%%Y��j�^}��`q�����J �@��]8���fn�;N�'����������v��ф���1�@pnR"�6���O����z�Z	��<f��8���=�x#/���?~Fޑ�����8���f]�۠����SQ�v
s:��%E�%���tF�.\:���I��/�Ja���;[=r$ܥ��n[���n3ʱj�/�hhnN���Ɯ����oC!*~��A.��LG�[	h子2�����Q�uj1@F�!C�=���|�ܻ�.��5Y��\Z�c%�@o�:<\���	kD�<�/��ikk}'���o�!�v��% !��@)t@L`C���\��L�V~�X<�;�
V-�z�Ȇ[C.�?��4�Q��o4�p���-�Y�	6�cC3�V��M��� E��{ ��P���-¿��=�6�"�M4d-t�L,���jB��R����D�����Y�(	������$yp��+3=�<;�Oe����8�v�����Y��Gk7�!7�m�w��i6��D퀁/@�!��K�[�mpHyP��E�i��B����E�#�Kz'�nr��>���W7�?�]� >�������˓���F�f�LZڃRG��<W�~j���
2���]&�I\��^����E�x�g_L<�O����kF���k�a��?�4�z�y[��&�?��9ui��p�%'����uA;:Zͭ)K��Ϸ��C���X���NX>�P�D�:�bt�����#�~Jv�%�4�S �� �.r��^��B*��S?��!V&�|����(����2�b���kq��%�s����^q���T*?#jjj
t��O,�fVL3)�����F#��#�)�Q �Iѡ;��#a1{a�%b����J�|��q'���>���H	���Z�!R-[)_ʡG�e�����[�kܧ�X �թ-ɺ2�V��`������'e��i���=��c��f(��E(�W��sW=IZ��!x��g3�|��}^X(A϶�q����Uabj�*�(����4P��w������~Ϟ=kpeWt�?2ӭԮ��{��E��Ln�e��uD죭�(����KT�3����^:S)l�99)� �A�-�{��Π��?�í�կ��?~���Η=���CP��_�����"kFA|(��˿����dXN���m@��|j&��ʦt�8v�����r���&�?�OZ���lqn2�"��qf��r��n��v9��r�{F����wC��� F?*s'DN�z���H��_�����2L ��-RE�D ��m�	��8Pg�� �S�-�4�M�_�۾�
�7P�?V�p`rrr����"B�K��e� ��T�eg*#����l)�YR ƾ-h���U��c��xO�����uR	�8�|�KlT*�\�Fi�A,#U��@|"%&n�rυ�j�.�Ifs���qB�6��X��vC��#�X�n޼y��M�
���7W>���[%�l``@͘=fɣ�ň
Z��IW�l=A?v=0�V��?S�ɉ�
J��|TR'y��U4�jSG�JgV��ԹM�ʊ��/_��2����pE���p˳�ޮZ̈���{��1)գ��գR��FR[��r@F>I=�M�_�:ܧ���S���CC�ww��dX��WZ�Q�8�=C$\�� H9R�S�I�^i��U荌����39��s���`�d�Y]L..�����I���M9lkR�d�������(...`��)�CW��m�����{�߽��Χ�H�N�sǧ�N�0�);�:��^��V�WD�c��������!AduP����zR
Q����a���[y�z��sܫ�A�ժ�0(�I5?)�[��b�eA�X�#��G3-
>�����p&�rJ�o����%ub�$,��Uy9�=���c��׍ǚo�R���]�r�ލ��e��Ӎӭ�0^�/�+�,_7s��e���+X���NzN({2www'��5>e%X~4�d�ڵk���C���G�B�t�������r��囵tu#���x:5##��&2�nF�΃$�n�����R�	��;�ϯ�͢_([4�=�)uGT�D�5<��Y��2���=d�|��2�:�}�Qءgx۵�~�̽��h���ԟ��H�K�����⤻IZB�8y���PEP�c4 Y�N�g���i�j88�E]��9�r�I�]��e�Ϊ撩�Y������婎��ojj��ۘ�lIK�Dw�w���9�&T�,��))0��v�z�j�}͡?W!=\$���57�ܺ<�,��z����	���� �����Xj�F�F��_-����h#���'X�s�,�E֋�-��I?�#  (��Ǔ,�q�9^�֔��/$R��4� ��?6>�*=[�8��&hib�Gxx:��O���M�/�zӭU1��ꇧձ���7d����|�� �`0ã���|ڹl3�֌T����sM���#�&Ï�HK�����T�>���Jܺtqj�آ��G^Jj**��[o�z��y໧�؜r�E���x�!�������\*�XGF����u�A����6QS<�#�w�S}[H�/��YlBn̤�^2$S���B��C)��1I�d*�f-"��ɕ*�nn�<d�S;I�G�W��?��C���z׉�2٨Zl1UϏ�y�˖���HJdu��1�~�rJJ������e0}ю�j�s-�v憾��ٚ�0=���iC5�c��s�bލD��"R^Ϻ{�l�a�S�e��ZFFm�yTO~sdnU0�������0/�����}���v]ASs�y+
�<ON�O��n��0�l�}�Νb�Z9B��x�����H�#�g����S2��5�Ɋ��v?r��*��6�5��7�]m�率�(R
���I��^�"��L����##Y$ڝ�mLVOS0^4Wj-��n�M6*8���k$�7�<5Wz�D*[/�q�n�2�87Ox��S�i2�3�"DFFVs��	���N����d�#y�����kը4�H�f抗�j�f������v��z�M�T�aU8�i����2.:j�*�Q�q�}���r�s������Ʈ�m�����3�v���3�]qBT�,���u�������we�_,3��r��ܦ�ӭ�R�Q�sb\�9"���y���Hj0��jL�3�pv&�\��*aݚ`L�%^�M��Ή:�}p!�cl�K?�K��z���s��݊�á����J����P}��{0���ȸ�UR�ŷ�o���p5���T�?xP������s�[ �	2��u�̦zXdm�e]n����S{� x?�Qov!��2�|QؒD��"����A,
�I�cJvuR?@P^�o�娭0?�(.���������Q�˟�7�
O�QM�A�Ņ0���  rST�:�<̿�8����:��CWW�e��ݟ��+�;�N�ZGRx��E!I���f1�����8��Dq"!����[~�U�$lb'�@�G����d�E�����6R������pȆ�|n=]BWH%�T�3�i������c�+_~�B6z�T�Unn��p����!2B���7m"z<�����s����!������{8��B����qo�06����ʹ_3:������'r�Xt���39��������*���,����o8:�؟8~�833��ww+���1oxsO�03��(�K�����'����E�s�.�aY�DJ���0v���q���R�Xk:���E��
����Z�0���>��uuu!O�x���C�^~����CA�]��@0�c�Ν;�&���{<�<D�@�7g�̰�9b�ޠ��q����!��͂����Ό�����h���w�bcy�N=���4�y0h�|�8a/�&�]a�:g�N�g�Йhkk��r�좙�,������i�����A�a|��a�����5�[g~?�OmvCfLsYqA�;s���G>;q�����]߇g��DB"���%���k+t����(]�t�T���Ј��xUp�m�\�E�g�'6������.��/�X==�Wyyʎ�ӟ{ݿ���d;� )���l-f�>+�����7����&1��l����x䞟g'�$2��0*��߆ey./��zz��%:�EǸپ�������,-���{aK�"M<f?��Q>��+IL����\�_SIM��s��21I3&���	�5�k0�]�}��Μ��l�UU	�g����($QV�V���rc�D���e"� ���C~ʒ��9�����)�&9En㘟��>?U	����8�:Ɇ}��Ri��Rdew��.�ˈU��n��e`����R�0_	����x"ɴ?�|��W/�����D���?��������uH�x3�\�qDD�����d ��$��pH�Kٍ^����ۇK歁1I��ޯ�v],K�}��+W|��� ��4���R����"��=��T�/�c��JKw�,u�tR��x�= lX����:�S���qpp@���o���!������C������B��0>u���OK�`����g����CȻo[{l6646Vf��{H��<�����{xc�	gE�K`u�_z�B�i���� �:!�Q����W`�3�ی���K	�pهG��A�K����yB��dŞǸ�?׊CA8��:��y�����If�ux-==0��X?�Ą�}��c�g��j9���K����(���"��Pd �J�7ݺ�-_:ܧ� ����i��J�����1���QA�)��֛}yuUԼ*�yZ��u����I[D���=d<M`�Qu�c[�w�;85�q�d�{���YH:Y�c)���y�� �m��D�:�aT\��U�vr�%%�ggg�}�l�����L[_�˗��)$EԄn�gI3sUm#�]���,�H�H��,]�Ƣv�d�A���	�b<
5��.����a�v_�kQM���H�ud����,�Ůĥk���B�� cCCN4����CYכ��J�Q���eܨA��K����Z�UZ�|�tqq1�(qGN��c!�p��˾��E産C��* ������C��������<OM�X��rnG�M{��--QMM����

(�!���i����Ec���5z�4J~rʹ�͒:|$�{㓔���N�с#xo\z�!�6�
T��9�5���0��7nެ)�+�N�%o����EJ���XOm����]<��QP.��^9���խe��5ݱ%%r�܊�u�����:�RN��'��2p���+KaBa)�%�\�����p봸�=�B�� �����cW�C�Ҝ�e��l�P��"i�o?�������/I�����,��T�<".�X�p�һp���*U'�Դ�ۉ�B���כ�oF��	%]�H`>~���F��k�ޥK���^�I�̴���Q�%e�uأ�*J],��2�����~u��q�Z�_#��X�Yu�Ȣ@R�}��C�/@�qF�:Ec�k�׈|G=I����G�Xl�y�:2:wZ�Y�*�Cð9�PL�٨g���"��|��B�!�Y1��u2vB����lVgz^�?�'X�9HX,:nϏ�Rvo�tyz9��u:zqF]&w,���|"�uzz:��ӷ;,�3/ف�4
aꋥ��X7���"/��?�`��� �mY��I�F�ʻ�ө�%XHgz1��3C<�z=�������M�/n[#��%�$"n��j�kew^�������X�#��v��8��V��WM�=J:_s���ANV�;��y���>-/.��h�B'�)�� p�t�7գn�UsK����)6LLlv�*��̘M��&;��]��		␨�
�0��aW�.Q�Y�'�6Qc%�L1R�V�ER�6��������CB�d��|с�=C&gg��z�y�������I�A;H�(���r
O�y��	�0l�u�R��:��P+P��_-~�����"ؙ���|�׾mmmZ999Z�f rv��͞�/�a��uV���)@4���.]\@�9����q���]ee7He�3�l��
�uR��������0d�h�����_��}�Ơ~-c�����7n܈����>w�-U/3x��Y��8�h��:.�#~^�ok��ez�L	.��+�7�@��E�ĹI�h+2=���tq�!����+���#��0��]J�?�vHFN�d`ˈ(��T?�4�Ƅ�ֲc�5݈-�d�3�e�"j��J5dv:���$g�"�k���X�p5�,�Z��X�:��!;��͌ҥ9h!x{ZA�C��ސ�ɫ��=hX���%j�	斏Ʈ󉘛���s,َ҉�K㨬�J��F&` �o�s	��Zbe;Y_"d���@�b�Q��0��:Z����An6
2t=O�?JC��I1�Vw+�pJn�l�BMZ���v
�M����$ J7Wo���_���O�>m#�Nʀ��	�M]`M���|��nSDqy����%J5E�2���>��@��Ȣ�=�*�]����_� ��^ֶXq�W$���n��⼁�6���ظE-�Pԉԙ��:`���[YŕBvq����i�<�6:1q�yd��h5�/�Y�<.��Њk6B3n���Y�܌��4 #�:P�hԺ��Mi�L���<�q���[�W��ᦦ��K�e5b;����~�'ʦ
�5�<8���=�AR����P���T��ػ�xzQ�o�֬d��)oɳ1�׸�;�jD��

��أcccr]�0���);˼鸹��� K?E�Lx�9�=��Y�bH��4Bg@�Y}~�����B"��ZO����w�ޤ���j {"k4n]H �Ine�,;	�� B�{ooRm���uxHˍqYwV��`�%3_��гx��FXP?�ۛ�+�%�q����e�Da��z�~t/��L���5�3��>�wtǎLL�[Z7m�LZu�1�k�5,������wd�������)bB���Q�$�~��%����LiN@���^!v@��-��ء�84�;w ��>�F�������Ɣ
:�������/�Ə��r�V2#�H�5H��m������ˋZ��[��x+��g��>e�v$=�8Ib<!�-&&-�:���у^ޖ���G�/Z�63%��R̓�!Z�k��P"{�ñ�4�i�g�S����M5�jt+@�7蜭
9���D�.y���A��ao!�L��|�F.s�D���F�!ȓ�N0VfzL�J:�����B�l`�]w�p�}S�����4�KD�����3ޯ�9F>�A�鐺�ΟgG D������Hۖ��"�qi{����܍�!��jnOv�Yt�?�)w���|"�kvv69le���������q��v ����C ���}�D��0!�v�x"� L�����cb��Y�/�yu�㶈x!>Li�y��%RY�Wx��h�'
�;��Jĥ�
�}���:�Aڣ�`faIҠ�95�2�n�4��ЗH����B��WWø_z����iS4�ĉ�q�r���u�+D��s��c�A����h�KK5<�D�^�=��z�OK�}�UIVbGC�	��r0*3�b�QY�wɲsHX�����TV�Qؕ�Sͣ��U!�]����Ͷ��~?�v���� n����d�P�̑n�g#j����2�d`SI�(��f��o�*�ink�B�r2��܂۶����,&n�M�,��Oǰ���k=���'�gGa蟀�.�vUT��&��X&u��y
<y�%yR��T����VN�}����P�1�1k%�|��46�ST�:V/��ǔA�A$j����2�QZ�&ɁFl��¾f��#�)u��i��K�;�Az6��:�*3�7�<�;�`;3���Y�s���uA(�v	��4�=8�ʾ��>Dn�
j�E)`�|���!Sh8��X����hD���
p�����g6 g�����J�(�k,֑�{�&���e#�HQ���u�� ̻0 �E*1��1��Sh}�wt 5S���q��t��]�J���cSRP��WŸ����	f�:��G�4���_鲐�?j�꓏��L��Gb�uO�\���r�M�)ӄ;D~�	5N��A:�����M��yT��ma�sLj��&�zz���Q��6G� 	4����MN;`"~ZqJ	+<^�r��x�����/���9�pw�qP��{����сO~�AjMMMX�\YSSs���ԗ{����)w*@
Tz��ڰr�R&�K֔�ԑ��fj�DĶ��3J��p��'"��l�q�`�P�|��G�^�H�d�б����ZU{������~&�J��2#���6����S	{'d���?�mi-�#��K���'V�>H23�ۨ����a��l7��DDDh�=����b�Ce1�}��0���^)�G�<fPhݼI�h6rL�Ja��xuW��.��Y"j ��x��2�6J���>)�gQ�V����r�w~�T>צ#����#i�D~���¼���x���w�O�Q�d�Mu{�+���,W�r*H>�� 3��c����
�XY���� �{
X��=�����f`���E� �@�.��$�5�]�TUo����FY��o���Q~�va,��&��<+K5G�rf�vr�{E�� Z���=n-���RSfT��g��!��j�	ʚ~�l
W�a(^ڱ
u١z� ���' �6œgQ���y+`k` ;�F_���񩪪�<��"%kc����Q
�)dط��χ�n�`ع��.��Q�8�8ر�hW���@����
�e_v�
�?�L5�vG��kg��p<b�O�W��5OhSxx�o�F��V�\���<=]Ok�
�k6�S���yFF0%˰Ə��B�^\>dH�=>�j:�q���.�	�̽�>�*�PB��ѫ�L��x��k&�L��O������Φ8�����w�i��<`�8�pSF���/y���Ѩ�J����J:�]<���,���x��×�1n�ŭZ�������A6E<Q2�j��u�O��h��J6�z݋���ݫ(�zO�/�/44�R0�����~=pP�hkadHU�`�Al��Q�*�}  5�+?~\GWm��JFb��BC�Y�.���MX���H9P
����<�XEy7n�hV��Ի��ⅈ���PH����%�S_Q��TJO���u��c�GG���2?(�ߐ�bE��-v�{B/ 2�L��'�]F�`D Ea��2S��pT�Ӕ�����X�3�J�c�~�@�0>E� �P�?<\���������I[J[ZX;��:��DT���C��@@S�%��9�`۲��Rۦ[4V
�	`p�H�VN�<ʘ��{'��c���^�խ���GU_�{::6\��H�L|]4}:������G^�.�8+7��r#�1�݉���ʼ<�D��^^�޻uF�{K�X�	/�L�?�ޏH$�IqE@n�G��!���M��	����&�o�ܼO����u���_�%��q�������$��x�Ow�����W����W�&j�VN@��WX�踞����U�c�8�>0���@�w�ct������7��9�\D��r~o4+$��kAlv�/.D	�E2�hyxx��O-����Yv�T266FZ�1�V@�9�3����&��J��L����IO��5ݔbP����7�����=��8n��-��̓���Pj��l@�Z(��쪁�ch�V������\�h���իW�5Rvya|�8��s�6� �r�Yݒeny�By E��>���V$G�]6�S6]�˽˜ঈp��21}�j�@.�N��Ać����ς���AG�a|�'�ƨ| �>�J~S.)��%��6U��ڿ���OQ�r��Uកg�cD���GI�C8P��P�/Û�/E��s�{�h��c�!v��v�#�N�b�@�no�֜@��9v�9�퓀��� )G5�3�ފ �Da��_���9swf�t�R>�'�)�R*�6���sb����

����&@Q ��8���Vn�X��(K��]@5���mG�g�q���b�{{�o��d��.���uG�ЅW��U��ܞ�,�Lj�B���Z�ῐ�?G'�ھ�\������K�X�k�`���8\%Z;�C�䂚�>�4ee����>�9�X0&$$��=cg����߁�{������î�9��2�{���k� �)W��mu���z)))�0�e0�@�����.��b�e��H��b�d*'Sѣ�O�Ao���	���򳪨���AU�njlA�˛�e\B��_R$0G�k�˱I2�ߡ��+66���VA`y�⎺��.�ꜳ��4�ѥ$t��.n�ߣ�c���:�N�����A���E+� ��S�n�r�b4����K~�3=���/�aFU�ъ��r��-���Ы���n�1�}�|�5���"��Kl>�a#�YhnnyIm |����*t�1E�'�r�x��ȆXH�����B��:thT�sB�w���K�_����
��BB��@���kx�.��R��U�:�mܺ8Љ5d˹���FFF��Þ?��7�.F�����(�FA��ϔS�v��E���U���@G0ԯ� �> ы
��7���6̼��t�ċ��g[��:��k��:Ŷ�J�Y��}���c���'��A��{��7����X	���`0��l�T�%F�P�̼�+1��r��,�T	��-,,�����A�:�42 ��뼎?��9����D��FQnq>�f%���*U�"��|��^��Hq��Rί��ji1�:������L�H�Ofz��<QX��Zzzz�ʅ�y����M���?%��m� ���x46fO�H�\�~ݰ��W/ �(�4Y�4�F?Iыq_����1R���葘E8";c�04�>�+��b��s6ғmvvivew��b�0�ʓw��#���~y	�{86�����u<	>��m����7���}jh�7�l�A�e�V)�#�}�Qt�k�&v�=8�SD04�vw5�.�ܖ�;BJjJo���)'�`����!%�ݽ���=�-��9(���!yd��X�mص#�t&����A�������#�fdϛ�麻���3�S�x�Q���/�H�dmS��wWh+ڦW��]�G6EGI�帖���	啃dr���<2Y����x�	:GV> èV�N��O�H�.3 <ѹ���Tp�'ORΙ72��+sEEE3z��~9�{<��|�$�*UYY��-�t��v�Ζ;��={v�g+qT�L*{�P_��y�a����.�O��	����vS.T��]:�A,�F�NR��qv����xI����r��1���(�u��;�v,�Dw.�����R�b����u����F�G�tK�T�~ѣծ�(��EҖ�����T�/}@Q$��m��eSZ���[� ��3H��H"�4+��.Q��7��
���@����PzKQ���1~aa	ۻ�#���ZN�m5�!��"�G;�
��tZ��_�Գ���w'̍� X/�.N�#�~/a`�N����εs~,�pٍ����j��Cg�讽����\�h�M�A��x'�1\@���	�᪞����Ћ˒���9���&Ƃ~BGP+WFD� :����o� h!R�{�-�#@� F�Q��;�y�P�Z�����D�|�AO�O׊SB��(����h<@}��8nE`li�s~�&3`�_//N+�R��m@���*��U�X�6b%�t:�%5袞��(� �#����r�Z����Zq�P��?�\2}��f9���.��_	���� ըe+����aJ� �|萐xc������G`�T`���0
��T�^�F��������o/�ɀv.G�G�d��?{I�V����ۇ+~��5$�P�<�H^����;v��>`f=��y_y��=B�� `������/z�:���9�Ά]��Մ��Jщ2���gm�	L����pr$����+��%(F�,6����Fm��@�mQ��gՌ�5�/���rFyN$���#@����]j&sg(L��%�&����Ǧ���u�?QeeT��1X���X:�Z�o�������Wj�i�{�Y�~���F[�AZ/����A�:y���C�����Qy�H�cS��y�."��}}}*����$D�������s#<��EZ�����sM�.);��:�D���υ���7I/we��w����G�~�U�c6��~<��z����6��ƛ��C�~Dg���4v�Q[{_�?�o|4�{�y��硭���S=�Mt������M8�Ǎ��$�bZ����Bx]�#��~�ć����D�v;;,�@E�;�x���{"�o3���'c|��i6��&�z��<ʽ���1D|���v�m~}���x��4mL+/�-��k�>f)B�|�� p�E�W�kʼ.?K����$�U-w�����b{'DnNE��Ћ:,�Ѧ��e�Ś҅ {�t�3 *yDA�Mt,/v����Р�ݤ�A�:��������4��*�/��K��%�i�2��өO��a�F�|9���J�Erl:�ҍ��`���:v��A�K?}�">�%����*��!�O1Nk�#�z��{��$3���[�][ڑ�O�A�loLs8�v��L�D0�4$�h@�4��9jO> �]m�����R �#-��E�Ν;MR���ӂ��0�@1����f=�]y4#�X	t�ϳ����������N)(����wov��=qx9�/��z��z��Lt���Pey:�+A1`����s�Nx<Y C�;��[`f�1�z�oo�3���[�n.]�Z�_2O���vb�K
�c���=77��z��_�}�?�؎���������7)������dքH�kld�ϵ�l��!m���Dz
lW7(8�|�1��dV
��޾ͪ{�1*B�288X�UN��X�Ɣ��'�;��Y��_i�ndccs��l1ǽ�o��.O�}������b��6��dv5[f'��2�ij6�2N��=Ϟg_�s���\�	~=�����Uv�ų=QX�@8�䙇r���ɲ�ȹ�?����SH���`fjqqvm�ŋ�5��;�|���v-??�e����� s�˗�X&i"[�]%L�o�Wx�}�I��f�~�z¥/i��p�I���/*xΔs�1�Ӓ�h�lIe4׿�z�-o*�������#���XmC�O�.RU5N���cץ4�Ь��V�Y0�Ž���n�x|zZ��A������w��}���1K���$�o��6E�>��Yv�R=}ݑ&g���q�o���F���4"�Y���N���;�g�����t�u�>ncF�ǲ���Mh_�d���Zi�N�cRJ�6����r~����hwUa�89R3KR�^��5biɣ�9;G��] �@d�B���Ǘ𷈤+<��		��z��uz���Tp@Ȳ��^$�_p�M�q�����+7��k ��q�^DH���"�W�KZ\\<���U}qq��?�h"�b`qM��`zZ��E�_��20�@�ƺ-�/�l&&n,�T�����j�AG~u��器�y*�s���z;]̰�w���XŹ$Ϲ�ꏏ�Ů3�R_K�Ù����O&���rȮF�ib��bbڈd���ߒ�T��0� A����0�q�ܚS4� 4ū�M�:Q~l֭I
� �4ИFdgA��$rt�G�BGC<u.�ᇆ��v¸p����]�9�H�8����X�5��	���8d��[��~�M�W ۀ�����&6�RFaa��/��7��/H��T��񦦦^M�8�M�~Ih�J�d����g�ݡ�Hh���a��{id��~�̅ό=f/��c��u�v��,�2���O㴍αL�%n�E�a�m���H�� ��{�f'����L1��I�s.���|� ��F��}dL���kW�f�ad���Y��q���a�4��=F7�?�d�dD����)A7;vip��1�Gn�DwTB����x
���j��2զ!�tI΍�,��&2�i�,�D���v�Y�ﱕ� �O�m��`[��ۅ�Y��YJ�=�\Br�*0�<p�|������iڶw	��z �%pΗq�mhh�K�K��Y�	@Jj zL�]�t	�a���		��tth1s���!'MLb	�,g�TPp�(7���Q
.B�LG3�u�oJ;g[@��DY��=ʯ��o2��	]n���S}=�j�;��e+%i��Ra�w��v���F����J��C��!���l�!j���:�O,�2�������۷��-����I��)�v�~�)��1��w�d2�����V/���8$Z�̛�2��x��֕I>:|��ev6��M��D���9::�&�c��I[X�8�Q���){��T�cWY�ʮ^b����� �ޕ����I1M����o�U%���y{��� �y�<~�Kέ[~���ӷ����@2�yp����7LT.����_D*�D��g.���~�g����1S<���)[���0}�����e�m�[���P��8~�̀.I����#22VT���	���132�6Gv,M}����*�㘽~�}VZ:]�+CEL0�H�qƽ��T�S�y�i!��|Ȥ��*�v�â~�d�ê�<{�ۣ�v����{�fY�@�eѭ�[d�u�s�1�,�\���ڎR�[����|��K~��xmmm����ׯ�2*�	����L���{	�a��5i�1����i���*��m��~�E��o���?iz�m�}(Z�]���CZ*#]e/���I��G2� v�DS^I�2�{�n��ӧ�B@�R�����9u
�=�Y�1ʦ�^��IH��D������Z����x�@�]iLѥZ�ʅ(	��o�w����4���^�{�QUS�>~�G�e0�V��5U,���6�i@��[�ݧvĢ�s��UP@���.h���տ��p+��!��	w�ڵ��a�%�ג@�#�d�t����2��2}?~���ƀ���`~Y�i-�)�7@�&��Wo�VE�[��J��6t@�����yрf��e~7x��5<M<��=h�{��ly+���t��� =��mbB��6��(��~&�g��
�.�=>��m��}l�s�Ƥem׿��"��pJ>ML�dp������Qq�%�����@��l�/�۰xy�v*��ZXh@!�w:;�����8����1����f�{IK�hJ��˄����z���'A�׼���OHH~�ܪ�ȷ��e�G^�d0n�Fd��.��7��l��عs I~1���ð
��{Eh�@F UW�Ux��4NG��A(��[M�X�Ƀ̄����Y^��-�J%A�U�jy��t���x�c��`��,��bbaa Ȥ-����|�P>Y�r�wö-ws �r1��3��z3��у&%�����������k8)H��Ѯ�q]�K�0�ͳ�9@�x����`��V�@����QU]@P0��+ `!���}���?��4Uo?P5���b��Y`�ɘЯ��H⹊�\�^�*��x.!!a�J���&���
�A����EkUqpȖ[�1���/z�1�"�b��?����a� �����{6��*�����}��s�U�h(��0F�p�V�\u{u��o���ÿ]�_�����?M����2,M�ѵ_�_Q��jaٜ����(0�9>�q~��zLI��_1L`DoJV�G*�T5��%��F(�'Ҝ�&���Ǯ闸�g�&��'�I"���_��6t�c��q��*?Y��+�Y{ěVYhY��q�s�˰��ΝsY�퍸��6�[o%J�HJ>oLՃt�
�G$�l��3��/$B��%���dΓ315�ĸ�7<�t��Oi1X��Y>$���V4���2�)�UG��I��ЍQO^�� AW~��.+�e��a�n@���/.��B�`�QWW����؀fF�Rwlp�x���j���d�
Y���,�b���l�C��끙'�g�<���3O������qtI��6+���~�p�Sa���{�8l��r���u2gv�����������-Tɚ�*�7ک8� �}�Qf<vd=H�4���T�#7�#� �+]�a��v�ݻwG��d؛���$ &VP"���4��*M�R�����87	_��X'Z�}�į�l���1�O��t,@��x��n�s�Nѹ@��z�h���>��$R��jH�;}�=�Nd<dy&dŉN�l�]�	�hT�.:G��a�Kc���a�g���Z��M��g�StS��Q=�w��irLW@@��M�������D3Z!;�J�Yy�U+AV���I��s������g��	��m*�A�]�e�s���X������Ů�����֛�S�>���;�ž�J�TDYCZP�d	�-�ز�Ѧ��&Y����-�#�R�PG�Ph!��?���������u�y���y��k��~fZ���<�3�kr���T��l;��o��ߏ��Ղ�������0�枚˙F�O_�U� x�V��RV�	.6/9�	>�G�IJZ�@��xɋ��o�u��3��sѬf�?a�����^!�����	׃���ij���U�x�C���9oE?y��*�0l�t��/7���Q`ᓮ{>��d}Xe^DI�a3$���dZ~�:FY�#�W�/���나P�[����4��#_r��N��S[���%-��[��%�o=�{��?m��9���ϐ$Y�G���{���;�������7�+N慞)�����)����c���p����D���GC+׮�{�ҵk0��6E+�b.b��Cs5/~$��[,d�C/v������k��}W�k����ۖ�R�:��s�������*z�}�^B�IFY(�F]?�n�rt����O.���0[�ߦJ���mlh�˺<==<W���(�꡸@�U�菋7_b~"��6�RG������$\��+��~Z�IT���I�T|����<>O$w23�s�, H0l�Ѩn�A�Ӥ�sqr�}41�:X�+6��G̷��޵.�"u���6M�z�bbu�E�n���ih,���>!���ϗ\v�065�-������}�����5;"�Xk�jr�__LMҜ.R�r�|�s#�H�<s����n[�+8�� �yp%�p��Ƒ+�J��K�#�:r��������lB�˺�;s?8����	��<��҃׭(��~,ή05���D�.�s�� 8�X�_��Xtf+>���ߴ��G�
����_��;�z��Y��	�(�G��T���F-����)��]�&:r�����p��j����@�����2w�-#��ѭ���.���5###f�����k>�_!W��K-U;��3`�~��#�_��|Ω�':8,C�

6@���E��R>�[��f�9V��Q?��adj��7L�[[gc�r��f�_�2���O��5����P�����毚���/�6��u���=���Ϫ���FjEDD�����0���NP[��� ���r�y�,�����.����b4\�|�l�3���;fo������4��l�k�wo�<GG�)��l$<���?��9�
y��@IR�������߇r'�����gՍ�����\Z�J�Pk���0��nnYR	��$6AN���~�Q�
����u;���]01Ȕ�n��D�7�WR��&=R���m����|�Eꍐ��DB
�0A1���w%�
�*{���H'B<�=<��㋄��Y� �w�}�$����;�\
Cd�Y�[X�||.4�I��d;��m�����r��Z�	)�!�eʆ �x�G��Ā�Ʋ�FT?� I��ם���1�շdZd�<8���م��ѐ���	�˚;�y�����7A��f'������/p����>����ꁘ�����J���LW8/��EQ� ���o߾v���D��4Z(���V�`�R"I�~��_�1�����Ɯ}率K��v��+�ظq��o�}؆UH�M�ɑ�\���Sʁ���:�N��C��g�8�[b�ns�˚4�`�˗{ �H�ϒ� 'w�8�|sG�]>>�$%�֯$�g���i@�?�c���Q�Q�D�qX\�����m���@3�ED�	'l�ܖiII���� 'e#G��ڙ�����GMì�~�{]�,���+���L������\}�w;�����x8N�%�dU��]���Z��3<�			Y҉A��,c���J�>;�{�)|��A«�p��R���o�[�'n�raQ�8'��K����J���V�wy�'�َ�_�*4ݻ��fZ[W�w��(�~�r�����j�A8 �8��V�	~l/<�ui���f�����/����˖�kη��x���gq��#���TY<��b�������\ s`Z����Q��`do��9�/�A�Wo]i��S��*t���*�.����gϟ�|mN �8�����1��������c��LDm���U�.:�D+�����uu��6O�)a�#����a�X��� Rx"T�
y��	ϴ�XS���6���Rk�s�yc9hm=:*i�
!�@xq�������|;����g|�㟜����#7�����Aj!��D��l���9���{���4��:��,8�1�	���zg�;Qc�?67nm�ȫ,��_��U��c�`z�azix�+/�	�t��! Bۥ��J�*�~�T0n��u�~-�ɐ����J�b�iچ@�m�sihmy�|6o���u���E���ʩ%��+�n�1[J|�
�u��*\v���_fuD�8�^��K�46�cW��:�2w�#�����;@k���"��>���;w�Z��ܧ%�B2>��7��M�W�޹��wA�elf�}���\�!�u���#vg7� >ڛ�L˵�$'!ʹU�b�*�N��� ��e�#o]�����+�:�<��'�<��8�v�|�~�j
z�%��� }��/���]����U�Dc}���oQ3���>������.��z���U]g��Y|��E[�e*H��>�Ƈ�ԑ�]�l�Q�>8	:s�|�O��I����~�q�����n򠾎�a�+XT~��'kAjj�*S�л�[��7�u.��J�һ0Ѯ0���<2�⣼�$ �h�����4�Ʋ��<R���1`㕕�w��%OX���������?K������ �/���k��z}ĭ�l��qV���;�*�Sς�j��t"Z�ќӾ�m��� �������#���J.8�������\��odt9��c˖-w��[�����!77ܠ�c&�UC^Y���葿��^齺�DR �~��-����6���L�V�A}�ͭ��*�>|�xhr�ם�,rwVx8�IQGWy������]�bϧ��q*F����QL������CA�v*Y�9�;w�v~~�jy;XS�������	��1V!�;�F����V��^\*��@Bn,��o�"�uiH��\V6��ikk�U����1ɹ�=�P�U���ǻƳ�4f,�	(���3[ݓ:�s��i��	| Jc��ywn߮V�[�:��K��O��|�X�h�Ft?Y���Ĥ4N���y�֌�#�0�S��?
0quu}~��V���Դ�H�W��W�%j"���I���o���|>�tr$;���f;�4���B�DUU�+[�$nܿ�8�H�:��pb<��H	�qrUD2�����O/�[�f)mؐ���*A�;7on��/�����9��L�������M뙳�{+d}����ǊO���+��L�򙚘�R� d������/G��a�7����(������6_Ȇ%��ԜZ2>%��r��A�����2Ѫ<^����l��n<�<���������{V�6�|���Z��Q�%������j���e%m?�;'g�}]�}�ߚ��ys)(%=7��!8���s�'h�N������l�`6�:�q/�էDd?��?Tv���ݻ�G� �W���fw�3�t2�����d}���Kw��	�?̴���?�����k���oK|�!�^�v--.Nt@�VQ�e�Ye�%"����L.,4el��d�fC.���Чh�����L�nMN��Ȫy���߿L�ulP�o�����K����3��O^M��O}�o�2��K����̋�	�&D���kK�o�4���eN��
[p-���M���A�� `���ANsi�r�<l��4ѽ��*�{����k�e�'����ۮ��ד�w�����|}Uל\\�$�qpH��'����/�w�����hbgle������'q� j�AII�w/j�� ���e`�u���6����SQQq'=R�b����7SQ�����	�5��f��~�u�4p]�9)��ش헥��ʖ��~����YS��6�7�����ϱ��2��w�j���in�HJ������`H�����$<��(���|w�K�'��_`���kͥ�0C/�x����C-�d���b���q`sCÍK��ܼ��ug����������g�i �1�!���H�Qx<���9�!c�;������`]"%׳��/^��d�	����[=����/5��B�����o����;�����2g�rI����><�����g�r�����e�VJ-�o����@��Q��c7|8(U�E�>��K��8�X[gǫ������塀�����f��m�%�ȃ��Pu5*��o�}�L`,��o=LJZ��ڊF�|�����I�5�#�!We�RZ?�>M�tUwk��Ϡ-eH�1����+R� ȃ7�⮂z��h�"A_�pA{��pE�ɹP5Øne��[r�j�����'�օ��)g�E��p���[���K6�[�]Zj0h+��u�2D���K��\��耬R�?��N.A�\ED����bbc�8�L��Ib�ǿbժZU�54�?���=�,��$�q�W��	r@�m�)ɋQQ�ǎ1ÓkTY�;�&�����}��SU֢e����0��<�4�z�W��ADt��O�̿.���,����/g>u�.�q��dWГa��OODh+�=1�"�_2���ᑃW�q�瀢� ��[���`�#4b�!i��xzz�v==�ւE�?� ϓ4�9wm���f\�;%�&O1��E�D�܌��GYoW�9 +Y��Ջ� D�Ǝ��*�����ھ8u�FU�B��̭���Ϟ=362JvnJ5s,��$���de�G��R� /Z���m�D^m����-s�	<]�k$����5ı����i��F.M߰u�E�3fy驩�)))xBə�d��9h�!��������̢��b�u,�d*b����f�҅����Up��tnTlr� ,�ML�b���ۼT��#�<n
�x~]�e�N�5k���Ӌ ��7R��b��V�~�������"b�5�IL_g'']���vo�~u��z2�H$������TTT<�L����m�S2������7y��<6+D�]��@�3ٶ�$�q7O�)��<��u��q�j�+�s�?ʆ�Ĩ����w"����EڒP�P��ލ��X|o���9E��L�H��@��,�K|���K�w��?m!߱..B�R �Eݭׯ_��z�~�
�r��I�xR������p�ӈ<E_����08�k<u��K���F��r���t9IP�=Eu���7X 
�Cʻ�?�̑�������y�Gw�cy�g������[UK'N����Ͷ	�(`Ïϟ��i1-���ҷ(t313�ο��6�Fs�q�v�2�8L�V9�+Ʌ����_�ƁO=y�y��{ZW�^%ώ���9�	a�᲻{1y zVƖ�;�h���׫W�RS��V�r8��ڮ~����������ny�֙IK�X>��6����?";v�(�4� ��d)%ʭ�8X!��̥�B��?oߚc%K0-,�R�d�
��ۜh�]^�5`��x6��$��]w��E���RJ᧊t}�y��R���u)�ғφ���������D��b�Tb}h�C���`�-���xYڠ@��Mg�ˑTކw�&�3���vH���k�e �E��;|�i@��׀)"��$��ϫ���\�� �m��'d�xpZ!rsVi����]�G�W�̲e�/�Ф�����׭���a��q�	d�O�C2K�B�°BC�<w�&a34Vœ��"&�0�Z���\,� �=�g_��f>�,�p�Y�PɮY��n�FFgH*���X�\��o���E���G�JnV6���d��ITrK~6GFFa�}�r�����!���\Z9����,,,o�d���FC`VW�\!O�u�Z"�?�\<�$%�;������H;��l"������?u�aA��b�/^p�G�A�� M7�ڌƂ40�/�W�Us
�W���<�=u{���OXy&�3eٵ5���͂(���4Enɴi�2�	��Z�����==N�t���g��Z�ǅi�I���rk F
���;�
%�>-�]Y����`�J~a�E/AY��Qܘ'g��Bۜ��X�����5�,<-Ԥ��A�T����HE�����5Y딕oi+̀���� ��I5]���+B�iw��'�1�=�.Ϻ&���hXg���g�n���y,��7�I������2�U BCZ�����nU�#�R�mʘ�MA�kq��Q>�[�K��a�S!.��򗭯mij*�b��sf�ׯoWVj��� �|������F��qk�	PGk�EN�����\�
�@s HO��L���hl������M�]k��������P,�(e�2>��C�28]�@���b��2��7�<0���rN�<���Y���>>>�(��
�!G��C<�Seպ408���g���e$��gWF�~[��P��y��ё�+��Ő��{���(=9�B�/}�a�����Ԕ!���D؀�z�,�nޢ�����o�ۏ[y���@��٦t6�����
���Bƍ8�бS�[2\_��[_�!: I��c˳n��'Z�� �1��QrO ��6,��o[��,��]��ѣ6"�����W@`�4Uǣᐴ7��W���pOv?>��Ԋ���KT�,F��E1�j(x�U<Z�Қ�|�K��v]L�z���O1�*o�8}����]o�n�0V"�'��B��W$�x� ���
[DeC��k`K+�s6F���~h�;���0bH��CLv�l�ڟA~�@n���C���zc�N�B���ooAp����ת�� �C��J\�0;���W�1�n=�=��b/<� ,fd�|���}-f�h�,���QB*oE�������lr�^p��9��ɉ��!!�DY�Ǐtď�b�t+��j�X�=� < o��X\y3�������*Տ̧�s�6 	*d��m���ԃÎ�ơ��^��Z��E���ڀ�{���OD�V>��}�ˀW>�����9ŏ���;��-����?0�pݬ=�������ON���̿}�Ύ�ܝZXh21`]|�Ӧ��w��'�����zEE�c,Ny�`�ʌ�D�km>����͛7�F�������<�ܲ A�m���[�GL��:�!'\Pa��x��$9rY��Ǐ�̥�R�]�����H���x~8�8�����	&�&��ǿ�9m�nĕk�/+�q*^W���X���?�f�Q���#,$�G[����.����ߗ���x��� �l�:M�<���6$M=!"*�
|�?G2,�.L��	~�W\��#��Sz�L~]#Q12:z1&D�f�+c����m����ݖ��P�N����e��A�x��9r�ѣGQ����7�����!��� ��'!w����|�E�����),�OXke�eKy��z&�ޯ����)a����9��^c���>^j�03�~�����Y�Z�u�l�w.ã�<�ٌؙ>��X�lYuA\�'�r�.#��$�5���������̡Y\�����ލ�g ���� /�2utrbN���2��,�
��y��
�qtt�Cv�����'zS����p�O�h=]a�!��o]'����:_C�4�P�R�v@&݀VM���۠ڐ]ɛ���ޝC���e,�N��N.9��1>����x�(��9Q.�k�B?�m窔�#�dN�W����Ct̗޺m�ggƸ�I҃�W��cR]����Y����|�6�c*��M.8._W������%KT�75>	
�?�iR��l�uy��j_㇂��
Gww���V��_�Sg�'��&����0Ǆ���fkx��y�t�O�V���{��c��_�{�Gz'>�hzz��l��,m4}�@�S:�Is���~�]q�?/�A�E�)���J��}�O�##��Iˈ��ѹ�lm�b�~�C��{_��J|���9c+Z��%�i��2�{ڃ������X����`B��TI�DV�5�u��IB�E�����x�~~�J(2���6Ѥ9a�]ݱ47]��)\��Pk #` [�[��m��X�sj�g7���&����/�����/�Z+Y|���<e������S�X�Z���H�W�<��D,}�?]��BԘM���!�ZQ���|+�b���j?�d������H�Bk9-?'�9�������A�)�i;�V9�4�g��QOu��Dk`���?�S���a��^�|)(.~; EٛNkN�`�_���A�Xק��Goc�CL����u���sm�������Z\�e�ݿ����`���X�ï;;�s�lx
N�yf���_e���Oה֯���-�
d�������� �0L"2����ã�Ѷ�X�뻡`%l�����p���*,���ӏS>@�ߢ@� eQw���i%��,�2�a���Ԛ�~���q�w�K�v``�8�A�W��SwRۑ���<��to�av}J؛��2���S�/�!�v#􌤙,�o����1�TG�J���[s��4r$�N���_�C�b�)fMg���^)P��H�'��3gμ�Kh�8ƨ2B�a"�\��q�RҤEq9 N��Thm��e!�|����Z��^S/�lw�f�9ƃ"*�`��ttt�p�\bx!۠�*��g���?c�|MP/|��G$���g#ӵ
�w�Oj�k��⍱����L��ze<���\Ƭ�E�k�A�arH���;�0�i����Jh�qQU3�=˨\8�i�$}���Y&��^"����$o�����=�j%�qH1�`o5��|�k��^�>uU�̯*e��R��1�VvEU뤞cL"e�{%�&�~�)�C8>{�g`&l ���5I�i�Dԙ��?2�'{d�w�~�p��b�rFk�l�	Z��xç������a<U(n*�o$M�+>��1�Y��E��
�������+��d2��`sxC�Ŗ�xC䎔K�Ҹ����5�.�C�N�! ̍Т�B�c�A�l$,�,��$�kAK,�Ԉ:_h�y�I	�ʒ]s�@�rӜ����+�LYմ�v�D�W7�� -U^���K���"8���tV��"N���rD����_�`w0݄�V:�o������2��;	j�`+�ǵ�+8����c�/YZ���rB��Z�K�~���lD\kK?6jR��k����+=f-�6���JX
4p�?~�������6t}7�\&��� ��y��t���U�u�����? ���*���c�W��v�^R����*��=���c�ب{��;����b.ChNl-��ݔ�j��f�y&�YTJ<�
v��݁�{��3*� ��'s/���$_Vq����O�J(��X�OIS�8�����L�̌ցt��fc�IA�"m:^6�(�ƎrbA,̚�č�uww���`�噱;v<����bߵ�)uԌu�ηč��;�_he8�"δ|f�ɋ�f����R����O,��b��F�ϬQ���O�$ު�`����w+�SZi�&("�t�g����GP6j���q�ꆏ����U�!0J��Э�:� F2�Ak@XPPwz˷��al1�3�d����{U����*�|�yl�ڋ'�}��,��̽�V�iӇ���<����P�+!� *>!!aŵZ��죔C֫��"�g���se}�,y`2ҵ�����♈繬��ò߉|�z�I[�*e0��!�ρl�����#�x��9���Ǝ��Z���%�i0i| ڕ���gdx9I��Z	E~��Z43�n%k��M��+ ^��9i�)��0���/��7Nb��0gAmijk�~�05xh�J����ʊ u�O �H�1�	=`�~��4W�:� ��Ev%{�7��f�q]k*�m@` �<�:ᒃ<d�Y�$Bn������y��'�����-^�v��j����iXrk��e��=��
�k_kA�� �mDg���Ֆ���T���Q���szPU�P̫nn7�����j�� $:se�LO,|۫�p�4Y9J���e�5�ˮ�=�t��qF�LWc=Ǿ�Rt��k�[::��	�!���	�2�s�f���zHVn�Q ؙ�r��(�<�c��=���,��		��A�,Y��bG��=?<��b=g�;�"��I+��vދg&2Ņ��LZ�>��:h���R�T�5��ʎ����9�Zq�:{oFL���Q��kK����G|[U��3����'�V�E��^o��]�yA����%��ep���~���5�"w&�xn��BEM�*++��*���++�t���>���V
[�����hG}N� �Vj�����s��s��/�z��j�ÇeQ~z3�MßBBBH�Q�aXB�(D�|���O��fDb����[?O��f�w�t)0�mϋ�V�ӊ�kxѓ���H�jg���2_H�!,"��c�e�Z[ooE�v^_�g�Y�T3�2}�:|7v��3��@^�����=�v��L~Fp�nan;��CCC�߸���p�m�ņ�Xu�׊	5y�dZ\�Q�ˀz�>4r'Y� w�0���3)���G�	�/�w���[����@��C�5,��Y����&@��z *˴�/~��y׌�v�2�:�`%4=
!�n����*B1�g�e�/Tg��B������Z�`/mpk����[�2��G�P��B �~�h~x���S$W���p��niQrĕ�����x��`;v�	�����C�3 �;���.�"���'ѠNV1�&l˱����{��9�^gpd��n�
x�	v�gcg���};��w��ࣤr�\��<U [��qq��a,�����a5u�ŦB���8����f�6�L��s���
��7��2��71�N;ԝ�?bk�Hql���X����ʈ�6��z��1'D���;�V[ j�A���ͳ�|{��`t,����l��c��y�dD!�Hp�������f�n�� �/ 
����b�NZ�n3�l�Ś���euQ�e�h��(a�� E�Xy��5̀}���P���B��c{�����'�	`�T�8$�?�c#�S\a`��5vAA�@��Ǿm��a&��1�م�J0C��K�9ۻX�c��H�ӟF���&B1
���n�ʳ��c���J'��B����GRٺhZ��:~��)�
�]�v�3R�ՙ`u�m3V�x����H9,�k��5Z�FZ,�a5���dBA6g�.��
�#Y�[�}^�q��:���r��)'!��������������h,܊�Ϝp����#Ǿ6
����� �+��mutt�F��8���
��3N�f��Ԩe�>���J6Lr�s_���M�'�Q�2W�73��P.NNl�����V���?'��m�"T^^����P�XvycE�ɪ����Su�Ũt�D�`�&^��+�Z�m�\FPo�&qU��xFб�_=ܟ6�`T����us�l��6Fm����𺀾xx÷]ha��?ݓ�̫�n���׶��`����Y�8�aI����ྰ���4[q��W���mٙ!O	[��N�FZ�v�e81�����Y��1ܻ�^��r�����S��p)l�3+���dyE�+p����w%���U��e

��p��S��l�f>l��	+�Y��R�"��:!�F�)�k���:)Ǳ���������m�j�m�J��l&"�>M��}�7


�9$H�:�P�0Ya�S�	mq�E�v&� ���h­�z�X�j�n$�H�	 v2V�D"Jjj{��5�gī���Q[��K��	�w�bo�>Lb�����`���-+�$��ͪ��zS�-�?��FivNN+๊�؁�FӚ[�v�;+ 0<8�B��=aIm��_�JN;����:��h��Q�'#D��ɐ��&&O��hT����tEEE^P$JX 9\dL;M�Kd���K���1pF+r[�#���-w�x��M<S@��j���Ә!}U@7�:8)��4�b7�(����h-� >�	����qk�oΰ;xP҇Mq`d�K�]�^y��x�����HL8�Cv]	Ђ�i�s+�A�A��@�1�n�2�<�(�ܵ�e)j�ۇZ#G�r�D�r��-"���s��It��֩�
3X�g�uWyn$	��-t�f���>�$�\8c��~�������]Re>��~+))	{�!��߀Φ#*cl��=}���6WVc�� ��zʎ��DO
;�Y�oӶ����^�0�3����\�|�5�_	5P8������#�z.��g�C*~��Q�?�O���z�G6>�j�bK����B;ʽ��j@��A���:���wz�Z�0x�౮CT�vtt�ąr�؛\�) o�'l��
���[ɗ�}��ϨU�iǣ@�{	`�
Vl�	��AV-�qr3vnę3yY��O�3�-H����w�X vU=��j�	Uە�6	��D�$N�H�՗��9�a�i\� H. �,  �)��F3�s���&̟a��֬��7ia׆-��w� ���ᪧ-v�255��&���1:�G�V�����ؘn0�������(�t�]`H���y�&Ҭ�E_�~�Ƃ��틲��oJ� �[R�b�GY�����ts�����oǦ�e"s�>+�9Q�f����23�!�J;BJL	�i��s�:��O�GV3��2��`$�r���*�p+�T�еȥB�KԚ��d����x�!�`j������!�1�
�>0,/�1��896ޫ)~�X�ts��������lق��Ţ�$S�2��=fv�����h�M� ��p��1�M=�4Y	�WX����㕭h����#��:2:px�k����o< �E�&ȭ��dLz50��72*D�W�+�H'z7�O��E!�׮i),�b���|ћ��%Nd�(�X�N;	~�_����뜕����1p���se������ p��h�އ�v����|�+\zޖ�oW<�^-��D���M�H[?��f�j0�zS�~��j�� rlu)��%,B��='����ַA���3�B�Ug����?��9����g����I4'�+	�ɣG�<����y����K�������1֘xm�w��_p��ޓ�w��h� � M�¾�I k��l�VN��� ;����	���y�=���f��MMN�+H(�ps��ϟ�c��u���h�1�1$�"���Ò�3S�C��<�b���������ua�	�cJ���t���ߐ��ERHHֻ����̹}�������3G�?oq�qf��@�1H����q}�z·�)�f�8�^i/��`:6��U���-5�6��&�/���X8ۓ6���X�ct�f1�-ja��%%�w�=ִH*����uv6B4���L:d`F=}cA��	~���$����u;��,Ì��pw◥����5�m�g���`R��NΜ�����dQ��(al�c�]��y��ͫ��g8
���� mX3~=}�t��A/y9�HU���»Ӎ�b�Ep' rs-,�����Ƈ�Z[����%��vN��~����R�2������T⹨�	�����ۃ����z�!G٨��:|��,���0e�?�5E��΀�0��\�����y��11���1�g6bbD��-����d���0B�9h�o=�D�fv�Z���X�{��(��\kjs�����䛃PY��.����w�4���=���Z������([:�}<6��>������[�Ӵ��E���b�J��oP��$��Bü�R&�+^�޽{�>}��~��݃f���۞Ţ��1_��El�η3�%�}��+��"���tɕB"�{��tV�<g�s�;� �N��7��k�}�.읁�M1�ZI�<�������V�'��1�71�#� ay�Ϫ�132��`s���^/[Z JP� �D��s��@L��K��},�o���g39���j'���q!!�3�A`pաء��u�ò�,I�!�T^\���I�Ý!���o�r��X}�֍3Ww���(�D7s"��F�����[���#���ۀ��8�h�J�G��UL�HtF:�4"D�	�� ,�e�����\YlɊ��go�6���q�ĈpZ�s0TAHÆέr�56�	Wc�p�3�Ȼ<
�kc��ao)�O>l��,��g��e[��A�l����ӊg�}	�]P�<�Ӳ� �:��e���$�6�sr����IWά�9V��<0����z���åd�}`��އ'�f⪦-�����F��J�Uf-f;;�AV��|�u�aXƙ{�S�Y����z��f��"�X�Ǽ�`V�� ��:��^��b�!���b�i6�����cSv�#B�p�<8�mH��i�賰��5׌�-Lk�J���^����Q�9����ʊ�l�Ӂv�}�V�y���$'� �ʏ��(.l�bx&Y�����Ǻ°�i�5G ���ʿ��B����`_Zƽ��2��_�V��T��hF��ꂚG��t��ޕĮd`�ب�\:�>�xrrrү/��M�t��M��z�?o�!�f]U�Ob���0��߅A�������bj�w_�r���Ǚ�̫�@� �֊��K�ut�O
X�&�m�' q�&E��ܩ��P���^s�!+{�p�ģ8X�̜���6�3����2���@'d�>�#�9՚J���{�d[�]����gk8'�1@H�!<�Z,�#�Q �i�q�/z�����ζ�h��|�x��V)\w�a�2�y�=���X��b��ꆆ�$4ҍaTJ `s�?��<�
�{1�����G����x��C��{���y̆���/px��Uk����ث��z�77fgY9Դ{��E+�[a_��(��khL>��fu�V���_�o�0�������C?��G��4J���(M�⺂�Ʒ�Ko�{��gZ����"�:ܲ�Y]�Rg/��bUY��\�Y�?�T�_�����iuLN�Ǐ� W�ip��y�)i��gx������`؛<��}M�**BxԨ��F��o�85�5�N[[��O4��*�2�C���L%�ōWg����11>��ގG����/��~��^4&�RP�9~5"�Z��&��e�Eك'�^��m� �>P��_���9rD�>�м��7/djOˁʹ�NK��W��*}�n}
V߽��׎��S㣅�z�,��h�8fH��>bӠ?�S�O�&`��zj������\o����nę3g�G��׷�RjU���l?��.-��qr/���(� G
S�_X���\�Htl
X�Ǻ����"�=w����0�;{J�n
j���x�\���
�2@Ew��ġ�/.��X�.݋0�kL����e��7o�#��<؛[��M���N��?�ǫ��yvt\���3��|�"�8��L�|��t�@xż�)�޺'s�]]��<�
;����� �h�%��rMUa��+��+���=٭ ɦ��c�;::�F�M�]���?i���V>����B���t��	���vUҏS^X�������� z����Z��[����x<�Ss�t¿� ��>p�Õ�����q?d��S���u�+�؁��+l�'���j�s�ʖ���=��I7�
��z����{R��"���>�!2Pd���HYq�⏄c�N��Q�kş�RqD<��ӧ'�Tk�4���.EW�sZ���-�>�a�� �p@"�<�# ސ���޺���,Z[qG�*�/��O�/`��?x��5��i�c/Nn-�w�0b���~��@��!���q����3 �x�u׮]A=[]�.t$�=�3hb	fb���<,��v���|@1:*��+[�x�>�l�6�
��w���^��Gz�m}
�*��@�)�t;j��w���G�Ѩ�@w��$�$��ȥ#�������@E"~v�h��=�z|�+ׯQ�Sʒ����!��ޛ����Ii�b�yĞ���,���X�k����!W������N�gO��ѽ4B�6f��d�$SO�+T*���;֩=E��[vD���Z���L�Q"�!_�x�/�Y�w���Ɨ�w�i�Q���W�~�J��C19���Q^��ٱ&͉&e���@��o�!��ʔ��e��
"�YH;��H����@K�6�\�|Y~������	։��⢢�z��ކ=�������̟,�m_�]�7'E�;�R�>�*�/�Rw(k�x��߿�G�UVV�����
o�7-=[�0����py���c��F�>H��X���hZ���ʿC��'��MX_P�R����z25�g���J��"7,9@��G��AQ[[�����x�l�hS��]��J��o�@��!P�79Ih8u�'*8�CN�ih���)����p��C��4�v&Sl���=��8nȼZ���R��7&ዀ�!��=>�)�L��J�R�y~�O�T�o��t�џ�H�xI��y9���x/�`�V��3�!M���gv<��N��U�����
��m�U!�:����j�>W��9gqK��ʹ>��˅����q������\�m�ǰ������v�������C��)��+1�$�cw/�;9k��� ��~�냶�Gھ��{3P����)�oT7�U������Z���6h<�i��%���d��ǚ~�G8���+p
^�.��3�ߪ�b�������7�zh�=\�c��={�<P=Y~��Y��q�6��2R)���D��8��Zc��>^��#bu��}���fY�C^�����{q0BK���'�C���$��}xp]zW�.NN'oo�}�ҍw���P�����mjo�������6�����/�Ic3��;wd2��3=��L.���CP�W��;&�|��X�$Q�����w�Ը��k�b�v�̡�CN�3�Ni&��
�,D%އ�L��w%)�
e���S�^<�BQM-��I���ķ�뮿z�:ܽ|���e�d��Vel��FAN�5x3GS��@�����;$�zA:}���O֓��8�*�?E�ˍ�u����7�����!������� �޾�q�\#��d�����o�I�{^�x��rM���P/e�T�,jyb}Zc�!$��9���I�l��0ܼ{�[�������h9�ʁ��G!M��V�K#��ŉ�H:'G Y����6P�zB,�|%.Ж�\�?4�J�� Y���|p���1cu���ʢ�ᇅkך=��`@��g�AOOC�_5�rr6 ��({��m���)4o�l9m1�V,I8:j����E].��6�� ���C �A 8��P����e��W^�QS���L[|�~��=E��H	��φ1u�o�2W��C���x��x���X���D�� ��� `� �@�z�Kk��d�.2QQq
�Trko�w����_���(�V�D���~�F`��͇2�T�G�ȶ���}��.��̒��6M��O��=�Ѵ���e�%v�\���4����*��M�\6x��C���ܬ.�!��{f���oޘ%������XZ�G��L�G�b��q)<�+�NMM�US�k�{�Ň� T�-�<�GZMfϺ�p�OYA�~vͱ��o��Pm~}���{�+�z*,�/����{�/��9����\sBΝ���dne���Շ m��{-7wh���,*���܍����s���ۼ�4��Ws���o{|d����c�N=R�f˅#�\��jdd4���oP��[E����o�(�K�Y>�<��ĥWw�a�2��|��d=�իW�=���M �k߆��Vbk�E����/�o`9w'E���ΫL��[S!��n�0c�F�
M��@Ugx��v�k�?C�#�t4/��\�
$-�1��l�R��6�o��b)ؽ�V�#���ۚm������
b>�}��<
7��TZ��ԇ%r||�cbb���<y\-611��M}pjN�<���(w�s�$�P?�ɛ�*
�E��Z:�a�O_�r�l�:v<JK�1�`��
lnmM{�rϋ�ϫ���e�c�z�݋NQ��o�1�؛���e��w�#�;8:�hN}�<���9�8ٗ���<��o
2�	�|�W���D��Հ6���@ �c�����哓�.������D��gVev�(��{�\|V[���RS��-��e�үk;ӛb���&�/7g�`?0�� ��'��6aϽ��։�������Z˗/OŕS�򋻤|F�MFFF�mm7���3��3���Ibu�
�ۯ ��.f��͹��#Oߺ�����,]I[��`��5��n� ������].>y�~��T枟F⇂tJ|�6��P��.��+�k����k�^9r���{i]���~�"���\Ǔ���1�>����p��E[�43���Hi|�*����A�azS�LV�%W#�+ tJJ��_zS�'D�܊�E���r��bq�;w��ǽ߾}����R?P>>�1���a�.m���x"+3h�~�n!����ڵ���^�&��� ;��/�~�d�~x�(l"u�l���#���|�R�klhx|K����C?E��B�w��7e�����ޠc��M�4j:�i� ��� ��$5?   !���нշ��~�㛚0���P��~|>"��WH ����=����u�m_�`d������X�v�<W��-�~��/�&Bb;��Fl�g�w/�;�P����~�
���δ�����ڌ�/ޙ��?8���=�M޷�/)2KypS?��s�m	.��������U��oѪ-[��V���pD�}i�1PO½�U�S,���s��X�m�֏�@/�c���K1����F��y���Jv�x�[�-Փ��ӬT�7�����v��I�}l3��G#QV���}8Nh[�9D<���((h�(�L�-֪���oT�WO���_}�o�H� wT$Q���~~�j���"~u�qm�t�~�:�F�������;��6<�����lx�U��tYi_�@l��=�reAs j*��.ޟh^�{'��'��7���q��)[�bU	��(wۗ�5�4�nQ�8qJG��W�үg��A%&��+�������C�N|�+0�Q�_Ɓ�E���������mZ*����+=9[p�U��s�<��,8	k4�۷o�cr����zn������~�"0�݆=<��9Xm�c�TC�̓T;��ي`gh�l�v��IIe�o�ؾC�2�/kI�3sW��F�/RI꼴>���!���ǏV�0�&?z��p ����f7����b�
[��j&6������
�[5��1����?�5���QҔٵ��X�ʓl�l���{��K;����%0ln��r]�0lA�_�����g��aٌ�V�֋�t�������V��~�b���/Gb�0i1�xt�RUS[��~���ڬ�l��.Q�d ����2'�kP9+l6n܈�3דU��R�˿��u_�+&"ף�-�-[���5,@�N��(�޹>a�o��5;�൴�lc�L @�S�[N�:��8�EP�!,]�Y�*�@9�X}fh��~d^v�贝*�V�2DWY	fXX�_b�u �wC����]'�2�:qH�AL�(�3�ZP�xb�I�9��<�'�*��̅!�����dSC���]� t�=&&)CA�j�\]I�~6T�z�
X��(l? �x�9��8H�*y}W����}}{d��^M
	*"mx/$V������N5s��(���C?4y�oL�hvr��ց���Y:b�[�\��0$d��k���`�.�8w.���"�]���6�f#� ��򐈄���IH��g���+h[��r;%e�cmZ��%	!��X�@���9P���.����M�m��ނ����~4*<�-U��P�ņT�X�7��t�K���R�<��kc܌;����c�;��L�nX�U�	J4�dQ� eH��"9)93�"�JIr���$�Y@�9���'����ǳ�Qf����n�[]]Mـ��p�坽�0H�jۧ�=&��휁�#@
��Dn��Y[ZBq{�a�fg�w��δ&���}���a���H_��j xm���JJ��[+P���������/
�j��fh�b�U��+�*U��?v��6����+Xmym��?){�ȵ �4���F���9����U�!]R�m'T�Wl	_
&�+U��y���N|���=�9��>���f1�kN��`�����I��W/�g"�xh#c�w�H!��]��Nyyy��i{g�'x�i1 ���]oϡ^\?_%����U�N��`��j4��U���/'�:�������`Eݰ�ź!��w��gK~��y�
���b��U�����ͥh`��]��G�_�Y@��	�`�.e 5�����x�)�B�Af|�0T@�F�nA6����r�%��� :8}4a�0b �e 6|����2�I�9N��J��E_\�������|Ϯ$/J�z?�J�� ?�J�ؔ+ @ި
<�lL����뱿(a#m���[{��{���˲���v|Y�� V����Q���}o�e������ 0C�����ǏM
��d�z����g�GPكs��)����\���E�������|	�s�y{Պ]�[���Z{z�C�v>@D��eHp_mmmD�C�����w��6�MOW|/n�ng�#���y���t~��:���2������N�@R��Pel���k��iUxG�S<�q�R�2�nDd���>yBaT��:���}y��ki;�J��cכ믣��p$�S����F��Ҟ��iMM�Ʉ �9t�]iQ���:�/����uE"���*�F��0��9#��ϟ?aC@���8��g-U�'���g��:���n�I/b@� �3�:vI�[���|�UFc!lO&�����4B ��BqدJ'=���p<�1�齄�P��~�/R���{��6*q��!���
i&��%��LNN���%�7������k�G�P0�a�|��q��)P�9|������@W3���)A%j3�S�JP6��i�N��.��8�~��;^:�y^h��~��HB�C.X1�C�i�����2��� ��ځZXc�[bN�� ���).�������Tٽ� �F�JެP>���iH�����6g(������vnT�@6C��<*ג�3�E"��4�&��I�8��N���-J �rO[;rh��Zg����g�4���^}|#�q!�8\��^LB�����#�������˗�QB�'���z��Z++,�A��&�QS�_vP!+G�vg�7� B����Y�j���=z�Cv"M�VW�?"3���}6�<�/^�B	

B�70�)������(���1�����֚o���a!hX���@Y�77�T\z���M���P�1�40�	��KJbQQBX�� ������HZ���F.VQ=���.&	
</�êCR���`�=�&�}}|!�� ����|ow�9�n>��C�*4W ,���dj��&����� !�h߉������G�,L�z�v}�B�c������[)�䴰�_��a �C,,,J��-āW�+�S&�����g�߸���5�u��cx���;������
�K��q���
,�e�r�<(����.� �x=!/������~�CgExo�t�Tո. �a�0�	@�fg}�-�30R9S @�����d��)��Wƕ;�֝$um��i���W�~�������~���>�}�"d��e!�s´���yN�����e��C���$����d	`>��ɨ�Dc���}||�߁���)*I";�0�����L�"��zDRw�.G���@5@Zα������QUh���C��/�F����oW�TÎa��Xd$!�y%�H��7��6��\����G�3�s'`{Z�K	f��N�� ��}� �z��������\u_���@���<H�ˮ��㳧�����.��uN]���� D�L]خ�اpf{m���˰�"���a2hJ�ӯU숣�DY���*���,~��^XЁ`�mt���@гk����*(�OP�����yRԢ����A��'�؈���� 
��z��8���M� /��"��PƐ�l�wmmm
�hR����I)�Q:�6	DR���,m#�XwC�}Pﰋ��zK�T���sG4����5 +o:X��a{��u OJ�����G~�ػ�N�		u�·�'�В���	,G���|��
-��_ ��l�u�����P �@̀��@J�������\t2Q�@��KT\��I�b2�,�]e��wuYW��8I�!�I
��A1,,,%���7>�R��na�Y:�F�;X�E0�`T�t�
�oÛ(���;�Q��u++Y[[kf�ק�Q����y�+ѯ3Ka/bW�.gZ�S�Q�b���Y�����,L�'�n�;:����5�����_r���q����� (]J�7l���$Vo��>���y�����I1�޵vvj^؜t����Ot���#�� �!1����$$FH@X7����v��"���'`+� *-�G���F�p���Ā�-D�����6M1b�bG d���C<��M~"��b�:;;��v@�������O�āG755��O�
 t���г��wDxxZq��z-��x��ߪ}0���>,�t���Tom�Ѩ+q&M�$������9m g �O��i������;����`�C:����|
P���|"�,������ ��_�|�����ݎc=��;�מ��\ȫ��Qg)���r������+*C/���t7d[�f����>Ϥk�X��}� ���<����]:�΅Ċ
������ِ#�'��陙�1E��X��2�q\]u���=���a_��A4Z�L�F��sڀ�Nt�1���~���<z���Ψ��En�SC灷�X�~�n(
b)B༯7���:��&\:hY�br'��L��5�yp��7�8�d�m�YW`��ɴ�

bW�8�X�Zs���x������?�u*�ב�k��<��h�R3����[0٭�BAF��&lv���l��X��.�/����ܡ���˿�P�ttTo��;�@�Ng����qη��� ��� ]
<X޻��E	�_�B��+L�@��y�K��$����%�Z �28�3S]�_�*�m�;vjdh�))� .��׌<&�@���)�vD�=��_�5B�;B%�9���<�[������~yy��Q�0�.|�lO[]�\\K��\
�+��
P��a.ܵ�Z��{?�܆|�*|�
}d:溓T,�-�AA���<��OX��RIE��크`в��R���-�&��bو�l��"��V����C²xxdπ ̰l���%���f���o�����Jc�s��?c|X��������(��cA4�ar����J����M4�ml!i��mӐ§:�ٯu���H��f�='���cR���Z���.Ow��#��:�B;~�WS������f���z��nʒM2��4G7�����%n"E��yy�d�c�Q$��� �P��}��G���������y]\]��Ђ �:?�)*�8�r?a�X��<K��fWN������g����)�<�F��*ĻթBB"�pKO!��㙙��.���ʤ�e��l�i(خ�����A���ߨԹ��Լw�>i�g��C�=|�����@�{�uw�Q:'K<G��	�/� R^��F�Pc���<�y��Y+��p��3�;)��Ϥ ���3�a���H@D�	0u�:�%ȝ��,滉7ˡɍ���Ȱ���#�BK�Pp�Ѻ@� 8�<�<�Ȟ4�frE�L�{R��p�&�@ �^������n&���%�������yy��*�n�7w.8��\������6
�j����kddT�`�v��y���a@A�7�c�VVm�M�	���o��x���7�F���~� Sw��Y�%��ж7qm��y����o�r`r{�,\����%
�V����c��2�E6[O�[m�.����?p�YH��< X��pq���A:H��O��Z�es�TX?�r a��x���A-Aף�����l'�v�w.7x"""Rޛ�@����ʀ�p��n���M�_8�R���D[�4%���L?�@)�K�$bIm1�"=M�u{g^���J�&E(��L�&�l�c���*kȘ葟v���D��@��m��F�(�%xP�r?�㼿��x�/2�	#�^|��ׯ'�6��77�	Ύؼ�~�3�m�r������骓VO��)V֎��ʬ�����Ux�a�����߁�]�'�B6q��$[-()����S�������h��,�����^���<"��o�ʌ��vX�/%9��˱3@"���tD
�ɓ�F�n�TNB7t'��P��{ L��/%�Z��ߑ^�؂������] {#��^�{X��\�Fx΍��J��f;	c0��x ��?�w��ϟ�a2|��`����yҺ��84�9#C� �I��۷W���VQ��V;r�d0� �È��[c��޸��VUa�n3]���D��I������֖@/�\4�K؆�S(�6��*�x�RC^�����D1��Pɀ83b� sss�2/ ��HA�w"�L����$@
X�F�`%�K?Xa+�J�JX�C��q��DpssC�TVV�&NM�@{x�VPP|43�^2�E���\(߀j����x�a?P�0�7��W�8�q�}��Pn��Ʀp���lⱍ�? ?�`B�\o�	!�(LI���խs��%�}/;��Xܰ4���-������\�P��b�.�FTF&n�U�
�L/��^jr��6���<z(G�A<<�_�,z�%�.3J�I�P��N �:��Ba���m&҅�ZzzV$�%sP=%%��ɶ$���p�27��U��&��0Q��x��VW����B�J0�23�@TE�`{��zmw���#� ���HK�����^CJ�+&��@�wi�ۂ��iiJ�(��D^BX8�%��˙��@�7;�S��#]jZ65X Gz��w�%��2���cv�U��M���__�g��T���6�� L�?";P��` ,���G��*�i�Gڒ�����qqp?���aA�S�ɟ�
UI��XlV�Z
q��uH����g0˫o`@H/ANL��p��=�a��#(0R�ٰ�`��T@!y��L�r����|�e'�ԫof�%����,�92b<��8���1`_t��񪦦� ����^<��Z���g�����wO�k-tc�K6����LtW�q�~eK�H!x9�%w�����&Y��nOG��Ȉ��B�H��F�l�_H>�� /�+�P��Y�P2Y��E(�(:DA%��R ��Qd`߂1*� �A(��e�q��_R�!9��!}�~���0l�
�Ɇ��ۋX��.a߳I߽o ��ȭ��=��m��-S��W��[Q|(�N�Lr�����1�(K{��Z��u����4�AQ3yI�Q�j��w�H�"yS-0Z(P9ЅK�|[���A%�>����R�wkO~٣|y�l��g���Ծ���t�`Z/�cկ=��U���������W\a�<�qp��a�����Ty�ޱ��Ur����G�b^�2���ֹ��O���^	ȸR;�} �p�W�V򨯐G�
h9�wu���,�z�,p�#�+��lTu¹8��jj	&j~o��P02oi�^R�Z��չ7t)+�G���š��Ñf�:�QYu~���n�8�]3a.v�UGZ&���������k�@����*�x
}���@\��z^*_�����4*	QϠg�c�_R�X�L�85�϶,%�!P&���R8�'��u�ЫW�Ǚ�O�h�;s&?�3)�j��֫Wc����ǘ��n�_Y"٤�:�R���#�L�HY�����\T��cv`���
�:��<J�<���ϟ&���y�h����;@O�w�;���n*��JS�qF�P?ф��c5?��?J8:z�N�4b��u����N̨�JI5���G�X^e��˧񛚚�#a1�)�8VDv~h�'x���#r��<��H��NZH�pce�`�k��ꨓ�r� cɇ�L[������� 3d��y����������Ⱥ��6:!w�e?������\�+,�[��K/�~$j�pp�<�)��
@�2�cϨ�`"�Zb@��o�9jhl7�c��>�����e'� Q��������|����2ñd.@�h#�8����<~�D�Ƿ��V�5ӧ�����ob�=��{A�*��W��^�-��VTF��gs-�K@���ʩ����Hy�<�+ѝ ��e8�E6ڀ2�����N{h|zC�-��z��Pz� E-6���3b���gu�Nǰhuwz�٠)	Ơ��dm��������:j����Ð�I���U�|!�H�kR\QÔ���M'�I�d [h�P�.��"����vz��6�!:S�Xi_�N��2Ӗ��G�����[k�����ݲ���RR)�s��?W�OHX��[hτ8e����4�����r�dUWH�U�0\(l��������F�%ÖsM�x~Zz�.3�����5��"�$�5���f�\�8w�}�a'GXXY�['��ݬ.��ṈT:�[~�I����jc�qC��n�L��,���> `���[F*�TKIiEF�]��>^~��φOL�h���D���������*�2�[��7��W�5�X�K����_�N����5�f��<� l���]4�'�F�I�g�$:�4�����xԘI��]ӚuM�Q��/�a������L����������E�Dfٞ�A���堠`k` �~Nj
����^�ee�$��5�D�z4�(*!R� ws��Hw�o��C:�fGT R���������5�X4�Р��#����Q��i�j�q֥�++,��]��/�={6������rM�U�x��XD) �����LN���:�8�$[WW�"�㍬>�X*f�v�q�T�@��n�ϟ���Y�����Pє&B�nX�}kVm���XE+Go������X���V�p�邺��*-"�?Zi���y�J��d��+�x2�%��Y���X9��c ��ڣΆ��<�@��7h���\dV���7�(bN��lh_�g3����J���G�B)����J%�~�x��������sjD��+��&�c�B�ވ�$8X�^W�Cwi{xp$�֑g��`(���AQKS'#�O��^��yTuG#Ͱ�s�"���p-M�E/_�����5��ε'�YB�x>��C���|c^v��z����?)�f�!�!�o�jo@�y�0�8�bicx��e��\� U֬d�)Փ��<�P�֪�Jߒg֘kۤ�I˦�JϾ��Q��m��Y^̗�w�����/O�Dc�[��,�na��:,�C��GS����[��o��Y�;M�^��±�*�:����;c)u1_o.�1��������QQ���%Ml��/��-TU*�~.�K{n�p��ȑ�B��.��Å����,Z�u��5�.L�nIz~�h}����f�SD�u-pu���XO���ڗ�(_����pA���L�C�]l����LU+�"l��������ѓA�_���	"��#���%��2�2Ӟ�JA�t{آ��),aT/W�,�������;��
V�b��RB����Tq�F�s��{�޺.������?e�)��b�������t!�D�1P΍�*?�r�(J�,���g�Z�=�����ɺU��F�~.�p%>�J���`o��Ʈ?E�¤%�!6�@Yg�"�jx��խ�G�f���Xg���}����Q�������	�2��J���S5���~���U�%2���^�����ʛ�hS t��*�ۖ:��*��ٓ�1m{_=�\[:"��bar-��NH�����ď���"���D�d����s&ǌ�y�t���v�66H	����c��h`�m�y|�~y��ܬ�oV('A��>=���"{���ykc�fD�Lji�A�o4�c\���kn�Tт�4���M���4xs��rx�4r�Sc���Hz���!� ��]��L�C�O�^W����b��㛥O)#��Q���9ؑ��Q&�ӓ��s�bģ/��e���"ɬ�'c��m�%�a���l��wpbS��K@�&��N�gD�)�w�k���V�z�/z2l8��R��W�M.�ķ�����'	���@Ȟ��8�a3{�9��ۋ�M��S[��-�WKǵ��y�5�_���P�Zk���VYi�*��W?1f���!��*m��3�q1*_�\;�ؒEg���X�:7�q���/
sH���9ѷ�\��6V\�p��Vʪʓ}����ˏ5�i�NIW]m>�� |��� 'N����sԃ*�$N�<�=b�;nkg��x��1�<UuY�X�V����oDӏ�dwť�pڃ?Q���Z��*�4NB��=��Qǘ��4�Tš��@���4�}��H%S�l� �l��lO&���њ��	��'~s���Ri�|���C�w�37�$�C���Td\yu�_��L����$3YGL��C���� �&g>�.�����)��&��0>�(�⸓���V����XM�+�+��0���5�&����Vg>y��o��*�[k	`�=��_����W�N�,����j��O��CT\�����Mwl�=�(���%��>��I��s&&�v�I rJ��U�e�k��hT��?�(��;���n��\���6[G4���z� I��礖[��4,�[�;������<��F�&Bi�.Gww��[~����0\!�fUŃ�7v�T>2���Y}�i��G�:�}��=�P F_bT�1��+��}]�i���,:�C��]b�����c�^�^lޑ�/�.������G���l;���4xm�6��yF6�܂1�}�@��-ik)�%/ƍ�#���O��S!\��썔\�H�Z�D�wG��/ֺ�>P����Ko��"��v����z�R�ԸH��D����%R fx�x��6ְ[,����ۢGC�xA\<���[�at@A|�EEͨ���_S�@����e2���l�ӯ����;�;>��C8\��5s3� �R�!���ܜ������_���w��}�:����SL8������Ot�D ݗS�
�^��Tϰ�2�w
�9]����T;��,P�Lc����,�BV�2����I�q�իW�o+&����b�4ClR��$�"�?G҉)�{�r��{Y�o��r�������IӘ��:�Y����Ԋ����
��1��R�@,�G �tCW����Q���)��9'�e��U��F�IQ��Mܳi�wnX��P�����T7�O��؊4{��x����qn{K�J�^��y�Å45Ӯ��:]U��Eg�@'��W�e'�l��2X�i���-杙��ۂ������9���[;N�u��}�:mM�E�"�>Tz� �����PD"���S?Z]��IN�W9E7��{nn���'U�
=�i>�J�
�����2�J�&�9�'� �J��a\o��O���y5m0�&� ��7���7JJ�p|���8P=V��^z"'��п���g�`�`%�(w���%��W�/*�",�rqQ�?��z&�ag ��ͅ��k�q)'��h�µ�f�5һ��K23��u��%[������|+�5p�{Q����7d232��v�v�/���[��)/��l�잸*�βQ��31�;�@J��\�@�5���ϬՏ�5L\]v�Y��ز�9�B ���Y��7�61���D����ۭs#(���
9��S�.���.�;@�D� ^����w��=ȱ�:$w��V������R�=���hص�Z����IY� �h7-!&-�(M�(-�(M�-��&�v�/*Pb�Ґ��C�1��^/'m��Њ{Yn9�d�����LD�R��R���/���w�%���1l��2]��'Mt9��k��n;I73�2� ��/����S�\f�x��_�]�M�������ȕ�"�l�$LS����{i��ɋ"�s�;���Ҳ��m���`0����2c�(�,� `��9���-Շ���������|�+{�ό,���9���N9$㞸t-�n�,�P]�zvv���W�	f�I���蓵��)����Ӵut
�?['�yb��hh ��5ͬMcS?����͎���K>z�S4���˞z�X���p�<�w]� ��5N���/���)�8z(��1��V�b�7YY�Q�B%��ea
�uɯ�`h�	�]�CT_��~�� ��U��Ҧ^F㫘
��h�$}��V�o���Y&����=<ܒBl�h�s������jk�^X}��C��_cA0Q�gK��{���iOZ�@���}��aɖ9�^\�p�Wc�P���QVV��	->[��(�|�gB�#����	�Og�����b7�ucгL�+�9��}�)�T<��uO�bN�sB��Xl�ᯒ��/o����1%�m!��
��;��[ȸ⧶�7]51�on=ۘ����,�Jc䳛Ӭ2����z�vR'6�34�;٘ +߂?5�h�K>n)�I���U�"�ۡ������<Hy$��]�?�b�*�V��/�Ԇ�G���4���#��/�đM���$x��x� 2+e)Dqc� `�j�� e� i��o����럞dm�g��Txm5�Y8C;�/��
�fs�Ԧ���N3]v����+�|V�К��s�<1��[W)�rv|ثG�ir��<1��~?��q���z ������'&��K�H��iӎ	tN�<���C�NJ����B�#���qx�l�:���W����Qvz��}��lE�~x7��@��d����T9�R'v��5�x�ڼ��1b��sҳ{���0�SA;��ʺ�Y���o9���0�W���ӷ���w��7�-滖{e��%&�� X��"�;���<���p�g�H�v�H?�->����.�o�ɾ��xG��RrTǫ�R��`K��8��u�YI�)F�9�ff���v��������q��,�ʴ�N�D��R�qW�y���>���r;������__H3����:V��4�ބ�~���6I�dO�-2$M�����RN��.���B�U����w����'ؓ�6���Q����zZx�w!vn�*����s4�v����fD]`���ä�s��%$o��zqf�?�o�`t�n��f�̅�5�U�.H����!=5!G�"6]g�"������o������^h�{z{~T��d�����T���l��3"�/����,�#�Wz:�Cf���+ր��k�1���/�n�,,�3*�s�ڗsm�--!���U�<R�EM��Yg3��Ɲ�Vwu�\/�#��/��B�trr�'dǮ�m�/�.R1�F�b�n^,������4�v�<����8�#��x���c-�d��k�4?\ln�Fk�q���|?��{���|�������P[�2�d�s�����Ǹ�_vu��`|%��`�b|IK9�>��`̵�k�*��TM��?.��XЇ��"���±O_T\+�c=�H:�N8���o�zSN�����\e&#�����.��(oc.C�-FT!�[k�D�Q�Cu� S�>M.6�/�Nj	*)�c�y+�fљ%)+�MW�bW�f'�'Q�S5H~0�	'm�j����=��[S������l�K���mOr��ƬV�nJ�vdA$ZH���@G���T=.k�F�K\�ƻ�d%}gV�MԖ���S:Cm5�
��n=�[��9�t�SNM�gнYgf��ga:d;B�;��%���b�=,:f��T��x��1i���/�LFE��_��~������?�}`����0 ��3�v���Ng_���ם�y�ʜ�dZ��cF�r��bP�@�����@�0��~0�g�c/���h�r�̌�t;V|�o�U�uq������A�v�zc�u�4%�P�!G#��gg��d֫��"Ͱ��g
!؉�li������+���60�k�3���gy����y��`����9|�C� z,-W���W���H�I/��`;��?:n=�3�e�h�1B��z���`NY{��6�9 *��d �`�֖� �Ǜ�h�ء_]�`vL��g)��SVL������3P�.��}
�ea�A��\�j����n��`��k�J.<m�	�6������Ϩ�؃����������'{i`�����өy����;��O��k���8�s�f��8��B�$`/[� �澜C��h��+\ݮ�y�N�Rp|�����xjwt+p���W8y��O]�S_����Qv^ǣă@���<�1sU���ypg?��Nޚ��$�6{���v�9�����u�F���xI��hifZ�]dpP�n���i�1�R��G=�:N[,���β�q�����a+绛kg���Lk����<w���<cc8[��;f��g�v�8Y�.,��(&*���j�5�!�D5J�l�_�~���﹟
㓀?.���3Łu+>L��=qJ�
Ӳ�޻�?e�QL�+��a-��әҢ烵Y���v}�4�`��F'J��K�S��*����8?O��.�������2k��̺P�D̔�P~qqZ�EUb�"�I-)^YzN9�[4�Wb(Ki¼i��}����=TVt
��b�0Q��,�?��hc��\85��c�J��M�*uވ��"��h����^����� ��#ƿ�߭��0yasA?4�"��y��Lp�1�t��|�M7@.������g��#�fL��ڴV�5��
&�/6����� ����9�՞),D��#`K~nq<��N�����=�Q��r��3�cH� ��v����f�E��0����3�e��<�nK�r���|CߤO��_)7^wI�j�T޷wޑfπ	,�9���VPP�@���]W0:QIOwBE5�t�ǯg�,��?�d������Ga�����8���������j6ݸ' !l�M�'V��J'(6z#;O i���δ���q�̀��j�P���R-g��b6)nҐ�KC(�e{Պ�7��������i���L�6K��y������)�g��f�����#'̵Fa��q��@���-�P�����a���q��ȇ���u����8�T(�f4�d�h����R�vܒ	�Ɓ'}}�v���lAR�F8K�D,���ރ EuN&�4�� ��72YN�ӳ��֜�e�)+��ĝ���l��7���1�)(�7��V�}����,jy�1{����TT˂����W3�-��9TT9��D
A憘!^c�Q]����2�`RI�����F�8�s���L��x�.��";Y�;O��X�Q����t��v���'�J3�b��ơG$�ZE ���p��E����ƫ
�pٝŦ�&�z��kٚ���{3�ן{�:��n�j0<8r��}R��K�n�4�P/�Z ��yx8�D6#����3��+d��T=d�G�2���^c����8�P�u�E l+A���z�Ų5}�C]��ʋ������C=��oő]�����2���\��xЉ�f����Mb>N��P�������e�C^�|��qB�I��StH�9_��\A:.�kR��&s��0��؀���Fk+��9"ɺ =Ҽȗ�h[iy�����je_i��l�����F{�+FH�*�9��^�iŬɎA+��$�h:x'��f++��U?�v���Ii��������I���Ur"/�r��zfM'�IM4%���e��jYҷ�e�7��q%O�Ctן���%.pCr��u��>�B�� &	�T�G��P�b�iv�����\A,�l�Ȩe�n���1o��}6�$��t8[�e����{Ϣ����Izr�\/2�"�3ѷ`�'����Zv�;{����7����W+��%	>��?7Lr�X�!V��g�.k����&Cfe�v��ۮMuK\�����Uq�������?���x�B�� a�?1�T�OL!�Uo?���MTU�lA��Y0�`)ջ��ie�o�!SV���kb�H)��Qs�D����ª���kzm�_z$+I#և��W"{����� �e<3��8z�(\�:FM����Q5fvr�����QK�tA׮ )��$�c'a㙾������B��������Ѱ���M&���{|L��I N*��n��Te��@��ʄ|\��rj�y�	��;�<�]�Q�1���ǽ��JpWۻW�$NĻ�.�,��hx��Ӑhb��HGJU�*�Kkp����g\���]8�I�"��������t����y�i�ػ�J�<��y�&�!�p�*+��BF�[a�v�xz�6���/i*��Tz_�f�307�����P'�V��63�ʳy��S�Oߓ��"����#���2���kpv�3<���3�:T�x�v�JџM/����A?À`�q#�E ��T���kjY�z������jI�t�*�>\d��
I ���o�3x��_]��B]j�-��УZͽ��ٹ���,�R���]�f�=?^�`���<���ߨ̓?e)��R�''����,��u�|���
f��.;�}�_���J�VQ
��yrFT� T���͗�X_<ͶQ�oRà*���W*�w������x
�s�&��	g�M��t����;7�!�R�g1c��n����M�F�����׾&N }r���@��i
�Z�x��N{C�'1`���Ϧ�95��Hym��<p�ј��5�/>�l�R�0�3c�)ݨ�Ȍ�<�� �`�����4 nIea�?�1`VEX�ɴKL�b=�]���t{RԴ�=�r�7��V��/�#��a�?���c�`4�����ܽ8ͦ-̶U_iS��2�&�geLo�n�g��Ee�����9�0�J�&�'B{��=y���Zf
��2q@T[�Z���lR�j���;�k�ǻ�dߗ|#s)�f���ꆪ���O'�m~��Ɠ��.k�jO�)�:��������k
�P�'�G�<V�ÿ� g���y��S��SN-SK��-�@��uD�W���5Ͷ�?��FW�r�Z��� A��c�6��H�T��Mʯ�D��a������͸���)��IQv�EH�ՙ�TpZv�����[�!��7�)O��
O��ʯ��x��u־�T���`���o&����������]�b�ȵ,V��Afw�o�!�⾮W��.]�
�aQ}���(S�EQ��) 5 � �����B�մ���

��?F;�:)y�Z�֮I�Ƽ{����&�X��ĩ� 7>�Y"�k���9L |�c�	ƣ	&�)�Ƞn�������6���n�Ɇ� ��ȴy�X��V�@�Gk5�)�L�¦7ަM}�c^�b�K�4�m��)�[���B�z�TG�Z�о65-�01�����Hi&��h�a�iB��G������Ezp98r����/9t��VL�U��������*D�Дb�9��7��=��69D�g��_��)�̀-��:n�!I���B�Cj<�p���s0#��9�.
��/7�L�}��Q�M�*�G�c1�]&(�_'*����-��{NV�o�@i�QyPN��o$��ef15����ӫ�M�k�
����s�Kmg��L����!S�4����"%�ͧ$!,I�
�I����Db�ru��=���g�w@z^0]�� J����>�c�B�+�e>?ʯqFw���[�ϖ��fژ=�� >-�G��S�W��oɓ&����K�`�NX�N���zRP���9�c�J���\���>R���;-Ast����wx('��Y�;��v��}�0A�s�ӎ=�r�FJ�S1�QO�br(<�S1��ӤR3����X�[��F�[�H�X��7�r'���n��`��.iSL���r
3%���w����	u!C��m��ÿ(4������pz��0u���gJ�F����R*�M��M�x��yk�j
q�݊��h�Ĩ�qV�����^�?Z�>��5��":��,I�2�۫�w�ϾT��A'�)H <X@�%���l/۴a,�h"l�VUt�ٰ�c:�j���5�~攐�����8>��[���V���	9�W��_C�x}lz�Z�8� /��o�U5����"���j�*��	��9�����6�j3�u���UC�mZ�B�3�?�V�9�=FwH�sڋ	��`Z]����ȣ��ڱ<�lt����i_OO+��"uo!��.��Ƀm� �K8#k��f;�{s�|j}pl�sX�JOM@��v}�
7�2�������K��c�[5�)�򌧜�]�������S!~�Ie����#8�p�sUaLLL;XY�n�x�0dYC��
uo����;T�d�m��l���k3�CL�5�����Z)���.�o�k� �T/����m���2���o��]�UqUa��T(��{.KAUV�<h)�l��E9�R�{L�:O~x����A��Y���,z�Q��[As,���O�o�
1�Ƕr���W����v�>pq>���I^���uLP�}��ѵ��������[��_��|b<9�Ҹ~bSyB����t��VF�`������,��T`���r�.��igx�4I�}�SA"���$�rg�� ��yUL����7�v�M� �����S��ՅŮ��%�D��Vc7�nKS�l:�jLCD��p�t�
�hpX�J~��Ì��C����<oG���u��A��/j��'
*|��L�E�.F�JA6��f�*�.FG�~=KA����M-�L�{�h�}��/�y'��� w��|N~ /�+ϱ��	�vn�M��	��9W��mzӴR;�U�Pf�lLJf��n���H�IT�f��0c�bBb��>f)�kS�c���,�w.�U��	9�B�:�>Z��w#̀@���b�q�E�M�J]�c��l��gչ߻�[��t�xٌx�{�M<�UK(т��1���8�2��G�$�:�Zd��Iz��T�������,�#��U*+=���)�j(���]�LH�o9�0�̰��Վb���� ��A|��A��}l�*�V@ ~w-[,��tFִ?3���U�lz�����:��:������R����$����D>���zN6A]�
�^�QIЇ(Ed�Y�aRS�i���7u�ƙ�5\\Bb��?kve<�Ol#�X&�10հ���@!{�=A߬����}>�m!��H�y8}�<�G�a���	-���熛I�^�1M�-)h��-�3�-��g�5�5�O|I#)w;l�� ��?u<��,��~Ӛno��E��]���� n�g�#�WI��������Ku�
���\Ӂ��I��i�P$I��뤠��;@,���8-ױ��iJ�v�Y..n?�:��?6lo�4�e\�=�hͭӾk�'�&JU�����6����!/�q��p���,�NG)"�<��h��������#�����jfh��Jf�l*�[!|A��� �*�wS&��>����I�x���tg���f�k��w�[h !��:��O�^�9-�$7J6�O��v�E}�Bd��hB/ƇormR�F�&9�G�<c:�ri�3p}/f�4#�� i�*j]��YX}CC�Dٳ찲L�����Z ��ʽ��Z>o}�Z���orr�i�!i��\��ߘNмD������+-�: v/�m�H��!A� �X:�{�]{QF��BO���-�u����'�U����7�RVF�PC<�o��k� ��ş����Wk���D%V�2�{ Bd�I\s��R�F(�Ó[��� ����7�L�}�nq�y<|�i(�W�i��������g\�����b�+��>u�����苫r̓{�ȵp��&��� [^f��S����:��$2��F3�r攺�����}7�R��1�G�����y���������je���a��#�8(M[dv>��s���*���1���ǘ�vw�z�L��ti	�x4*�[XNc�u3�M�h�Q�f����	��;���%�o�g+Emi��H��|���J��H��p���M8���a�G�k�C�G!
�����������~���Ht{P#����V�|F���䯑�R�|��[&����%�Y�;	6��@+X	LI�� �_�c� ��j�q�qFKrP��_���g��Y�������/M�ca'K}�����u|��u63������ݯҋ����^o~v�"{p��w�ɞ`b�$���	��Y�lyt�L�Y�d=[z#]X0"�>�S(;n���a+Ol˪��=oAp?an���Wt�+���q=�b;�Э���TT8KI���Ǳ@���3v�qU�)4��o��n�c� ;��-�\�j�\��D�8}<��d_ܴEURP��\JW{�4���U��=�9_2�RK�@���������j�����ɦ���,=m#�����m��Q �3�w5�o����<q�R����Y�.�L����*v,�����h%R�a���6����Z�E7#X�mZ���.��p��Ն<�4�ns��N�!�0�M�`Z��0^�0���M�r� Q��n�������������ox��D��R�z�B��l�'�z�8�.��ND���z`{[�hoYd��
�1�=���/��:���M��R����(
��BM�D�$�%�d�5M�B�ވ�gYBeI�d�ٲ���;������3�y{�^�ܳ<��{_��)�y*B�f���K��������F�l���IIIFj�ed��߱��ח����Htkcr���X�^=�e��.|��� ϐ��e�ofX��Lz+��x�s�b݂gF�%��;<�ڵ��*׮��H���PMM�!��(J��Wod����0����o��&k�^9�?���Pc0��{<�\g�,��W��}�Ҫy�c��j�ո	�lƑZ]�u��n��Ƙҋ������>>uib�1���� |���h.ޯ���y�V�鄔#�I��r�u�᳻4D�t�T]k3;���������Θ1���v���ҥ|k������Y���u鴤۠4n���b���%����}�z�#՚����B���� [�/u�.&&&Fmd��}nӍ�T��d�l�k��4>Z�޲�%:�bb^$'>s�v~����������T�.��/�n���ԥkH�~�������d�	6�#_i-j�di�L�~���9�PR���࣫C-�&3�dŗ��Ō����Y��1���.���\�LS?�k��K٩<�N��h��z�7�Y�h��o��M\j|m"��%7��vJğ���y��Y�ً�n�)2�;��������"^7�:������g<�F�q�)~���p&�"��'�Z\��<g�6��1�l�����J9S�n�����W6�j�Ƣ�j4�_87X�LD+���tkLOO4ۅ0��y=�Z��s���t:`�m:��t||���=I�Ul���.�����_��s����ӓ�����o���ï��ދ���w0G@�.���{L��q���W�D(��=�s���/���=���];~6��N��/w��U,�n�j�d`⯕��.�Q���r�{zD�����9Y�-vx��z6 �%~aҚ��9��RJ�� _0��|+��c��]Z1#�w����5L�Xv=zd���B���k��,�v�P�Ն���v��5�w,;l7����*7#������q�y[���=����[��ol��X�����F!�4���*�OT�;����2��ܻـɩ*ߎ~�H}ˋ�]�@\J�<��·� Y��J��wzys�ߟ�ΎU�d�<rƦ�V|��]�j���dq��i�l���u#:�����M�ͫVX�V��Nc��_�����*/`��}Q~#X}��3Y��f�l n�����w]^4�o,;�`�_��6)8�:����@�L]uL�^���/Y0�J�~����y�o�bzƇ\/>��� ����=Lo��!.�=&�-�����+拄{��Wy���H�o^�`�ӿw�8~�g���6�:���/���Zt�*>�\����*�\���:rݰe�|����c�E2�j�.	H������ᙙ�/�}g�9�M�/�t��L��,�En�2���;�&!�c�3m��@�v�O��y�s\�t2�o�a�K�2no��-g~u>RNf^�������m��y~hP��������
5^�������%���/�S�%�r��mL28��-�_S�-}`5���l��\��sms���#w,��V�[V&B��Kt�Z'd�c��@QF�Pѡ���?d:�?R���Qxd>O,+��k�[L��x�8���,y�n,�h�i�!����~�����ꐐ�f�a9�n�yќ���,K6Ez���ױ[ ���
�\�xHm�Ȼ%�

���q���vC-�w�`�9�������(��)�k�~�L��|c�{g����?�׌��Ͳ�O�j/�tx�����=T�	����F-ZC�9ӆ�>���Ek��ۜ3���-�r��\߇aןM��\G��au�G�-�7��	d�ճ�ۏ#ڿ�i`zd��ЏG�wx��άʙ�'& 	��#�k=�dr<ȱܠL[�*=ykD�,�@҈۬�����~Y)W����.r�,�낶�t��8;���ZɆ�S��^[!7�'��?7ƒ��a�V�.�g����������ٺ�+mQ�v?�8�{�;��}�ï����*�X����W+3�W�i�l`z�L�S�%wy���������7:\F�rOrΙ�Y�cY]�A��%�IF3�2�i���<#/h���������Zﶁ<.�o�s�jD���SAY1;��s��f&�����"8 �&�*�8�rGw���Rg��m>=���]�-�-O]�9�x�i�SwG��ɱ��(h��p��Z��%�xf�~Y����_ڜ�·�bW|��?�<=)��]�Z[��M�,�"�BdɫrEO��aW�>�c�� ���Y�_�.��:J>��z�
g�9����tk|�my`|���\c����-��ba�M
W(ᱶr�cꔹ�7���S4��*� ��E�N1ky������O��>������0�^S��yӛ�Lҋ"_@�zmj��D����j���_[�V&���}}�.ݬ e�쥜����?��h$.��8��*���:A��;G�\�g���K1��*�U�w�o��f,~����Cf�92�-o��;�q��R���(��e{�E#�k��*�ҕN*]��t���9���,��x���&<=/O���f�]��,;�t�jHB��G��4�>m��O��"���HZ�,�]�Ƚ���v<�5##���Tt	�e�6;5^g��\��r���x���M,9�ԝ?1�w���B��H���RR܍��Xa��8�����������{m�m}`xFZ�G]�u��,�Vqu�20)�a��fYܛ��^��,���h��{F���6(���Q��rؙgZ���DH̓C�a�]�R�t˽��Ѿ߮�վ�O��E=�y�2��1���1*��:�#%�����6E=1(�$���~��ik��3�|�@� ZO��/�[�9����չ��rS)cm�J��M������i	�1j���"����of����
���14-�Ѽ����8v&?Sݚ�n�%<�\%X:@�r��X�%K ��m~Y���q�wtW����d�/p	K�i�c�4~JX]�>(d�ޝ�5�~W(L3���9�X�dĉ-��ϲ-��:9'u��p?X���Af�
I�'I�'ܷ}��(��`Luy� ��d��a���.���~4[���aE<|������I�vF�L6�:K�9��'�@�G����/8?�d��V�&S�Y��,	K��@#�4�0'��k���u�lw�	�[��}ť.s��GF�x!��S)t	;SL�V����)3�i���g���OoD�/hL'�F�p�xk~�A̯zg"����z��3*Jp
}z)��Ѣp4|�ڋK�w��S��1؜E�����`j0k��$scQ���@i�S� [y�s�1����5Y��|����(��H@����J����g�r���鐇`�bo�Q��5G���p^c�(����h� 7!�E�022�oL�����S�?5�S½�k|���i��`	��;._Xf�WVZ����+��GWY��6�B��ɓ�z������i�o����x�8�/ϼ9�}zbH����г��@�x�1Hr*2/���O��he�X�$�� �ffJ�'����h-�(���VE_���"��^É�1#S�*����>���6Z�:�.�,gn�o�g�u�(�Ýa<x���d'��lAJa:?���%���j���_ @�+�z���'�W���gn��N�(v��$��i�O��W��9���Uֱ��׵�LRz�L�SR�����u	T�-�5�w���I-�9SLФ&��l��`��_rI�4��+K�y:w����K�kρ`\i����P���p�f۹k��:��i3���"��[���W\��H$�3^Rv�Ȗ�"����&[���V��n5�
����P����m�	f,a݈!sƟ'�`���Igf<���$�"(���{m���7���[�(�4��_�c�Hd2rt��j���6����S;� ��D�H���G�=8!�+�!���)֜��Wn���J�cĥ�<���̕��x�^UUq�^� xD��cl�����r��>�����[�)�;Z�}�m5l��x��]�:\m����|���z���H8�OE��������O��n	�~m���	r7�E��5�>&Wc�L���JR�n��rc�W���u��6�/6��С��ڨ�3�;@���#��2Ĉ�A�J�I�ٶ�6���aT�UU#����r�>�sދ�	��vt�~UQ�v�A��?���Ul�qLi��6h��[�Hv('���%�_A%	��Vy�:!��[� qT��ы�E��8�%XE8 �E�;���Ȅ�Waҿδ��;��cvf&�_�H����K����;R���V�6y�NOѵ�Zl��{�Nl@��u"ٸ��U��샲;��o��hGx7NRU��V�P�HB�]��Q��Z/��Rp��Ԏ���{r�W��㾭���Ub�B&���H�!�����_��Fw���t��!��l�)�+�rg��R�����)ہ<</�p�ۅ���o��*�L_t<���"nU���#I���w��� �(� l�����@_�~Y�y����Zp���Lk�S��Q]>���=�8��~�צ�U��ik{@&:��x�h��'�����=Z.E!�~Հ��3�[	��x� �$��0��e{����P��ޏ��'�g�5R{΢��V����8�
�=0�E�:u��X{$Q�b�^���S�!a�t���n9�k��s8�NP��lB�p"�3� 8�̔�llB��B�h_'��IZ�+�dZ�a�NB���-��h��.nt����{�����"�:�Y%�8���0�]`�/���5������{�?��)W��g�h�b�ȕ���@�h���p�u� qm�W�Q�b���;�	&�?��J1�P�+5�YMU���5���OJ�m��Tay���������m��<M{oJ^?��$��t�%�@:ݛ.eG�|u�CT[8T-��9������<�.���T~tو�3Me��:�8��G���i��`����w�m��٠�>A_����R	W���&8��Q�eM�� ��γ�u����U@9��u�ƛ_�hf�*#�����h<�	@%�*!7��-�d=������T��?�Q�6����n��qzfB\��W��D�N��"�}ޱT$���s����bBP�UK �����.35�`�dީr��w��h2����EP�?�_ߘ�W!�,�5!B9l�ξ둹��E��9�9_z�l��@}���y�C*3��Ӆ�ڇ�/�L��#]����[�NAݺڢr�=�����7�;��`��Rs=;�H�4� k�z�E�U���x&a�G4�j{~�5�==���J��?	�����q�P��\ߦs~��v�C�&%&�'�~n�*�C��S*k��uN�[iЊ���AO4����H7`cERCُ��It����o���j�����q��\��G��FiA�
��p��({�0�l�ך��@�d9�j�
fH���]b�l˥48�;�]Q�u�ŏjG�ȷ�ŏ,;?�$|湚?�y)�A� �|P���"_�7�Wy��W�@{�[1=7=���+�B_�k�l/ ��Ϳ�*<uҪ�#}��Z����R�x)��E�yL,�Dx��g #(V��h�������T����6XHc�~�S��	@j�:,���/J����E?;Ĝ��;>}S�:ؔ��+�
F��rJ��S����k�i�����m�W�_��lGF1]����o	�.eR��">�������]���� y}H�
Ņt��wKx���{�Hl��Z^�K�I�S��i����*�L��@�5�ހcV.8�&>���E���;���ہ ���*T5�	�-z�`l���Q\N�7�n�Lz�����@����,L��Y]�:M_��2�y&�b�a�b�ؤ*7��${6��X!�^��\�H�����"\+:���m��f�n�sl�L]��F�� 1-?֋��xl7A���ȳi����J^5�� ����$��U$C?�r�w�oL" ��Vޑ�C�m�Q���t��_���`��YH�AM���H['ʥ��lX&��x���Rrc�|��@�Q�m�j_I��أY���B�= ��+�w����7����e��}}�~U���F���4���l�4�@z,̰�g����H�17�R�_��U�Y],�9k�Fi���JΎ(�^����#\뎊�B&U*@�M��O��[��̄#�*|����ͱ�1f)$�}8K�J��U~�5¡1�o��^���;��;�@����_r36��ƬAA��l�e�2,1�K	2���C�%LuY�7Z� �]J(��d%ˑ�PRV���}5>�"dJ��"<#H����WD����b�W�M�&vkm�g�+�L�2�T-;��5q&���N��D3��vg�T����aP����bc���0_oU�cD��j��D�qe�v�N�2���n��/���V3�HG�����f]�v虜�,2R�g�!�'@KE/�?Z�B ،�<�&�ylT�i�t9�=�it�cEe�(�ȭ�$ mF��졄P�[5�gF�a'�Z�q��Y�ϳ�5�o_��ӥ0}�Ɂ\�1��, Zb� �dL������*�4drCqZ��w�[?"�����.���j��'ٔ�h4�����Gp�ȳ��[t���'>�g�����魮A�L����x��=�҂�1z�ǳ��{7�� T�,D$md;/2?�]��w�ژ9D�����觗��l�gtt�x������-�>'((�$���n$�ð�"�(�]���{��0߻ʂ������[�g6e���ת��&T��Q��`�8�[e	�%,�+��񾺎�hu����Hv/qP�£�|�
�C�M%��[��.���^6������Ծ������QA�!8`���?P�ʑҲ��y�Unʙ6/-/�(w��$K��G3�٨���w�v��I̔MV$ e�0�H'%�L��s!�$���%ؓP"MsZ�^�ƨ�\�G��1�"���R��BUI�V����XO%��r!�4�lݿ	'L�����_���/���d%<ܞo=8�y�+���D���񮝩�+L������Q�ǳ7��`���v{�`S�x8K����I��@��4@�r�k*�D>��|KX�fV]p?���6(� V�T�w��M�CI&� �Yv�-�,����i�.�<XS+�Q�* j�D�8�G6[�����L�"~�pZ�`f��{RSf�+N|`Ү�W߀O�(�%)k��[ۃg�6�\gF�@/B��̞n�,!|�6�����%ȱ?���Q[k���i�T���������>����� Ly�X����"�^��R���k\{ .���� ɝ4�B��&>���}⸼�/4v�DF�����QZ�5`�r�� �#�;e,�� 
��'jD֗�O��Db���*X!{�hL��bv��X�RŹB~�B��2?񐔼-1O�'Yf�B{������0�;g0q���wl`r��D��;�l?�b���Ͷ�����,vV��9��\<��r��-��R��د�qߩP��j���O���>�/�1�,Ј�M�&� )�)�ǧ���ԏ��4���j���h,P�O;�X�wy	Pu$Yu��ʿ�Q����=;F��WWO\O��y?���v�$ڦ:226V7��F�Ȁ�l7�fLd"�r�H�ҽw���m���-�6���{ ,��jv$1\�FZ���
`��Ϳ�sIX	*�8��s�˖�N0��ig�D�ς����\MT ]�nÚ�x��v�anO�����ݿ�x�>�T�X1�@��'\_2��\tצ-���Hd���h����喽_^��Lu�����͚���0\J��~�9���7��&�:g��S���3fgj|�fNA�]/��q��{�'lv,t*V&X���߿�hI�w�_��la�U�����#��6��${�f4�&dZZ	�'`�N����1l�����"�J��!E�|�5��FFۑ��'�`ɀ��Z���4jPfo����]�g����������b�5��B��5b����[R'GM�x���R����&�0�x.���h¼U�?K��^�>�E��އHzh�#_�Ep}��p�6�}�S��I�N���߭�&�������8�L��uI�a�5M��~5��9.$W�w�-�Z�t�(���4P��·���' #mu~� ��s�]�$/.Kފ���W��qS������Y1�!�8��W�v�z׀j.y�y��W�g� �n�i��Ͳ���V�x��=3{�G�ǰEZ��0��l0�jȰ2�Նr��2R_=R��������@c���f���ysm3*;�w�災%�on��*\nPF�^��]��O�" S!#��8�h���:w�bx�
i�_��]N��	��/yksrb�%�	����q��
~{Q����Q���ݐAmX�a��?~v�`�L��wF Q�}��A£���;��g��6��A�Y%��e�p�Q����k;�$a0ʢ:01��`}���b�ױ��Ó��~��@���K�$Vs���>8X��M�X�&ڋ�LOx��ȝ�O%3c�}�-��I@�S�bWFt"(�e{o"������LKpYٟt�X��T��ǋ�~�[�ل|����+����3����U��"����>V��G�K6�)H��h�q#��8���l��ɩ���*�}:�l�dD[v~f�hm�au�{�vG7���dS�b�׷N���k�P�xı��r�tjD���>��G@���˷B�^��2�F�Ǔx����+����� 7�7V�٫f�y�@�h��/!�8�;Q�}��?/�X&�6���>߬��Q�#h{���>�wWߊ7a��ގ�rTL�@@}`����4Ǔ��I��:v�=�n^@*K��*!`̸���+xӪ����b\�M��	���x�>rc����F �#E�6:	vg��DLKV* ����+:W��vI!ԏ��kWi�o9�C0<���{��BB;o�:��O&C��9�홹|��k���զ7�3��b�V4g�	�v0�(�j��OQ�ݡt�+1t3��$D����h���� ��8��)�tVhcϥK�?ho���≶nUU�p"�F��k,	+q�n�z��:��{���mb���5�f����q�Ӡ��h���������Z�����,�h��%#���l���!_/p~_b��j}�Q9ܮ����s���)�� �u����י�rX���)�����ҟ�?J�Y��0)����<3理u�I�^ml���y��^��n���'ˎ�6�3��8=��P	_�f�XrR0��$�}"%k1��42ĕ�n�	w��dA]�Jc�_�P*��3�� x����'G�8�x
�}rrC����Vt%e�
a8�r�i7�`��+�-Y��(©49:�gK�ݐ�,Xn�8���R^&�lQ��.c�<�7l�28�6�C�O���| 4
��������;��
������4)��:DM6�n��z)�A>� �#bv:��ΚQA���eE�!ޗ�AK��$�����i��B����eSު��''>����e�Lj%�?�A���:���Ew��/���Q���]����� �<rɖ&�& x��ߚ���b�;����Xa��ܛ%
sB=�,:���ju|� ��Y7�:��-�9\��#�2Y�J�o�@��$kT�����������y���7�$~�jH���&��F4�_v%`����I��`JFת��T-�਄�9I҅����!��'�m���ī�)(y4@��pV��vk����/U.��;��7��-L�s������p���C�E�W��Ԑ|��F��QDF���"�����H"�w؛�M���Xh��Q�/�?���e�t��8�F,h�����"7c2��"Kִɡ@=;����� ���@��t�4�mw=�r��1�V���d\���c$��L���dg	p��_?Y1,s4w��7ٍ�\���g�Bo�-5c�nr��΃(��i�fɺ��WTdj;��L���*����ȳ�+�3	&d�SOȷb��4�}B�j!;�]ƨd���e�,�y�2Nd3S��.�9��_�:�ʖcg�-�W�{�#6�3!6���ur3Çѷ��y���FJ�`͗k+�i��z�x(9��qW72V�n.J�}�1�#�&������g����1�p��
�i��H��¡\~ҵ'^S9#/�Ӝܯ�8���Oӿ���ʳ0w�Tl���Ti���������w-�¼����MR*w��H���y��Po���V�&�^�kK!��j�h��-���&�^��N����k��[g�E���sPb)��,�!^���A�O%������g)������!%�󀾴�����VPk�?_���I֖˹m,))i�>��,�טq״I����;���+�-U�;�OC=�t���|�O�z,�Aޓ�3�$�_��kW���S�]f��?�Ĉ�(൏�����8�\��bdo4vC��H��f���7��gR��o���7$�O��T�S��9��!�!H�ɯ��~����v�7}��p�͙V�*3@�`���8CJW$���oN��m��r�{�*����ߓ���P��<�h�� ���N"o;΅h�{�9��477�
��O���H�N�A��oM��2�ID=���/L�������`@vٮ|g"z���ޚ�wDfw��;V^��8��< �q���@���X��ޞ�����󘗒c�~_D>0b ʕ��P�O"55��q�(=nj Ge�v1��t"�Y���TV~�y	����
��X����vv)0�H��.!�Y��[�J��ّ�o޸ͻ�m��W���226
��J
`L��H-?2�-��� �$�n�F���?6��{��ڜcֿ���ݫ"��k�Y��ח���c��">�o.a�74܆����G�*^���FI�: ���I� ���)�%*z����[�zb��yLv��q)�.��sr�ڣ����D�u]��\���� ��<J齜�U���V���hs[f}�S[[[�{f�J �"�,.Xs��tP\e��5R��^7���"bsy��%��.bN��"pd��hV�����;��d����\܀�v���d4A��\�J���߂�JC�#êƜ��j��o��CKpA��I�(�����a� �u�z�߮�R$���2�,���U��oP�%8��(�.�@n(?�_lS�B6r2d����J|@?X�g�y���!:E5I/�� c��U���^5fFĻY{e���'��?7Jۯ�r�
���+�PA$��B1G�t�Z��=/�S�m/���{����jO��%��M���9�v����7�V��N[�����f�I፲�ļ�dS�ɕ+��������G��bY�njnQa��i.�B78�����O���24���8 !VSB����Q&����?���^ݭ���������G�mNڼ9�<@q&$|A�J���mYK3.���TRo�A�{Kwi�4���˕��mETVH5pV7UE�v�ӥ�¤P���T��\�Uf��nl4E��'�,��B�e�wY��L^B�f�P��+�}�w����iR4��^^�輯��<�|�B��.X�a��`sI����D��Ŭ �$���5�q�N���0�)����ɒs�yO9lώ�S���h���Yy9Pk��~qq43�n�a9Dd��?L���.3C.���ޅ^E������/���b:�ҰD�&��������骷O{�(�w���r��9�N?�}��UܫI̲� �
$8�S���`�KēiNc#��gW�~l̲ѿ��H%����)����V�U3��?����7_��M�HT��7ֽ��h��W�:��~�|-���w+.:�N��O<5�%�<�j�'(p��`�/�����,�q2Z�8S�,$u������ �I��ԯ6 �#�#�EV7{����o(=ۀvI�u�O���q� Xs�~Ă����MDN3�Ej�Z7]	b����`�����$H:�.�m�?!qC�LU�[��H��MQ˿#�nZ����'ݎ��+���e������u��7�W
�"��W-,�L򐘄]SK��ۇ;��:Y`锛F노�k���v��n���	b���ݗ����S�6x�V����O$���ĸ���W/���7,_��yq����TF��TK���M5�����R!{�x������i�O&�𦬉��㛳��E����������?-���D�����q�m˺p	`�.I�ɑ����4���O�$��o~�y	��9r���N��`5^��Ϳ�#ֿBk������G<d�dj����$�;*�M������	o��^��sϼ��-č�m�ߌxn �� }�4��l����&E�ͥ塷k���E~)ѮTE��/��F�'�m���PT���l�m=��WC?T�Q�ڞ�C�h�m)p;|�`\t�T�����aH�# l�"�%cA�w��N��K��r�|[@����Y�C:��f�L����$y��6�^.o2��JUZx�S{�����C%TU'��&�+G!��VS&MPoZ��� 
�4�{���W�w���j�i%)�m�#�����ߜ��ͣ����>��i�K{B~ۆ G�� ���`'��*�&��'��z��ojྸ��K$=�d����V�5YY@��5 |�=4L6pPI��Iqߍ2^0̮�˨��F�],�k���	U2����WJ���`�ɂA9Ř��jr�P�y]'7��wHu��^R"5��8�ZJAW.�2#��ܣ��>]����RO�-r�|���פ^L��cCN,qj�A��7200 �ٵG岓i��Q�e���l�55�G��t8��&�T,D�?!�FF��6�;�&�#�� ���*�B� B= P0 �()R���H:ե�Y��oA�bV���Ѐ��/��h*�5y-"�qy���f�������*��w�+�=�a�v33�|�7�8�bU?��n� o	�~p�V�y�\d���/8����V��g��8�R2�
��W��*5�u"�e%yCs�!�-���F'\��{�W��=�Ž��o^�jr�.��`�uC<O�wc��:(���$��W���U��9�J�#��i�Zd\g$6�8f����R "�n}�p�.Pq�BR3�B"�Xl!d%�U�[�~O��_��Dk�Ϟ�*��s�X5�Z���8Gf����UBos)�Y}``���h�w�С'�b�E.a�L�d*ں�����_7��}��K����m�l/o�$�
��!���_��˯��R��>e�{��Y�nK9���P�n���n0��0�5!��7��撥�GX�h��t痜���ז@�rO� ��ᷚ"*'��[:2�!�u�y�))�!�(�=��Bj���s�.���k+q�k���� W��D�B9ڏ��O{�G��'����ɇ�6�?�����_d� �&���wE���,)�s9(X�PbU���dvR��˹�R7���w����0@7p[�ՕS1��:IW�e���L���_�P��迅��%O � �Y��P7I`0��7��C��'�.L��� ��Y�����ߠAю�u~�e�m��M$�]���V+�{L��1�o��M�/���������I��J ��з��wp��G�ӟN��i+�c)��C1�����?
��.���n)Sb36ұ EYL�^�7��u���?}:Ff���������ƌ�wEՙ�'�Bĵ�dv�Q����0���CAU���V:뭔-�L1}��su����7�����#��d�RX��a���^���u�A�~���n�Ŀ�`�6T�C`����#����`�r"23�M
?4!�=�O�p�dē"�e+�z��'kNZҕ������m�Ů�O�\� �i#�%��J��M�_����ad/�/������,*>�$���
�-n]@�klj����o���?�n���<���c�k^����}��������{�D�/��>���0�0�<��Ҵ��<�Y`z�+*�=9���nAA��p�7-+)<�>����ĸ"�L�K_5��Q.�@��vu���+5�g���o�e��i�#e���L ����V��|� �F��Q?.��4G/IH����J�%`&ޕ�����'�%��3)���t1/��4������ȇݿJ���T?��+܅�#��Z-A��3��q		H��G�,���!�\���ᦅGA��t|w��Ne6�E�#�S�z��lFvxz�rH!R,b�n�J�H�hf7]�i��d�zۡ�1")�֟��F��`R��X-��Q�W�^i�96��<�Y:1{B�p�`�_��@ 봵�?� 2����sӹ�R��F���y�/"Т'����s��HGQRNN0z�eZL��'�����P�����wzI%�Ԭ_C����)��g�|A�ս,�p�	�|>إ����>5��6�ih�i�ȍ�Nb���n��.痳�hnn�m٤�IMJMe�|����&�O������(ĸ���V�K��<}0�h_�sG�z��Y���;�|\\d�u��;@&,W<ȢY��m��#�����9O ����C�����(=��j!*7o*荎gڔ�e�1=D�����^��[�O��-]�M�s�&TKa�[�w�$����7cy��2�A�ڙ֯4����u���~'�`�����7D@=��Ө�t0� ����P���Sdg?�d�02�H:��

�r�����rvW� �ǜ��APxT ��N0�a�y���HQM�Yvdڷ�����.W��ICCܖ�fm*�RK5��4�H��漉0b\��P.�l�/�g�� _ so�~͵��2���h!(��X|��$f٧������һ�ZSSC �"�j��>k���E��Dz�5t�K�8���z�!9i��+W};��Y���L^�3.�K��X�*��z����dɞ�lK����2�s�W���ՠ� �ǅ�Ї��%��Y��B����aoQsy�P��c������E`����|X��S�fޅ�]SM:�n�QϾ�� Ϯ*a<��H-����������@����,�i��v1{��Z��&���������OB�%V
�:�������8�i�Y��e��`J_��|��[v���|�P;��ʧ�Y��O�.��jS��UVH��]�1<p$�g�QdA�7$n|xq����}T�o5�����"	�?57���'��k��Z�B��Zʵ��"UI��|)~�Cސ�2ˢ;�=��ב����*��r8�3�s�,Al��2��$xv��-�YK�6/)!| n;y;���`SF���!y�3蹞�����FQ�o�P�Z$%'?D��c���p�#�|�[�,�i8��,�Z��C��]x0{��؛���'����8��3�2�!*+�V�H�
�wu�.��!T��A���Ch:_�|������7�C�v�X4����)o�p�ᶃ���k�"#)M�HH�2���"�V	�1��!����q��:(x��z�|k�͟�S}	���&��"�z�1p���������B�
�q%�/&������}���t?�	�v9]�Q�|7���F6���@A5Nn�O�D�_^|���}�z����+��GG;|� r/ bYA}�t���d�������>�k���B��L�������/�k-_w{I�b���l=�nC
�i��h8�VVE_䗺��qj��U��'|�ȑD���ux��XB���) �]�%��Q'�h߃"�ׅ��F��H<y!�vI��j����M����A.y�g�ΛU�s�A�[j�"O��Q��b�Ή�2���i��°�u��KTBߗ����B�?����Oɸo�Ƚ�����*�]15&�I�za���p��@\U������#�WY)U9VC*�M�!=���W0UF�Dxu}]
���C�\ޭ7ZJ��[��xIÆ@l"A�*k�B�c��M|FRe=be�&��Jo��'��J^J1���9S>�* u��X�+$}����9���J&7;�}<�����Ѳ��//��#���V��m�=ڍ ���\�eQz�c [x��~kaCe)E���j�ܢR�jx1��9�Gn�o���n�!�p��?�B�W,���D�j��o4��8�]=�?_��p��,�̄�D�dxbL�}��� r�%r7rBFi���2�YP�4\��%++x�3�b�o�k�vus�H�#���B�x�1���	YY��eDR*܉���w���:�_hΰ�GL�K:72!������o��7�4E��]�/N~�8�� ��.�_�?��z�1E�)Ù�_��{dg����ri��[%LŽ$��P�a�afH@�����X�s��"7<-y"T�����J��a6⸡��۬u,�C�A������#���O�<!))k���a�4�-0�L��T^�F$���"I��t��n��C�C��1 ��>{���|+^�Hm���,�@��Һ�V��z��߆v8<��Saɢ ��̃3*g��Y��@"l�Fi����𸝧,nuSs��G�e�I���`�,�Q���A����!����[(A�ȕX��H��Wx�Ȋ'!Qkq����;Hf]�	2 D��n~n2K����+.Pg�XЉ����T !d;
\��7��[:耾���
�G���R�9b�Z��smz����|6/����Ka���R���Y �� XX8�J��� ��ꅈy�u���}���	%�6�
�x`�Ӱ���E-Û�Z�{����;(I|��yU�N��5���i.��h�r�|9p+�'v���ֵ]L%Ԟ��3�įh41c�h TIii�PO����h�$����7ϳI��WAꕺ0�&C���>R��F��R,�9U�:i�^߿�M���g?E絿���w��#��E4yoģD!\7]�T7�-�<�(�1�=0���ȍ-(.���'�4֣ffa����������>0G�'K<`�(G-P�(���E}"Y�������V\*������.e�r��T�y�H�Ql�Ic	��V��i�(WF޻���=��Z�����[�y��H���D<iY�$kѾl�c�j�ȯ@E��?����^s��W��_�R�>�Y�eW(�J���%���d�QO;���������Oi�s�Ο��ӱ���L}dS�a��WHGd)F���+��䑂R��ʫ�FD�� �*��K;��@�8��la���hl��KUB���O%P��V��͸)x!ǻ/��4�r�"�pƦ��V��g� ��sɹ��ȕiA�W���;����R���w�.��ޢ%��Vi�.� �b3<S��')�����=^w|?�Cb�(�x��qL���4��4YZ�A-vv� ���)d}K0"
��t��i+�ۃ'�gsgQ���=��4]��+m*De�AU�T�7��e�.��р\��ٹu�h���G�F27���]��g��O|k�v��a~�[`�۳7A'�����k̀���-o1��21hǔ��x2/�t:C	�iR�G� 4����hL��p�M%���Ӏ��� �2.fq��ݶf��E�Dq]V�Q���q���dhE��Wl�hW��u9T�"#f�/�$ͨC�I�˴�(�n\�ع�Np:�2��fͱ��k��b��6��D����gb�h4���L�{om����2���|~}�q�yn%��rJ���

�_q�U<�s�rh��ܙ�������]�����w�"2�2O�"�o$��(J���"w�8rQ�����^��<=� ��o��r�P�҉FF���\1T"�-/���Y\r$[�v�U��+�-��oi���͗��+�,n�}Ob����h��k�Rpe�8-=݀Z�q�"ДJpX��zKҖ�Lk�

	aK�
�]�����M��E���?�+!|��Q�������z:�>\C	a��|����F�1\�[� �ߌ��\q�F�f���`�����M�	B���ke�n���j�����QJ�ѩ������Q'��zd���C`��c_+M��k�O�]����9��l�'�h�����|�s�q�k,�RO}I5gW1�QP���ƥ��Ƥ�T,(�0K�"!ʗY���uu"{���dn�d.�/|@t,\��.���
��w�gv���"�:"am˯��Q�u얯��Ă��7-y�Ѯ��4�|:��k׊�^9T��M[��9�9�h��]���<����k�VE�.��V_k�w=���s��"m��C�i�i_�o��2S�IS����י���Ɵԡ�_��V�H��5��ٰ%��n�ꥯ�Z3Y��ьށ����\��(Ϸ����f*��[���n�3'hY�����QVsD�);�M��f�<����t�2i}�4�Gr��#+f*�gT�Qc&��*?

��Xrl�%Mg����ʽ�c�,�t.4����5���� k���M�]����ў-��+;�k���g����:�}���4$7�[)��P���:��{�T�`2T{a��O�1T�x�4N��fY̩��֦��ϼ��^%�E���������<k�cF0_��A2�C89�ɉ�y���-l�ظN��1.�olnv���k��U�&�Fh�Z��`R!g���Y���`��l뼷�Γ�Ƭ6<:u��b���sJ;��=6�p%�_L۴��=�Wzyv���0:���H#bܑ���&Vֹ��4d�>E�?c�/(��DB�x/��ʽ%7|1M��&O-�U8�ƲV�A��'���&��7���ivx�Ѕ�{ 3��[�Oen���1I��'K����HK+��QUn]�]�,$���?��7E�y`���7�,����J��~�t����������͍��ŗ2��1���y����u�FC1�:�{����'��c���~5�?l*�9��!�DpL�W/)�|�N����`��Gw-Q�f�T�o$�w��ѐ
�ӧ+-���Hs�!����0���E���󎮏#�feeᇉ�`����NN�-g�]�VW?����u	�������j��0s�Cn���V�	zY�,�ޒ������3t�#�_������,݄f}������~�s������c��/:Z���y�r(��������:{����T��|��k�!&f�Ċ������m��V�~�-���.��)�U�=>u�DՋ;w� �T�F�� ��
�sL��$�흛����������oު�;�󥵛��ieF)D�8ў�'B�`��T�8/����XzP	��8����6��h�2�58u��2�
=������ݼ�u��^N���i=��w���� !�#TN�k��:ȆD��,�����MT�"T�k݄p�Uf;�X��Py�YȐE�)���(���<M��R����'-�`2 0���`��J^2Z�N֒����鹭`��W���o���X-��
!%�!**b}j�f�J36O�ut���Y��T���7p���Z��\�7���;uu�<�ǘ�>�}�"��d4$�y����[H�Q���P��ezkh��h�1��u�\��M�e��2+�Q'`�rL%7��[l��'Y�=���wp� �n̞h^����G�u�Eut��F1*c�H1�(E�� �(J�"�� RX�^ņR54�Ra�.E�^E`i"�KY`)��ܻ��|���{����w�̝)�cd��W3=�f \����JR@��F��Vr{ �ˏޞȃ�F|�_m���qZ�V�SQ�:�`L6�37ڂ���w�%u��뭇���Y��.'�bHv�-at����U��nw�W|���nrQ6)!b����ݽ�y�J"�5��&;8}����Q��P��4��Z��1Gu��9< �9� �W�c���!�D�b,A�} �b����4���].-e��-LO��0�vZ#� �o#))��2�z>�]�\K
���r� /��Wc��m7�+q�"�wpvfL�y�U؏"x�zl3ei�ee���;F[�U�U�����|��i���R{�������NAy�#OMo�����5�R,N�xX��$�^�֫>kщ���Q�Ϋ4����@T>� �Vr	�{2匈j|I R��4�r@�EH�5p;�_��
($17�nw���9�-�Dj{�~c�_��ɖM0P�ج�f��)���nt�R��y:��]s@(dW�>ή��w�}i���.*��'�F\T�j/�z�Nl�,���ܐ�+� ��	I�{�\2
��&g���0u}lsn��T�e���js���>׶?�M��[�D��8p�;�����z͸o������&��� �* [�u��7�5���9-퍁�%�SQ�DH��'��)==�x&N���:18�ޓ���ڶ�ኇ�G(����ӊ�w���������U�M~<6�ڍcQo:' �n���a�0F�6�\�;^N)7i���a�M��!�:�5����/	L:4���~���X�<�_{�-h�;�h�z�`�l��ԥ�ը�����%,�W�?��Q�cSdH�}z ��=@A�[��ňX[����S�p&"Q7+�
p�����I��Q�Z�D���xZi_�z~��%��� w<(^^�i��Fx��J  8"�f $��,��'S�ǪD���j��d`���֯�	��b�Q���0�P��?� �J�H&�E�쎂��j�_&�Ey�F���"m�ѡ=/���2�y��\.�I�#60��̏c�G2���.yt����E,�� ��(d�j
8��#�p�D16���G����`����ޱ��GL�v�W���DTk�9����?Ⱥ����1P�S/����Ťo��2�5�Y?t��x��~�mX:/�U�=x�69Jb�\�$N%�
Ċ�(B�c�4S���C���G�����l���v*Tq��T	x�*V��{�J�	�0���L�f �=T��,__|� ����,���q#v��ΐ˟^¾�on�; =
��<^Ŷ��Ch�@M:<+��*䊠��[Qa�����%�*�'�;`܌�B�ؐ��6���]t��ki�;H�9�9���z,��a�@����^���z��~z�	_P^�t^d�F t!߸����3~t ��rS���['g�V>��hv*D��BPO})t�J�m��s�P%r�(�x� -�� ��N(ŏ��q��}2+�v��%B�BK�����@X��|��?��_�K��p�%(��=�
�D/3U�h(؀�Pmv�3 :��F.@��G�s�-t�ŵ��ʵ�/0�����y� .xTe'�},e"aw�	�������������6������.��vV���!�4�L[�L�a�!��&O�nG/6�<0:���g���f�}�<��z9yoZ�2nk��F�+a|w8~G6�c6)�G�u�<�"˲�0�QQP3W\�k\N��+l��9�r�؛JK�GOgI6�F$�!�E�(���w�ϖ�2��>�� ¾�R�7��!Z���xb���*��J���HN�C�m��=4�����E>���NA>�y�MXo������ �BP7^�>~����'pѝ�6�����]]	�:k�kH�P�J�zO`�=��q�zry�����6��!��S��Z��GN�����m���D�ku�L{S�$��S�v�`8g;�1��A�7�zR�Q퓟;�����O���Kn8!�d3��E��^���s*o��������`Q�`@��G���C������#W|
85��OZ��P|4�
�c���rP��S[ےl��h=M����z.�q[� RֺT��m�o;o��F�ah0_���A��oT�:w�X[F��3o��AD��7Xz%�7
��6$�=5�R�^d ׎E���9���+q~tC��$Du�E0��
��Զ�����Ц8ަ��oTP��|�M@�D�^��CN�����5��M�w]� 2�`�g��x��ax����(�)�$�����_� �م������{�aVݾ���&�9x�"P�	��S:��VOp8�̃����WIT��C�˲yqd�Q����\^7e�H�E��[ͬ@���ӥ���wN�3�;A�c6���mb*�۔TO�@ �������}^�fSU�LDe�cy����={G,�� ��c����I� �[r�1�n��9Iϰx����*�8�]��.�q]�	�|xR�c\��A�3��׬���2���V�N>�F?#���c�06��!��j�����c�ZA��{�G��!ѐ/Ҡc$���U��m,4
�����=�¿�h��34!�"��'��P�P���e���#������������q�$�W�2�.^�:��	ňXR������f���^�[*#�����	S�� &)2���/ρxF1��F�� ~�M7�Gg��n��x�mj���&"�sbGs�}����*���߶M�%,z7��5�)�W1�X�>]d�3�.���Q=%?�J�; ��p�"�[�\|Z�p��#�F�l'�+����xӥD�r�@��S!��A���]��czR��DJoQ���َGٸ=[����|ja�-�C��D��� ���W"�3�2:�5��c��3$ :=á�j�� �3��Մ�g��@���b(�LԶ�<=����ٸ�%�Bȓ��[�tZ��&�*���DoonN�}��b��!)���c�� �6���0|�����V,�O[G���X�}�Y�S�b��	���{7�6�Ю�8�cF����»�l,ԍ���t?`v�����G�'�A���Ui���e,��`*\E��<�@��/�;>j�PN,�4~H�SV����dC>}�]B �M��R�Wru�	x\�Z�Z�F�@��c%�E�UP~��F�a��:�����Uos� �P-? C��S~�C��l\�(�h�y�ײC |Oڱ���mA�n���x�>&����%�y@�Y��}	��A=݌����a��9n�����'�'�6�i�&2�����V����47�l���a5�̈́��D�;��#�����y�I]6Ρ��$�����F����x!��w���S���0�4������)�/�qd�N�FJ_� ހ���s�m���XL{� cZ�qy�+�/�"�VJ��}s����MT/���	��v�4
1�q5��t�8��vOJ��~��Y$*&5��A8��I����P�������)}��j|�[��ST�ȿ� ��D�@[hQ�� �c
(~Xh��&? �M�?�$C�!����&ئ-�혗(���V�r�j]��\๼��Z����Y�,�B�6�!T�Wb�~�8Gao�n2Aױ�ǧ$��ۭ����Ș�/���n�-cv8�s�h��J�����������Rj�l��C��/*���>�;ji�j�>����I��M (*n�+/��GV�����^���.��5v������^f_��A`x�G�%[��v��=�Ї�1|[bX10�.�ur�Z
rJ` �ʫX��K��������i�8�rA�: C'��D���*RT2�#��kk;�\��ޜ\-������U1�'8m�����ѨY3���}rH&�N@&Ƹd����`NW*>P�'��$
e�urU��mRz�t��:u��C*F��a<���s��m�:��#z	�^b :#���dol��h	����:8����~�J����a0��V9]�+��2y�4#�Ţ,��Y�$��[A���	�Z�����4a���kA�������B���33ڮ��/��"�h+Ȭ4��w��W��x�mwP�v�|�'��a��f����BxU��p+��NN	�d����Fp{X��)�����q4�bbx��~(�����P~,74�Ȓ�"�q-�r(�z�r�OS9��h]J����g�iOY}�O��Xբ��U'��ɳ����2�0����F�<%��1�����Y۬y	�#&s-�ຓ0Ћ��}6��t��9�1�������C�W�6n�"y냱Z�qۤg#H�  Ɯ����Yn���`�2+��� S��3�bj.��d�B���f�z��7al��>=���b��(��Pu��"M�o�	�μa��RTq��*o�vOG��妍���"��NM,�?��ۯ�EׯJ�6@����
`3a�`{#���ް�l�| ��ڳޛ�u!*�ʣ'�h�p��1ٲ��A8��]X9v�4.놧�j@�Y�΅�Fο���Wu����]	�6���X���VS�T(��ܧ�����Y�N���m�C�~L�߂�%�%Zo��H����H��L�dX�ķ8K���}7�n�C���\�k^�]�y�mр�>|�X��(&+�H�� �P~���|k6�׋����
�>�ᬄ�م.����>[�:]0�4n.d��k���F=���%�����	�X0�!N��8|-*��nY"�Lfe�/T��٦�!թ	�'�&g~!���}�J��8ݎg!�o� =���`J6涖�.�1�C��eC/�(gi�|�Ri����z�ꉻ��o����d�+|���o�	"6�L��(�̻����J[���^\��"��wo"�
O�R���˧x���``�i�bY�Џ��r�^x{��
H��[ȃH����	xC�k�e��v-�r@2��t�|�M�~�����i���q��on��t�oY�,��~�睅�8���H���L ��?Ru�@Ner����6��2V��#�&t�� ��j�B�O�С��"�)2�˧�5�e�B�ʳ(l��ͯdc���,�����;v���o�,��k/��6y��B��0}���~`9%��In?h"fU�@f&:�2���L�4�z�������h��&�%<�����\����*�!`T�Ȩ��	YD��#xL�B��yc��gv焴"��+h��zr�V���`����
�[u.���l��+�
?w�̷�̫Vb�
Jq
��MK����ծI������F�O�iH (�MH`���r3L�:wS:S~f �jC7^����A� {��q��PJ�f�����|ł���;�a��w�c��a�� ��J��R��[	��W�(�F���6��.{.��F����n>Xh�M˥�)�C�1�f�� rVrr �[B�AM[\XN���R� 1	��i�oy}7���Y��Nt;Gx�I�õ��m�����g�>�lh���� 6TI���ۍ�Ehu�7D0�����;��"v*����B"��)�5������	&��+,���{9q/I3�����އ�/��V`��6a��@r5_O˭��I}�{�n�^�@�_�<�Zxj�R��N�������(���}�]�<6Qu}�~�����c�D=�Ѐ�8{]�l،�/"���X��z�P2����h	Ovv0	�q;L�ݥ;W�F)9s������]?�{���&��^+�2.'+����¢ʁ��-oz�})Q�WJ����׬��/�F��2e�4&V�FO�f��'M7%\0�d��ؔ�ed�6�誂�cOS�a<���]9�XJ�T�x^*/ ��d/�
����t�b��ls���6�g6i�;��"�y'��Յ�=^�$�fp����v����ۧ�`�L)��hbd@���ꮔ�E�5�e�j/q.�V��Pd@���a��8�mr%UTWl��$�D��������F�]X�x
�R&$��z�X�����$Dૼ@ �~6x(߹���c�(���f5ɻQVm��!�(T���"zc]o,��������&R��b�zϲ�U��D��Y��Z��К~�ng�FS�S�����+���(���&��F��8�%:��q�K�.ho�V�������\	�O:�����6�x��Z"�+((�KӀ�J��h��Ou��>�<r�"j��=khcʣK��S.(�FG��������+��n�۰�8��zԵ	�]�y�����Znn��j��-�[.�jw�F�eN}(������WυwD;,��g͉�+s��5�H[�#���WB����!1�{��/#:�L�9��c���i���fz���n%s��o$�������m��=��.%腣n�S���-�ߕ���>���@/l��]�j�<l����;x?%V���$m�z��]m�)խ6yPtD�S{���{��&�9�1M����t�G`�,Y�1%��؋/S�Y(jJx��[|.I��_c*��w#C�� ��b\jʶm�[��`I�N�������N3�����h��Ѱ>�);9}�2xכ�[�n��L���T��������m�pJ�Q��4>t�����iW�u���Zp����e�O�>o	��;����>�*�I�'c��tf�{�>��H�����n�|��w��������/^����^Y�.�	[+q���41uV���(c6ЯVJ>�u�\��8\6m�Y}#���۲�F��%�֭�����"��5�[5� 81.~0��t*]}��낞K�J�dk���$*�8�;<{8H��KDҗ&�i�N�n�q��Q;n����q���gQ�aF>����i��$�<��ކ��l�./��N�;]��~e�:��Ʊy�����𳌇	^�y�_��4�I5V���u����8�=�T�mQ�U=gN=CY�\F��&H+&Z�%[��YSq�zd���/t�����ꗹ�0�O�����k�~�.�;oE�٣,`�p�C����}ʞ�!��4/Mt�4!�[j�&j����CC�?G�
~���Qd�e�z�))�<",.���C�1�-@=���#�����Y��*�"�H�c ��ܶm(ى��0@��"�T؅6�0¬����:$�y��q��>��,ا-q��ˮH��f����z8qdC;]ch����!i�Q��@�qg�YCBB���f�̧�A��#�s��u{��@8m��z�#�&(p7�|�t�]����� K���=��H+hÌ�!M��2,�x����g����I���2ܶw�OP??���>��U'�c��f��Ð ~b^��Ky6
?�P�y���)�{�,�UkƤ� e� ��5��.�|��+zj�MY�hw��|������,�z��Q�!����s4������W��.(�]���KS�˟�7�v_�f��o2�f�T����%ϻ�Axo-�$��.Ι�n�-s�"�/M�e;L��ͦ���+A��L�ժBDAT{U���`
RK�:�����P{^E���7ڥ��(}Y>`դ��^�'W����Z�e�`��r�������ǵ��A��6�&��`������H��!J檞S�z�&vL��^9�&w��J��؛���)�FOO�,����ƥ%+�eJ�����g��Oc�q��;|C���|�2N��o,e-��3<�܆�����#���:�����r��J����B����T0���O�u|�
a�\�|vM]����x��˶�]1�'V�%(��Y*A��ʕ���n�%b���v�^}�9�ZY�Z�����?�#;�W2�G�@#5`�`�4'�/[a�O�Թs�w�Ǐq��W�h��#���$7��7�j��	�} 5���VO6��N9�`�m���N���32����vl���˗|Td.;w�����^��<읱�r��:���OXT-V���--߾]u�}�8�}?E���
�y痧��~��-�?,�D��C�`�=x35R-� ɇ�ŚJ�Bl1/%녇��x��ִ�����U�/����o�y���"'��^8���?�����f4��<7�~8v�3L8��r��.S�~[QJi�{��K�ю~θ���s��0��~�0h��B*J�*2�p������.Qڇ�o�a��z�:!**2�o�����Ń�ū�2/���.�߂?�=�2U�2qc����n����DU��-��ƤܥpR��*�n^1A����Oo�j9���W�^{m�n`iްM������s
K����G7��*�4ͽ9���K" Tg�|	ʑ�6YY�˱�[�;���h���Q�9�k<@����d�u��҄5n%���ƻ(��mch���h�p`�9�����Q9�LA[q�e(���O�epO2A��0!n�f��8~p����[��P� � �A��)(�>��o������=N2��"�/���Ԥ�ƅu��M�́O%Gy�ρ�5__��<Vd�溷��>\ER׷)�J3ٝ�Ln�m� /+�/N��#��A�qV�R�%$߇]$GJ�7Cl���<���h��<��B��
��{��u½|�g�j������u�w��X�1��_�F!x}��[�z�����K̞�: �y�" �A��ƚ��@v�JV�w��+',� Y �yfD�!@@����-/���l�
v�F��<���VnJ�r�({��B���C3���Q��o#A���J���������X��엡ܦ̓�䚹9�Pu��i��˗A�tt�ݗ��C��1�:J=[���ш��Q"���:���N��E�$��6�j�xe�����2��Q��>J��	��/���7͇�q����@i����O"+����oHQA�#�����7��/��U.1(YJp(V�l��]��G��!b���3Z��W�a�:��	�C��.
����_��������guu5$�P�֥����qL0f7��8ߵZ)(���O�̳���P+���vx��ƕm�x�L%M����fR��&��D�xȡ\y>���KzO). �Y�z���N�z��ϟ@Q+3�A�B��\t4�V��n�r��'f#���]~B�~DP�A�8����!�K;E. �h�u��&�Ck�����[%7�j�ع?c�Ƙ���zf�3�x>A�g�V-Ŕ s �o���\/�)�p����?��Ck�z���=��̒���ȓ=��OIC���f\�7?ko׋-�U̏e�|o��U�tm欤, dv��;�D��c:hL����	L�;�B֓�C��1�L���%m~�ing'ũv�!�˿���@v|�e���Ok�u!��9z��xez��h�JxD0�Mz�.�u�wƱ�ޡ¼۴V�,���p{N3�􃠒ݻ\{{8{�r�Նz��eo��8�;��e�Z����[�2o_���Lq�\m���"��U-4�I�ݞ`j�S�8����m�����is�֜��g=n����S���7y����m�G�2��&���ՙ"�K��)���?�n@�W���ya�7��B+ֻ�KWG'{��� .���DA_���[����O4�< $���2O��#���-Ŵ���J�k#zR\S�r������O�78�Q�)��	� i6�(�2�`J<���Vn\���=2�8��7Q�#cc�a��"1����{Z��,�Î%�H-��T�j�#������|VN�s�����=�w��ۅ��֌�LԽB_8��NvL��<��+��;�!�;'��]Lj��}�,� ���a��R�R0Hy�}��maX+7�r�[h+�,rw���Q��{��nY�.0ԁ��|LNQ+�N�c�׬�.��i{{;�EPq�A���W��CqO��������{t�8��˱��kv!��P�hZ{�g0�kB�*�&oNu�y��� _�.�Ր7���SX�����Լd���_��r�HuR+돷d��	>�2�ڡ����57Q��$�<F�@&7o!4C&SM�Ug�����f�.�Ⳍ�P�ڊF����7��CFq���9���e���9qD}Kx{i���[�{�\�C��"����~W$�Kʷ򅷓!���\���*6['#��}���;lZ�ӨSJP��N����X�y^�&+�QɈ�f��@�^\�"*�7�q<����wl�B^����Ug\�: {�ŀ�{(8�L-bv�:�"*'�����LE=����2'Yށ<U*�:8سs&�	���/��S�0u��鑎�N�4��;��+˯�q<8���R�T�mڀ����R��e�J�C�>5�D/��;���:e����hy��0{�:գ��Pٻ���]� ���p��5wsC���]cR`'��`_�l�����;����;�ĝ������L:Ȇ��G{e��j�_���9�d�^TP4�<��r�I��aC.:���u�6�l�g�W�K*t�RT���v#M��1c�h)�<�p�d��k����0��R����'�,&�!Vc��F��a�\��&�Sa4Lk�]6⎅]��|�47I��:��i��UPל�y�w����];d���4��L�8���Cc����D�Au�ڧv��/R�&�X�J붞�l�L�t�P����%XB�l���(������+)�uJ��D5�bf���SB��K7�ߺ�n�7������ݿ;�Y裭�JroW�Ā�Aŉ�&������KWg�ȆU7��'�*n!��:<ِ��yG�㬴��N����7���S8r"g��*��M-LtB����WPJb���OZ[�����Fљ �ߵ ���|���w�R�}<�~t�
�8C���4�=q�h�pP-5u6 ���[��ؼ�E�[�PPV'�bH0�Q��R�=mȱ���3P��D1-p��� �ݟ�r�WW�����%K�v+�X�z�:10�6<� ����$J�*��8�ʆc&�ݔ�#��1hX
���"�Tr0�y�a�6��f��r&a��� f|��`c��VE�X!�۴n9�95eo��_����$� HCb�?�sB��Q�.N<��;%�dw���d9���o�1�nNY-�i�w轢�o�A�OE��=����F��k]�r��<����� ��N��q�.=�u��l��YB�ؗuho;�~eks�*�F�J��2q4 U�5'G�&���N���b%�3{Z�~�r������4~DE�-yX��������- {dd��hz{�D!0�w�l��L�q���~'_�_YA�Ǿy����'�U��Ӛ�/:&6�vȏX礆�'�.�'KWMPL�g� ��'�J�F���e}����㊡�څ~������3 ���x�n��Zr��Lo��OY�@��Xz̷6��4�$�] �&��
@��+��&��Ç��e�l����7��gfϞp+��Rl�dl.��R�I�wZ|��������31(�ʋ�;���5�"_�D.i��w���#
� ����f�����]�I��_P��:��xnC�o��?�Ր��rAy�"�W���ݧw���W��|��!" ��%"֕*�m��L���W�7b� �)��ĺ����.���- a�蜑j��n�zDn&_,E�3_��l�v�tu�Z�,*|��s���@�5k�C5�]/A��(�U:~QT5��9�)����㰌|Z�60Z�%JȠqWN|��T@�? Z�;�8{��K�577����UjQK��U���/J����t@I�UN��V�%qz���)�� ��(8Y���F��..y���<� �ğWe�׃<.�(�M�%' Dv+$�p&j�����r�5�MZ|"�(:dȝ~�e�/rl#��H	�����0�+�f���&���.��CՊ�5�Vko�Cc�+3�Hy)�{��P}]��h�R�b�j��.���/\#��I�>��j�bd������#��@^',K������㦓qg�l���_�Fڃ�O�F� �����luT��O4X(�es���b�Rz�K꺛;lӨ�E�"���|ʸ��(�#V|����[=v���Z�-��۴Jx����E~K���e8�\�{;�g]��c���Xeݠ:i��_�	7Y���D��:�H"�d5${v����[=��xų�m�kЛ��s�m�1_dL�*����f9 ���\�(ˍ<J~f��띜W�ٿ�*�oF���oP����4ǧbګ�����鍊WL�ԸB%��p3�_x8�����q����x�fF��{�8���ݘL�=�Zy6�VRd\��!2�i߫�\7V�ekM�|ƣ!�2�b�^��T��[�tUu�� �TF3��<��{۽�r�]W�?)=Ǿ�wdⳡC��W�k�p��ʃY��e:$�6���[]1��?P�������i��.��X:�} �
�^}tN�O�7��O>fg�'���؂52���4+�b�!S�x��z�/� m�=Կ�d�)�;�' ������$��^�q=�^?�!A֞ȒL�l�ך�ܷv�%ߜ�;�x�/UM��e���̃x(��(w�)�' �6��� M��&��Qm��Ǘ�[��U��Y��Lʞ����'**���v��k`n Z$����T�ou�G������>��g���#ܭ:)r�V)�vS�G���Hާ��)���+�,S3ԫ9�m���^�쾱� �<��wCnl�͏�K:�����BO��y�#r���@ x�G4cҿ��KoU�M�(���@�x����`rt}�ۭٹ��L���c�0��N��R��k�P2�\@$>�hv�4w]�B$�������!��ׄ���&��m &�6Qsj�0N8���<�89M�'L�i�g��1/<x8L��B�/�� �QP�:T��@֫!�q����W�Ѧ��n���5nP��շ�T�e�K���� P��-��3|d�/n�1C�<b���p5B�ox�?��.#�:�7'�O[P�{�K�!�F�s����d�0X�4�4n�F�����S�Es��d�Yy� m A�����m #��x2죈:��YkE�l��Y򶟣r�c4�N�j�ơ�0܍(U�b�@�:be=�8 km7~��a����z?ȧp���	L�qBF����k�(� G�fK-��Afhj_�'Yq�LoP �=c� 2����&KS��2�*�{��������M�	0��T��0��Ғ�� �\�46�פ�a�8���|R�a��mb��2Rjr6S
��o�)�_��Ю�TtH�������-�mp=�ybH�\ ��7�+UAa�`@���n���	�i�w�F�Ͱ�O8�����[��h葻���E�^_$�����ט��^: �rJ�Y�SG����rN|��R�C����w� �j3[4i�IU��ܞB�GDh��E["��V�|�_Je�A�Xt�%�͚u���9
�|_��`�Q��&j���-�NfI����'����^��$��@��w=�K֍��S��_�,��3�6���u|��a{�'�}�u��ѻ�e�̉<b�1C(b��s�m6>2[�Vil�_M��9��	<\*Cy��gUP�d��@�Z��^|yni:��j7'�i`��|R̷ɋ�\�@	$��Ʀ���X�o�K
�Lej����OS��1��y�X�E#,>��y���Zh��O[[[�|t�ʖ�zĩ�o�;��7���ʔ��zES�?j���#���z��}��\F�]��L��FY*/�G����� ڂj�$==���SP:G�G�������ny��7R�K����M��W��V� ����N����C:yS�<wG$_�Z)Tn������"������Mn5Q̗F���wl�"5�����(�^kd�����70B��qZ�ܲ�a�T4�)���2:��rj$�KB��>��/
ܡ��4u��F՛����/o���go�O�9 �T>��A����i��U�8Sp��0��iW�;��_��y��~8|�A5�l��8	��'�)���s��Nj�ڍ���|�SF�s�Mޥ��'���<n0[��N­����!�uZ����1���(�e��c��+�(|R����J[�������yൈ�J/�8;��ZZ���m��p�68hG��3u��@��0�	�E2$[�I&�׉�g�q�4(3j;���Y@ПVW��=�
�h`&�B��
����D��l?�]X���G��{��
��T�*Z�=�d����WN����e�t������rQ�|~r"1�Loy4��Dz�4�Ɵ�{��_I~T9�/:�疝0+Ss��`g�Ǐ�q�݂�a�@�U�@��?�JCí�x���1��r\Z�za�Z(��E�����L����%�̠�Fض-9Cv��փ�_)�oLZY6t�2\yd��1T��F���XH$�.��k}�c����[ԮK}<���ԤYuS�;��-�9�
�#��m��j�;p�۴�R�&q!m�Q���<
S[��*N�ӊAx�Li~�-�*�{��O^��~�\�Fa��O�&��� �a� ;t�CU7��5w��91{t�fB\B�K۔5/��1)p�����w{�6�����Jg`��^iud���Fݶ��R��3}hJ�%AOl@�介�S�ܜ�����Ef��7�L����J�B�P.e��Õ^ �;P���B�CIm���se��Z72��!������"�'Y�6�[`��rs}m��V�n`/���"v���]�U��Y��xm��(�h\4}::S�>j����9�Id��(���i(Ń`:00 ��
�W�/�_����'��{S���y�Ά��{̔�����qބ�����`�r��>D�q���e%29h��^�a�:�q3j����ԯ�V�xv����+�����P��e~(���:�b��˦ nɆn���������b��뺷�ˤ�$�j}}s��DS�
�+�f�}��q��p���c#��\r^��viD����S�����&��A��T4;�Cm���A}�x�����߰딨�F6Lb1_���y�}DͶ-�GK�¶I K���v�"0�@�G�PBSE���T.�	n��.mRt-$G �j䩟U�ޑs��������7�9ܭx�<Z��m��A�^Sw�_,s��'�-��F�i��@e�m[�Fx䱟�L�g�s��s�<���r� ���B�q?���w���M�6��#��/h����� �`G�N��=54y��������M��Aզ���g|�z�c����%Wd�I��3�h` P=ؔ!n����_��)TZ���P@���v���,Lt\�<.��w�����f�
+׹aq�|���z����[:b�3��R����F�9��)���Q��őZ�A�;� �(,8g�~Ě�CKV�I�yN�p�����^Ya�Ǩ}Fjx{{��f%j�����H��z���A2��&pK��D�+í̋��]���¦&r�k�P9hR" �j�T"W�����֞%鑐�?Ev�.e��s�5�ޅ�ل��-7
c5U0�6�m�ݺvݚU���{u���������9SC�g�	��r�(X������Xxb�t�;A��+�b%�f.���N��q�g��T��<�*��&**)e�<��+P<'��x4�f�N)�������3���@�I=}���m�f�۟_�ȟ��CG�����7�d�uW���-����",�S��G���9��/i l<�GTDD��62���y}�wѶl�!�.kKC��7����
��_���N�Ww[��+z��q��#���'�J���� �Qj)���C�޲RW,B�׎G������^\~�*>Y�*�zo>��u
��-������K�0dＯ��+��W��M7��.�_D?+��z#^FG@�r��r�����9z��nSS�v�S�bRW����g!Pb��L+�).u�6��K�=x�D�7��4n��P�k��=E�����jF�#�ժ��$�=��ސ��#�d��oViT%�]`�xC�RzkU�Ű�l�M�tN)QF"��٢�?�b��e��놮����?�rA�/0���hd�?}d�A ����s�U�$h߆$s�im���sB�c�⩆�S��J<����AHs��kR�㭳���֖'��Go�u�ͻ�C7�|7�<��u��FQQ1AG���	���KU�(8fl������B��*U�![���)[D�����~�f���E�MU�����l/��L�^�G��y��%t�]<����)_���,��0�޵�F�;�Qq�En��::YP\�mc�<y033�lRg�I��Of�`�pO��³_�X��@�����M)�8PI��U��NB��9��Ř8%C��v�yaX�6�f`@���Sn�/��NjpO8�X���X����}a]�=/ܐ����m�����ݫF�ۼR".y|�����o�2(
�Ğ������@�ߛ�1;��^#�D)���%[�EV�漩�K@?�G�vk�dK����{�5�;?��j#�a}�Ő������C1�t)#rssӥd~HI����.��y�:�>�_g���%f���.�v������~#��A�~�-#��pC���x�\�2��� ��yK,�<��*0�W��B�D�w��K*�;�ϻG�>�r-���<	�AQ˙[֯:o��;Ք��W�1��5wAc�5 ���k��kwq��rny&)�4�#�xS�0�)��k"�;�nu�$�
���e�����ζ����g�l�4
\ťL{�M��9������E�/�*���b�cR����[1v�Z����*�|�w�ؘ���>K�����u}_&�*��w�jxxx�ٮ;�/?ž?(ix�n�`w~H��_�����Jd��C7>h|�Q�jr�4G�Aː������Ðf< �|��x�����q�#$�<���b-�@��U{���&�g��'�Q����X������D��;'���4��K
F���R[M��hgx�s��u1�F��,��7�X/z�]�
d˧jP4
Xg�.��𐮨�D��"oι��V/={�Iq lޏ��:���&���/�0}�_ж��� �e�+��-��6\����X$:�s�-z��#����&��L���hV��fo���>R�h�%��Ee[�0�����D��*L�۹�q��:gay\Ո��n&3��S1d��b|彾6~�J`,x�ȅ}]6_v����ʴ������5u_�
.6@ GWI�A*Z���9@Y`�Df���s��1��ͯ���v*l�#�໘H��]jU�;B�V�Ɓ��UMyo�,r��Ï����@6nb��㮱k�Nj
�S�S!>&nY�����{_Pt)�mS�3��o-.��7-�E��k��q�Prr2������u@��$�Ҍ+_��M/���@6��\鳐̇���z�އ�W>�`�Z��7�?�4���YΦ�Z÷�.]�"]3�5�����]�6�6x ��PUx U�W֝�O�<�X��2��f���2.oXS��Q)O~ ���FKk�gec�D���v��9����C�1�c�`�{�ۦ/�D|��+��*kf�B�(� ؒx�<��̘�:��*�W�#?R2	�tx��zɯ�˄�=oo��Ĩ�����4tIv���1ј�C,��X��~{�\�s����1�@���v�����ݟ`^t4Ee��G~�n���ZU��۪f����rt�3)�q�e3@w0@ � �ן����FE]�T6��͜��� �]aQY�Rr��I��7RŻ]x�k�eA�q�<F�zP���!A҇��t�;�t��r�����:�i���l�u?�!��b����ɋ��� r��ҏ�=�0ԗ�O�WuR�^&zE/87��>,�&+��c>~W>"�5@X����=,��~�ر��W�~	620!�.@�M7�O�X�胸ۊ���E�^�WOpe��<	>'>u�<T5�5me�'%�K:<��2�����H�&dÕ�<�/Ͻwp:ɧ���~�B� t�BQ�U)��~�RO������1!##�����x�m���&�$�yP�ytE��W�#�}$��~�Э}O` b�B��h�5�ҩ�`����*����G����O���o�T�AH�DM��¯�� GӅ�;��i�����_��4�L�@��?����{���0�����H陪LJ������m^$m����(�(�������Ϡ�_	
v��ߏ�||4�2�i7�#�*�T���#eZ�ݗBg[4+��~E�u���?�;M��`��m5v�Qɟc�6`u��m�ԉNt���:į��t��]e+z�)t�i� *�1�3 �s1s�j��09�&�B����0XP@Q)��=��N��%u���w�g� 	j���w�n'�;�X%�ߎU#��������K���f��mn��t��ټs��v��J%�I� �y�$\���[�uc�b,��5[��4�2���t�/���~�Qq�f�y��ɖsF20BFa�'j�
J���iMew�%��6�w�զ�\K�1=��/[�Z�K9d=$�Sq�k� �bc��. �D��.�l�މ콹���˻ޭ	R�5�������{�3�:LR8yO%R�Vz��r����g	�	�#Wa�rk�^�ZH�W;Rs�`�~b�`n��	�[۵�
2��uF;�X��V��;���E�Ʊ�nǑ��|7����Kn4�0qx�2�
3�һl*H��8p"��#T�L��\[G�Є2��^�3Sz�hhz4}�s��8�!��!��=ExNЪi�dG�K�r=����1 7Nv����H@��uu��� ڍT�!&���ݏ/�za�T�q����u�&���9���x��CR���r ��ҥn��][С�|0��b�&�n�Owv��Kъ<i�
��C�lV4�_��nY��u�p~�10��v�L�P�Щ���q��n!�?D�@8��1�R�N���Ӱ�����P�@޷�����M9��]T2t���]Q�o��'z��,e��$x�6"���ͼ����K�{R���^��c 5�6��W����A�������M]�j�[�-7�W7N��F�j�Dj�{^�J��s��f�䬭KV��6��\v�ҥ.2D�	�Ni;>m#�L?I�9��nyOCHtPKu7)_��J_��9qFS�fF� DPċo[���v�)��9�N*�ZTWQQ����c��t�%�,��?�K*��v�%>�]-�E��{�s�L�l���w�0{۞���k��u�w)�˜�Ka�/37�8n�����_Ż  �{������^ߊG��եP��Y��Y�}nV�	��˽{�{���5��3��/�S\y1�����b�N�0E�2%���ۏ` y#��PT곑���HIA�4ȗu_�${�yy/� t�m�ked��I������jr�o:�JYY�'N�9Ȇ`�/B�>#��ư��p%|�x��Q��qYf[��p�����R*�*H�c�"!! ���� ݠ�`Q�H����t)!"% �t>R�����~���}��Z׺�����w{��ğb�/!3(�4L�J�rq@��Ò�,��YN�/��8��~P��+*��R�S���>������#���C;��ɂ+Fp��YN�b�@�U����.�]��0���f�$d��C��i||y��Z��`+ *�W �og`\u���}=_F������y3u����^����f�v��ϼ�V��Q�ٹ_=d#r��|d�BO/	��Z����$�' ��}�\���mJ\�A���&5U���9A��D���)*)]?�3ښ����tt�Ed	g �	�<
�B�ɦ釩�zƿ��6e`�Zp�á4���.�i|o���r�#]tf���uDx�F��8�\d���,L�P�Y�eA�ys�~��Ă�!^<�����է��n2n%���g��y��(��q�������k#���F!�i���a
����I~���*�U�.R>^��D?)� d��o�GK��aѹ�?+��dd���}���١i־Z�il�X��q�Nq\��'�"�j�����d�Za����I!�N���!���|����cB4VWm����Y;ͅh#�Ј+!��y��`~�Ҝ;u��C�օ�n2v��`�c �I	G��*[���c�?>]������~w�r쏍�8?�9P|��l_7�caL���.e��o1��hEj'0�$%���?N�/Q�W�A���2�
�
�:ζ��^�&(s�MʾfǬ�Q��]k�lԳ$vxK��9=SZ���Ņvj�q�#A �����db?����l�%��^U���&f%��+��x�a)��+n�cw����jq��f�9���ȱ8aINi� �:���=�������Ǐ�4�2vX��>���m�(���R����F�T��|pآ�c��<�\�3�5�<�M<��yR�M��|n���~_�����ʺ��%y@�ǫt�`e�T��k-���( GL
JB�&�ivL~�	:�k�vK�k.�^^�13�t�-e����Vd�^�.B�����4`"<�]��)���!(x��) ,5y*NB�9R���!��e͉�[L]��|��y�ӑ���滪$Wڠ�x�%��{��Hy��?-��V����u�Gz���_L����WڟO,NV�ʘ�౐J�sC�>x�ZPJ�hct9��fmm��f�� =�Ԡi�]�o-"�r��R����ț�'=�����VS��(i�H�E��[:L�����_��@�;L�c"�t2@��Б�����_�_`U�wv����ؔ��J�����<W%(h�U��]�����H̛_Y���$ux�ή�������/mY�ب��p�f������>=>HpJ�q(6��H�(�Xk7�V5f��l�P�Ԋ9`!�CBC�(i���̆��+O��f�h-��v1���]�9`ЛfW��L�#�\S�Y��]r��!��fO��d�;��|b�u�l�UEGGwg��WTq�A���hg9福���6��=_r��5<
�&>�9l����S.��g��D$�T�E.t�t����p\!���hcŢ,xO�R�b����܉@���Ts3��7Р
��V�M�#���Ę٘f��&K��^�4�k��۷��3Z�;"��즳�gk����m���ϕ��8�ɢ�4�b�����0��?��qX���uKk�9��!�Q1C\&J�`� �ņ9�ք����ރ���{� @��p�Q>�F��GHw�Y+
,������/4QSX�k?arD҈[��qa�='��G/��5����HT�O���y�\�\��p�` RJSEq"��Ȥ<j$5�|��"�{��o���wwR4�N�P(/���prFdoYr��$g�y����α��a1�`�G����j-D�)r�[���sK�T�����LWs����z��4@+��mK/���Z��k[���F��@S���H[��dd��������s�/��ݝ����,>ZX|=���̯�2O%H�CNW��*(�AHb���0�����F�Q:��2B
0%e%O��q����I�݊aFFF���+�ǣh� ��ўc�封E�����i+ݨ�ݱx¶��yp0���篸�j#�Q�Q{s�rᜆ	M/�'�.:^}�l���ʶ,�cslsBn�(�:�-�2U�L��K�ؒ2?��������8�m p�������.�꩝�����M����\�4�;6	kn99�!y�M"��S�\W��*�@@�9�o�///���{��D�`��DV��� �
��~�r,j�Z>>��m#ZePvD���,)��/����3t���0�E]$��;A)f;��K���fJRCva*�I�����|@̑����w9@l�v�{�,�^�=�88�K�en�ΰ|F���'�@�"ɲ��%�Q��7?�����Nေ�ѻ`��og|�N^bۯ~5���He��>lt��oNnk��V�m�=�\����R��@�'W�����UHт�r�|����}��]��옃K?�޿	���H���L��?�;EH5ygD�j���f`^��r�����I� ��uʯ��؏瑴r��,*e��I�l�a�6�nл�+v��46+&]��1@>q��Jڍ��v ;H.����Oԓ�6��I���~u�F��h���4o��+��il5M�f�u�"K
@4�xWS�a?&G!�X����m5�ZZ�������U���)���[x��m?׀ڍr��Ò���7У��|eh��TD��u�۩�g���L ���)�ݛ��o�iʥ,Q/'Qk�ٽ�E�CfN�N��-!YV�J��9F �t��/�$��ʲ��eJ�~xz�S5,��y��C��yh��ڰ$�dG�������0���j�\�IB�ל��tD{�k��H��UR2�Wh���-B���ùB�9��"6�;�d-s�,Yrs>�"-О��!}?��3�+�/�!H8�f>r.���w�̷��p|� ��v�X�������L�"_���B��;�v$������{�<�2ov�O[�"�����f&��{?�Dه����q��2�ha�4�ITc��N�k�]EoL�/P�A�bd�n�r�q�F��	��#�����l���/\����Of��l�)�� d��ȯ��A%�-y55��u��u�u�;��S�1V:�yO�9)��EeFd>\��Fz�,�b�x%_��<���wfH����|�h��3��0&ܑ7��H��l��`_?/ʷy�Y��Jx���2/cs����,I��9�E*�J�I�E_����� 
ncc���KI���������y`L��^��IW�L���}/by*F��4�l��g��S%����<�g���CJ3O�[Z��5��$h��:LV�Ի�W���|�tX2Һe�늡Cs����c��-yw%��,26E�:�0Ҝ�
��7��;*�	�wOyG=�!� k��OxY�-N�^ݦfP:?|���c[�QՔ�w�i������1B߂`ZmWD�C
#-=���ѯ�֓f�#�4j�Ә�~��&0�2$jd���"<�ԑ�d��I�^t�Z?�\G����q'3�e�*�uk��u��*E;=�N�6��t�����d�JnC
^��Lz�+7ė�����I��<=-e[��CǸ� �R���^ W!�V	feOpc����v̚ۂh\,��%�ڄPOz[��d�yaF�X�����	�zVSy&���ҝ#��gee6o+�-i����`_��ƽ�b���wwfC��������������o$m���X�Հ��ҥ,�Tn��')��I���Tr���&���ÝƲ��cR����hhtk�{���(����~ץ����C�ny{R=[=^=�\8�T	�����n�L]Ĳ0V��ba�Q���2�_ř˟���Ӛ�F�c$�Z�mLm??���DL����of=]E�a�U��09]��0F�Exz��n��ݘ��]�Fܳ�X��[9]�Wְ�����4��pC �YDh>�]_�XN��q3']7�`�옷�d�U���za�����con��Gޡ,p+�b%)���{�|����(5��ח�4S��G���c:?�p3��=���@��I1�y��f�j�?�8�$w7l���}+��}��G"�`M{]�E�cܛ4�
:�L3��L�P�A�q`b)�>.޷�a��Vk:S��\B�(Uܡ�E�DT���م�A����xn���Y�iۮY!���T~�>������	X�x��\͞�*��b{�!�z��!D��u�<} P����Z�;�-�*o#��#\���/k����ܘ�Z�!�X�*�GqY/aʑ'X-�x�.)'���?����Zy��,Xj-�f�L&u�ؑ	,J�F���	ׅ��c���
@4="u����p��x�ߎh���Ǉe��r7�s���ܫ��&��$a���1f����.Ї�UZ����{�ßo!��q[�u�Ѯ<���s���u��=s��
���NW-Q�݃F6�A��r�FF�6<ɪ.���߷۳�����i��VZޝ�p���M�Mm �/��Z%���?AA��}#�Wԛ���H�Y)`d�v�+��ӽ�N`/�p6h���ٔY.����u�b�r����KY�A���Ʋ�P�����.�m!�+}�$�h7��ܨ���9XៀqX}��kcN +�'���z�d��1X!��k���m�<��:PWoc��4�g���N�y����̡��9�k�$]�7���#Uv����m�j\W�^��,�JE`��Q�T�oW��A,���'�|=��'��ChRK�denњ���8� �]`a=�1��:������̗����������k߃�ۏe��a*�'���U�^��9�g?��Q�>aR�b�XYYy�[e;]f�M�w�ߑ~B��r�@��h�����Dc�������0��ɫG�_^&��Pv��ݻ"B��R|�B�F:�o�+q��e��O�\j:g�^��<[^�����/����'C�O���l�/v��Xs���%/�'%v�©� �啾�n��@y⑕ҷ;Nod$�ؒ[��{��Z"�
�X���3M��2>YG1�����#,+aR�ķ��]�P]�˅�����b�]E<Kwv��`�U}�폖�����]�ew�2s��̕i��+}�����A��E$=�P����������M)�Γ���xu�y�D�N�#8��͹�0�@�O;�ߣ_��V���$�A��+����*3혧�쵦�}8�'�W���_��9l���U]N����a�)*(�`����@+�����׍�} �@��M}�ͱ%
��S�����W��.N��4�1YB/��vP�N��[������ޠ+TqG��
f���谰fP�ll�n=^���4n�,/��	X`V
�e�{du�+��NsZ#F�>"gr0 %�&T��T`Ӥ5�|� �/���ϡ��/Q�r��Ή ��7=�Z)�}��.�C$�	��z ����-A����\mz|/z��{�9SZh*����Lڞ�q�iA��S���YH�H�b�!�a�IH#������Tp�09=�	�h@r0�=L]%nNbZL�#w���l�)�S����H޿ؒ��d���m@r�"hw�i�)�̋�2Yo��jk@�{`�������1<�L��l��$H�nT�vM\���y�My�Ie�@H0��Vҭ\�k'H�yOTF�#A�W22�խO���w�e��(9�Rn�@ꌧi���!=$��f"�7�@�!�5�4�8\��ԭ�a��f�f��ee1W�߭��>�܄Fo�q����|�TY�+�*"}d>��Fms��f�Oa��B�����%M�t~�ޭ���8Hkl:EM+
�+JÝq_M���d�-0"�M/�ؔj�[���VCb�h꥿�z)���l.�}��<�G�H޲}?�f;}�+�⥥s�W�y�h--�����ZF�(�~���?�n������Џ,"o?�Jk��,UZ�x��v��茍�U�N�k����s� -�Wօ��.;��Ӓ�J(TO�����n׈j7+Ò��o�;�`��h�5ګ|F��@ui�f"��lي��*����]��>��-��y�Wfq�㛆/�#*E���xN$f��d�����ׅ��
Jj���_gV�5ԕ���
��֕�땪�x��������b��i�)dyG����u���v>�Z��<!�)��_���Kߴ�����^��n;$%*^c�2B/���,=�����8Xq:][1����/��H=���:�|_M�����	r�b�4��"�����	(T�&N8p6&&�gE)\>��6���L�D����]���blC�y����g�A5�4�d���%0�2Z�Ӿ�ʪ(ڀ܁Iե���=�A$�u�5��	�M�}Q�d����NY������B�-���׻����X�j��a���)P��뿇�&)Eˑ�i��an���+�Mx9��tN�M�H'�0���WJ�9���vBt��!����u���6#,��G
�j�\�vm��@LU����r�sq��ߵ�;*�cb~K2�������9mgg7�������ű«�yLxKFW���ƞ�K~G\�dl�g���]\Ssa�3ɿ�ߨ��+p�LX��|�~���(���j�k��-�Y:i/Nz\O2��Х��}�7��V�.�����zX�3�LF-�^9�ir_������2�4�,�f�U�4�ǩ����ScI�i��y@����Q��NHvNN$�Ʀ�Q;��F
��6�b2/�,]}��O)|6�C��>���$"o;[.*�I���Q��4�t�b�q:d�&�PE
�Ν��(�<���2�nrfܾzu_�������	�J&�+G(7B���I l^>�{xG�r���"v�]��&?���v��U��S�J�+�X�^��d�Y��X���ȌQ��7�������[��Yvw�`}}:��,�v|�8R��ق�%[�h��:ٝF�_]�~6;y�١l���i{�N���A��޽
-َQ1�%7�8V80`r�R �nC�ve)_\��K>>��F�:��S�M��
y2���koW}J7$�<m����A^�ʥ��.����=�w��.+�bUC��}�I��f��� �`�8X,��hF&��h�#�������2U9G��YlK)���^�#RR��K�E���	/������1��/����r�7�>�EP��&�R7x@�p���ano/�s�xj�#CYF�t�f�zc�жc�*"�[�B�x	��1E�¶dIH2��Jn;_1]O�<�5W�C�=��G_�
d,{���Sڬ���-��mX�K޴iSI��0�n��{����
�TE�b|���"?��0�����|�	w�g�.�F#V��&�>��l'{�7[�]9m�Y ��%����[�6��Qr����,��2�DZ���\�����_<F=����y��۴�=(b��Vbx�F��[u�����H��\�c�=1�@{>�@_��aJ�'��!U��q8�al�ȑqz��W
s�v) J��9�=��~@Ѩ�~��N�p�v�)6�}T��f|'����`�*:��R25c��>2�&C��*za�`'$�̟�v�Ŭ�����A���.��,,�䣞�3�M|ؠ����	w[�W�}����
�B���a�"���`#�S��Ĭ�ج�;��£���0X�^�HiYq�ۄ�g�e�c�TI��
�4�M�+s�M���8IZϨ�PDr��ў�����K�w��d���Ҽ P�)%�\)���!��/**�^��}$�>/���G��;�l�v�˶SW�6�������D�w?�Ea�r"��u�K���v,e�HD�:E�tݤ���]Y�M��.�R�,�t��'�����n�|����^$e)N�E,�{��8���-_����;?-�4��߮�q�f��%��ڳa�%$Z�Flww���5H.1m��{�r��I�!l��;w���7�;���0L���O��k����9Ӟ��053#���<�)xLBb����:�) �)^��7���{��г���Ff��8&d�%�3݋Ǹ�n���$��I,���k�a�E��(��-X0��=�g�s@��8u.�����n-����z�Ny����� ��޹��G�AR�)e���r`�ᙃ��r�>J$������CO��B���~��Y�|3B�7'��t��1U�����54�pqq��� ���OOPaxA�t�ڳd^ }}�x�6�5�L��� �'&n�F�hfE
�� ����<��H���>5>&��hE���4���Uss����j�'�c̋�.0�ќ����L��B��;��<q�̈́q�d}0&B)��<h�ƍ���@�Ѫ���e��6�! #�w+&|�1J�9ި��/���Y!xF�X&(qp+P�,l������"bV�
I|h�)��ՍQ&A�e�V5�T�X�c-��f�g.�O�����F|�!!��@�xf��4�����Q��7�2��s,{��f�>�pbeeg�:������a������
��NzT���Z���x���@���-��2��}^���]�h󪲅��\�֡�1o�V@�7qq���uј$B1���d~��
~�F��y��#;[��x_|��j�hw��v�+Gl�Ϟ��k'@�� L_�a���.�I��)�l�w#Âa�c�O���8��-7X-�g.�BCp���nX8#{�9� ���HE�ջ�28!zޖF�{::\��+c�������h��ڪgnn�]E=ѹ<��S{�S!~�VLW�7��$�,��s�wtt�����\�c��{h4MVz�\�=s����6p�݇��===_à�����Փ��)���M4'��i%d�t�D�tyQ��d ���Ъ�<7�!�H��*�1D�6!M�d�ک����=@Y�e"|�#{����۱?�5��-���T�R���|��cf~aA�g�祀��y�> K�I��¾>&���#���jl�UE�h17O���vWtt�	3y���C����;x� V�H�G�Gr�����[G��J�op�m;�a�g��ҬR��=;����8��B#�@�c��1�o�n+�+҈u��7�b��8�SH�*k�WN�G�����d�q�����14Wֱ��lM�Vɢ��˄�S�a?�]����>�촶�����*)I�F�6��fؼ�4�hn��N���}�\+QT5��?�:�6��t�Tm�D�F>�v�3$d�m�V�fb��<1-M�gv����]��������JryW�:hh��x�UtG�?A�"���3����p�6��\h >ؒ��y7�j� %�)ioz���6�i��K���+�c��Qe|B!�bء����*����Փ��B�Wh�N����K�������'0ݍ�6��L��?N7m$P@�1&��%�'�FT�(��	:M�?��2���U���}�����k��� ?%����U�ꂉ�����������*TcҰ�R�/J�\��#pB�1U"*v'��T��H;~������-����0����=@}	��
ВA���>����=�F`rF���1�E�|(�SE��m�@����6�C�rtrR3vV
��|��sW�;lX�|�	_Aֈ]�3��i��?b���q!t/��[�����m�xs<�B@o������zu剷�� ��u?�Z�L��[����?E�����"f9f	�����A�8W5���>�jH�޼���y��h��OW����P{^��$�"�:����X�p�`Oqo\����`dQ�Ճ����C��6I-'�bd�-?T�e$���##����Kg�b�iy��چ���|.�!�m �ސ�wF���{DpP��q�%)��V^�́ժo��XҚ���:��.���w,�#A�<� ��9 G҈U
�G���8�0F�{d�i�6��J�0@^<�>�O�LA�# 6�����=�U��r�?��Z�?�`c*\�fFR��v�A%����� ���zК�;6��?.���ۢMS�(3c��%� �*��-F[�)���g�hy�f3��Խ�6}`x��/��:lO����Q/���n�w��bn2|��2�W�1��*�V&�Tَ4�Z&�SB�!x�{��E���b.\�t��r�;�%�N���m�����A�'T,��$hhG�=�y�hܔ�]��������rG�ٌh�_J���^����.���ܙ3�Z|�Fb՟ _>-`<�٘YY+:y�鍓�'_^0�j<h�H�[0{���~?m��7�g��I,ި���������I���n<5��1�����2�.ށ]��_�����
b�,^D�>tE��X�,�8����3�����Zئ�_jeq��4]ᤠ/��C0����2釉�;���V҆�R)�]� ���0)�d`�i?dsO2_������)E)�NI0w�%Q#]'�|�`�	��Yc�j���eה;�3I#���e$��r<���x�&KW)��Y�Wa�+��B	�;<+vF&B9�n��'ɽ���&���{ϕD/�����L()�hG�3;SE�RXx�WY�P��k�g �M���\(/	N�W@�`k�2xz�{�&���=	z{>{�Ī���x3]�DnS�5��4�VQ��R�m@ං،T�����4�`L�&���{���i{��S_��a�W/1�O�]�`o�w��Gц�ڒnj�+�D8HX��'f|�v�'jj��>p�5X�M��� ��|U]�B��K�6rG��b���F�0�#""\Y@�HU�����9�W2�\[��)���1�W�����梩f�ٙ��D��¨����m�)�����
�Qs��+n�זC2���������.?�aw�B�:����L��6,��w������x�VS�O�C���YԺ�=f���[00(�~Orr�2K����L��X��{�K�
���cOR�-����� * �֭�4�t\&�]�� ⛅O�
�ذx�4��f�(�߹uk-D��)���� 8x���͛K�*C$]�ª�u��}qNN�L*ku�\6�fJ�#��=(5����Z~���WBq�����/_qv���d�y4i�RD�Wp�c^�R[�T��U�q���ۏ�F��	Fb��ѣ�\gÊ ~������7.'�~~��3�1Ug� BQ�n�/�i�_`�9�O�I�[q�yR�~���H2tv��/��	�e(.��E�6�!���Pr�L���,���v��s�;]�b��z��0[�G՚��U��z�?=d��-#����\�2)2?�N���ÍIxM��s��son�[��a`�c�ð֧�2/�L�����7zA�Z?l�+H[�vv1U��۳m��W`�'o9v�ϝi1%0�k��F�b��zϟd�qzg�N҅�{aU���LR�`�`���7@��T���M����.��'D<yUR��o>�=�Em��?rL(�L4x~bo���(w�����6r�N���I�NEr�B��8m���<%��[��'��p�Iw�/Y'7P�%�������x�e����f��Sw�и������;��Mu����X����Ζ^�l���t�ȕ�����3ݎ����,��R��^GȪ��n݊�/`104�_��k2�Kx���8�n$%)|�Þ*���m-�"�zX�R����.�	�Ô�2��u]����v=!�`0������ß�c�l��,K��i����"�+��vc�I��\�4P�:3SϨ�ÞH�L,������"r:J�8_�Wd"tfEF>�L����� ����p�����$Yq����$V
�C���2 XՄ�)�t?)1���B�B�b��l?qq�7��V�>w1���n3O7�W��@x� 嶤-Ex�*��\������[&��7� xE�8D��G,�h~ZNP��M�SB����Y������� jO�QbN�e-���H������ `%��`��8��d�3$!����}*A��;@�G�l%\�.؄k�􉲜�<^?W(~�
�m.��<[�	��i|a�.S6nKӤ^�T!KכvڢQ��YM��a�y��/���$���������6r�b6�7f�Bv�'��í|����v��A�h�e��š��4֍nÌQ���K��G��,�Pc� ���ާ�Aߪ�����`>��q��"�Y�� $�ԩSy��||"�rHp��vb�@`�1-�����|����ĭݟ �xR;��c����^����;X]�����%��D��
�MF$mdl��~B�L>��&����&��0H�a�)<
���O�W��׫�5��*t�=? @��yk�E_���욨�+�q�uu~i/!��&�}K�`��m��ok���iʴ0*�΅����{�f��07��J��w7[�t�C?����,lYdAp�s��I�ֹM�F	�
,|����=������6���.�2���5y]�֮X��Tj&�d���*��:,�ȏ�9<����%u�.j�]�v�e����a�g��5m�N������jٖb��_�� ���:�2�=��@\"���g���KՔ��%��|}�fh�?FÂH��'\#'P��4IF��?Q��ٵK���<��)t��SXTTt��<��6[������2��a������ק�] SB����a��A.)z�9�p���Czk��X5���R�:����Ae�]���7p���
g��a^���C�����7�?�J���_��K]�W��G$��t�6ƪ��C���槭xpU�4�ʻ_g��ϱ./u�Hs�w�{M�����ux Q+��Ex
�2)�u	H8� S�
�t�/�7(_�����SkQ&8�Ç�Y�\+K�Sj��d9~u��\�q��VG�8ѕ��sr��ج����֔��\kJ B��
%�ӌħ��u��[�-MF>%v�y��^�ڗ�<?�4Bb�c�����aEz�Ios�t<:4-7�_lҮ����!��Mf�?��_;<Jp��R����x�w5��/��{� h0 �AJܙ�C�H�%����"�y��$� "�òt��FO�q����� �:��(�����<����]�W��>��.�LSK�,�|�o�����9�M� ��<��*g�N6Z��.���	����ծ�|�f�/�{�t�X��?��6»���Z�.�w���tϮ�.��Uu�����66�%� �Dn5�3��tU{�g�T�{2�D�E�2y��؅m��MN?u�����Q�U��<���c1{-�]]�!��t�zuz�U�<�5V�������R3NLL$M�"i˙!�ś��2K�� 9 v̆�u�r/�zI=H��u1��͕�0�т,���i�������b,�$*W��=�@� �O ���q�ͷ_�
�I�8o�z�VK�!�/М�S33���0�od&ӜMZ�AfھZ�G�lW�5��ķɥ;��V_"�v�͆��z�~ٹf�,�}#����ov�WZ�nd����a�������Ӊ/����������arP���,Tc l�tf����`�r�4ʋ��QO�ż��b���>H�6>->���C@j���,��e�}))�������o�myt��~�$dvq��^KP�L�'�ج�m�W��b�p�O���Y6��NҪ�-5���G��NM'����j�J��J{z���%6��r|�r[����f�����Aڡ�,���f�C|�y�w���/o����޼sl+�L�� *^�n���2��%K��)R#�4���2X6��֏�}9ߤ����+x�2.�abZ�,`@��4T/V���%]c(a��7<a�f�邚ȶ�S�XRK�QG��a(�3�MX�)S�č�:qi�
�����R�v�ik��rt5�*��'��v��aǘ�.�]�/ΑNL�C���:����[ Ɂ�sa������>а�5��0׈�/�*֫��M^|(\?QH�P�`����Ç���R&OA�cͰe�5G܁}�eD�C)�#6�o��`T����l�����y����@�!����x�ei�5��v�lW.����
���	WApG!�i֦v��������L�"���6��Q��ӳ?�-�Gn,22RE P͸�PӲ�eݲdH�K*"���c�����C�E�v ݸ; ��]�[��?�~�R���nA��OҴ� �q?"�thy�s�dn���E	iF�hrrz�2KM0:�@KeW�3���3LȚƋ����?.V�Bp�x�315WE���3r�\��c�/z�~>`F��ggٽ0��[��N`���S��P��ʂh��>��?ءw�(Z��h0���)Y�399�{^hrE�������%��"�������ץ����٬gGy����j���]Җ%&�	K��MCq�ef?F�c��_�빟<�4�����o�0!k��վ�2�7��2�s��`��?^�J5Vx��J�c��Y��lI ����	=�@��e��!���o>*C�<r��?�h�-Ja>r7ֱr��������S��vE�m�h��9w�)�{��]��_ʿ��߶la.׬��#�UbXG<_���d7�h[��y��7����$�rcQ�3���J�q�d��:8k��n�Fe�� o>Q1�HTR����z��ʪTzeeէ�Ƙ�߀_����b3H"�yg<	�N�%i�Ƶ����A
��lŚ�z�"ۑn��{����~��Ƃ�*1L�򆽎�h��YDx`��Y�^ܴy��#X����w�B����ğ��mt�R~�r�����+��y\����j-�#��oE�q�yze<�q�&��DJu�Ԙ��� &y�R�,f1x�4"��s���29vb-2u�ϗ�kע�'9�v�vt�]���G#v����4����	�;+�Ԟ"�_x��={��H�c�^��Xﾚ�D�ۀsC����>BySS�=5|7��Q7�R�����i@�'+ӳ.�g�-�BWE�ZѲ~�,�9�ng���=:\�2�;!3$k'ç��ꂠ9�Ֆ�硝�툛~~H��kݧr3f�u�8���^���jO�{-��o��v���@V���C�&d7���m�]����ɑ��Wó/����qi����W��d�nza>B+�e9��lm�bz@�;��o/*\����RO{� �*���"�y;�HY��t�I�mq��T"�K��t�,�:Zl�dd\�ZZ�@�:���콵��$t$X�_Cҫv[�$͝��@@��"���U��`������odM^(n�V|hx�j3�@E
���Z�IiF��U?l�{m�j<����+�~0s>&���q�R�yk����P'D����Wc��7~��⪅`I��ɧ�6��'NDG`��>���%NNe�8$`�x�$˗��� �Ng�ö���px�4GG�վh󪘪{�a�xyy9:���t�����^��O��_B] ��7��#|��B��˿�W���2-�����i�31�0s����T��(��u/p�`	3�G�[�Ҙ]����`/��o	:���	��Ǉ����rz=�N��N`n�P����j��x��\��ҵ{u�W\��މ/����v��� ITh���C��� �1[Y��)|xϞ����p?�J��d�G�n��&��mYV���7�8�B��l��4���T;0�����~�ؚ�Tx3lV(u�?4!����f����V����
?�=@���;u��e��ؑR���yٌ�kƶʍ9m8_a1�A�ѳ����s�� �Y���9ݤ��6�f�T�d������a1����Ax_�����^�i/ͻ��s��3���@`
f]�Y^���q3������s�~f�����8���ǹ^:��_k֮7is��sj�)�|�mq���Mw������ռ�}Z�@<1.��fz����i���^D�����R���rN�Ä<�[�M8��f@��_���d�� ��t��ޮ(�����_���_#R�O[?mgcS200�_p4�ʺ���m-)`���D����0̰3���i�F$�uUXn4pk�$3'}�	w�}���bڬ��rcmO�'{ܖ\��Fg� 5�X�P��?�l9�FUj�Ȟ1;=M*�Q��$:j�QUA����x,�mH�~�+ى���сr{'@%	*���	�zp X-@�8����C�nq���#Z�����C�R~�L:
��:W�ֱ5�����c�3�?��^A�1�v�x:��x�E�r���	F5��X�.�����8��'ؓ#F�qc+�'�" *� ��T��~�V�<f-'�:�7(]Y6qsv�Gs�N.ߠFq�`ǆ�y�6_	��c��9]�D�ښ��{�Z4��Ar\1����M��ã�6~��l]���uia��l4т����9�]v��=�ѕ�7�k�A��JQtJ���|ie�����l��ů�ܾP���D=^�D���,]o�dQ����)+��řV�?��[p�hZ���o���Kc�Q�@�}��Y��P�����FU
��h�2���xg.ʄ�p�R�� ���gNoA���+�����g[J��4rB?���X�Nf����Q��7vyɱ���,-����-�q���e��:������xX%q�;:XCfaayT��+x[zYĲ_��J���,c�t���1��]�(W��} ꖜ�Y60`�V�ø�:"�T��Q_H�o�N@�����iǡP�hX���X�Uk�AG�<���V\iC��+�kp���)+�z@ب���e�X�^yNN�!����[�WZ� �)s�ssW�e<W��&���,l �ucc�t��-ȭt�����U �.�g]w��e�Z%�G�l�IN"W{w���jQ�xL6*���P�|w��y,�~�L��Az���zÇ�lj'\��;v��m0&�%&&1
.�t0v�ZRE�]�䴶��6Ņ]llؒ��׀W��p�[a�=�l�y�Ȯ��X�|8}��@^�*�z��ږ��
sW�9a��̉I�����1!��%i���� �ϰ��1�4ܯ�V�h�����8��ݕ��Z�\$i�����a���缼pزߠ�<p�N��g��<pK��{��s���x����E[g3o�Azz�pS�
ox��\��[��Z���}5�w)�&���=���9������ޫ	x_�^�>Ӹ\��$��߻A؝�j�����k�I�Z�mڷp������]㛛{�������ݗ����;�R��~^���/����&�e��z��Go����(�Cڕ���4�d���+�m"�����B�Q��c^|���J��׻���BB�`�����ɰ񁮢�\��A�/�;v�<�å�������sp'{��%i�����tZt4������?8�Pe���>lQ��l�樯�M����&�?��'L�g��Nxz$��fUد��z�Å�A�q��ә]
 _i;��ׂb��r�&/O����g���K����9U[�j,8���Y?6�ћ���H�E�]s��=x��eJ�ȧjr�-AF��i��˯�s3Z��߹�ٿU��9��)w	a�-Z��ˉS֔�i��y��x���V�wG��G���b&=n���j*o�tPTT�Z���J�w<G�w�aL��s=�A����}�Z�2d����ǞkE�d�W}���_�ҡX�	E����t~�K����#���*akN^ay ��i��O՟����q���w�|�n�ڷ�3&?�p��3L�M?O_pD��ʥ�nJ&H�b�9J�ܥ;��'$�Zw<�}������c�~��s����Lѝ~o�����=���c;85X��Ln��d�o�a5�G̛�q`��`\�������ԥ84sڿ]>���汗Ns�]ͻL�U�/)Ӑ��1&_Y���}�(���#nǦ�=;�+�X�_�pџ�?��K����O��8���w�w>xI�v����I 5Xܟ�.N덜�b:{U/�o��9ⰵ?���>�{�A���9N=���B
L)�Ռ^3���wa��gnf�5(N��v���-O�s�x�=hI7�rf纏����W?j�0>������/e��-za:�b����{�k��������5ΘG��5ȍ��l�vy�V�7��1&�_���j\'P�����
;S?�m�k�gbb��4pu�{�����8u�FF\#bMk�Ӵ����7H�H���J��@���٤������`���|Ϟr?��̣�����-u���g8�K�D�]A��#v��_Ue���+��y8y�,�k��f��l������o9[2��%EWռ�7d�j���d�CSk��w�9̤�OoR�]���\dpD�C�tD�p	����_�s��I��kM�7lؐ�8�6��z��܇I)�G�v[F�O�2;�����*a����g��fh�!����p�'�r�˧W}�UH��>�rwE��cU���6?����0��qk݃+�Zo5�ut6HV��L�n�������Mo9�x���1��^��?dF��ҽ$ey�I�i~������G�!p����zS��)KO?��*��/c6��� {�y2F)LU$�Ar<7���� ������٤;����8��<=�����w��eFe���[�Ԩ���M߶�%K��(o����7}�?Wi����Y�����3�b��W�W�d��9mC_�UT+1�}*9�奤l���'1���Й���aw��g��x�x+h�5��uKD�nc��$��W+�z���K;N����r��
�g��A���D��-��k�v&q�m�-Uˈ-=�Ƨ泵�,cy����>x�-���~:���yzp:%{����gk	韖N�j+
��=��b#O��*��𒳡N\��w�4j+9"vҸ�=����uG��;"��/�V[['���	�&I����s��ǫ��6���`lM���zIQY�g�3�iv(�?��u��˻�i��.�R@���oUcM\\��9�������C�*:�����a�+��z�Z��G]���(�LO�tsVAd�id��L������)σΪ>���O�ˣ/��>����
�L�����=��e����ۼ�,3;�j� �?{Eo3S�p�F����7v����o�Iφ�-=����/������4ڜj��0�.�6�����R���p��}	z�jit��_��$ ����!Y�������`~P�m<�2c���8�$�k����x�n	Q��޼3YKA�Z� �����\�յ�~����t���<mӮ�<�9���7�x�ݹ�7^j�F����|Pz�9��{�ii�+��T���:��>���r����t�qю��M���A��בg|�s/p��!I�Y�G=~>>��'���&��g���Zh#��\�`LؽyE�VU	��SJ/�r�@k۬7���v���&''S�L�cZ¢������;�ͫ<�*˃�lb/�b"�1
�4�����=�I��= 䊨����,��ߨn�D_������p,����T�$IFG�
��le�gvvFh����l/�+�!!��MIVFF����}_�����s=׹N�����s>�w<F8DM�b���~<s�%��������Č쨳�S_S����"֓ٓD/����<7	��<����Q
m����hC�=�K�~\K� Q��7=e��{:����*-#�iA~���}F���hD~6Z����>��IG�:�������/�����b�2�ѽmQPD$�������@g�@�ӹI� [+Oi��L�� <��L�zg��S)ޫ�G��=��o�����ks��T����Mon�0{s���-���Or��h�X����:������r��N�_�
F�sTA�9^%���f�	�슌���zeBu����������{�K���oԉ�B��=��H�.O1F��`��Vj��~G��T_OQ����/�[(�NVp�b���+�MO�w�/<�Yj��C��Z�����b��ϓ��n�.r�"��"�_�$�IJb[����߅�����Ӑ(\��9�vs��P=����oԅ��F�B�kK�n��L�P]Q����>�}��R7�
JK �x��?=%/��V9p�'�q7z�ɉ D��Wo�{���B�}�6!1�B����)��|���)������mm7��4�Oy���5�T7��`?��8z�<T.^�(�}`>�m�sm�.^�"���_�!��gzĚo`b��־_��Z�������c����Vy�-)kG0�x��,��fa�#��	�iߕwB5~���^�Q��-�8����s��P���S�"��c���5���Nc˗��6���q�}�����pl����9�i�����n�����h�b�2~��'u�Lt���@�h��q��06��Y�H��R�zg&�*����)��1��)���	��o�OIVqfLN�%���v͛�{�g�����i>~���"�{��彩A�נB3��5���k?��sO����f �L�����I�����kP��U���������U� �Ag F��C�k�]���M��������s?�kfr@�:3_L��W�'�q�B���`T�@gg�6ɕ�J���G�D��3I�-^I}}�?�����
��jL�Ŀ|��#ÒjR�i��؜a����z����/7�gU�6��s�,�s*Y��Y�<��:E��W��P���{�����賓�����߬�!p�C$Q�nN�W�j��Y����aGʫ�ˣw����{��FMvq����Xx�E;!G�^A9�p�<�_�mp0�������''�B��|��!R�eN���}u��_	2�Z�p7Qx:1^t������f�&A���,q�ש4ҹta�%����p:����߮��<�
qz����bu퍊�D������Qξ���݇�޼��*��K����#��:$�O~{�ܽ�@��!�ԏ8hC�������{F��L���Ui��k6�rZ�7BЉOc˶|=e]��Cc�6/�D�H��{��s��S�vΏ��~*ė�*�����.����aA ��C|\��Q1|��9K�e
ܙ[�2<-[O������=�BK�����^*,g�;��;�`�����T��cK�<�Q���D1��t'vxH�߯��j6Zhw�`�6�-��P(���K��\?�.�����{�K��4<�Ć�,36�}6�����2'���y����������|q�}�&�ϼ�ӦW��Ry��lB���)�	��p�4I��/�c��g�M.���&k�(�?(N����isy���Ə"Zn!��{���:��Ӹ�����yj�P]`]r��O����$^B��+�A�C�,�iѨ�o�y9�$5L��#�	���zc���_��`�����_�ec��W/��1�`�>����$�`������:�
O^�SG���������f��L_�����f�4��H%v����/����D�|�F��k�89S��N�1��]5��:m��!w~6�_ ���q���2�MW]M9LxAQK���l�0G�J7Y�I�~]=��CJ���p�������Rm�D'YG��q�YT������6'7�!��f�Kh_T��]M��|{�o8����EMI
=�����_����_�4~?�@y�%lowp�c޸��S�F;���=�g���z����m�����w_k�jre �rӆ�̷KX�.�Mod�s�r'�� %ѻNb^���0\Z�.p������en�=AnR�lC<	߶���x��LJKο*!� 1#�U��M�cHW�9q~��qΔ����Զ͡��L�󝕄7U�'2N������Iݺ�"B��(�Hcؐ�cI�}�R\�C���f�{��t���
\�?��ü��;��P_��QL��X�{�ɵ��j�i D��,�[�/d��hO��9(���؟}(Â�?���uʸh����N�r��a�����'�����sE�ox�:�[��5��Kr���i;��;��;�)��w��G��	�~U{��9?�Sx��v-Ƿ*�p�+ �0!�1��묐?������]��ݿ�xl���G�|��bhl���Im��� :,�q���$���_�o�
��4ϝ;�,�9�O�0�JjN</|�^ۄ�\.��:�ȥY�B��h�L{�����1xE\.ؠ��k,c^�������V�7�^o�/���$�{��}�sR?�h��*�����Y�<��\��d�5֗����7S�>�ct������m#��W'P�p�����z���TI�"~$�C��~�3>|t"�6Y=U�nʈ�c�`�h����@j_��,���`\���X� ����c��qζ���'Z���6�A����d�6�o�=˶����&Pz�,Y�⟠�����P���Sh%*ɥ�Kr��[�xب,�J*̚�����������9h������v#�<�%B@�{��鹶	%�?yT4!%E���T�h�V� M�J8�>һs;3��I	י��鱵�t�]���ӿ�%��cup}}��Νݩ��_|�!w�����"sߌ�{����'t�8=�;�a����h@�)bzi��u5���J/yT��C��A��8�!G�Z&�*��<���7�Hdй���i������O�l�����'�ۯ���}�;y�Vi�M�b��fT@Eo�Mz�+�d]�v��d'��<��|�&�����W�v��W�Q�TU�{=W��<��ɦ͚9A"�X >����neg}_�{Z�]�'��e�0�#�^�r�#:>TS�co<(Uy�QP5�c;eX��,�B����=Ē��0	��P���9��Sd��_Zڨ(\�W~HR������K=�CRW'9g�(;ز�5���^*�[X�*h��Ə���lm$܍��ƅ����w��8��q*?I�bf#��
R6����ŕVT�XW>Oq5^I~=FA�v���CGnj�,��[���-���8
W�a^�F}/��z�MT�d��㕸�Z����OD�3����K�LF,N�9�
(t�o�'���Maˇ��-n�D�	�k�.�G�Ug_m`/>��v�)I:�$E�Qfއ;͆3�10ɝv���NZ&ݬb�QQ�i��i�d�S�{�	��&
'���ړX���@�J��U6��u:!�VYy1�����
���֥�q��|���o7�.�R���㶍�����p�T�St��Cn.����ȇ6���Ʉ����\��WJ� ��^�*)��e�����jGЕ�@��G�3N��{"��ݸ��ݟko>��|%�jw\��a26���l�7�s�J�6�]U(6Yi�:zݐ��/[ƺ�V��m��$�_P�NR�+���1$����~��8K}@��(���L�=�:Ÿ�FE��o��:��u��WD�B\�I�/1p�P��ipSnu��u#����Z�d�Fvj���ŵY�:�N�y�uG��|�j��=B>����$�mk��D��V�� ��[���4�;��'�h����#�� x����.̼��K�]U@#����vR*��.""R�RT�H]69%�5���$y`ʯ�����G%���^�/�7��rȰ��q҇�;99�:�^�e
�<{�ӱ5=��|T�%�p�`F*�ϩ��5�_�ܴu���!K�x��N�����L�Az�f	�n������_��o<d�&��[�y-�455˥qцN��>=��J&?�=���*>���+/+����-�3c��&�֪����s��E�v��l?3�k�PH׸o������(��c������z�C�$1ϩ�|�����2һ׼��{�4X�cu�A�ʜ�[v�:黎�mVn(��u40������H�uu�)㹄�� ��}.s�j�L���J-v{���ч����:y��os��-R��>ny�v͟>�*�U�ua�6G'7lYg���N��hP�]H�uU�v3�_	?���~L�k-zeU�A��ӽD�;3��"���	�*�	P\���x�pQ��f=��I=�mY����$qo��Ռ�̀��Y�n<���z�sdt"��dUԦbo��N�v�	^���&^o*6�ލ1�^�-����m_�����q�%-vzj?���j��ێ��IM13�_�u���s�-|uyhS������������F{8���Ƥ<�������=�?cވ>��yû�;m`m�u�qi�/���#Aq��kV����j��g\��7�ϱ��'2,GQ[gm����u�֓��2��x3�x2�ʆ���-�7n��AJ�%n�Qr&�ۑ������}/��Ctr<���K���/=E�V���?o�<�u���V���O�I����w�����E��ͼ���̕��=�� rvlل���蜦{6
�*_���]��ݳ�ؠ����I̸�����m$\8�~���&��e�Q�r�N�DҞp�-.u(�M�n��I�	��ڢ��`�ݜ�y�l$m��-�3�!�7ؿM�B�|vݎ��faeL����w/6���pr2.e7�۵������h쉼&sV5YH�b���X���K��#A������+b���;�(��!����n��Ι��:�7��&(�վ����%��îD����t��b�0)�t!�&mllB�k�g-����	�h;ym"=Τc}���{���bC��کjj�F:Ž�A�/��]b��Z�_պ족��D!'�s�U�L6�D��Pu���C��T
��d�K�/���:��������DH� ���5i't�f�4�
j�_�8_�L�9��Dr����L�b�~�'�z�)
���X�ʪ|���^�K����ָ52*��)	���0RڄN�ٻ
b�϶-��y����:���+N09m׌29�Pc����D���H�Wzhg�Wz�_�3�d%w���Ҫ!5��W���o����T�.�g�jRn[�PE�.t����iY���K^j�Ƅ7����s��� |岃��MTM��N�r\RU,�Bq
��IZ\����1ڪZ9.7J�R�J=�O>����這�C�4 �1���	�	�������:�Ie� �#�%�s�b�??�D(��h݌u�5(p��}���OYaQ��)
\5�'�0=�kd�1a:ame%.7��1�V(��Ԅ��P��j/���0eL��s$�Q�'x�@�|&-N������E�?ST� K�BKo��_��Q��ڐ����P����٭&A����{|(����5�m|�j6�'`X#�����>%V�CR��'�;��fAg@�p��t��ri�
�ͮ�^~���������IҒ���ȕzK�L@g�u��&;}���).|�ϑ�	%eeΨ�O��:;n���?%�2���,��&�m�)�7��R���D��"�}�4�QH/�"�p��+�x��6���}.��
&ٳ�������7L��Պq��i���˜@��$�g_�����L�M[GOq�	m�{����,4s���*Kb�o��/�(%�/-o����C/6�����ͪl��*�@7��dt���(���V��S�a�G^�Hlm.�Snm_������O 8f���[�����:ۿ��S��|��궷�b?D5��:�[�+�(���-��P�C���U��i��恱��E�~���Kl�)h���Ռ	��q��s�%?��R�2F�("�X�$����+�m�	 �+���L<:��uks}�xK���8�3���e/��ۅ|@WkS�i��Xp2$5[O+�����g�U{e�2��?���&3��)�I�h�du��]E^��'yau#��ln��he\S�#��<Ċf���7����'gʇuꆩ�;�57X�c��zM�,����:���V�S/ֆ��u�+Æ:���`�s̑=w�f¹�b 
���{�k�AH���	�4Y	
	�f_����<�vUa��'�����`
ϟ�O"�����Q0�v�6�� �8 �����u��*�!��ԝGQ�D�������.��Vsf���x�+,c����L�m�`��]Xm�]~���<��ْlP�S���T����EM(�j%r��9]Brr����/�#~9�{D8��U��0�*��l ���������I�JA�A.�YNql-�ې�������??\��i%pRr�W����"��PS�10�,9U�2�3�Z8���F���#,\�||ƼǾD.��N�ۃ��
>�ɹJ�J�pZ<\���(:�x�ȍ4�6�W���u4#^N�+2��.0�����\�-��+�l<E���$���c�ȇO|M��;�[RTD��\�ͽ��)�$
���t���O�K�c�Vs(���!���7π��7x���{��onڔ��46<��T]w¹��eEd�x���9Ӆ ��� ��yⓟ�����X����K^�ڼ�_���`q~x�r H���0�[���2�n*�|Մ�e�8c� Gm�Q��|ǃ&��Vd��w싱r��3>Q���}����͉<��9J��d?J�̛�A�,�ϔ/�����1�Ӛ.$#3s�'Y!�)�ZFb��2g���u�pa��ӛ������EW9��.�����.��v�e��K`�y2��}}}5�����T��7�W�HQ��j��@�3‧����i��� ����
~�����:��8���x�����9.VS<�~&|j����f��.�ȭ�L#޳�����$�ʮ�K�H� R��p ��we����Z����Rkgj6��O��~;��s$��,J�h����8J&���5滨��Y�§����]��Y�1�1�3����p鯿�Zq���KIu��^q��S��&�%�nLHH��>�?�ArQ�!R57�Q2���M��Pu��w='��x겇 ��a�������`��6� ��7d�ڄ���!��aZ�)u��jA�=��$$�'&�����@�&2mK��h�0��P��Hm��[�H9쵃��N�;e�ϡ����7k��`��!�r�w�D`�S�S��Ԟ�������a�d]����eLXYp��D��P����4L_�
 <÷:MJ��\v�nqE��1�Ǎ�ޒ�hfWb�	K䧝���t9�ʏnen�)��L�R' ��;����;�]Cè9���H��SKk9B�k��ݺ��|c쉰O�b,�ߝ��8�z�2����+�I�U{��M��\���)/S�ou6mU��:���¼�a��n-pR?�Sy�
GJ�Ebd��ZA��&R,�������Q��ĵ�/�
R�s����+ks)��/���:�?�Ҭ:^x3�S�<o�A�C��2��������{V�{�M-��4[����u_L9�qq7Ƒ3|�'m�`�2�}]賓%~�Xru	��>�9%�y* )A���������ǐ�1���]#)tk���>CU}���~�Q�x����b�5����2����3��o��5���J���g���ůt1Rt�,�l�1gᙳp��:u��?�)�[w e7�W����hjjB:(/�Q\���� 57�KjP�?�yb$��ai\q�r���̝(�<���� ������#Z�e���Mf�Oc�@���<��� ��ϕف�ԏ�l�R�(;?��k�۶�Q��!�b,'N��^�|m�?��S6���T�������b���0U'#�� �#�no����_�G��iUM�Zm��ˋ�9���VC��4u���i����lQב�����L^�Sg�k�V����լ,��m����E<p�E��e_ӺT:?=P��~m_B�L��W9�<is�+U�Z�<v�L��dʰӞ�q�c"���Zw��5P�w=�z����:�����w7	hF���~<D`�dChh�yc�S�4�N�(�u����,&��{�v��Ё��'�n�esi�8���� ��Q�|ß3q��$���a��B4�	 HG��O���ku��:^j��K�,��i���m�����AZ�����W�1�4�/e���6��S�|��}A*�6��ތMq�B�K�ē����z:>�l�d�"�zV幚T
�e1R��������l��S.���\ް(Q��k��X^^~=J����`�M���e�L�9���7�4�<�#G^[�Tm���y�w�K�0Ĭ!�Mԏ�C��t�:��~&����F���kN�W��,�{j�X�Bvz�=nO�^l�2O/���.��t9
�۲D>�9>�]�����hsH���%v��V�݌��-c�?h�}��h�
�B[��<�������c�AcA÷-jek��"�p=�A������64����V��|2s�A�s.�旑E��js붖nK��f��?�=Vȉ�C���)ᴸb:��J(�W�9��|Hh���4�!%�p��ʰ�B#-B*5����=�_�{qq��.{�H�����X�������/���5��%�������K�5֗��~H�խ�yl�-�3��>�a�H抃�C_O�~��ˠ��arP2A
3�V���@���&���:�K�x�����E_�_L�a�zU`�_F��+���8����k��5^�:���($�N]&����SI��� U�j�±�k��h��J!�66�Ї��M�	�8�} �O��ϟ���kg�i  0�_��n���l�˰�����k)۫̄�m��?���.�ޅ>s�a�E�M�co���**^3}B;�\�G
|~uZZZ���˛ߨ��͞�=�[��h�K*�N�qb~�����@Tᦣ���
�W�e#i�ND=��\c��GK��7�<ǚcΙzx3��'�hqY�A������Z\铓v'C\��3���9՝��%E�3��i��Z3[�#��-�;��D�&�|___,a1b�DB��\��u�~��T��d23E����9	Kn��c��%�N�n/��VU��k�Y�k��(Ґ`�%U,��)�鵅c���=��R�P �G4�;�۽�+�Y��[��~u���Ի�\;]��]��v��U%14����Ǩ�y��	b�뭭�ϖ2V�vd(�>2���.¸ۿ�J��UZ�ײ�@����C��)~��{.��g׽���sT�����UU0o�?��8�_�Z����UnQ�LNN�MǧO;&K&��/h�YWV6������E��Y��G�e�B$���zn���K���l�<o�CF�P;1�U����yK"���<�,�<Fd-E4�i� ��Y�j�� \ԏ>���ٱ��x��u{{��~��B&�{hԙJ��ȕ�ohU}� D��?t9o�Q6�rii>��r���/�qg��v�Ѝ5�������U$�b�Kf�|�(�x%���w�>66
�?��/�"�v�yϯ��de��2�е%��@���qr���$F5�1	z1[����e�]]���ʪ�����֜ԏ8�(��~� ���sysK����&SJ[�SYvv���]�x���s(�U�����?����n�Q��by�>5'�+��?aaa��9P���Z[[�R�8���V�6��CR$�_��tEKQ�S���`��e��A���s� 3���c��|@�/�QD7{�ױ�7�eL�ϯ�����E�{���`����ٙ�4��,�m�k+�}ܧƤ������dFƟ�����uy�min�SYd���4�͝��;�\�#�@9��W{�:`�zx�Wo1��վ{��Nx�M`K��0��z�uȚb��~;U�:��G����y�>�y�A�8P���ۋ�l��6Ŝ��G�� EEEe(̡��Qu��畼?ޕFu5�.Cm$f@KEb]��I��nC��/I�]���ᜉ�	��^��111`��ri �H7~�d���KY�:%������7IY��ĵ�$���9�Ž]Q
�Lz@��y��R���
��w�WDcZ�K�~kk��sR���T��(��2��WVZ�U�p�ޗ�0O�R����YJ�h@���oj���WR���YY�����)0���ͥw���S��a�sW��(�=Ĝĺ�+��:;9b���MV���瀨�)��������u�I8�I�s�֠4�ځ]����xJ��skj����0���Z�^@�o��;�"pl02x�-�gve-88gZ�f�~����/2�ɉ�\NLLLPH�Z���.6��i�M zK<-�:����s������Z����=�7R<F��A,���IO��a"CjL"��E�R)p�����#p�YB�j�}��{�h���!�G /X؈KU��vB���Av�9W�g��uujri4�����^GaH}x�&�����Ǐ�}�� ��G�C�A�xΪ���ru[U�l��'[3.�>]7\�Ǔ����u�>��������`��T������|�9	�{z��M'�N��\N�|E����%�1�'�)��f��/�Qx�tϔ`R���MĊ��w�~Lm�f�+5��CĊ�l��*�mi�S�e�I*X���r�8k}Y����p�p5��sݦ�O���M�%���|��+�}}�<���X��g�uPH�6�'�أ����g�w���y���o�Wh� �����|^�6�¡�������k�4'�$"�b�X���<������9�g�����]Z�=0�lR�^+A(%�,�]��_j�_�{�Ճ�j��~>>�h������*����AyF�ܺ�Z��u&���SQq�|�r���3$5���Y���3��n��� �������6b# ��1�G|w���� U��= دP�;��s�.�L��.��M���ʻo�(�Cg�� �T��L�yS��@�|�'�~7��`��Aon`��wȐ	@wM���ߒ0(s<Iذc$���.*ػ��Ƥ ������%�2�F��`�-	�A�~��j��3�������%u��[	H'��s�a�ڵ�f�9�,G��i����i����>�ַwpЄ2����X�a

B�댸Ujik�Ր�7p!� ���m�:?]�]
<\[k�ض[�����O���v�f�jVu�a��G��� �p[@Ʀ��aH�'�#�}H	*l��?�*�+RZ��9���-������ʱ��?o����YS�u @��z��j������A�h	:��*�[3�o7�(c\L�59��>|XV�A;���2p��2a���U�M���A�o&o<�.�pd?\��n��ek52��1B0��)��p������q�B�;�Vj�ف,��fe(P'Ooog��#��?W��ϟW�8�v�ߴ4⍃���(�|E��[���ְ N2���(>�?&a�f��Dt����Ç��zMJ��	#��oIpqsG��W���&cX�~��գĞ%�E�{
�A"zx|&��������cccP�_���]@k�1som���Vr��x㦋���kk�Nõƀ��H�f���#�`᪕!?P���%p�����8+�:�ekvv�h�Le��^�g�k��P.2�ձM���90�wΰ�"�Y"t\�Fy�w�����@�w��̴�p���h�^	�(�� :���f�&&�&������naq�X��N��/n:
.:
�5Ӟ-EZ��و���4_"�8Z��#�)����+��g��@�C�l]Z*<( �2F��e�/�{�N���q�*����7p��<m�t�D!�o54���k�wq!��YU=謭��Z $±c� �3�n���~p �M�:?�z�bY*�Mcf����rn�h	{���%j���89wv��5xh��W����y���������q��Ou�5g��!ii(��S���3��/�9�5�J#�/⣍��!�31u���>r�C��ݣ?yR�=�<��P�R���\�w) ��^(p�����2���9~���t�.Dc	^�щ!�=zgz0�8\3�v�Y��u*�����9A�}39�8�ר�Em�j�nnnNMOR��Y���mh�[U%���M[����kG��n�9hkU��`q^YI�#�%>�S�ҫ��Zr���
����g�D	�|���g�޷o�ǟ_��KKY����_�4�sRG��ۻ�����ghz9'?_�['����ܝ==Y�-��[8d���Y�?�X��Ç=㗑?����S�;~0���7��,�>����أ�:�L�2B=I*����ZO��������U��oy�2�Uɮ.�)�$��Ii��CKa��� �Ǿ����
rgsw)�"{:Y^]�s*ZL\\�9Ǐ+�І��6� ��0���G�}a�c+��˶���SSS�SCP��"`
v���ay<��!K$����fp��&JVb:ğ�B�B���Ag>)L�w���� �������'/�xH�4��Y(��便Bl�TK`�h��:��*��X�i�|FF3p�������q�|����*-��b�J��|} 'Q��號bd<�o��ȷ����]����;Q������i�!&h/:��Ǭ�J��ݞ&���:�Os��f�?!!��DDr�I0X7�$B<c���n鹼��%E��Q�AL�2��*�S��zϗ#�����:B�7��>Wɤ?u�s�U�e�7�����F��o�^^^^��yS�=}��ȋ��xZ������� ق��*I��yH`.=B���'�,�r���D{����ث��Ej|KK6}����Ȏ"몠X����0U�$ǌ��޶7��+�"&ְ<'#����K�������Ի�C����)�*t�D �h���9PM�ܪ3�va(���f*݃��7E���t�Vx6<��������;���j'�;�p8�m����ϐ�JSGL�򅱒t��U��NN1���4Kl�q����$I?HUnG$�Jؚ�x@�e��^�`��u��=`,�7�\��6?[��!�E������{���t��4`X ���!�<�NS�~uV��+��W��d��Q�̭�P��/����� kD�%?��ohٶ%k��F�$��kf������ཽ�s�TWn�E�A!!��o7��yf	��Ş�k���v��҄��3~>�Ga�,�DaD�U2q�j�b>���Ô�\��<�Natx�J�k�"�]]]�..��o�����":���~t��ڒHJ\!?91��*9tgUV�ࡀ�FE9��(����(���5��������H4`G�`�����C�[�h���X���a:EV��ϭ�-0��{����'��v�:�H��hiI�pcHJ��Ȗ�N.��Y�����Mԏ�O�q�n)*�_u���9��� ��0:�IM̌�#��F�����L�jռ�G�s��aSH����4�ݍi���@���o�.L=�����^ r4�����έ8,Ouӎj h�g��߿�]�a���rre)G{;;u&y�g�7�=��|
�n�ۛ�h��''�����V+I����?[�����$����Yp���Х&}q��;F�y* I0ߏ���d���Ǵw�.��c=�A����E��[�q=]CM�1K�A�߰����ʃ���Н׾�<]�:*�����a���J �	��'����y������9<(��FJ�6wK�����F?��]�S�-� �7X� 3F!�i��L�ݹt	#��w�''=PU����B��EK++�puH6PC�xL�km{\z�c��]/�#�]DY<3\g��gF���#���u����3?>�sEuZ����s��[[�E���Ԋ��0z�m�P��P��}��J������eX�������bԷY����,c���"Q}a	z�҈�1kB� r��M������A��� �6D Z��\�H�Uշ�04��?�ԦV�81�ʖ1of*�7S�M
t�fw.��_��)�el�mM������,�($j�	��Qƞ��ݭ��a��K��1A����kʘ�Z#�v�cd�WQ��O�"D���,
ʰ�BK(��&^m�f(�����v�c�/0v�����ۺ���g�ߑ̺�����|�7�09��]!��LPkOd�#j��D��	��A�*�/�9L�ǙX���A��/�3��)':�"g53�KKˏ-��F*�d����Ff��ؚkT�&��ֻh�D>��7����>��8���ȣ5[k�hyճ���6E� ��>�6(��ԑ犿�e��=5�3�9�����f���X�]IA���C0����_�@�A\����e-z	����/Q��� �|$����:��+W�i\ �uMok��k&E�=�7Q��ϋ5���`��i����~.��&��f�w����>�\E�Oz�z;�.�e&��V�j����oq��G5ѰWkz�cx��|v.�>��H��[�2O�ݽXk`-�*�� �֝�Nr1��!�'��?7(s�Gqk\��Is��CL{�1�x�a�Z���ZP�a�w�/���h�q��m��}qt���e�������j�`�p���+J�fDVm����p�n�	(�0�����ç��.b,ht.����7UPb��[�{Ṣ��䄺@�N}�-EJ������`�h�6�K�v�DV~~7��[�	@�ܤ !�+x���]�w���u�&K��@����ۅ��ۻ��8�r�@_��b�ȇ�	�i��nG(_mV�p@�߃��8���C��]Bc֔��%p��E�H��t%�_�e�AO��o�{N��P1�E/6iq�ߒȇ"�*��g��7&slQ}��R�#�� �E<�GHJ*�-�G�W�R��^G(?�C5~]CC_��1������+o.��u��6��ǀ�K{�����41�����:K$�X��M�� ����t������5&��d D�)��CA�P�����Ѧ1��8W����i�hU���ap�-�������|��]�or삂���W���v@��ywJ2�|�W�, �6����l������C�@h����c�n�����}���@��j�,����N'�)���{����Ԗ�Vj��
��<t$�Y��_��x������B���H@h���MQ����~���!�;��O�m���%��<_X�9�"�!F�zD?6��u4��S`�$F��F���(�fc����4�d�����h+�P�'EQ >���#�� ��A�P?�I��eU c�{.�.����#������B�^kq鴙��V�JKK[[.�B����S�l_3w{�1�ԉ�J!�P�t{�v_���0`ǨW=x{ep�1z�y�T������n?�����&h[�pXt] �h�I�$S�pKKK)<(['�{kO���/�)굹�-���";���d���2�~��~(#�3 �zP'�	h7�\\ 9�����ugT� >��Y̨�3��`҆lz��*2{
F�dU�ߛ��	�.���l�u��r��b��
@#��
����D�)����\k�H
��MF����u}hEjf�&�v�[�A�� ����E���0�=/'G�y��|��P�秈F���+M��s����ǏOe>��g�F{�� �e�F��(1��B-�|�\��!������!MU9��{{����������l�\7�|�+gaD�2ꐉT
�¥li'�<�2�6*�e	�-1��F�7N�ҁ ��qvg.B��J�aI�a%ǼX�1x;�m�7MF	�X$&ϝ;0-��6}p���!��X�q�-c�]/�؛���53��w�Y�T�h��s�\����U]@�:+���j�T�<�QM���9�����
��)m�j� ?�z�w	qR/�&��^���,��_�T��S�4�
�F!( ��6�9� �ޠ�@?��|2���P}��J$, �;/,�uV5��\�0�?qҭr�7�l�Rs�Jhf���n.U,���)����Iw������*M��������+uۛUc��
�����#�����_��Ä��Q����~���7*��p��%��7M��b���^�rJ..����H�������(�"�����ꘑ,-� p�U�f+�i2(WUs�����1f_��yxyM��&��Nr`:A$-��4j��a�Kp#�Z� n|e%p� x��8�{�s9jm*�s�!���7���y�H�q��HzUj��`�az�+�C���ZÄT6f�Ez�,��|�ׯfb1��.
C##/���@<�x�`Y�#µ$�$�_adc����ը�ӧ����j��lS�t�V��#�}46��ꦁ���3����(��E4���glчQ��%��IU!4mE�cS�[b�B;������%)�$wb���m.dT練IU�F��4�C�;Qxٞ��lm�(d���+��W,٣8�3�V-c�d@NqVT�^I��=��+F�x�|XlH�|�T�m���Kx���1��?�.xr��]@�*�$ IV{�r�3:�k�ϸ�~7�\5`!�_ -�z`����������S�&���O�F���+���c?wa\�m3!R�/����
jH6�ps�oxbD̀|��UUU��fz(F"#n��r/�N��!Cfac��>+����L�aG���/��U�a���Ч17r���(� �s�ږ?6h%���1)�?�1�U�WG)	+��+�����G�2��2q�[����m��
�1�q췿KQ�Ԍ#�s��~�� :� I�=�7���Y��2�7�.�9����d��p�7R��М�F��y��@�o\"�r7&�쓤��e9
���}������P�Wi��%����4�f�b;Hߵ	y�3� �Fh��GtF,����W�(v0��޹|:�z�}������188853��C�	!3��I��9@�y��;��IG�ST���[�����`%y�/Z,hZ��NM� ��~ q�s�u=�+�l��5 ?�9iiW���#hB���?tvuM���VQ��,<,<|jidBW�^�+�k���x%�*���Eg�3yB��9�]V��:+���䐆P�(L�ʻ�����ZTPD�i�fl����O��h\�pL ����{��ҁ�{�o�����e�Y;�3��L!�G���&_2�燆T�ˬ�`oN^jΡ�T��x��"�E��Ў�D@;��^���^�RK�TMD��àD��1o\		�b��ξ���h;���r^�Z	�D�A���I�L|}�
!nA���\��!ڛ�����[4��W� �K����A�L�n����m��<,]]]�#w�;;:,�1�@k�x��F��~�nD�Х�߷$�T�B��<ף��0@��k�g�*��+���M83��XF� �e#޸�w����JlZ靆�Zs�h<۹�Ś�R��HIؚ�(�5aɼ���%cE���!�U�%Y��h�{�p)[��B@ݰ�7�����jHH�S�B�c�%�4Hj��LN��Tf�7Œ���(=>�]b�c���zF�ӈ�E�3�Ä{*ʈ2t�-������H�4�z���Z�.W���ʰ�-Jo����&3�U�}�����%(�ă-�"��i�*́�\0�T����=EO_����8mF+&&��Ƽy-�|��.דQ�>tB�s"p����@4� �� ��c}�|zk}.��7~�r��VRQ��X]�����<h��Rmcn	���KK�K�*�1-c?7{0�*D�x�ҥ����]K�H��@7�@H$�/\G�	�ߛ������堼�?[@
?;$�Kz'�I�bCĪ���_�ҹ		����?@�9��q�D�B��Zً^bI��C��Z�����D�:NNX����y���0/fg���Q�����<��$2K6�y�Ə���N�����<~�?ʼ]���:A��mCx�|C(�S�/˙2�V	E��:�ќ�Z�L'@P:�u���)(�k���x� ��cn��!��&�UU����׫�S�R�/�{����'�k�Y� I�֙)ņ(0a8A�JH���a**#�ZY����$J���IEa�"Zx��XE[;���k� � �*���}3GV]����<�1��04[1J)�Oef��,*���EzffD�~jCb
�kN��/����u��� 4A&=|M"�!reW��59�a�:��hE[�3q�f�Yp��Q����������^SU�i���
m��b�DY	�2��8裷1h�֮�������H}���gO0�*�ٳ�PSR�;:���̱}��}��� ��`�;�\ �����wq��/ ,��^WW6PA-�,��O׉�R	;%�iv�
�4ik2a�<��k_x�I���EX�z���:z���+�ߒ��Ё��F�C�m�3jM7>uz�|������������|*�!�=0Ѩ�b�NOF�Fx�)�ٖs��[?T�U� x��Mc�/g\�'!�WOq鶕Z<�ScBL��
��vu4i��u��1�:Z��#�n]�e.��QҠs\��Sªe�0����G9`�3^đ�:���e;����%�To��c%�2�QR(�Ch�"�<��)�H�2��IHu��d�L�#!eH�B2d.Q���C��߿ǽO�:gkx׻�^{o��n~>��d ʮ��u�� �&�����`0����u6__�=B1�>��2\k����v�����p�@D:Gj�oŮ�گ��|(2�2��7߾=����'�"�e�A�I�K��@�Y�����`�qf�YY�Cʱ��i\~��&�_1o��Q�t������\��_����{䨪�<�QDx���ȿNnT ±L����6��?ξ��k�(:��^�j�Z�Z��H�~�9	�����9�~O $���}���š|7X��Fz����>'�yc�b>�)[�����]w����pt~�/��?�E��|��n]�n~QӏO&
�(w�C0<,Xq������\�"tk^9Gc��e]��{��B�/1�va���x�oh;�7L���ϯ�a�{qm=�3�Pm��`g�|� �2�8:�y��O��1��E�8�2���_s.����1�\ �~{�{������WRi-��;�O�� �*=,C/Ni;��j�y'��߽Gߜ�T�4X�� ����\��~����?ο�~~T�oq�o Xஞ?Z������l�-�]��Mk���6\�Yl���-�/`��¡��v"��z/�+���1^�u�!�r��	��3��(Zs��,�0�rL�=��-�j{��u6��y6Pd���f����$�g�C��J��>�+~�C~zE�i�w?�~��º�#G9o
(m	:�2=��ȥ��3����Ą��rS8��Eb�R�6��M/�_�_��і�Q���x�Q@�qq*+W��vÎ�1n�;#w�Uε���������r�^j��a�!�5��=З�dR�ҥQ��ĝ`��A
(���� ��I֊�.n�ԋt+r����[�XPH��+w� @��#~oU9�	���4���r=<,,�I�p����M��׿[_w��n�=�z��b��#u��#�m�_��f+/�	{.���ayG`mO�����&�e���U�M]����GTT0(m2���jd�H�,m=�R8��0�� ��|�9/�r�i��v��{��&#���a�^����c��=Ƶ�cƖ�%Me�l ��!�3e��5��SЊ���T�Q�\ �����Q��!��bCu��̻��¹�/l�����:���he2�2�x�7+�GQ,�����\��|ZȔ���_`���7���9�+�:r����ߖ�"�]����Q�yY����q##�OȽI+u�v~�6����G [�^x���X��p��-��m��{���z{<8�p��sO� ����������p����B1d, ��0�*@��ó_��f�@��4?�V�qz%IU͍���j�`oi94 &���D����RG��|1�X��.*�@/a1�m�D���eהk�$覴)����b^)[/�:���n��(�������#���
�Pz�Gutt4��6t��?���yS��&��2F���� ���ϟ?ҹI2��U���C*1�&?�/?��B_-n}t�-y9�,N+m���:Y��Zt�`��&x_Z�������P�U><\)���*������9B6<i���^XT��It�M�����`��G�_��{������s�]ʡ`��X�ƃ�ې��~6�6U���������v�����|b�tXm���h�6Mk뎴7i�e�1�_'s���������
�>^v!ݼ�av�!D�
H&�:?S��Ӄ4�OB�K��z�'H��]{����fF��+�Ph�z_�C�d]n2A�__��W�j{�h��8�"��r�o�����}A��3��Q��m�6l��7 �p�/��'�]�g�a�em���n���Y��{l��yI�0o�}��̸��&���o�kd�U�`����E�wYVF��b�g���싘��j�*߾�1�KdR�D0���e�_����:t��r*_��Ҽt���ކ,��o743���Դ�W����P��@���W��� L<��G�.�&'���	"�p(�?J0���@t�	d,�?��+Cr"|�a$�BƤ�8��ɚ�ˆ���p�ݗw��Y4jjk?{�����i�v��ޟ�x7y<�,�E�m�Y�O�6,�/y#˕=�Z���n�|�BB����.����ĉ�0Pp�-`6�:KB��7:�~<��ڟjQ������"}!�ئ�7T�5Y"���
	�M9�M扺 ^լaa�T��o8��M/،T��w���놆2�y'䖵��c&�,N&^��-W��M��*�q�+m|l`�u�ǏG�u��J066�����%d<��2;����nA�ϐ��ٔ�LF��#�ƪ�� ;��@,ܻ3�
��5x��K�`*�m�����4���32R�&|� W�t���܄D�6�g		���Y��#�4#�:]����lxvGv�����*��Pů�eN]j��/�~B�u(�����9�D�l6�khkG��jI[��x�L��f`]7�I.�����p~o�������6-��X>k�Һz/�8�YE�ӧ��c��4�͔2�<��]���ǚ�����~L4J��
�r�Hw�H���X[��q���T<�ܐ�Pfr|���(���{#cno�s��;&�n�wr�������*�z����N�AѵL;_�8�������Fr&o��Vsf�ǥ��_��ʲ��Ns���*�Bׅ�~]�/�tL�������d։���B�v�7AWrr�w�z�GeUՓ���@�jsv��p������l�H.�9j�j��t�=`����A�w �p�T�u��H6����p|����^z?���O�t�k_�Z*�:9��ɉ��5ww��9�ZL1�J;�
2�����艺o��z(��'_^� �p�4x�*������s~w��F�P��!�d:��G�M�����¯�]w�J��B01�����"1��&$�z�����6(�Ι~�S˛x4�(�������79�̴o��Pr�
��g�{�%�M��rĐ k/E�{�#\ggh�j�g�iQ7.��5��kn缩'@�|llL��`����"�@G�ɜW�Ź2���E&�MK�M��?��:�����A}�'~�;�I`��R������h;��{R���888t�?����^���ɱ�ɾ`�9jjiu���E,�������x|����rSM��Ǜ��k���e'K�P�L��y.�0^�U,P���j�U�����ɜ�Ef�N�v8+���n�[L��)+���p}�js�l�R�����C7zHQUՏS��)�����+B2�i��T$�� �=��UP���*��+
j-�Jz�v)�wl�������b��>�X��׮��ݵt�>�w}�a�9�5�)�1�eÆ}��K+ǆn�q���2��[2�&�#VC|۳�=t�Л���A����2j�j���6ۏ���]#�c�0)V�2|���Fp֔����,?'��ԏ����1ժ�~E5��Ɇ	��?�	4�2����}�`��T�|}}G��'�����(�'{!y���F��Z�j�,X O�O _��Eb���	Vk�D��8َ����1R���bd��e��w�T�ģ`XR������g�T�P�}$fQ��nk�@���j������h�		5�j��#���/�p���M<����Yk�yv��%R�n%�g���U���ޑ�����)��(���2|��]�T���T��ѭ��Ј��\B6䓊t�#1����[9!�c�&Mf���ڴ�IN��-<���t��󜤶J�l�xSW��u��k:t���V��F�K�n#1��߾}���s��#p��t��X�_��ű�~��:K��&.�S[�G�jq	���� p��T�v<������G]��k�l1�63��U�d��6^J�)&��b�הzQ?x�#���ֵ	Z {������3�f���D	II�H.J�K�5�?��*a^L=��!oN#7k	���M �p��,xeޒ�/N_�$�G3���iڴ����WQcc.n����������}�f���@��ޗ�'���{�]@��A��=���˛uɚ8�N�������K��`��|�B?�X,a�׸qe�-}��*��j�����)�	snY ����=�s���W�+�5c�P>4��[ׯ�r�W[]�{�#ŚF�����V,�8�[D*X��9H���ɡ�U�l�:�>���������������g��}ddd������
P���-x'�=	�`�CG���cV#������ݧA�:^ �e��`��K��5d�		)ӯ3<p�S�����g��;LZ��� Y]m6g�w�y��%���nZ�p�YCPx��� �����"��=�@&TƦ��G�eFD�{�y���Zy#���1��n4���=��Ku��F~�OƝ�9W�w��~qJ3-Z�î����/پ|�Y��	�Dq�����[�frVX��5��C�y��O���]����n_��v��]]]5<
&J��B^:���u��Z��$�L���|���{2N	�rh��ƲiP�R|a�"�����@ ��V�]��ȹ��R7:�?�a���ۛd}g|tT	�5��ԏՃ��ѵ�U����V$�g��`���4�
* V�y��3o������q�_B��whA�'<n��Ө��v��K&��#�*H,\M^��F���;{�g�$k��>\
�s㤢5�ߊ�5�{m����>��>�N�Ie9'��&��U)��E���#����3T��o��]Z��o�G��nDMH$.�9�?��i��2��\�p�H� ��y�y�*ס��5<�0�������1.��ц�@D�]�+�����6�����h��x>�F����O@Nl�Ui�4-X��3�^^�]�^GXL:�u���X)�4ɕ4��/|O)�O*H!���k�b��[#=��[H�}����emR~s���N�R���#���='w�.�'��4�w��D�����]"�����"y4>r(�k�����$��E\�		g�j���Y
������B����_��𥿽ie�WXX��yi=jB���Q�@����V	��9�� �l���0������'%���x��#��> ٳ�b�aӏ������u����8�<S-+��j������ey,�y|�k�f�!���\BB���`m���u��c�]- �C�ŧ(/]�x�cﬅ������-JR����a�=֗��j �;���Ѫ��n8�.u��ߥ�8TF�K]]B[��'���V��.���W��z+�}b�����B[���K��ן���KKK#.iij��^Y���P�5��OS�ֳ70��c	����ۮ`ۊ���Aaa��˱����{�V�M�5<s�A�z���_����t�O�������p)��;!<� V�P�<�'^?���%k��ȑ��uN��l	��V3����g�"�H��2Ӧ�6�U��C�?�v)�;�):R{6������X`\�4#���U&���&�8��s7Y��ϒ����Սq Nv�r	UF(�"6���h��>.[|�#��R7�b 0�K�ܼ���|1Xb��$99�y'/9��/xxP�~v���7��ߗ��_�!ر��� �^GȦ�/	�8'F@�7iD��h7����c����F�%V16��D?Ö:�ɇv��}��gz h!YYY�8�xr	��'Q��A0�81
���3�q��ڼ5ܷ^@��%��[�"�(^h �8W߹zI'=��d̩�$H�0����_p�ׯ_0l�7���m"��R��X�7xpX[Z"+��l��p���q����l��H��ƾ�Cy�쀛������27��wCI6��[��b$G;t�uyrŴ���&D��`��CDt��2���DF�_���`t� ��������IwVZ�QQ��u�^��AgXH�蛬�G�D�!w�n��������	��3����}��$���M��}����%��?K�0����w�Un��ԑ�.w�0�~<��̏�4��]	ET��cX���X`cҰ��(qXY9�v��#���g�%?#��� �a �n�÷����XƷ��� ��IE�MHa7����n<$-l�dݯ���/�:���DA���=����g;���Z�u��E&[���V'�8Sm�D˭�؁�`�NuC�������)���y;i��KǛmR(�6.�Z0Ȑ!���Ԕ�\Ν1�inum1b�Н� +w@S���~�`���С�����*f�o�_ ������ݳ�Ȃ9���<u�N�"�X�����'j�l�v� � D�3+��	��+H�(���kK�k'�Q<,�OS�&67FI3FJ��9�b	�|#~�Q���AT��e�B`�׀w��g���!�PH|������L]��뎬>˳v0w���.	���C��� |��0pi�b4\5߹���(hC;�RL�$'��9i���L���L�p�DP� 2�s'HK�gnB��Í㞆,���s�G����YDs�D�v<%Vq��+@;e��G�M鄼��""�\��g�X��=WX���i/^�H	ω�Cx��c�u=�:ܲ��q���h~O��m��XOJ_) r
[8�	ȰZ���_*lNe�jR`u����v���`���k���2Q.Cd01][[��U4S�p���X�h���i�w�$��t��UR�2�yP�#�l�F�r�yv g0��Y�mZ~b��j�����>��lf����F���j�C��2`N�[BU���G��.~�������5�D�E�ߗ�{�Ҭ�GJ���?���2�P��2	��{عO�29��J��K�.���r�+>y�R�&pA��Õ�h���o޼�O��
���ڪ�7m�'�����b5<��Q�}Q##��
��M��
�� E�X	�Nr���̑���&�y $S�����3�}<��˗�%GBw���ɂ!�K�����@���������'���7
�c[ed�pKi�ȏ}�;j���aR~���HC����i�Q4b~b�G�}+q�O��_]�S)�~�Y������֡7ϴb�jj�g���Ǔ��	�V������0� +�.H��s��0��l�J��<�;6Q����%n}L���~Uy��]�Њ�֛b�)>���.�7����V��j��$�22�$&��n��H��8@Ӵ�L]�hUjr��
6ρ/?�t������&�n�5!����m�c��_�׳��v=��߿���"�)���J�5iZlx%=}W�^J!)�
2M$}�M���E�+�����&dd� �0N��|��B��ӳ��,��/��iffV�C�Mț�:��:_�ĉG�E�%͢�C�g��ӗ%fER���p�3��G��Y��%���,�?Sx�"��`�f�փ?����ſM�CDV���`���0'Q�E�cz���㫿��T�hhh��i�.�K*���}M[������o;%����m��pVٸ���Q:70�¼Yl1����� ���g��c V�x��<o̴���i[��2B��C���Ϗz�V�$��OF��e�3�9w<	YS�=�2U����|�lJ=�y*�71�1~��72:��sr������ѩ�1t;��#s>���]�87���oV  w�!�+���(�f���Z�RF9xuﺶ�l^ o<p�ӑ�I`EK�qi��.7�,>E
��I�F!VB��{[��֋vE��d����5��x؁7:�.�x�0P7�Q��˗x�8�Ltٴ]���F�Oj�)E^�/�9׬Y�I���	�_���G���2���`R>~��~���y9��MC�3g���l6/�_�b��mp�	-#��}����OX�RQq�zb���?@��C�-P��4��:������iȬ ����M�r�[��b�-�F>4�%�@��&�v1�犾����Z>*������~�� X��=���)7�v���������n��o+�ș�^�Z_oM=qW���ǉ5�H�Uyt�-�IA�>�>B__�G}LK:5�̹M�! tOO_��ˌ=��eۻ����Eݥ
@��<��5�u��ub-�T	�B����x�=55<&
#�Rd1���
�i��JBN��0`[�͢^J.$]������(xCn��9�:̇�+D>i�ֵ�T)��y�Y{i:�y����ԅA/�V���I�K���d3�]}xs���C)�ׯ�|�soI�o }���� sC�+;�N�B�OO�� #������[@�h4��:����dރ�: }w�|�se �e��zhL���!���X�t�ҥm�� ��Ӭ���jj�D�����\^��Y~���L���Ԁ�H�8��ׄ�6 o�$i��Ջ��q�s����$9N6O���Ҷ�������������<����wG��ځ�� X޽6Z���Gÿ�|!�f�q���]Gbb�y��GU�4���Ŧȏ��wT|���~��� d��D�5A\�g��V�gu�����6��>%%%�E;33�Eܐ��?c��H{j�,�"c��ͧ��{鿅?�,>^KO/��4 ���S�!��].$��}&�KAwvԙF)ρ�K���Z<i��;�k��"4�����Aj9��X���k��sg��[�f�e=�O�EI�x��9#�x��F��۹��S���OLO�nkk��g�/���<�o`�D����Yk`�*⫴pה��~�Xё���ӬC�/�,;u/�� �gΗ������ƅ���%�&��a܄��@��w΁ �޽;\]S3&��x��A������MP+�o���:}�	 ��74�Lc��Ç�{a�sO�����i�����=��-W��t�}�(��!�ce%�37���\�WcX)�/��;26%-�4 >>P �T�rz�������x�!l�����Ss�˚��M_� �Ά0���Ξ?}� ��,6��i���U���NH���(�Wd�n��� �&iZh[��*�V�Ķ��ŋL��hoN�)	&#�2�k'Տ�7-���3K=>&���Ke��v��%�	�K:�[�bKEm�R���M���n�o�=����?>9�J��$�my�������iI�A������}e��
S��R�E�w�� �u����G}F9i�����"F6T��rhh(���wIH�� ����R��b�r�.�>S|��`�%�R(����݃37 �m[P	�ھ}W�'�z����P|{���F�OD�G ِ��HL�E�����p��8�$����Iv�)�3��H�,OǤ2����pIl����"a����C��N`\Dث�}}*`�M����;��׀�������������Íۍ����(I�!.G��hL	�`�QDI�m{G�Z$ԗ����9�ӴӦ>�����a�_k��R�@h`鎌��T�@�"0�������+^�)�潸Q�ބ!<OK_��d�]�O�N/y�h��O�t�O���ˊ}�K���q�΂��,"���=5#��k��U-���N���*GV~/���?s'sM�`ֱ��^���\�깐�׹�x50.�0Q~�3#�&���v�`:h7D@��Ǐ�.Z�$ X�0?�Y6���54.�i���V�^=gI�� �?}��|�x��*�w$&)y����=���###�E���v��<�v��6_E[����P�?AF�ٲ�a ���S��=HMo��E����]�B`A��f��u��=z��s�mii۟�F��T	<��1|���8;�XT�����HC���f�wgg�z�H��7,S�O?�^&�4�ge{�����/y�s��u��i�sg��^�L�#0�C#}�K �c�R~��e�"#�*����[��k�瀯!�R�A��Α�D`¨`C�7/�SE�|��W��(�����{&��<r���R9'}�����2-6�u�2�>\l�K���b#sY�� f�VF#^=o'�'H'�*�9��n�Ց���a�Ϸ?c�O�q��*�#S�������^F}���#h׺����K�g�P&CO�0�:r>�ii1qq%�Zb�����kJ3;uʲЇ|y% pPv<j:��
�f��m�ٗW�#X�a������ů��1m�SX��9̲9�Ep��*�]�:��<�Q'W��=7�pd$���;�DcHKK�	 VU|��sC�,�4T��Ĕy���P�X���f�Lu!���)y!��S��l���O��� �F� �� 	�Ωz8�����Ga��(
H��)��ɉ��4����E��T�Y�p���M�=�஌S�@k�v�'��̮�*�z����\�I�V��{a^��*�j�@qկ�<��U��<7��R��:	��%ȹf�Y����O�JH;p,���[G��r/t�?�Ek�|I	��S��ZSw4��'�{ׁg=��?��J����C��ҀSXO+�k��w��ie������0�u�%����OwW��$�2n�U与�Y�cl��KVU�­�}�����ѪT|�������E�����P�*X�dA�^�禔377ϖ�fX�>�~�L< T	*�!s��VP>.���jJ(��D�h*$ `ٍIj_���3�]��^YWW7w|'��v�B�)͗OF;������t kb�wn 1(-о��j|�����7�ֺ<��F�<�*�dFe2�GC蔊n���o\�(|z���0��L����I��wt�Da(���K���zD�~gC<�e���t�eй��C)%ϔkr;�e��`ֆ�'��O�fFm&E}��/�hg�p���[�<��,�����/$��0�xb����}9g𔨇�b��&�X�kC�r���n}S�ԿDLtai������kj����������RƘ��3�����9���P�}~���uS9Ӝ����h-c�(ط������
d>~���`�u^�6m:}�L�*�Ģ�;��3�����x�᠟��T�=>D_&�����jp�,0b�����ɏW��H$�&�<�/�j�6H?Hes|
qP�eͬsQ<4��9�R��K��;�j�#�����',��ڦO���(�ǎ��6]�k}
����]YYM�U���?6A��р�I��<
�]Fb�,���y�hO�q'����'/n���75����.�b��J�HB�a��8�}ۄFA����w�ϟ���N���9� v�]�1\�X��q�d���o{���|OO�±��S6? XM{��(U�3Ȁzěn÷�|Z� \Tf_��Aa��~��Ã`��Cŧ~���ߓv�2/��K��)�L�{��,!s��Y$�S�	j�1Ϟ�c��5��ꘄ�Ւ�Uߊ% �D�b�H�"}��#��A������� _�w���`ݾ�+�WlV9
#g[�0����O����ir��������s��s�!��0���yE����-C�8 Rn:,:S�
:���ӧO��|�x�1�}Hc�1�.վ �A!!�SChӁ�1��l�`o`0���RWD�ْ�>_,|a�q�=6�,&������D}N�(-qѵtk�|wA�����b��H\���Ш�u�m6��pnb��}�Ԥife�ڽ��G�z��-��t��b���ׯ��Ret$�#0�\�8�1I��z��PaZ�=̡Fό����x�YP@�	*�Z�{���P��|���|�w�ڋ����;�^rs�1/{*fq��u5V�
/b&#�c�=D�>&��2 4��(]p~�+Ȋ���K*k!X�,���A_a#B���޽{��ٽi�o,�Z!�y P�.lV�����d��ƅ����ץK/!��kP�4��-������E{v��$ǭ���t���h��\|��5~v�E�Ԟwj�K��K�����Y�VKHa�
kc�����C��P�/�����s��B�I��M��ÿt�ط*	��s�(���2NY���|r.wg��&Ar���s�IJ:�{���l�z���F�/4��<�y7s���ظ�S�>���TFc���? կ�B+Q
PzCZ$XN+p���_MuZ��`^FNN��Q��b�'��Y�yY��C��\��N�)���>�ym������;�T"ы�K�s��5�5��tp�D�/�X���N�\U���� ��a��@�ކ��[�</�\Tpr�Ԣ٫�F�%)�r" @�&ا@��s��=MMՄ�A�=v�׊���������}�����k�)�i�O�7|rjgq�k��@��R��&oo�̆:�˄�T�7����ƀ��c����]6w��-y���D��=x1|um��P��ġ��xf���	y���3u!���߂�0�z��ΰ��|J�w��4�'�ݕ� ��	��Ί��~2s��lć��
`��ҀI���<�|�_����&���\�|�1�K���)_�hx[��Y�V�*J���>��@��z�Cw[=�F����L��xtߑQ�����߿K s+��c߾��T�(���	n�~d�6��qL̡��x� �p��'�)���+_ZZ�UP��`_�(�$�Ű4��;\��2fyio�}�I	�������c��s�%�>�i޳kh�df�dfEu.8f���57�]G΁���U�1w����y�y�l<S76N,+S�a7ܜ�|h+�9=��x�O�8 FX �
�L��V�b<r�'q��)���>��^�"���� ��8���C'���O�뾸L+���QMh�����'��Sċ9�c1�l /�~����LPLLO@�W�]f�I���t��˗+���r�M3��=Q1l��:l;���` �X�2�A���3�#6��a��T�Wޫए�K�����;��-�o��� Г���p	<s(	UG�=�Ԣ�lܴ|A��u`����Kxf�ˬn)m��'�}��O/ߺm����k\�(�8��14�0`oh^����'��i
�>���z��B���w�p�pN�v�� �m<�>}���ns���#)�X�︊���=W�E�B�qW�Cc���L���N��;��|����lD�ٖ7X{g�	�IO�!1V56&�?��O�1�}������N�$]��r����:2~�������3�z%D?�B^'7:Y�k���� ��'b<��l��S�U#��q����@������EC��!#��C��'ΑU�*��ij�k�4�i=�8���bA��tڿJ�KZ��� ���MSȾ��9�H�RL�b	|����/���ȿf�^zo��]j[_�H�j����½]�q���N�'�2}�i6��c �rǁo�+)IU�׺Qp��3M_�k�y���̰�:v,���M-]ݧ�M�:�[�7:Q��!1�ͽ3� �½vVç�I����G%�����p���_�P>22R&��?��P|�)B82!���df�g�ͧ�Ok�%�~S�����)�|�����f�����>&�|Y[r�������C^������43sjǘm#���ϙƾ��OS��%9
 �⫪c4�����dUWV�_9�'���H�#�e���0':����y=��@IԦ+w���#�Ꜹ�FΛ;�����.~����� �VS]I���W�;S���591zo��7��J,���qjl��*E��9Q3ā�z�P�W��c��pU�L�x�=	嬬��!.$���X`V�����O�� u��)�z�\�#��E�@�1�GkZ�[tlG�, �<Р�M������]��ծ��Ճ�^���4��u�j%��
�z*sC�'����)=|c�!�]�~��%B��|�Y�zW��ĝq��p��[b}���EZ��˵����Wd���*c=cUF��w]�Lg��>~���<���MWel:	�`��S�l���`Π;w,���=q�)a� ������@X(7��#`�a��z����{��5�������t�]߯���+�q�c9�oii���,!1��7�
ֆϝ � ��RO Bifn�=l��x�ڢ�Qh'����6l��̭Ӛ=��G?�
�C
�s�����	Z�l|�������l�j�'0��K�cuM����;�Ұ��_iS4�cJ[��ǋhZ  j�U��d������M�0[q��TEO/75����XS�4��.R�gJ(DOo��������5��I��TjF4 l�ܹ�[��}�����k&-~��$�����I �)0�[�Np�Fn~^��G��_�~[X��\Fo�'y���{ϥ�T���թ���=�\֝��X�u���L��c��/k8Ԙo�$�tܽƉ��7k���ڞѬ�o�! ^�u������V�Q=��*�$����<<^999o��9��HAf);�����ʰ�&�3;pz���6ױ�"��x�.[f�ݯ��?0|l#�y��Ή1
!	��5]qn�iI�5�	��wc:��܆r�������D
��4,hd�5��%s�����l�5k�=z���Pw�	�ԛ�<Pq�5PM��Qs~8��H���&G��k=�V~��%k���Z�*jk�"""pN[8�b*��	��,/��t�p��Ȟ����p�5�uRΑ�$��� �1+L���(��}���W��i���;w.�40&%�R������V���/�x��T-��z4��}��W�h�`l�SO�Q�[j��}r���(GE�%K����⒒ѪBBk݆N�ʹH���AdR� �M�T�x2lm"�C�3�}b�yb�#�ի݊b��10"ҏl>y7ٜ��E��H,O�����~u�Z�5�<��,i)����5x�'�%������/��F«tAL�I��
.y`���-xuC�9����c���'��I�^�Y������z����w��?�c��,`�.�'�3t2{����Qk���p]� <5*㷆�?sVC$�w�^�����8��|����97{vvw{WTT覝�*�'!�XWKT4�L��eR7,=��/�X�f�*�	g��o�Y�8��r���-^-_'~|��tU�����h``��qWM���Fe*!�[*���}$�}j������|���S�gL���;�:B�DqH�_������Bϟ;�������Ñ�ݩ�X�/��_;q4%
S��̛���*���e�r�6���S*��Wnذ;|�������mt�Q%�$�f������[K�^������jM�8؍eY����	���sr�'��=�ÿ$;@%�!���]�}���t��v�n�H	�ft�-��ڧre�{d�Ђ7d(O�(V��Ek��c��ݴ·0�����7���@��������,��P���ɹ= �P�m��[���ÿڎih��.�;;6�!��8oi��tDޕ���]�%G��@؍��<�����*��o�!F�kǚ�����8l�OD���7tfzWӓ��&1w⢸�D��G}||�<�v���&��?9�CNN.�x^���������ud/x��r��&���N��:��t��.j;/��!s��IU8+feY)�-1�a�xkME}�j��Qѥ�{O�˭�wk���+g�\��O�t['�]����F���J���h�0���?_�U�] _
a�lr������v���G]Z���/�ǃt����m��&ɐ�����͠Q�
rs��<�P<]L���U��}h�|F��P
�+Dn�/�j�-�"?��(�����vq"w�;Rޱ�"����'Ё�}�~�Fy�OmY(��j��lrc����������I�u;��
�	G�
��FIػ�߾��V+Ry�!�j@=5=�]���]�V��<�!��D��HEc-K�m,s�0��fů�i��8�
&��߉��:���������ٺ�Ŵ��-�E���ƙ������W��d�+���8�_4m���<Ϙ�N�M�s����':��V�7��xr����C?�����y/8�o������Ԣ����@�bd'0�M���w�ΰ/^\���[�F�1tL{`�<	�C�-�`�R�'s~�#�������g��Ƿ�>79�[�;�>�Ym�R��%rw�[�~�N2R_�T�E���g�5���|IFfr L����^J�p�tG<����|�3�9:�}���u��Z���u�GF�ۀ�D/��| ��z�*��8�������|��h�&�D#�I��6���f�)��I���</�.�lE(-Zsi�v�!���iEc���{���@���� ���_o��^�y���+�d����r�W'ˆ�Z�[�b4b�� e�ޏWz9���HL���9�}Yפ{Wk�ހ"�Ы_oI�#����d�N��)��#$_[�Z�U?��i��1��,������ϯR��?���C-̟.m���%����x��s�T#fy4����kݸ���ϡ��bA����ɿ��&���֎T�C�n`�x�LQ�|= iM�?����/}n� �* �,������osfR�qп�5��Sq�I�GFG[�B�U�,K��q��	��L���L�Rt�<��0��.���J�po�QX�R}m��,D��L97��Q���|v�?6d2J� ��X=�r���d��5�t4��3�V�!h��X�SP�a!6���6�"Lf\B�.���n� ]|cq���o5���0
�iu����?�����A��<ΒK�½��	���\��+3!u�7����^0�-����s��A���߸��K��<�MYD=��@9�ļ>dz�3J�G�풓#1l.X~�p�p�~+�O�nW7�V���iI�2�	����$1+�WO���:3���-ɉ��ʐ�Ŭ (;[f$ɰ�gӯ¯�gct��5�t�̙�`Bc%�S��%��IXkc�>R��wf ��i�Mˣ���	��3-������6�d#��m�xӔ8�e���;,8�fz�.
�м2��9Mgr�^��n{�Gm�����?#k>�O�:X�ŻThsٌ�44-&TN5���?��孃@~pG��.���NL�����1�Y�qM~�m!��٘�ɷ�'��j���8�r:�X��N��-�m�8�6$te��*8�c��FAo�m����� ��0�6�XAw �?�?��؉���&�R�=�>h�cin�8	���>TU������9��C�2JvLq�t�m�BB��?���.���.�E�S������G�SI�0�L��o�1�?ZH엚^~P
�<���@�UZj*�@h�~��S�J.f"�^��Mw��N��5�����޸v�Z�?��@�o�8�5�8]�
@�N��2m.�Q�G��ZM�*�9%A��\ܐ�}d�1k���3�Xڡ�>(�R8[���%�	�u����V���:{�0�>�i~��a�;͙���������刍߶MM��@>�5H݂ �.t�"�����GsY �p�C.Ғ��t�^�M<�-�^�5.)����JD�"���|��
�[��L�3�m۫�*#�N6�	{'2==��^��2ߓIwILe7������y���`Fƴ�H��2*8:p�cF���Q�u�uLBB�Lt{o��8��F�X,�<s�L���bH�+*������~�.,X���}���OH��RQ ��U�s��)%��|�4E\�oC#Qm�k�;%�!օ����7�2�K�Ȉ.��6oR�M��8���Be J��dN}�FH<U������v[<}���^VB+��K��n��=߿�`�M�
�<��8�룋�ݳ�KXe���������*�Q��8u���kl����_/!V�yoA80*z�5�ʖKz��Y�g� q�hR=�����=�{cc��NvO�.�P��D�mZ�~�z��23�a�_�P�}�_2;����|�j7�#{&?d�>aaa�1�n���i�ijr-�8���!��;χ�ڐ��`�z��0Z�2A4���wV"Ȯ&N/����jz�$�
�L��&�M���眜������{bFL+�w�}���I��ro1(x���>�`��Q}��tEC���]�`dF�$(I�7�fJ�*Fjjj0�mF�R��*���zW�&4w%N7Tlkj
Q��Y�^���u}Dq�[���g9tDMk�-udd���ɽ��Aڂ'@+�b�t�F����ψ�l������қ\"�Tl�tT,�6�|�hu6Ǐ���; �@e�_��L���0X��zw�h��<�����+���M���c���] "�q�_H�de]ݪ���(�uK�O���.H9x�!��+�ٶz�� �F�������߿�  *FFn������ G��r����͞�?���l0+k٠B��X:-S�T��"|����D�=|�s�/v.;m.4���i8Ԉ�ݦhllL�hV�0���U����*�]ӟ*Z�Hջw�>�p9�������'����ʜ���b���9=0� @xA�ϟ� 5앥��sgZ�O����Q��d�{�R�VΛa$V��W���[b%�hق��B�W��9���iS�t�t�fP0õ'�"�;��A��z("��P�THj����7-`�T�ȝ�����-�M����߮�6w����/�K��8)1?&�˯US�<���\L��.�8�笀�r��g���}o�Vx�����!u�~�����L&�s!������h[�\�rl�Գ)0T	1{| ��>�aqέ��K����D���c���V}����!�!e���`�LN�.����w�]eZM��[j_�|���� ��@��ݻ�-]j�ċ��%o􊔼�n෯W==-{n{�L������*������/o����h C�TZ	tٴHX��J!��Ȣ�(d	�BNjZ�'''�6�웓�cim����677�ئ|�ĵ��7�OFc�>�Y�����8�t�>��D��<�Yjz�N���ģ�`�[!�E�K���>x��V����������@20��@�f��6��py^n��	���^��0�ǃ+0:\��o,\��ld�������t��.2�,-J"�#1�_��Ѳ���B�Y�ظ!zC�Y�B&���i��u�G%�\bH ?I.ÿp�̫%m��O}rA�qn�q��dkkH���00�6K:��_XЊ\~��[����n�;@Б`������o@+��s��n�A���&e�/����V��#���zմ���@}l'��K2ՀM��T�]h���O�N���d�v�a�" 
>�� <�M��]]^���0��ջl>5q.�r��-��-"B�q7����P#`����]�adOOߗ�S�&4�X�D?�����|M����>}�E�_FP��B�l8<�s���u ;��e�>q[�&����x�A=��"��í��o��ˡ�r�\Ļ|�s�mK���F0P�B��������bw�������mWˮ��7f?D�gF`X��*`��l�Rg���:x�D!�� nr��6�7�[�~���g����-y<�a3[0��n��>���Ba'k��e 	�.��\	����I c8���L��<g�i�b���zj2��́���2A�b�o��6NhR�޵?FDX̝��4-��)�MgO�?o�Ic���7���_��Jy����jժ�66��R�2N���v9�PyT"a.��k����\�����&�
�B�T2;�S���I�<ώS�Dʔ��$���n��3�e��3�w���������/g��s�^�Z�u?���¸�vsV��0]�jK�=�qp�p!�9�����\��$r����� ( a�{Q^��"�9J`Zg�WM1�UeeM
v��ia�Imu�A�� `�/
�X̢-�*�C9R2�>�2ӚW�-��r`3sss8��o�'���]B4Cv�^^�d
8~��OY�cT�)���y/� ����h��oݷ�>y�d/Á����J��-��X���MB�~�ԃ!����u�Rʏ�J[�d��OP����)���6�*�i:���|^�Ao�|�c�Y���ӎW�<�ry�-e�Hi	�ŔNH*6t��;���A I��>\�'��Lu�&�@^���-�����wu�u�I�a#W@-��34�wY�ms-.�6�nhbT�jaT!w�3�1�,IZJǡG��:�Z�v�a�Q��k;�I*�O#S�Xhw% ���4�CSwc�Xx�i��x(\���Ҳ�j��ȹ^1���
�5,,����w@�9���1�8�%!!KΥ��j�Fr
-q�%�����!�:�_�F�W��)Sdɢo�9�������e�e�s	|��W��k����,�� ��̀	d�$t}��5��]Gk�����D�x���|Ȉ#w+�'�!++�OmP��ò�%����16�\�Wu����R���S9����0��Z;(����y|ͪfa�Yp#���\˹~�$ƗqdM:zzy�ڄ��WS����7cjkϓ��Xr��� 3u����G}�Ʈ�Q��x��ִ�tͅ��=����l���~�@�Lk1U|����GC� <��.-=�e˂���?e``��(ר���]�lvB6ݼߕ�M����rճD�q��jvߑ��!�7��(��T������ݳ8+I����	qꍖ={�����ft���*�qqq�x1$���8��r��EY��+��`{��:�:�q��&^Im������7���-.,���@+z��������t�+[�J�$��a���'wRT�BU�x�:.·w�&�S>�Ҥ�˷��kt�Y��N1㗅�/*�����K���9�g�����\c��Q�eEL�����M�g/0L�#I @�B��!j�OIr�Ww�������M���N��^
�#����h������I7�/��|r��w�L�<A�*~~
�YB^�͐��/G]�6�^�b�l7��ހ��&k/��Vn���b�uh\m0��4D)eO����[��&o�hyww���Rn4e�UW��xU���x�w��ˑ�%!E�G�� 0�`h��Z��XA�A�".�N�Yʓ��k8�tB���餴�a�s/眡9 ^0~��w�_�6��3F7+S���zr?�)���⓾�l�<A\��ek��g��Ţ�����Fm�]��0V���+����ԥ�5������gl3����HW��;7��9�). ���/�E|�);�f��#WUU�_Us�^���H�E�i=�n޺�T�IyM�r�����[�eg3::�����I�㫸!��%ෟ�(���"\���P�,���bZcT'�Ny� 0�8����7����O����Ʌ�,5�(���!`��ٳȶ����&*	R���ױu66�=��q���%�]�aE��a ��7�Nn�~��l��^p�]滇�b\��R��Fݥa���m��\w'���$/�} /�H�1ta���ج�f��O^l�5�|�^l�YS�\ t����@�cR;�Aoˠ��T�:ʚ�1O����--O,�����q�C����ݔ�S����SP����"q����a����~�F����TUV�ƒ��o� [��i�[@Bnpὥ�]��2�����X&Ld)S����,��/�5jи�+���Sa��--���\��qǉh!?���C�D��C�Qv�r��7��{M�[����7����.��s�n�̱jԨh��?���Aު�7t��3&���w�#� P蔶G"��@� �a�v\����_�(��"ۦ��>7g��аPW`�U-�`�]ܖ�R��"OKؽ�yX�.���L�w��z�|���o)F������5��-5�EFզ?qq�f���<1������ |b&����GiC���W q���
q������Y:�~?nk���hB�235���4�EȺ����0.��o���`@�}��$��quu��y� u�d�P0lѩ���'�1;�*r{�ې��w{z»x6��J8�����B����(TmC�	+$���I�ס����� 5�a^o@4z������5333����yy�p�3�zAƅ����d͏?��&���O��3�Z�G�[�Y��k\�-��Zs�Z�N���,)'k�b�Rz�毄�dPu��ٓ�
�8�"bA��$��	�>�%��i'CC��C��ۉ��� �DA�^�elll�+4΢}���' xV]A��j$���b��)u��-4#
�%���^s���U���*�5�E�j�7��fh;#�Τ۵ ю�)��m�=K^���-�h،����(�j�}����-�B���k�T�\�y���^�~�ݘ�m�O��!���2V��G�#�����W�I�M�B�d�+��E�p�M�.���^W�3~��n��D��dj���?:
M�Țȼ��Pʰ4j���_^.C�ۈpxP5�(� ��f�f;��.�d��SVV-=�	>� �H�@��W�7��D��:�4;9�6�󤘘�<"֢�Z�#�"{�����	���f�\�HY!I����������y� �,dl��
�@7i/-�,W���?&��pp�Ɓ([ �-;�w���d烇X�`�e}����P.�6�$�����.BJ�CI��@࿦"�-$GV���5*K���͚l��ic��_8;5��D�~��D!�=kћr���O�Nۑ"\�����7�����GmB�w�G���P�^��*�(��,۷C��GE[$	,��i���Ve� 	0j;�r������5���``N�0� ႁ�<�Z����D�N�iB�p�%�R�^;;�Hy�[��'7�SfV�҇�yڨ�*!UNQ�y�Ĭ�3hܳ�ewvv�@�nyz�y��/�y, Yʏ�t��n��
�����@\^C�Ӌu?pB���ID!;����܍������b�h�3;�l},�����F��Ƃ�'����(����BhZD��A���D��ᖁ����^��A�w7��mも8GCk�Z�g�q�^PXD����Ӣ��,v�����G�!Qÿ�t+�zv �sݸ^BRtS��.B�H\��+�L8s��a%W)��I!O�0����$ ����=Z�E�u>���9ȢI�aq_lEhl,�e���l02)�}.쯿�"�\yBE���3�H��ʲ>n�0�a^(�ښ�h�̶�R<�1�v*�.�#E`�
�9'׋1Q�p� Ty+����Y���Ť?�Mc|��ڊs�Д�ɔ�ag!�S Ehs��� �	�����ؼ9"*�S������CD����m&�g��Ͱnjg�^����6���yӄ���ڹ�&]%}��O�HJP��W�������:��[��]�*��p�^��a��B��U��'=�k�^^KVڹz�L��>N�s�R�:$3-qf�a����ؚ����
l8��t��$�~�4n&x�̸����������;�HJn�d�����_�˫��O���653�DK��B�	y��͛n�PfoμW�1�d]�L�{������U�zzhi�b���|cpA��7�O-1 ���/υ�7~eQ�KJ�L��A.x/p*ـ��o�k:fAL�'�����d>az���_��
p�4&�L����׍�࠱��.��S]�A��J^6��P�]��4����~���YBY���˗!{B������A0�|k�<��Md��틻�!�i��	a2�[�����K��K��j�s�!�F�3yS�@�[:��y��9{ԯ��Bl��7멐�l3�B��_�>ыI��W[�j҅�F������,6���4i֕�oa�e�s��Z�����օ����ߵ^|RS��E��8�o=�ɵ�&�lVW_�%�SJ�����%�CVRJ�3�.a�j ����)�������	�� eO	����.[L�S,B�Z�9��>݃,�5����ӳ�F�lS�9�/����ޛ
�k`p����t��i�	~|�ۓ���(�J
/[Ԛ����P �<� �ŁB�DO9�U��׃«�Yy�{v�G�r?�K�ý!>��� [t�|���( �-"##�{�F�a�h/*a��Gi77�pj�o�/����Cv���>����������;����S�����k��D�����`��e�4x�y!��3�����Pг�v�_��D|$rr����4�ir�HS������;uOI$��'��č{N��g��v-ҷ�
���fgvJ�l��f;�t�G{�ns[y�:l��+�&�~Z���~�:�����ނ:��إ��D��"�wڜ\AcM�VT���o�� {tK�?ioH5$�p�����{K#�&�X�������fo 6�Á!�9�����t7���W=��+"�^�����p�1�����	e�[`�~!�5�߸'�vm�a��;Ӈ��Nn��#e͐�\ٺt�֨����_B�ۏ�>ccc���{���W���b�#AP9|����4�?����٥Pg��)�d s�g�"���v�>��M�o|�����/>>�v�"�8B|�Kym��*K
�j�)~�;L$�<:0e�󬰰���x{U1.,`^)&�����1�>Pboo�-y$������Ե� ��<���(���s~� tZ]�ABF�C_����O}d��,{!�\6�����!�]�^f5j�,:�������H0��"�wKE�,��wo=G0�����F�[��+/>F~9?B�PPP`�i��0�֭�?at6&&��޽{��D�� ���؃��F����|��w�D�����S�4���4s;��g�����_dU�:�1Vp����D�3r�/E>U6�<6ߪ>�!��a'�+�U���T�&� ����Y@@Ey9��0�|����� ?Sè�)�b�}2�6�"�o�q�b�~� ^Qm\q^0\������n�=��p����T�5MM����A����<<&�l�^[[�Lh	�o{wP9�`WIH	�`n��f��x?ga�`l7��c�!��+(��R�A<���Fq�Q�`pk���OL�n��r�x���uȫxf�جg�O֪�qH���l"IP!�ߐ��,�~�T'vAgvrH)^Kz��ا��HY\��Kb~
R�����O5��^B`����=�|)b��è�T������&�4?
���%,H����/E�����)y2+����x����D,u�3@^M�L^�0�=R�
�;
L���'���oH��Q�o�q�@�sI0�����n��r��&�	��@�0Q���4Y������xw��9�/R>b���3��_<�=��HoTl'�N[x9u�<#p������>Aj�N��_�S@��W���v���<�����D�^��
�1�_b�?���$텪�Rg��b�� ����!��=>�UңL�LO�Q���_6XEk3�J�V�����&&&�����oU��cV-N��cU�?�a0\�Gyno&�!o���czv˝�A4Z`s�Y��旇�ώE}ݯ�F'N?��K,�%I����Z�C?�qx��R6npݕO�F�W����?jѼ�
��8��e` ʄ�;�~$�dAU`���l��>�,P%м������׽W�S#�$���H[����羢@���|N`���`CJ��y������U��V��U�t[��y�c�pT�Ƥ��D,��غ�С$��Eqd �Ԗ�D\��޺�)��v�lllf��D��6��a�����VC�嫄K���v��X���3�Px�Y,H� �U��⩥3�@�i��"Yd i@D1���G��w =s��
ѣ{�]�jR?�J@r�]�Kl�U}��m(b�s|��XlG_p���駿Y��5�l��]�3���oZ��'�4:�@y�Pk�<��i=֓��xwŧq�����%�JĎ�Y��X��G���3�r��J��.��/ y��B2>Q���v���p
���:��S�_lH�οU�&��N��fVo`���n�ϫW�p},$|�tSiIUMM�Z�ɿ�����.]4
�.�;���+P�!L�A���B�C>"���R��h��q�P'�}[�	MR����Y�� ���>x)�Č��At��Kn!�q������5�G@����p|ρ\C�1����,���;�531�0C����p�0��fL)�8'%%e>Ф
=Z��#�^� �	�g-��T.�{�����d-�D�"�2 �lOY��"�0v�������d��h�]�iRn�9��k��\�&L�y�?���f
�\����ʪ���Uʹm�v����vN�<yY1oJ�v����-T�h�VJ��%h��ޞ�޴A�c"2��%7�+���ӊ����ۯ�=	�6)d��c��&��"�B�����#�T��ROT40�222����/{;˒��gjKn4�A���|�͠�M�Z�jk�qE�G���� 0��=y��jbLMM��^/���1�|6����!~RA��xG��Dnh
��(�@x�TZVSS2���[}rW����aFډ� �%�l^{�6EPI�F�'�H~؉�PJL���o�h���|�8	����sD�,� i�6gcc�)���P$�P��I�yMڹj�̧����|�f^J?9�sE9A���`�@O����o�>��yyx�b��b�7���m۶�o���f&��&p�U����O�O�4�)�@�����d3!�@@����4�t!��jT}���p6�
�Q���$
��OdC�F�`�e� �>?9"��)���
�7�yTP+ ��V����n} �G��Bŭ�1=Y֙`]����.,l�Y#h��s�QMooo�Tcmԥ�Lđ�6�al�Yq)�� �`^�P�?FR����^?�PZQ�Ѷ���}�.�rU�!S�o�,��|
dW}�em�����q��H����ʤ��V���
��y�" c�p������3\[b<d�2�A�ݾ�8M)����>���K25���-�+��,�;��؅����T�8cc�;?����~q8��\�x���Sȴ[�LZr=JB��.tv��ܔ�}���E|�S��H����f�ׅTVW����Z��[�6i!���ë��p�B��.���鯯/���j=z�����R6�w��Hun���\�=��X�
V�폌�.p�6�b��R���c��7LSi��	�dJ�Y�|�/>]��p���SD$ip�W��I=ڑ7Ԗ�vao9��q��dd8�1<<<�QRb��c�Dtt43y�Sٜ�;/d��9�@E"6f <���s��m�st��O�w�����	2��V.���� K�mO�7�56k��<����W��!Q\�E������L�w��	�����#�.�h�b��8�!>�'ۉ�Ɨ��n�����3 Ԏ� �@� g1s��\�>�>?�=/�n��-�z��'s�w��&]����R�I� Q{w:��@@b�X����i�jbe�tK𚇡֜�o��><��K�C�-89q>�x�c)v�������<�O��o(�H2�*B�:��hW�JG"z
�rqad˯���
��8��g����$�FGl8�h��R�$�F����y��ā<r�!�0 ?x�j�z a�o����@��c��F�<��OVS�#�%Z#�EPK�\L�t/V�����#���ő}�3�qf����C"O �	����5 �WJ�u�J���D@I���t�D��a��y�S�Ne{Ǿ��!нʴ���)�K�I��G9zo��W�-<�]�/yK7��{֋�)	>~vWȤ����Uk/q{77u�JjL�r w�L�06<i�@�Q.��K�Uf�_�t���+'��Sa8�e�\⃮z�]D��g5^�3�y�l��8�S]DǑN�6�t�@����^�k0c�3�i��#^������O��N4�X�R�f7��@��Px���VEA\#"�{lԧ -hP�UsM��l��mhr,p}���,��=�>�N���'9��(��$dV�ӫn�aV?��_װ��v�7�.4/$�����	�~R3~mV��UĎ��ԨUG���d�2ż��>,=]D���en���92�4�GP�����mO�۷?�E?ĂlSN�/zvLo�O}^S�zH-��8G�����Y4����q��.+6�0�_�h���
@���c���H�A�Y��!6���"��HM��&�~"�s
�� -j3�LԬ{�q˻����Ǯ�@�0\�Ϡ�����!ߛ'h�QAA���*�d� �F�#8+�y)���NN�o���� �I7h���Xz��V�Aќ���fͅ'}\�zյX��& �Z^�/vٺ
R�e��\����`�NT��zl;|�o�	��t����K'�7�S7
��ޜq��0�/���i2@لX�*� `c~S�M0(�K���x9`i��
`,��X�\]�>��Ԯ�����m@"}��F�JJ@
8�gq�1h%��?�(�ع"��i'�ֳ]�!�?�W;��%h���^t`� ��1�],�����qJ	r�����H�>_� ��<t���_��͋( '���y��=W�����!�m)�y!�y!Z@K���9���g�l�
�C�I�5j#F�9��q!pK����f�t�sF,PK<����]f��yr2s�Jf�U~����m�S�L��o�+j�=���d��ma�	��ܞB��B����z��^�%]PP��usyMӎ�%����vf��APǖ��s�|߂�C��x��=��t@O��:�kY��)L�0�x	���o�fpQ�����}.k�U���D(pg�THB�'4�T��-����� �q��6�w����)-V^�W"��|�1������x/C��	r4`�����^�\�wI̺���von�<���6"�	��ː^@f�N��`p�bQQ�UbM�f�#<W��,oNw����s�AF(~��p	��ϑ����;u�N��^�u% U#�|:]�A��m��!0'=~�U\\�5g�^�10��� O�k����P�^���1ș~�H���X4���Z��5۹n�*Uh��Y�e�c^�QJ���{��RǪ�M��F���WG+WTW_1e��I�������q+R5%�I�s�Y%V#ͅ��K���Grc���ZGr(@'2/�Б:�X\�[�����M���8�%DN� ������9��O�AD�W�*�j��vs�XWI���=ni2�,���������|��a�@䍍�����L\���<��J8�= �:r��@��?������3����1����z�������,[^GF�M��.��5�G��������v�k1�C/]���ZgkApiiF�����W�g$�<�K��8�E��X��\�t�~�Q��):0�8��'��H�~��#�]vX�S6�����\����/���逵��b�&^�sL���2��!4�cѢ'�h;0�^]����x�I2�cйZ�o��O�S�Ĭv��!V���m	�}0�g�����^�*�@f�A)"�~����X�6]]]��w��M:ρ6Y3)bi~��.�[�wcmt����E4@���qڝ[x��:!�NaA���_�*���3j�g]���r�*�a{���I%1s� �\~GL��c2�)� @��-5ʻH`P�qd�� 낂���E�L��}��W		𿙳�c9�UA/B����3຀`������A�+Wn��DFF�^VUm�?��	��U%%�����i���^ 
1Ԧ[܍�ٞ��@� �Ԭ������g���:ǂw�Y1����6y� ��5����]#x�~��A	��K-���P��t]}��t_�Ns��ρ�|�JV�0�D�����@�O������6��M�J�DP7��'�B�k�Q����Q��H �_�Q1�@GVU�;�ׁD���:	'�\�G�(�^�O9�~��D<	j^�|đ[�����j#0���U����ٌ�P�!0������eho�eHp���y�j����~C�Z�q�� @s /�7�.s�'k�kHOK����~{5��X�g?	�`�4~�� ,�']�l��q!(m��~꺪��g���<�����ׯϜ?_t7Z���
z7�Cڸ���d4멯/s���d��4k��	�֣˷;8������<�Ĳ��g>vg�;�:��a���2�.�=����#�˗3;��E�/\�|���
'� ��w&�QVq۔�j����Z����S�tQ�N���׎��y�3h�@\���d���v4�˃�n�]�߆�?s��Z��g�(��*��?��ϐ���7�oKA� ��Ѿ���#8�0~|Sf7[���,�~o���w,m�QCY��(E��g�����FG`J[c��4v�1m�5+U)tN(��|��֋�ڛ��P�����ձ���*'��h�<�Y�G��/�ߔ)�(�G��Wb�{����3�j�Ӵ�YRt$�aЗ���T5�h�$[�^�}���7�f�TY�eo#8�h��%.�K�t�9ٴR�1��x����z���9�a/��GM��3�9�؊���+�8�V/?#)Q�9"�S���D"��X~�t}���q<�C%*������(�f:������MOOo����6��/�T��JKKn";�m�Z�����3�t���~�J4n\�X>�	�!7���p�r��$.�L��u�k ]�VwP=p�'
!�������H�:9>�w=U���G�l|�I;�oY�&�^;�����ˍ���� ^��i�v���7��`0�l�XT��!@XD�f�8�m�0�Mu�x�ML�@uZ���Z��C8�Șiܯ���3jB��TM���b�V��I;�,�ö����L��c��uc3Z��%@�C�TL�
�P�Ĥ��<ΐU6��ĹҰ�H��{͗�!���\��љ���S8��r怣�Y�P=$
��7{V;�9B������ t����C��s=��~��&z*�l�p	�#��'Xv����^���'6cS�9@�Lk3���9V����<$&�n7Z&>�}��.B�0��W":r.�1���F��"՘;�FˤLȳS���h'�NՖ����>ק~��:#7��8�Y�|�#��؏'��S�C��n�3u�AYV�C�&��v/�N L���뛙ͺ��PjÅ���W�&�@"�O~��j<�~��s�)#����!/<7�6�@}��-����� �M� ��Y]W�,d���nc�:C��@s #s5�����M�M0�	ҳg�Q�PW����ꍌXs�[�v��L����e�3�������"�`����ٿ�ĥ���|�^KSU�7N�Z���5((�)����?�0��moWF��'?b������%��$n�q+�z����C<P���e�õ�����}��F�~)��
$<5�ŋ�O�91�+�jA ��~�Ձ��"�l���\���:d���Zl`/�����/������޳����@�+����\��`1�_�̄�pc}5�AC��爙�m���6���i��/cx��is�j}��ky���)	!�a-x�$ԋ��k>�z��%j��ުS:4�pB%k�� "!!aiuei:~�&LEeOG�ZX0��� ���_��@�<yb���G����!��&b��awf���X���܊S��S�b��KR��)� T�x"���dTF� �>b{�M����֡ͽ$R�E�H�k�q];<
$�	��e�/i��X�=�kq�^Zs�����_�3�-f3���m^뺝l ;@�/���~���w��xrvD�sy�ZG�;�&&& ![�{]ʇ�К1�	+�~�fD̘���藪�$����\�)��?��Q��5(j�K�!�n�i�p-���ˁ��ƥ�S#]n�S�<~��͎�v��
��¸����s�b����9}r����_#o��YV��/�=� @��b�K1��4Ϩ����aI2�.�ʄL���~�.p��9nj`~.���_`Y�`���^�a.v��YX޺0td�)�1\7N�	�~�5����0eO+Ld7{i�z�+�;�4.��"�e\T�ub�o��������)�=�ů��E���`�����9����p�}��@�sy�'�=���;]$f���f�(��|��)��T�
�_��m�#�v<�ي���aX���O�P&T�,?M�g��.8�n`�?{D���cf?��.��y��Pw���_�S�-���U�C�<��M3��؁��o&�S��l�\�������|��� 
P&�R�@���`xv��9�L�^�j��4��kl���X��'��tEFs��]W�dv#�ƒ�E����C�q
�>$��������y��.�[���s/�zJ����w?|	i�ܶ�G=T�/�~/hQG@��ʂG�ϞH�l����?
� uCX�C@>�����H8����mm�w~X���Q�	��o���f,G�փ�����8ÁgS��뮀�Re��!wʤ*U���U�d�'�~����q���(�<���7����g�j�[�N����NX��
�}�����t���z�M�6nz�f�|��2�x<�!�EKϨ���]\�ݵ����j�5\d`/@���Æ���A7Qkk3fPq6�f�C}�ϡ��B�/C�G��:����H�����yj>�\�������
�f��C�,qf���P=N�^)?��@1SPy,k����i��CJ)��:]�	�}��%I�aLS�nZyU2�^c��k�/���}��������J�P���t�_�{���\mv�]���K�rgY����(��R��H{X|g��2�N�K@jXW���XI�	n,�n��������zf_>u^�}bN3�G����J�����20���O��l!����ƃt7ˊntww���xƐ3���{..2���V������^��W~i��1*�����?~\.c�ӌ����}<�8H�Edd����w:�1�}��ܾ��#�bﱟ��EB� n��%�bTC|��Ѣ�}nf"��]��+��8'������fև�K���U�pch$d^�UD�>q%i"���P�����}��pHto��C��\�/�鯫n�w�Z11��JTN�|�uc�#u��/.E>��ˢ�����a�!p4��#�4p8�e��l3�Ɍ',LOO{�S��ٗ�\�y�\f���]��x�Uz��+t�z����)1j��Цd2�\���i��v cπ�w�Y��"�J����
7�М.hλ����|���DϖP�����������#��� 0`�'+I�?����1?���nsQ�l�[�W3��y� ��߸q�l��#}�$(ˎqMʶm���R�������Y�mR�vp�ioN���}9����ǫW�~����p�8��ˡ�=\#�3����Ƈ����Kԓ����2ǉ��:ũ�N��}�xN�ߜ�V�l�q6��5��Ά�U���]$>8�����s��mLa6e������ 
�����)�۳g����c�aX�9٬pvv�3�)�mk㵩����{�Q&-���LK�g�ka�3 δ��R#��BT��T�o�b���4���@��-�_�1E�g����w-��;��9jZ�N�F��e>l�b�?�Vw���f}�9 ��=�Q��3ý���Y��+&^��F'7���|K��\	���Z>ˠ�*άn{�����CY�ǻk�|�o��2���R�_B����E`t���w������]�O� ���]�d��+�W�pZ�3�I���#d�������W�0� �^��ō
�z£3���b�������K��0�[��w���}�����W��:��7���8�5#�3�n���GO8e�X�ۍiǶ�P���#'N�H�ԖPn� =����0$����o���Ϝ��>�#���\%�"�<���T��׊	%�7�������T�UWo-**
_��� �1333�a����Qn2��GC����X)�;w�|��EԶ�<�^����ge�����b��<����<��ێ�'QWF�5뭌�̓�߄GEFU���V7t���1����a�UR�Qז��͎'���b?,$�d�8�hǈ' =~���[��5�J1�)?R��,@�+�"�UMS�ה:�Gj�O�x��|�n��x�i"�O��b����n2?�=,*�b�f�}�]0�3���f�r*�Ң�30��LO.�����������:�t��OF�=����8���s[�v�/8?_] ��ҙ�hl�<#Z]YɄŵ�
iii�x��� ����?�)f}Wz�D�^a�*2uNtn�b蛦�w�20E�DU�N����-x�Nî�����N�lV�b����啨S��qP$�r�gZ�������� ��/��il��n2:1��׊�>��[{"BA8���l<l�aVVV����[���Ш�����y����	�A�@1��Q�M�RF� ��J�6<_�zv5����	��E���~� ��@��P[�,(8	�U��	���Err��N��i��R0w������ˊmQ���|�ÿ��u���se��©ٍUY��MȔ\�j�,2q��z������O�C=��m'g;��K����]Ij��S<9]��Σs�*:�h��/��H]��N��v�P���ÍKH����R'����9�Jo�8a֫Py+����J�(^R?��g��Km���=D]��i�wK�����=��BMx�iݺuq��'�}�w,$��2>*{|�o�n*+��y!𾿿?��^3�>�t�F��N����t�q���K��oH��ܸ\�0@�Qg�?��E�盪[=҅{VX\�'��)[�I�[c����r����]�^?4T�l���-����>��L�Х��c��:��J�ˤ[Uo�z���w&�rܘ۾�i��ֲB��"JlL�������t��GT�z�.`!���x��I�m�9�wRn�ō��QWN�����L�޽y��A*����q�n��VT��C�\h��f�!b��'��!r�"mGݨ��7;��3�:ϯF��
��d�a,�$PĂ�{�F�7�O�RMt���渭�[F��y��VP~xf�	 ��{St�u.�ݼy���z��v<)p��QZnE�7� ����A;�����eJ�=z0%���8�����������cc=���9�Y~��]��@�����{w��IWq�ؖ���y����H>�	��	���ު(̊W����Xu�u��?oK�@�Jʚ�9 �w0���W��ek(�}㼼�Zx�3�s�n���_ܷ��w����ϟ�X�K�������U�`a�S{H&�''|�_I<|H=K��իxH�E	���Snge�%��g�]���R�;���K�Q˴N=z&*l��w����׵��B����f;5�O�x^0��]ӫ����oRX~lY
���p��Q��'Oᰜ�@~c���G�wv ��9k�D��@�>	�K#<4�A�C@���-<��q(R֎�#NM����2J�����fx�4�-�Hr�����S.��T3Ѯ�y���K�>�zeB�&�g"��0�	lO�=z��)MM̓J��$������^�O��o����2aݺ�1��?[��Uu����C�%P���p�����G�3�B1e�?0�a^^� 0����o=�J�Zu��ƻ��H=Dp[խ1�6���\\����}i��J�g~܃?�p���s�#�2g=Z���� ,�q��@����BɒkVPٽ�!�J%z�K����ȴ�
{/wR飝���?����w����]��*W����U���w����]��V�8_�V�����A����׎$�OLW����ΩǤ��4�+�61P��������$�_j��K_��@�ܕ��-ZMG������w��+�]���
y���!\����+�]��
W�������w��?Vh���@zL_����=a��pqպ�߈"��M�-��IwB~�����G�p�o]߉�)}���1i��� PK   (}OX�Ɍ�� �� /   images/53a6c856-3ba7-48d9-b0a2-5ca2401e7b62.png|�T\Ͳ:0�M�w�$�w�0�C�n������������s߽��^��kWW�׵�wuu՞pEyIt  �.-%� �  @i$����N�4  M�RLLQZL�L������ �
OTG�P��Ҏ�������I�+hJ�BNU�,(��D��Z㇮�A�z�ᣑ�ҩwMNNy|���z�[����!�W���fS�"_7f����*~'�L�숒9|�#�E�Ƚ����M���m}c�oc�rE��u�M_.pp��O\$cb��@�	��	 �pe��*��F8��G�G՟�C��ئp���Є���!���wb:4�ڜ�(VOj$I�@'�Q㦷aB�g�N[��O�[�	ě�;+K��g�Z��Ħr����3�6��b7:���_$G-CDD���|�"c8W��!�E��H.Lɝ�7L�k��y4���f��0��$ɠ�{#`0��EP@��P^�;�?b�����G��lƝa��!)���Cn#M�rĸ�B�7�슩AՈ�,�Bak��Ra~�B_2��'�����Dk`Q�o��u�)TF0�-�x��o0A^�D��!�Ĥ�GZ9�:�=@M��}y�U��}x��j6�2�*=,�b��)
s���D'�%5�.z���W�A���nq�8����e���T?��at$�͛�V럓_�����A��z�f�PZ��P�{
]�>�s�]�j>N���QM)�T®�?/b-ܶ���±��v?�М�ݿ�{�4���
������5ba����n4ђ DwT�l��y[�l�AV@���1��I]*h�2�y���b�-D=�q)�	�z�"qqHi�<��L���T;�|�AZC&]��'�=� �Z���-v�i�i�I���˪��𡜴t2�p*[��˒�)�+_4q?�ت����4�=����v��=�D�����Tf�7�͚���ˈ�*?!��(���c#�o0�ȝH^��C.x_�����c;;6�G;���l_I��h$��u��Mt�W�M+��@���O��#<:`��� ��?L����|�wX�w Qa�0�Ř j�k
�Y�G\�����3�� w	���}�y�{|D��cfa!wDAJ$Q�b$�i����}�xa\X~A�Rlq!&��c���C_M��J$�(冤��g��$H(ڇ������|���WB��v�M����?Rv&�
>�L�}��]	�Fd�3�MA6�fe��	/0�O�K�L4����-�������:��h�y��rˀ��pG�����@�\��=����I�`�!�`�cć�d�ލ �!�"m���s���r	�&���@��;�s�La�Kv���� \|�r9�M*�
��OUTKaE�;�.�K��G�O��x���>"'�HIt�D�ޒw#{�Y3�Z�L2�c�x�t�l��ڑ���@�/�y}J�t�!�f<�FFF
G�G�G`��G 	�t�*>�/J_T��ĕR(i�֪���$r���ǝ����(&+����IU-K1J�ղN��Q���J�燾�|�������w�y��ے�y�y����'r'\����W�I��U���3ushS{�LSk�_�Y��S�5ؙlm���+�#�M�F�gW��s�*J��3s�ZE�S\�1
�Kz��5��C&�0C(S((q���L�<�c[:Z�֕�y�!-�7G`0����9d���i�I��8{Ⴐ�cƉ���xHy���Ѐ������� ��"a����+�N-����S=�5���J9��cȑ͍60� ;|�[<F�d�����B����fh��~ϛU��98�>�<n5v�È���c�8���XW+[�c�l�l\`��@_[Z�b.WW�e�k�=b�[=\�lᴌS�R3^[Q�n�Ҽ�|ʹ�E�ӑ��H�㤰���l�T��kn`�X�X�X`���A��D����$���Y�۠E2�
�ǘ�6m�J�l}�\����O���ԋ���$�q�5�\��Quu.��
���f�4�U��5A�[燂���%A�Ѱ�@_����S|s�(!��A�B=��
=����]AA�l�l���M���1��!I��M��{�����P�\'��g2A��@�ٮ����W��|� ����Ov���:��B}�&ߤ���ZX�LI6�Tس�Sy�=�#E ��Q��HV�h#5��A}"���K�B�d9����jnlYo�6�q���Ƶ����������	�r05R�9��)�?I�+!(�������<�ӊ�YbO(�e��].Q�KgH#�"Y�[��v�S�e�;��M�B���������W��'��ؾ�ݘ�M+GNǯ��'O����js�wN��-�~NIO�N.JHNZ��{��JC(��٬bBK��"w�Rk���[���t8;fS#�wo�z!N�
�ڎ�	EHV.l�6��]ww�0�������*���D6>��L0�?�ޅ����B����y=�Պ�To�m3�8B�33����;����FF.�{x�ށ�dp:�v\/N�n��e���q0�`�U-�L�����K'Ӹ�J͘�r�~�~�>׷��zec��������*&�?��8G3G��
��ϴp*���!��C+��=Uy�39��ϑm�꜏����M���E���6U����kߚΎ���}�_����J.GU����~/s-�ܰ���Dע,9^�o9��{k����׆8����{�yO��u:��CD�W�pB�A������g�Z��xB�t�4�t�t�w�u�����$�""}{��bӭ�#����hm���D�-mg�����	�,�$�������C�	.]��#pM�z��S'��Yq�k�e�����C�`Ճ����I�թn���E�����\�n�{#��p�ǥ:q��t�y���ީ�ڵ%2O��;���J�y�V�G�4�5�9Z������[�d��|`��3u�p��#��q�:1�M���E�q�i?�������Ʌ��x����o��ӆ8���t�~x_@z#x�4��~��Sd�]�C�y?`u�8ew�p�����U��_w��	 
�̙ ,�}%�7߆�b/4M�^h6)G�>�i=���#����V����x׫�}�@�ӥm�:���OA�~�J���3ݝ��Yסm�������/��f^��9��$Si399 �_	 � ��`�� 0 �� �W���V���X  � ����-�?�߁q! Ŀ��+(���ar��E������I�C�;���:Y�9Ӷ҅�e �Ki: 8��\0��Tп�EKUg9Y^c;&C;#S&w���w��Kژ:���X�:�P�K��/�����_*�Vr�dbv��d�L,L,�(ddd��&f�������	PX8;��23���1�}f�s4gf���afacfcc�����a�l��h�D��A�kqS'cGK{gK;[���Fv.����w��!Sw���d���i�� �?fV&���li���G�o������W����ZC����R�}4A.n~��S�jN��bv6�΂��������Ӥ�����?Mj��&���������?K�fk�,������7J�催����O��Fh��������ߩ������/O`�_��o?c���	��3��N+�rZ�V ��ET�aN�-����
݌F~�T����X�N�tH���֙Ʈ������%�%z���;��:�_8�'����#"ۂ���t�Z&���Or:���S��rs�ߦ��ϟ���\]9�>^��ϫ�UUU����U��<]�=��|��k*��d���&3�)dV��4�45!N�xP/�+dW�+(�rG���'�N��@Z�T"Vm�!�+@tǜ\b*��N�?�/��c"їB0������%I�ᢽL�����;�x��	�ǽ��N�]��D	�b�`9� t�v���F���Y޲���XM���q%�	~=F�2���r�k��T�P�r�E��hݫ�_��XǇ/�O�ݖA�H�i�q�c#��Jy�X1�y*'E9������Zڗ�.���1��T�*=S�f��c�;�����lX'X��
�-k�]�\g����$�OȄ�귪��U�6���?����[�߈�j�x��,��(,�~�א��V:?���@�h@{���;~|�[0$о/�a��N������[����g㋀ռ�Z�E��~ڴ�`��a�F��(�Ǎ5�wAK��d�'sB��T��1L}n����Lci�_�a���no#o��,E�_3R�pPԵ���])��"F�q�@�B�X�,�7�Ԃ:u{��{J5�g�Ç��9R=e�WV�G��@�Ö�ٵ���lT�4�x|L��V��*�aR�F�M�{?1����<߿�b�2cqr�HyB ����"Z��jQ��xC�r���_U���CPx��i�����f2��n Sl�:�l�I�u�zb	��M)�7��:2(�B
q�4` ���1ўy-��w�
'ͦ�3i�~��ش��)
#��?�����
�Qk�|֜dw����<Z�zl~��⺡s<��r����֙����H$,���'��I^kK:�c@.����}Gmej��o4���'�r�]������ �T1%\޳�p��]���[/��d�q��]j��^W�m%Iߙ��s��~ �9�_�?I��z�Ǒ��b�������A��V1�u�>��=ʺI���*&�88t0��8Do��Q02����!�n�b�^���]ge�:�y�$�:���8O��i#�h�Y�F�wh+6u _�<�|E�;�6 ��=H��+��`p,�z�޾��%�V�x�����m gV_��/aZ�1���+���?'�o��8�+!g.�ǩ�e+xn�K��j�y؏+��G����M�[�@r��z�p��0�O
�m@'�M:�ĳ:�44��)�o�V����8wn��C�u0�c�n�L
���73�p�c�-,Vm |G[�$��
QY-���\�2�n��a��:0�*�{}y��/� #�����5����lWɾ �U�/E��|��''��ʥ|�{�\;-�7�`�;���J(R�L���WV�{��x�/�}�e�+����/U����(��#�����_�H`��:��#MM�l+�^��QȋU~��W�泒���k��P�iM��q�����%k4!�8@�㒟����(ċ8)BL��K���	t��_���I����P�|rN�+�4�4�5�۷����R��ucc��y��#��SƆW��٦1Cq�\A���#�Z�~N�Psj\*W��f�����/]����| ʽ���Y*Ы7�;�����]� B������&�1�=1�0���*�v	����O{|Ϳ��sa*������V0���nQ������3�F����q��
��5�*�R�s��)m-rX2E��eI�Oc��9�q�@a1���u@����,�ٵ�3:�T���6��&T��"�:/{م����;�2͵/K`���V�����k ���M��rT&mc3*ܸәN,��
M8ޫ�!�f�64<��g�'k�P9h���8�1�{�C%N��	���lSo4�ã�kB7EP/�E���,�-E��`"�s�.b^�ψ����u��/����[l��/&>y<���~:^����>�؍�RdX�[k���H>7�!j49Y�"�(Gw����y-5�NRk�ڮ��V��$�!^��8/1ߞ���D�W&����T�F�Q���/*|&���\kXSi�h����� �m�1a�H�sx�f�Y����f ����:��!t3T��D�Y �"���wJ�����Z���2|m������M��,��V�D�)Q��ǹjb�C6�BQ�Osj<�ǣ��%��ۗP��S�\?�0�T�4���3�n��]U�}�#�I;�7H˯+��Ir֬����ω�Q٬1b���s�m)��o�Y�#I*��'pd�.>��!tJ��;���#G��j�r51�L��`q��|}0>���v��v*R���;܀f�D8�l%zZ#7��s�O]��;e��V�ǵ�gy�zcmz�H@!ڷ��uX�=!�'�� �U�w�B�y��iy���hC����ėK
�٬��g&��<��������u��A���h�>V�3���E��.S��z`fF�d>
C�ԭu���b}��=�����^�.��T������
��|���kS%�u�CՈ�Q29��$K�X�h2�w*l���~z�������w"����S�A34��)7&�~%�1�5� ��9�2��ң�_�LH�ϓ���4=%�X���+}$��Z����
B_���3��"F�8��F=�M9�bd&1�{X�K��ȓC�Q�+�=�_��!�eΆ�6�SF��*�K��֗�|���A[�Y�-�����60��P�v�[���}��ȯ�6uG$��:��B����N�,�K��@og8]8��[�$]��w"d��_�a��+�%��&5�y��Iԗ�?��rΕ��}Lb��V�LV�X�=�xO���]���[S��qs��#�;M�(y1���y[Rgdx#��z�I}\�*�"��F:�ڧ0pζ�ۑ��(�=HY���_s�~�>힪
EMq�w!9�oLѵB�����jfSo����V��=���L{�ʞ� a5Nvk�Z��Lhcx�V+��L`�s�.�����b��������n����S�`�;��e��ΩلX~����
��{
��N�H����:�nn+�I
A{���揕��3p����񭏫J��������؇�0�Ao�wUs@H������N���	��0#�Ct�`e��볻B��I��=>��$�>=V��Ê�c�K�w�,3�����Y���QB&n�O�������p�T4�8x���:��x�]���h�i������X
��O� 3V�sy�@�W֯�#��e��EyYPB��d����y�J"���o��
�Ŕ�m�A%<��c޹�t�SXw1��l�*�߼��U1$8L��Wy�k=+M�r*�E����N���i����^��;{h����b4��U;��z�&D����V�R�n�׉\]H�S M04��C�7���Ca0I��r�k~4$�Ojc�j,|:���U��W�T�G�K&i�J��%�B��:��5���&����;��Q�
	L���������8T-��<�#6���fi�ύ�I�gI��7�ۑѰ�)����55��~����Yt���>V��ϑ(*z�Kd.�SĶ�s��,���K�'��H��^��H<	$K��P�j�6���-��p�Q�L�`���������M%����m�t�n�<Q��t7��B�f:_D�.!��r~xr�����W�1�h�F��Nzv�Y�ǭ
+��6�yB&�A���l8�8��{|�z 2Q�?S\D0쏐���w��$�\��z� ����@�(Y�9{�:K��8|�82�㗰��b����d��q�R1����~O?�N�6�]ݪF�q�� ���Z@.oA��E�=U"�K��8�Wx�X���8T)$+�r��OThE��Ɵ�'�lKE.���ġ���Ô,�sk|��+�����M��h��a�ؙ�P�G�v��| ��q��e^`��FtN8��@�]�(�S��� w���Tg,�&8��}�Z��~�H��oq����BѴM��~�E�ܡzK!��k1`�(�n�l}A}Ae�|L�1�����v)+��-qG�M}�}ae�R3j�� �H�� �r:��(Յ�a�ȱ.^�� �D�EA�r����/C��+x��7�*��뿔�j�bKѻzm�s~�����u<�
D��ufȸQ�Q�a='IQ��B|^�����3�x	�������/�RY�>Q�G��QU]�1yG�K�]rT��F$X	�Tp/��J������:6�-R{��C^�8���}^.F�8��P��R�݌��5�-����,�|�~t1P޾�
�prT8uA��Z�\��p������Zm������I��dɦ�
�)DA���1�ҁ'RB�d�b+��]������2�#�?��G��}�^���8��^�"��;[�I�>T���r�
�c|LҾ;q2�#��'��8g��[!T���Kv�����e5�r1]��~B���^������h |1�k-R��,4g铗2���DsD!}_�$!��RϷ7M��u�8��#���P���K	�p35�^�* �K�t��9��3�0����y~���<bx.����he�.�֝��z���ԧ�\\|z�w�>O����fo<��x���������t��x#]c��-���ݍ�-��~����c���h!a9��{�����q�xw�EX]4F|B�̑ob��\�~PȨ�
�F��AFjk����!=�]JCrAәw=q��~̒\����q�0�I`�>k�4"�~n8�<wص3��#��K����e��tI��@7�A'���ǜ�i]p�+���ko|��ZSEx���4 @&D�ٲw7K҈���Q:Y�����ϱ������"��%7��o��9�K�����]�?���$v?8vʓ�	s�:�������@4`��hU��@�@I��oer�Ew�<K�6C��U�P�iU�S�W ܣ`�e�(��W��l�l8�wn�M�͚�9P��ƍ88��6���U���
D�y��+��v����vy���%�g���2C���?�П�`|�c�Y���D�"�)&u}�o�8j��²�3�}l�D�h�@�������;�Q|{��zZ�����'�ڦA:0B/T�&��@��%����qWE�Ʃ9�)X{mso���B��;#�����ވn���jϵ�9�1$ME�D%b7��E �s"-/��w��4�y�D�0�J��BI�Ns'/d��PZ9�x4n��4Z��\~x��m�F?XM?� ���9h�~�;��V�Sݡՠ3[��Ck�����- )L���-���9t��ɇ�A6VQl��-#��Ul�'�"ЊJ��n�뼛G`���M�y�����RN-X���[C�l����	�+�EJ<��k��<�u
�Y�֌�r�"��V$| D�,�c�n�S`K3�#!У�Jak"��q�W��<LZ$�{D]�{�^kԙRa��gqH�HmJ�!�<���c�Sz�v��.�ul��`�8�K.1��� $����|V/���c�N���
J����X�P��^h�1��)�)�03ޒ�^�0:ϲ��Y�st�kZ+�R7{ԭ����4���� 9E򇢘��۔�@�F	��]�Ko����8	�S�o�R�6B�����_����Hw����J43'"{�io�|����?�9jä��6f����j�ɉ����G�W\^[/�v���t6e�y;����/����1�7rg�����o���_ɃqaA����L����{����PEi����ԜщgWe��)��M�u�s�)D���Kc��=Ü܍��;O4�l��8sop7[D��-������KVe���6���1����*^�����n}vW5G"�ۆ�Ԇib("��s��󁟇8�E�a�1�Cqp��\�E:v���i&BZg�a�G6:��Nn��
[�e����3z�a�c���cz�?�-ˉ Z���,Oh���i�f'6>��`~��[-�8f�?x�pQ�X:���x���hզ�r�s�3�#�W{��ex�����(m��m0�v_nrjb#q��$�r�j̊'�ĺ�ԑ�6/�=L���1}O^w��4��&���=ө�G��r%��t���o������z�4Fu����D�ޜ�a���阘��Y�x|hRx>��g����م��|A��R$Oh%����(�\���dڛ��\�������X��~��F2�o�^T�h��c�s!��m����b�8�{��bo��`�|O�s�۴�*z�)_8��q�Pd^+�
��G+u�&^;�Y�������n�.}�'�!�dG�tL_��'Ay����U��c$�_#T�����%o$�El��v��.��v)��L����hG�����xuFB.�Q�d9���\��H�q�[{}m������ʛ�g�%��t�L>Dmy�Œ3N�!ۺ���,�[Ou�V��5�2�.]�)�WؕM���d/�f��}j[�T��J�%�!q����T��i��5��P��1osO��u���x���u����I�I������G�:�47Xdĉ/��]VJ,S���N^P�¸�}���F$�v��F+DQg˄x����opN�2;3��@\0t��B]��2Śߩ7SȶM
q�Z��'�f|F%�� v�`ƲQ1����Fu%k1��2�e�c�j��6��?��M���d��i��NVy�r��\=�,�-(Y1��i�	�� �U������j���I����O��J��6va��ٖ���_���$�;��7�}����>{�ɻGBR[���G��f5���c����톏���j� #��]!��h�@ ��Ez��K˅�="P�C��|5зc
{-���W���iɬ>�$�ͱ�͋���X�v��²�j�����!����Һ���d3�谵��F�� A����},`�!Ax��\�uA�Z�
���@^e��HҀ��{�;��"�ӾȔ 	T�,#|&���֍��X˶���Z��!V�p�3��k��m�2�����|s愘�� �0��Y�S���.�]��^�sەA4��S���B#Po_����P�`�?��<�"Ъצ��[Eϲ��]�D��&u`|������"��,L�>=v$�{�1�b�N]��au �V�`r��0�T{�/���.�ރHho�N�`\g&��Ky(����V=x�h]�W��������e�C���j_���\�^�O6�%�H籄29^���̓��I
������Ao�5b������x-n�Y�6+��3θ���gz�\�>�rš����k�dQr��i��z����t���xu)�W���.���=�~�9����-����GN��e��������$���S��EԊ7g%ůY��V��5�g3l���3U���,�YmQ���]��%�� �8�?1��P��_G���(�Cv@��$k/�H��f�׭ln7YZ�e��' ��x ��9{D|��������{�~�$A��eU
�M!$���~VKb�#t�v1ZW4���g²���`��g<�)��氘��	�h��=��2Hu��ǀ�`Q%�
JD�h>�^X�d�ܤC�+�[6hLғ�H�$�xƷ�E V��F:ۤ�83��O���	N�1���n��7c��W�Q����c˻(��wv�5N�c��ȳ������N�U��&���^��Q�͘�{Uw.�5Q�Ɖ�!c�s�'^� <�v[NӘ$at��eo�銒��]�*��0�,���L��6�o�Z���G"�V^�5�rh�3c%�o��5�܅���4ND|�ũ�sa���	o�S�R��,���y�-:�r\�]Q�l�~T�wh��y�!Rp�]��t�<����$�����=�u�}�6����$��[�}F���k�L�AFu "ɿ�D!�'N!=���RH8�gFFDD�'���K������������EebҬio�Y�s��-���@�؊?�>;��8�[���)���ry�z���0l>b��{Xx�#��f���Tq'w7wqN��35f��<�F1�u͡���V�_5x��U�8��|T_���+o^��6�xo�#�`˹6\�v,�E��7���{|=Jum� #�0���g>����$��!��M�V�	��p�0%�ϱg�-��ZY��OO]���|���]#0p>�;2��$+�*�U���U�@'�y&}�cr2O=������6G?����)�oz�21\�^O�8w˞I���J)~7�8�A������m_&Mj4�Ą6�k���o��,�׍�O���L'�/�>R�N��E��Oe'"l�������9��o}����yS�������K��X[��fD�o'_`�� �_��ݜ�
.aʾC\4�tFf�z,`ح�c��O>�����Gnۜn���) b�{�4t{LZyOx�SJ��i�q(3$������i\�}i�Y'��}G�wH�41���{-gݨ;Q^��Or�\�����:�l�Z7�2V��|i$��u�u��� ��Oᶾ����a�[,*�M�]��Yg~#��[�[?���'PQ����G���Wj]�(�Z�0� �"�A#�(,�G� ,;"�����rp��y
�J�V:6�f�ǨW���f�o���'>U�e���4�I,`3v7��fJ�r��mKݐ�7���\�h�F#�<7�>�
e���̱��� 0���ę2Nt6t�H7-�_~��~K����$+?&�Z~@��SUiL����bo�0�o���@�4�3��5�zy���l\�s����Z�2�n%E�auF���~b����0��D6���l2i���tzۑ���5�`�U����2���z�=5�˜��tV��'����㰞-�;�]V.���n^[5r��Gk+:�L:�aK>�D���pxP���Do�!��� S$��U5-�H�r�����~���+��z�-����③Ф'-���?��'v��?��g���[�ٟ���l���?�kI>[����D�1ʉ?߇�`-*�T����jS�G���0[�-���%A>��܇Sqh�ZY��Z\�H����[�&-Yf�����m�l*����29+f�0Z&�OX�.�\����W��{�.��.F�Z60z��la��ɬ79��~�Qd�r����~�K}��H�����H������5J�8�o��h�3�z�3�̰��`����'�0>vA�;�s�Np򋞏�A�)�Q��`]���5����g���r���?-��1�U���+�S��`�E�+���I������[����x�x+����'��N��lφ�yc� gͰ�j�p�������.�"����6���O}2�]���rX��Z�����8??:�;/ɵ�l&[e�f�[U���f�Fͨ��?e�e��Uܜ��ap��C�;t�&�{EM4�jqn�,���3��{�/Z��4?2L6ot^
xi{8IN*���<�u�7��PW�|D��Pq�������i�:��T�	�������V�{2�i�`�'���q������]��gu���Y�qF�a_�b��Wi�����Ʀ�yU��o6l��/��Z�Z�
��E������k�$�5�]�9y�a��wc��I�VR�}�}�F��L`��Pk�I�#�mzπ�3R99�2����y�d��p�m&"��sr7H��ى]Z��ٍv����g��B�~�}r�p��&�9ӛ����*-�p�D�M���w�A����t�_B@�F}t�O\������!�_IJL�9Gd�4C,��~6ڞP-fr.Q��r�մN
3�Y�.����_7�n��.nUu��g�t��ܓ�����cÛjze��N������-br5]��$8����2��֙��H�Q��<�R�@�~.Ůk����q����E�嵦J_�Bd��C�Jꊌm���	F�(t��'��b��1cz�/ȟ�y�Nϕ�����m<.�u$��G��Q I�4}��yo�D����(eW�dأ��:�j��é���n�$�S����U�%AgĆ��)�(�)tG�{�'5�b���^:D�oP\>UaJ��AN_��iTY#��� ��z�3H�B_��$8��ͅ�!>x*��?q@/�}t�;k)Xg>
��
�
�D"ӫL�/�%3>��3�;�|7L2~n�Ez�X��ˎ��Wo�o�>25�-�x��pX�1�r��k����D���*s��~̕��mGh��n�t�HD�j��&4#�@o�]5I�l~���[�VY��UƗ������֟��!����I�M���hfT��d�SϞ4rK�Ͳ�XZ��q�=f_3 ��`#k0�1���B�d%�Ç*��E2�U� �\Fb����x�GkM㮗�o�?L����Y�Ԣ5l�v�2�A�A��:�
T�:����v��맨j�%J]R7U�L ?�����Ֆy�Ox>p.C5+����!I�rDWw��U-�:ϊ=�[�6�J+�.�M0��uܖO�y�OK�U���C��w�Ϳwt�!�	�e>�c�w,�����:N[�3x�Y���ʻ�bkJ�[NZ�NI�"��m�!��sVP�����(XQ�U4W�ȡ���F8�k��U�������@����~������N1��/t�߽Qrh7Rb��(���5�A٢8u�_��6š#(�&��;�]4��a�8w��[��B�w��s���Z�������N=�t;�W"F��~���Z'Y��@k�;c$�՘��a 
p�o�Ԡ��k�<o|u��Q��`���]���Xs�×�CC{��^i��q��w���-lĠ�Q��-k&��f������H�+�9y�=��P���$�d�Q(d~w�=�_I�����Ac����I��%!�=��;�_���F@��;���O�g �ba{R��5^ �={��-kҪ��X/R�5��""	�.IL�"�O��������$�r���+n�P��*�E��[D��܇jr=G�!ԟs����4G5��%4�w6�.�7͛Ș�����9q�y���N�h��K�U��=JP����d�z�H 	���8c΂�fG�!H�^|\$����i4�ۏw����Y<��\����'�U��2MUyn����@�]�Wk_��5\��v:�_�B��6��$�R�oqs&8��|����SV7W;Z�j:�5��;̚&��ƹ��;"�C ��Y\_ȇ��Z����d�=h��F���K��HW6F��}�2/�
�m�z�
�蛣�}� �*�bO�v7��7#}R�a�҇1�j��J���*E�l�Kv�CE<����2sK��	\?N��m�x+�O�K�#4�҆WvUk��c{������te~'�_��2�e�A�������&�2���{��\O5��Wy�6Kk����������;�UI��f��%�Z���,�-����e����d���.�F�䈡�'yduoE�(yl-̸��}��tV8�o���;�!J�Qf��M������h���a�'�Q̭��+W	����}�"-��\����b��⫼���h枀a�ڏ��z�{x�{�['��/�1նu��y_>�ׅ���F�5q7�ȋ�&1˥�8��s��,k��M�r.� bC�|��r�,�H��Z7��<�[.�n�2?��Fxn�8�P{at�_��Gx�g#׎���>��,�e�^��0(�&���1Fa��1_��/c�+� ����������h_�]k���Z�axP�I��l܆��\�D���5X��E`B�S(���ow�.*���I��ڃ������+"W˭ss��������NK�>/yPr��
��<!�"/n/��*���s����޳m�G\9�\�0C�M��/���^��v��]��305x�������z�`Um/�eW7����j����G�I���)�ઍ"ڏ.p)�{w}fM�Sa�@�2:n�R��6Ȃ���v�=(�'k��z	v��H���mJ����maE���{"�(����I@�wA� f�w�N=
�V_I�RFƑ�Y�t�I��aZb�#<]r����D�%A�����h"����'��<=�;:�e��s��ÇOv��~*��6G�֝����\����ᤐ�m����ߵdZ���hz�Zě�K�4��L�,�Ϫ���*_B(��1�����V�j� fC�E����G�)_������opDYt�^����Dl�6��r� #�KD�8�o/d�n�b?��%����"�m�Ւ��"-�	Q�7Cb�����|��w�
�"=tA1p�r9^%o�Ѕ���[�3��nL�T��.����Ib�YJqer��~��%�6'�9����Z���I8-����
���`�kIE_hNI�;[�Ĺ����O���Sм��U��R�1x�:G5�I���N��ɬWS�t,X5_MvO� ��m�=뉂��N���8-����F=.>��K�{[j��LV;֩��B��=|p<>f4O�_Lߧ0���ŧv��3�:�V~?*���R˲�<[������������
i`���9����9�"I	e���i�$��?�-��*^��c)���a��2-8�h��y&�ۚ�)�<�K7N�8�%2,�����5�-V�>�.�:#�C��$�雪Q*�g���J�"��㒏3�!���n*
Z����� *@տ֑~p�ڱ���r�K�ݔ����a�o�VÑ�e�^ou�s��;`>��y\�w�cR/��Q�vK�(�Xx��Nx��:��(@_���;l�Ei*[���S�ǩ�WU��V��s��_�5�r��0�m��Ӕ��9�u�m�n8�z/�x����]�^��������v��Anyc.�:�z�Z�����{��G�T��B2sW�<�/���w�l�v�ҀxM9��q�<Z�E�rl�%�5�m���u@r�Lj��GT�J�:HT�����L;���ٿ]�}��ɳ�^���������T�s�#���z�|�7��Z1)�7�m��t�|� ,1t�̑w 	��96�yb�{|Omk��T�������
n�[���M����2
��8c�,d��.6O�W$�>_�]�KOm,�	 �}�"�T�����s$6H�D��*<�\3e�ͿK|����p�3�:j�6XW�Vs�+��s��/�\�����ޯ�5��9�j�2vV�IoN��2F���:n6�(ӷ�]��]_����n׍�v}}�^^^�,u��ۜ�`G��Z�r�G�Ԗ0�rڜFu�@�J06y(�6��R�sFry`)�)�6���Vܮe��{+_݉��O��4�Zc�S�-Q��5B��F��K���Ё�t�$6�MN
�F��pBs� WP��Ka��	�F��'n��>����Hbf$�E��I+����]��u87/�I�#���)��C
�F�MSy;�)ۖZ���9v�{���k����V���_2f�t�u�{[:���T�����t=|��6=���g:��G���#p�_?m�����?Ƞn��sBǧSh��2��̢5)�D�>��/����<�ǋ�m����d�c�ܠqwM��d� ���b40�B߾�B�1	ɕа�
�8䍘*�L�Q�,��B'����� n�)�7�� eřS�|%,u��^H�C�N�Q��Y�$K3�a��hB2r[��f���etE�Z�~��T��)]o�l�ېk�����`�R}V�=���/k����6��|Ju�J��[}xSN���ӂ��y�n[]�a�&H~���g킝�^��F;R�\|�ķ���^5�_���d�`Q��u��8�4\x�+ߛ�zwat�x�Յ���dC�$k���Y�\y{����6�1jp�? �
S�%�{���u/a;2�sηՖ9|/~M��ui��\O%�?�ˌ&3�|��H�;�OLLS�o��E_z�خ鴈�J��Z��D@)3pȂVG2��AX3�e�
1q�j�?�,Z`����5a���$��mJ�$gM�HܛaLaI�F�|�g�r�5L9Pc:]�˺���R�7(n�;5��?S'��#��*��d��淼f� np���z�����",�
e���=0���c�9����F�{�l2���0���V�������n�����6��;6�H�'&O*#��R����:O�:r�Y�H*%Ϣ�5��E ��%q'�]q�g�F��f�����d{@m�;ЪMX�-jB�Ȗ�A���?'����������m2�'7�s��l:�<آ�j�h m*X�i�$��)��f�m�׼���k������*�r��ep��x	ǭ;]q4E�̓Z�͋�Gz�`Sg���&�9�$[���!yM��/x���rlRj���r`A]{C|]Byʝ�7� ��B��TXS d�����>���6
�h2�єG3:�AN�i{��"w���i)��5�S:_�i�x� h�Hi*b�GF�!-N#̍���$G�ڃ�6a ��+2(��
���=0K'�j���1�قі%�$������^�<���ꁇIۍ��f7��T��!oG�~�\��z2�N�E�E F�DPw�z/,&N�.%�=O\R��B$Ժ�{��r�9%M�%��NS{�X����{��^y���X��*{�̊��%])p�p�����[ᵼ�_�}d>�;����6�1U�-hk���&�Fa������hş1kh�,�-����֨6�D['�e+�_Ji5}$EEe�A� �F��Nkt�p�	>�N�74�aI1�Wv��i��M���p�k�Fz�5I����r�iļ���:Կ�##���!��#���2 Ey��=^B���,{��uJ'`��.���V��gd�U������{C=��-h:jHj�O�ؼ�c=n�Ju�bߊ���&�v*q�i�������>=���fnN��bN��}*cW���<٦�c���m�I;s�����|A�&�;�r�`�T���"�e�]��|�P7��
�lڊglx@���c�tC�_���mĲl����1]�o�ʫ�%y[it�p	A�����^ 2a�*M�a���ן6K~-Ҋ���E|R�2q`[\��Nڍ�!������P�\#�i�)�4�Ib���b���76 ��n@A�4�bf"tMf"�p̥A�(C�I=�d)���Rף]��,�2�}���#�T�#t,U�uTVܵ?C������9�J�hQ���e.�� ���}i��K��M��mI��R"�ڰ��!�t����ޒ7ȼ'��}o��l�}���y`���G* �:�H]@ �H�R����z�������3T�:I�[|����p&%��t2l,�e��A.�1��F���y����l���ܛ���v��&������}}Ip���ԗp����6������oW_<��%�<�|˱���=>��*�+u�[�*���9�8�2�r��Q��;�2��$�oa�w��5����ͰХ���(��z�N��|)nc4�0B� �O�Ȕ�N 0�q��<Q��h�z�m՘V�;���7}�hS�&)���c	��]�19X�B��l��9�V�Fڑƥ1GkR��6�d�6ep7>�L��)�k��IļJ��9.!�������U�/�I�m+�����DC���Vа�$�<��S�]���P{Wm��E��-
{,彜m�{����M���n�V5 P���X0������M�-֓�|d�w��I]�)������)�ar,�َQ�it.,�%�#�㔆6q�$9/���&~�ȗd����wM�@�qy�,�l�9�����և��ݕ�:{z��|�n��mrz��;����������E��^狋W�$�\��_ou��^_���8��f�U�7����T_�z"o�����s��<)�)' ����/�'JHʣ�*M�%��k��>�e�NG��fd3��HyKM��t6�6X��� ���}���
B�h_�'>�����&Y�)���`BNh�<]eZ�,�O�*����U��I���7�b;���>XG�4KMq�zJ,����f��A<�H@�AP��\�Y�pN����D�2�Rٕэ�d.�;��*|��^�NHս��^�C�՘%���zL��w����&�+,�]��,H�p�s�u�)z  @ IDAT�����'�F���o@2�qGz�@��Y��b~&]^mR����G�˅}\,�bosB�B�'���!YNvkU�:���L����t΁�dx��J[�.��t���o��岿*�=��k�ߤ���~��}��_�~_Y������|]�{���5�p6�/��8
��Le7
���^�ť�[��� K����.�,2���>���|]\�aDZ�o��%6o�#������Z��ă�����Wr|n�N�Y�ל�k��@#|!9��EAG4S�c�ɲuR��<)��YP=���$�I�c�Sʆ	�d �6!��tJ��4֋I7�Ѭ���>j�lo�3l�0�%��?�9g��F�s3+�+֕S��w�5� L����ld|�kY�9�O�EӮ�q�L�6R�Εt�NRG���w��'�|1�^�6�CT�ESlC�r�h �o-A3��=��N�qn���,t�A2J��`�[�
�A��;B(!)�%��T�p��I{lG�����������ɦ
RG$���j���R���?S\EZ�@7A`*I#��wz��w*N\�́5�w�LB�|�Z�q�������ip����{���;�3�<�ŧ�lC�L�uE�D���~ޕ��[5�>r�+~[��[�s���F�uT����M_�M]Ѯ{ӭ�M�J��aQ�nl��\JLS�yl�&�S���j;���.4�����]��f��<����{8�Є�V7�.y��H:�$r�Z=ۘ����QAB���h�xM;_7�O���~y�.v��Ξ�|�z,��SXJq���4�>r?�?��#��NV�(H8��ǎΑ" �2�|!/�Y�@Gڮ�Q:�YO�!�:�rdd0c]X��`�T���E6��#Q�C��aK��{�K�r��Y�@�Tm�lA�-o�٩� �5%ۜdi�v+��"�+~|�@߲�d �ƈ�@��c�lrr���'OOWO�?y�|�aG�����4��V��y�F�qܸF�H�&>��[6�N�&���t��׿ M�7,��T�f�:� �[Wv��lX��@ih��K�RJ�[�2&�j���M+r¢f�۔~� P'�ߠ���$��C�5�cg��\��	z�?<I<m{�#!�s��Q>Mq�����G��Q��T��N����+�c"�Gv���ְl��K_���������&��"b"��'w��� ��J6�OM���т�֌���O��ѿј&&l�"l�C���NV�6g;��h\�y�#O9�> �r�A%��o�P7�敮�M?劳L�s��o:rh{y��o�S��~��g�a\�nI֨)��Y���mi �?���ۻM�6�ۻ�O=�m��26T�{��4�Gsi�z�����o�s��<d���K�JUˀ��,���E�7�5O�>�5�nF��ˣ;�Q�u� hut���f������y��_ba���^�kG��?t�|��p���G�ў�$3�2XFL�d ���:�;9�qJ��T��{�呾p��ˤ�>�wϘ;�kAd���T���-s/:��r�)�*7ѭ��h��ٕb�^�>���>�`g�pc�Kݣ�ҧi���ڠ�	{SE����7�`m���H�� �����!�C�o�o�r<�t�����o~���w����͛W�gϞh�R0�~��Us���QD�Kf[���wҕ��ty���g��9M��(6:�2��ą�mT9!�EE��v\&��.���)q��<Ў����Rt�&��p�^h�-c�2`��`�$m���6����Ƭ'�t@� ����k�;9���}�v���޼	eRg�\8y��Y��=�HL��kTd+%��a�K�-uv���b���4��y�&�?C'����q�]�`���v�p�����I!*_����X�=�N`�ZB�4������Jn^iv-�r��y�w��������و��4�<�W�.�����o��?l��8�E?�`(7<J�'D�4G3��)nW�+]���4K>��hyHU�$��Z�Y�d���f$�(uM]�k�%�v62�	_E'2n�D �5�Z[`?��~�����߮~�����啂��՗�s�QZ�c'������" k�����Ni�X�	@4_^��_<&�ǐ9�bo�e�b ��ud��y>�$3���3����H�Te�̯��\8q��!���$D����#��2�#�%�? �T�Z\0�ώ-��Mij��Eò��º"��;W�RDP���� ��V�U|��5� ��A���\J�~��nיu�֫��Y���#{���ꕎ�/_d0Ƙ
�I�����:g\0���8m� �N�N(�$�Q��@����-����:��4����М���`Pс܁����9�lӲUOy_��v��LY�~���������f��oЋ�>�׭3i'Ib8sR���d4���X1���'����d!$iO�� �ic�hF &Kd
0<�?IP_���[��9	��={2����./�QfLgjG{7"ho5�OW/_<_�^w��q��>�G�Bkh�w�8�G�U�.���NѪho�\���$6�����Ǵ)|&��y�����Z�\�w�����O�[�(Wڊ��]�<��.;7�\������,��=�&�SZ�L!��`d,����2l'mٖ�_��.�K�-��G�]�|�A#�^i�p,ޱ��T2&d^��;�ҫEY�]���jZ�<�ؕ7����;C�N��ڍ��/痫�y�z��/��?�>~>����2wƢ�Z�����#햡�V|̣�<��c#c�y�v�Ju���y�tr"+��1V)��^0	ଣ�uT�4���c����>�l[��MǑnn���
G�bLA�e�x�<v��t�_rD;�$��l�|���[~(�X!!������]Ҩ.mA&q$G7�faw��?�%~e-$G*}xzz�z6߬ο\I�����"�/����Փ��VϿ�q���56~��߬���߯����F�b߬^�|��l��B2Z�U���}%�is����r7���N�9e6���RKmYr̕������Bw1�P�`�Ȕ;
�XdZ`����c�W7�1U`�q�(CmyjwEW@���ľL��1HL�:_���<~��v�R�
|)�A܈�U�R����<]@�b7�ai��::H@!�0jBD�2m����en�ҩ�+�#/�d}m��JE��@Ή ���n����9���&�~T]��XļX�\� ^j��oo�����2����~q��T���G�(��A���f�L�;TB!>���{����;5(�J��ęҧ��k�����z�3~�Ǹ�k���9�y�3�f�u��p�3�<�m|��\i�<�ɗ���eh9�����6�T�'�ͣ`��m�u��S�#w�z�y�W���8�O�i�r�k6����C���ڐ?\����o�5U� O�#a�Ac=��|
�����I��N9�&���5�\ػ��V��`���V��iM�%�ܱb^�Ӛ��:P�y�E��ϩ%�3�+@�ʆ���V+��L)ЁR��0S"#�1F@� p"=�a���-�����Ocje͆y����haR�/l��?(����sa	��A[���tCp���7����5�����bCZ 4tǚ!4m�!S 6����C��Λ�\�B�֠�bY(A_�d0w�x��K�e�e
Ԟ�}��~��ۏ���|^}�r����W����v�^�^h�����q��g�G¥���e�~�����{�6#� Bm�S��/�5�Ϻ{x����Ƿ��~��O�����<���Y�Xn���8Cs���j�L������QC��F��� �N�$r�
}G'���H��<)1�Х����X�bt���#=��7I�5@���~��Sl/c�|����px��
���S������H�$%Izq.)X*�j璱�{/_<[}����ǫ�w�uGq�����w<_��zc�N�!�1q�fp	>3b����GN�	�j�@���7�9vRG�km����R���^����1�i�Cc΍�s�s���:�v��y]��.;7�R�9���&8�u�n��8�������*����|����N�&�9����k������5��R�~J<�w��|�	������q�w+���B���m���)��f�@اO������»^,�l�>����G����̏C\�O�0�F��	r� M�{�Ad��hVTt̕�B�o�Jف ��BC�!����$�+�s?�	�`�ARDz�����ɞF��@� ڃV�	hG�������K[�}p�v��톂[�r*$���C}�������ñ���v2էײ�N�7�b�P�x� �v���b���ϫ�ߟ�~���������׫���߭�������{�,�!����/kQ�H�%�9��_�E �3��F8_Ç�|���vyQ�˗��Ǐ��N��߭���'aﴵ�^����vN�p��=� N/���#�r01�Q"�:����=JѺ�d�#� ���@�1�G��
�1XR��O���m��)Oڈ6��QN�jZ����1����<p:c�#
D��eӁ5�>��S�Sj����\�JT��\T� Hw�LxW��<_}��߮�������?�]}�r�R\꽊�ᓄP#�q��L�!���q@�K<�7#�/�_jb`�>�OL�EB���O��u9sxÜ�����M�9��߹��^� �x������r�m��fS�˯u��#���VM�T?g����:�R�#���F����>Gn��SsD��: /,:�����<��v�=�i^֊�iE�0������1�0�D��|�N��Z�x:x�ȼ��A�M_���� f3W�b�E��k�}#n�����j*���h���7�j�E;��5����e�E4�砃ڑ��D0z{�g6��=-�R%랋������3����Gc��1wÃ���R�X��G��l_�G��e� ��BY5p��)y-@�{m�ZE���(��a"a��ϻb'�ǉvC?�_��:v�x�s�5�_)��rq������
��n��Ri��;+>C�')�sU���0>��7w�ZX/Vo�h���ᇷz��N?���z����ε��L�&۹��j�����n��?<��-W��z�(��Gg��pc���luj��75����R߄�a{����Gwpq>����f��?$�0H}�,��h��c��N�l3��c�!�>R Aa���1iCD��L@�Dg(¾L�]ip���ၳ�M�� �~��ͷ���?�/���?���~�:��a���?D��V?���}>�!p���;��$dF�R�?ڗD�;g�9G)r�ʾI�K���|e�9K��ky���`���܆]��g=�eV��iz������rӳp�d��y��o�L�����g��~��;��<a:�sΕ�i����k�ql�|���o?=կ�xL���_LW��x�%�0�iSK9�N���S��ãǒ�2ë0m�+���k�ebde�#�`ΐhl����Y��z�1gHHȌ�58s/���5��#��w��k(yΣ�$0x8�/c9�EI�,� �!��ǭyu���;P�w#[C6���@��J�� ��#=၌S�	B�F�@>0�R:�G��oZd���a|��*}F�̣W���x��@��C4���H���ձ�dG��ֹ�_����Y����?���?�^+���v\%�xA��-����mA�i�C�� p�-����O�_�����?���ӟV�}�C`��|�ӧ���xq����������j��:)L:M�`M;Ơ���`W�Z� ��ДbR����v��V���$2��D�D���Ζ�=�Sy1�� 4>�c!M%>� ����6��D�.ʐ+:�	t�O��a�l65�):m�͘P��ە��m�J���+58շ��g�)���ȽQ ���m��w.�CL؆]Ͷ�&�y�F�������@G�3��j^���lJ�cp�2��驪�Z6�y�Q�4�l��|��8����Ǚf.��z��z�>��^6�ϗ��ηY�+�&9Ue�����>��D��m�,��e���.t��Kb���89�dF�Ï~��I�Յڡh'_�S��l_��@�;d���{�J�#���`C�x��ZG�	���Wtb�IaZ,��X�̍��#��"	�2�H@�x$1x!9-�o��\�x�
^��6��'�!�Lq�i�N ��j�*ic�S��%�	;�>S���2(�q9>T�H��H�N>�b/	��H)�� �J�I�C�Ru��i�d+fw�������fґ>%��	�>|� ���T��V�����7߼���%B	�4�R[�>m<ugAF���ǝ���9��\/��^�?��w�?�]������~A��볶�.x�x���ė����Tϓ��"M@F�EkӘ���T�@j�rӐtr��O��'��H�"o*
!Dm��2Y��(6�TNY���d�ak"�,_ƀ�I��ѩ��x�6�Ȥd��,
qj�j�<��Z�=l{���|��<�$M���BP�eG���Ԍ�"�W�<��/��?�X�w�{�y'��~�i�J?��w��m\�?��� .�0~k�r�$D0�5Nc�e�?���g�O�sҀ���¾F=���`}^�K|�����2=劯pp�vB��j����<x{�_�^��M�J�I�����릭z�Q��X~�8Y�s֗������7�F����N)��~�D��R��5&mD%k���|���OtN5_���������G^:j����?$#c����Z��.�fA�TV�lc�k
�|*ꡊj����%��	S�#�c}�9'�m%f䄘��� ���g4��,� }���G�-7I0	\�33�<�ҷ�8����!W�A�����s��%�4
�'e� ���6$Y��]�n��%l0JN��e��|C�$OcW�0��+<�Q����J'�X/xT}���������O�>��>U�T�
{�a��b�6�
��Ф�َ��݋���.���������w���IA�?�{^����z��7
�nl�3W*�����K�]5��y*+��'���&���yJE>�&U�i����J��=��>�a8"8t��lM�@�����3��VG�7�A��B?p8�Ę�g��T��%chtg_��lscɬ�+tʉ��l�r��W��#a��V�C�#�ȋ�o���Q3�y�����=x��	�_��W��Y��C�Nۂ���3y;�e-K9[��q��>	������f����%�P�ÍTciv-��6O�,��<'c�9�Yή|U�%�����Z�v���I���s�8e��������mm1V�
������څ'��µ��n��gzx��va7��E����5�/X���j�yVu��̀�<��k4�z�s�w���.D{)^��H_�U��D҅�_����Γ�K�	��T�YQv�]�eJ{����� �_D9y�7�+����lhS� c"Bi��B�SQ���u���ڴ7�����/���PE�N�iS�Z�i�!$�'x����0#e�sKR��f!��b���/�I�X��	ۍQ!�j�D��ػ�\kҢP=��X륟M�k=ջ���U�a���t�w��c���� �x�#لM���\2��G�iTF���z	�>~�O0��u����^����_V���;�)���F~=r�z��9~�K�u�<����.��7Z�6��K�$�h3N�Vg�y@���+[/���($}vTk�(�@�|�h'�B��;����l^�A<�=q'�̤c��W����@�iղ�����4�!O:`F� ?� �	� ��,�]I1�@��6��/�5y�Pt f���=w<;!��N�&8~U�?�y���	������
�~��	�z�\e��(cW�勧�Б}�m����/��I��	�����m���6'k;�<�}m�4�mO/k�ʠ\�s�˷>���->ʮ���1~_=��s��'�Ǯ����Gw�٥?�e�Α���4��^y$�T��:�;���pT1�����#� #봋y���/����c=��O 	��/����~	��]�c1��z��E�<_��%�ʛM-[Z�$���K۫��=_��",m��@�f�T�v����v0/'$��G�J��N���v��d�*�����Hy/m���0&Z��
�pH`'�}�TJcD��
a�H��(��@(ARM���<����_�'� 0ͤ�f���82�K����Xճ1^�Х6*�����(*
���~b�!�T���������������W����+f�6b�b�l ��1;_��������տ�=����v���|�b��vƾ���ݔ����	�b�V��eW6��/���.Hg�r��L�B9y��_v���NBj|�3�8J���X�#�l����(��9����x��%hUD��� U�C	x@�� $�Hi���Xz�8lR��v�	BK��ť�م��:��,�������� ��◈��������mA���&�&���纃|���������ۧ� t.����,����~E��9��@�X��6�m��������d��>Ñ��k�>���Z�EnO��6g�y��� �u����n�5�]�m��G������s�zY��r6ј~��p�(����m^{h��|�!�ٟH����V�����g?,�|��`+�R� ���52O�Uz��~��O���9������'O�i-[ō#߶���|^
������aM�B�B��2r�T�C��:R�b R��)�s(j�e�&�g<�k�k~f� 6�n���>H]�f=�H���ܩ�܄�Kڑ��8�����G1�g���$d$.�OL�"��X?N�B�l�&ۏL��ܴ�`�p^�ɵ%��G	��1*Ъ1�<7.(���ŐRYh^���^^�k];ү"�z�O��V�;��C
9؏��҃<.0	���g�k'�G�i?闎�߳�u��k�:��v����+��s��{��謸Qcr0��QAJ/�Tg�&��t�ʲ	��/�4mz)�Ă-��K�xV`���#����5�4��lۘ�t:���(m���[��x�O�%`J:�>��J����|�V)�R ��|�?�0x�n��m~0������W+�^z���#�)�bE��՟�q�����s���K�қ����ўT[�u�H'�6�v��QҴ�}MTь���B�/��M5'˸��!���{������_�=�<g˜����̳�������s6�.q?J�v�1����zh�@�l
`� ���q����e�ߋ�����9�j�ST(�u@�$�9F0D��׌ϟ�l0v�nӂ)�[� ^)�Rp�V%��ߢ��"g:�~�t��9v��m~#��B�6�]����ե>�ğ�c	e���4G;��n 9��k�AD�ri{��PT$K��Jb�Kc�P>�!i�d�!��x�X�XX3�(���(7�A��X���p�ǀ��X[�gL���Kak�C�:0&5������`I�B�Y,ޒl�خpX>������&"^e��ї��ߢP�3�D��&||�K9�>ѓ�՝��';�z����3�Y���?��UoVO������-�Y=��˪R�����~���G}b�Ƿ������z��\_
��9Ջ�-���e�r8�����,chǰ_�΄�MwX�2"�YcGed�}�i��(!
M�ȳ<��kP���n^��q��>T��A��n��N]�i�I[r0�3���`p�A�$4RFo����4Б�����`�BuP��� 4vA	�������Ԡ�����fd*I�)u����SC߼y�]�g�IwNfLh�;.P����n薞��R���M��&�u9 �v��s)���f�7}��f�%ے e���|ٻ�]���9�)[O�W�Kp�v���ͳ��<��Ȝ�g]Ȉ���9�^4���H��������<�k�)W8u������x��Y�a���3Y�T�8o��qB)>��=j33N�c�.(�,jaԇ1O���HA�7��D%�?>����)�s���zt��o��o �V�h�6~Qy~����K�S���~p�I?6��C`\0#bS��̎��;b��|�~J>��9&�N���G���$V�S2c�je}՝�+���m>F�	<H<��G�ݳfkֱ��Ȳ|i�ϡx��Vqd[�hc�	g#A6�A��DP =u����ǒ�f��L�G0�v����Am�Ě�P�k؋�t(�«��.�2�ԟ�~��ǻ�	��#j6x睝����������_�y���Z�BO���vM8����|���^��Q�|���^�]�+���e��k=e'N<z�G�,P�bqn��~	���� �{�3΀�ϟg���N�H��p In��>�ΡM�=���A|ȉHD"��O�焜�,�DX��_�����G^�N������$�}�#�کGw�q?鏦`2� �&9@98��H�F�0��&�^7vac\�p"<�g��F�ح4�:+��M���TUȭ~��o�U���w°����F�z����1�^h��F/�����'v�d�����+O��|";���w|�x�G+Qj��T����9�Y�sld}�X��釼��9�ek�}Vrdה>M}��l����*n��&�����Y�����/���_y{��;GW-3�d/�ٞ�.�Es�����,<��93����ڥ�\Cϴ���`t�M��4o�Oyۮ��/��z�5� ���5�y�����]��я�*����:����r�W�ޱ������a�z�GG������5�����'�����7�������߭~~�Ek[̈���oO}ԙ�)�r�a�I�]%�1�IF�C��� �b���vy�T����X����J� V� �?��@�ݴ�'�����q��f���0���Wډ�06w�0:�eC����й@�,K��G�\挅���M�lك��m��@2a�����;`�h��'�=��X�t�����9fF�����U��B!���=v;� ����\��\0$�9�j�W�̬����,�)���d��BY�X�Ѿ ����c�{[�y0�1&���1g����~�o����Ox!�/$>Jg���j�כ0��9�#;_���w�����+��]�e��a�p�TFO
��T�(_��IzU�n�٠V]3�JX?tB���3��~�*{Z��&�T�چJ�Kx҉�敻��&yU�O^��z0m�7+n>ʺ�Z(�pk1nk�Ҵ�F�T��e�>��NQ�T8�x�~�l<��2���ͭK�)��(W��#���<���F#�v,a��J&|��)�t��Cs��£!&c��Gɖ����t�� R�39jb���p����շ|��w��-��_��x���ϫ���Wg,r���~'�7�șp��7��_zO�Z��-�#����>�W�7�����L���4�m�}��������q���渥�6��Җt�
7�K�&���n3�M�7�ϸ�GՏ�fL�z#�m������i��A&<�N'o<Im�>75�6Z���}˹gƝ�-�9n��L�T���)m���G�t���R�[�El�4�ht�����c��}J!(Ӡ�Xc�/��=��$�{�O�܀�O?�(GwIw�z���d�����]���C���5�9��ѐ>�\r���v`o	�}X�p?��Owp[�����*;���3��k�plLYT��T¼a\�o��v��J��P��8V��~	c�\ë��bHTX2~��W��88����L�<�U��P��;�%���?S�7��2E�Y�V�6�E+\��� �Dy*}H��4Ko�a��,e�������I�P��pF۸@?p��_��V�'XOOVw�Y�4_��m�3�f����Ϟ�ʺ/,`?s��){n��^�Ĵ��[qY�C�5�2$c*7V@Ș��Q.H��ƛm�Dv��E���>huG �H�Z2��68��ے�'�t�p���c���4 RL�2-2���	����7�#�#�Jȡ&oʎ��8*[*]�ZȎC��r��9]���_N�l�Y�G�3o�T���/!j����@L%��9i��x�5�Gx��!�(������d��Ŧ�EWvȓ��c���M>tL*���	<�,��o�^�����oih���X����'��!�!F	sz����,��a�g���������Ro����z�G�6,��}�)����A+u?\Hv\�]���4y�;X��p���Z۞@�4n�ӂ���Ȭ�K�9,�}h���⑎�۽	��k�&���wyt�{�６���o�n�\����ؿT���<��$d`q����4o�n��~5əN��q^�)\��|��N��OĔ&|�;�KZO�Hɔ�m��[2O�����3�y�:_'B<��C3�I'f���q������g��[�m���
��O)�빀��,�?Ǌq�b���9�A�������$��X�����?V�R�sɐ
�GS\�D��=��5����0���Mـ��j�j\�م]������g��Xm����7_�#���?�p]X���� Z��α���)@�e����d�rD�RfFpeNrJU|� @ￖBD�
J��T�(���l(���G��"��с�rlNDNޅ+��-d��;��%��%�Si�<d�hɄ:�mB�$��K��g�P���!;??����~��!��ë�3��_����%�Xm��Kb|t�ǟP����5�_jq*`�*\4(�:��U�U��3!R��qSHR��"@-<���T���?���ě����0F���U�43�Y�
m&��,����D�CW�(�(��5�hU@�@���.
���.��,���xV�'�����K��Z����F9B�1�^QI*a��)n)a��#e��m(>b}7������>5�]
��� ��_t(�H I]������9�W��aR��M5���m��Y���1����������z�������]��8<���a���w1�;e��bOe�n�C��xƤ�����.�L��}�
P'|��\�����Z�B����@#��yx� �5�7�t��3�N_����םq;|���Җ4�[^�����v�x��p���{嗆6Z�u<�0����n�u�O՗��j��<�%��!��kjb������9�λ�i�iuz��5>ퟟ���i�xa6�i��kȯim
`��<��b�7yy��Z��z��w������%0� L����x�-_��8���~����>����ӟ}�,S�o߼A��\��QL�;e��.��W���`��q鵣]_4��i;�Hf��蟠T[�}2�, �����`��®ϋS�+���V�����!�=�fl�a�����"0��Y�K6��-���z몈��e�"��5CX7%���F$d��!��4R8��7�i!9paV�]�S���@	�ĩfRv�gPL25:���p�yq9�1/k�Pz�CPD�a����	�JuZ�=��}ҝ������1|ʮǿ�i����?s�S�?��̫���X|a�/���u;�˟�C�ڐYH���U���_w��Ȥ�:ȏJ�A;H��*��r��NE�HZ��X!���F=�����V���������=,u�#�C������5ӵ��o�_�\=y�lur���.�)��%e�am�t(�nK�l-�o-%E��OS�j����jl�Le�Z�!�dn�%�
��"<��B)_sHIi1N�Z��(��~�`�{ �<#���t��>@����W���ob�:�`�u��x�"����l�F!;Ps%/��9cm�1V���6�����%���KI�ߝp�F0?�Iy��wM��트�7�g�˼o#Y�ۧ��D�sh4�/Qn�j:Mw�k�/�;�ϸ���v�q�O*j���]�k�5�F�퓺C��;`��9�����-����"������<�bSZ�uZ�\�Òz��:LU~}����oDf�a�3��Ɓ2/��ު��>���d��ɓ��o~̺�+�k~��^>������S��X���ӟ��5@~����m�j/��N+l��3�O�,��D7�(���y�)\۔c!媺i8eC��>`pxp��!��ӟ9,��Z����[�{K������뗫�/�Z=����!}�����Ɛ��d�y��x�\���Z����	J `�ƙw�(W#�z�1��%�wh�)���a-UQ� ���X�!����d�NX/�H9���zS.y����K7-\~@BA��j�w3E�JE�<��s������K}�:0ۢ��� ��A@�����s���?g��S�/q�ӎ���puHy�/�Bj
K���p�B�FA��樬!�0>j*p���6LF�9�#�RQ�7�D�)�QF�
ѻZF���Vj	��!\p�p�iu��;>��6�p_�~����;����N�����)1��[ގޓ��JLY��F1
Z978������:�=
����eΆ��s|će]�Cv_�X5]��GjP��xȎ�L©�0��ޖ�~�2M�§U�����{������'�ߣx�|}��7��t"�{�rR.�[��fr���\�o=X�TI�!��*�A�����k��?���9?�<�:���!�k�����r�'���2~���ĝ�� �,�V����&�o���qMg�3�>W�6l�����q��%�e�i7|��ԝ�i��-x�iS�m�M�]<J�i���$��M�����"�Ϩ��[�9>���hى�Cgd~�Qe�(T��)�t���X��.F�v���S���\:�̝o���Z�ǟ�^�3�o�1�ȋ��M��C#Mྂ�@�T4���/��fl�q����qGy�`q��e�b͗���p�xu�Qg�1���׋�~�v�:E��s��N�	�dc���[B�Y����(h@���'�an��L*��=D�4�¨o��H����cenHgͱY�X���xj� H\�j�����-|�+�g>�r
�
���#���,ڔ9�r}�g�y��)˻��"-0\�UֲJ��3C?0_��Oo�����J�uJʉ'�z;c����l�%��^aq�|�ɠ�@�-�>
i��@B	'PJ�SM�*�����aJ $�� 7���7l^	�Aj�\D�r�$ � ��7!���͈X��x��w�)��u�蘵lc6/ץ=z�d����2�_��z��+��ybQ��!4�Eq��OU�L+)��:�Vi�M�o2���}��a��������9�:���/W��㿮����S��A߇�l���||��o�)HNz��l< ���ǫ��]����������b����[��j�2>
W�yە�L���dA�9���R&���6�[k�L���Ca��J��o����EO��yk���e|����>�S��g���-�2�v-i/������h.�ę���M��9��v������Tx�[�=}��g`�dp
��k�,3��������֡�xd~"p�c_�?����1w�[~B����7��(RX�=,��rF?;hJ���aA�ZQS.�ۣ_=��E��%Ӗ,��������3�����"y�]s�.�0��O�M�=�a�T������k�sAg�*�o��0`;�b��,�g����s�v�z��1�����.�.�cl�a�����n�Wnj}��4
pIw0���L���q)�`$���U�i�Zj�?�\�>ק��^Jy��(ʋUe�D���F�!��~$�,o�H��^��`��W��ME����!�EG���.Ey�ي���$v�������w�P�NV�O��v7����ߺz�71Kj.�re�>i��ea�yv
����Yp��G�*�6:b��]7��	���+T�LV�B�*a���"i�B�d���Q�7.���5R�7�O��F���ᓟ�.زU޻��F �{���a��b����J�l(eѼS}%4��Rf����
��7w1, �I#�V�}�o��  @ IDAT��z���������n�}�x�Sy�;��x�7{[��gsA�� [��	��抿}̩GLu>Ą�͋�~��7L=���]5ʡ����6�6��7
�8S��9�4�'�<������S�jE���X>�A���)DF��M��[�A��ԏ���U4�ם�]�K�ߕ�}�n����ʧ����a�/�w�K:��n�x����L�-���-��w=.-�zԖPӽ������v�Eh��fK�wFI"��̃�s�s����ˌ|<}~�������5&�taY�(\�iu��9N��m�v�0-,Z�vv8���Sr���N�6i����Fa��?��J�-C���@��H�h�lעRx]v�'��VEj�Ld�W>5zeq
�ʑjK���f��X�X�N��W(�=8���=�i?�9y�k�%P�+����ߟ�jūr�n���X����1D��l�( Nx�@�<�c���x���%#33�e?�[~�Ji5>�x��[��A'Ҷ�4��}�� ������f��T���"vu�nu���՛Wǫf�VW�Rv�!@5J��pگ�d{*��B��\���`���s��wiF�n�R��fh�Rl
$�.���G�X�&�k��P�5-I8�o�,��t��' h�&P�0$S�������+��~��THǄ˴&1�a8�ŉSA��e>S�z�\T���{c*4g(�*!��F� ��
.�~��&���ld1��t�̷e��0 A�?�$N^Tmp����ի���+
����y>z���C��(?|">vP
� ~N=�}���^}C�}�u͗��#�w}�Փ�o���iǯ�G���B�C}$��PIOs�o�6Z�5�S����R�Ҹ������Z=��?r��	�r����a�փ���hk���\+���� �y�� ��x/sC�E7/3��kg�����������M�4�M��v[z�t��2�K�Ҕ��-_�Sk���g��s�i����ϱ���̌g2�s9�������|���T_]Ho?dڛ7��b=���|��>���իwH��e���$��������s��p�斸t��:0�[E����{+T���U��q�B���$�׼s۷qo��Y��W�~�����9f��!_�B�%̝�҂x�ܠ%�����Z�k�3A)��c�S�P����%��9w����&��K	���R:����[Â�r�^�=�ɏ�<O���꺛sDkL��2�X
��z-=�|�CKb��Ƭ��
�ɴ��%K~4^�.h܇���O������kxz�jRǜ�GM��y�3�~ba8��!	47P��d���B��3mu�GKW4>�����\
�F� L� ��	F�fa���HJ{�b�+�A2���&N-VK��@-�Gx��G�R��+~��DV
�2g�q���4��]SZZ��ЊT��.�=,��ݡr���P�R}�iM;J��2�gq5X-��_CZ:���Nd-DiF�y�gT���`#=d��1��vv4N��i�c�Q�x�G�fS�ͱZ)YN��u��5`0I���껯_��?~�Ɇ�"iɳ��,��N<_G~�̢HKU���U �R)Ĺ�ΰ?�kC�v��\�w�a���p�<4����]��1)˄���;��w�K�%�e�S���_��.�鴎���o^�]�g�ms�V�#�2δmq���m���s�%~���-��7x���x�o�5n��t�o�6�eZ��G_jػ���������������ױ��MN-� ��A'>�d�Z���z�+�j�_���Y�ό?���A��Ґ�z���X"Y�u����BovY7�2���$�{r���Ȍ�pg��?L��r苌L�0#8��2_%�`��DO�ȅ~�	]�bo�m+�f��x|�(c���Sh.�y����3%�t�rf_.^r�L��Q#+g�KMsX��π��2�!k��X���񁏡@���B�a��Q�`��(��^��*� �����(Rk'pI�c�z�rV�ƥ�S?�$s\ŧJ��Q�_�Z���f^��Cn���R�G1�� � �]#�����د1��T�A�2�^qv��)�W�^�H�:�2�Q�4�9s������+z�s�����S�!z��R�R@
75a� F�J*�%Dq�d��WK����aH^ai�z��>V'��K�x�Z焠����8�b�(�F�2���Q����d�[�?��'_����K������Rr�no�/�Z&��
Fx��@����Y���*9���`������#�y�!TOc�K��xyM�b�
��Z�T¤�����Q��ڱ񆅀{X�S�̬'/�yWu�V��v�ս<;< �����g���������x�%�-�J��T!�6��e�z����p����ʖ�q��~�Ӡ�s݆�n��M�Xv�����_�V�Є���=Z/�0���K��F���P%yN?�E�w���o�c�ϋ�i�۱>.����Ԗ�2�S�>�7�ϕa�/���\��pX�o�g\/����]6af���n��F����LCvYG@��-�w祐>v����]�$ǒ��ǳG����zŬ��'��R	�s^5z8�WA�������`��I^��dЪ��㥀����+�M�>��?�A
S�H%��"�D�ߴ����9g�����{N���7���x���/=`�/���H*����3"�T(U꼻n��k�w�X��4�;k��!
��t]�p�|]��Ԣ����ɣ����T�P������2��b{d�l����3A^%c�v|TTh<7��w��)���7<��a��%K;���#�~���V���V:3�c��o��1�c�b��;ŪF �66M}�O_��*֯}���]1P;{A2Uu��Q�(��1�#�beT������[���aP�4H�-��7�����eA�l~�ae�g���ZP
�؝?�&p��r$>�;���]a\�Q���k��]��Iږ��!#}@��/_Z4/x�xρ���!IS	;���C�Ey%� ����i�ew�)�c���:��/�88�ٷ�$T���,�|@�T�pJvc��nG����Ό���ƾK��Ž��dS,@�d�z�8�T�=������8S��,f��j!����c�������p�\�?�V�G��]��a������%�\�� ������p�i��*��	]w�zܶ�pMs[�w_��p�ǌ;�o�_�%l�-������t��a��;�%N�7�n��q�﷝l���wJ�<���8[�ш��7�܆�<5N����p�n���c�gf��x����X�k�'@�7H��
�~n��歞�"���K�}��(�ꅱx�T�|h����ǟ/���Uv�_�%*V.59d���g��}������g֎2,Sw6�����=��m�[�7U��qV�ę��*I� m�B�qZ��*+��b{���=�U�}Y7��,���Ȯֻ9VM����w�g�`�hA!;�����t�Űz���|d�٤Z������0�r9LY�T�Tnz��Qޜ�i��Y�vkg�u]r����r 0�[A���>yW�q�mxL�ǚ��0��>8��n��9�	�/��0ֺY��u�oC����_b�z���9�E��v����v������B��#�;<�Z�а=�U��Ge�*c��4�1~��x�Zx) GR5́� �i\�w#��k]L��?5E�0�2wT�Pz\�� �� -n�C`��&���64�z� J���|���fI��3B�Pʄfn�1?⣭�>A|�S�0*�?q��?��T�)
�|��Ք+e�el\�d@�p�/Q0���i��.���@���&s�zKyOY�w�Bt��.�OY����,�%�U&��I��"lۢ��)�4���=�x�� �Vf�������u��]�eط;��.a�2 �(_Z���!�Zw&�&�_|��7d���|L���P�7y/���Zės�.� m~�k	cx����]����o�e��t_�,q�ѿO\�Ȼ���C��}]�ϧ�1f��nC|N^�k��J��>�g�����,]**T�����4?_B�v���s�ݟ�^�z� �UǹXA2�V�}/]_����쁥�t�v���9���+�Ҝ(O�l���G�bY���M�KV��߬�_�Ο�}�²�I[�Ӳ�QS����违�p*�s̴z񎎥�CZ!��^�U�kl/NSh�u���b���/2���ŋY�����4��.L`|�q�8��A��C�:`����hjȸKţXԍ�Q����]yn���۟1�V�0m3�Ln��=�`�c%Z�v���D�gL��2V"�]�2�D��������f�v�l� ?\`�c�6���4e���r`(ݑ�V�¿�ߊ���2�뭬m��U6LW�je�b���H���AU.�u%h��S�*2T�"\--*Zr�e�ƃ�I��]�N��B���A*9�"�R�0A[K���x�)[ɲ�)S��+M��C��<��.�T����Ȣ�}Ú�3 O�Z�?~r���@�sd��֡(h�dT���IZ�H�f|K��lg����-T"1�2-胲s����.����{U��9eIQ!��Go�\uv*'6*��C��j48doC�A��mY�G���p��v� �����I>�T¼�P�^�$)���K~R�V ��V�$��}\A6W�	�����|�q��O�Iﶫ���q��|�a㗸��v�6��,�0l�2~I�����^��}�g�.Gӻ��T���uz�4�︥{'��R
�q�FZ!�u�E�?�7X��Wb�YJ�z�ï��&O���I�M?�����K�4��|�6�0�����.�c�������Ef!��#��c$u��!�����M�V�-�<�G�U"E古q�|���*�:e���'0i�g�~�`�<v3�T֙Xx0 0x�g��Ll�����l�ƌ���:��S�Oɕ����TJ�֮+������(^n�����,���GߣD�i�#��ii�x���q;N+[��
�o=pY�,�i�֭c�u/��� �*g��!͌�Կ�.����:2�8�2j�alv��Ǵ]��QxA��ڤ&�ُ�b3��K�2�v�7�<�)�W�f�+����
k�ʴ;�V���!��5��>[�����7�T���t�0l�؝<�
�����D���~���d���~H�&Ӓ(c;�����\�\���T�E9��P1flyQ�E�3O�O���`��T��e��36j-N΄�G<)G�g\n~�h���F�Ez��l�y�M�}5���lV�OQĞ&��X��?e���������u��ʼ��ʥ��4ʫk�h7�]>F�K�'˔{/S��(Y?��NǗ/_Dq�`�V^�sʤ��&�~;/i������N���Y����S����&�97�]M<�<���ך����y�Ss�6g����_�b���Xl>��������K�.�2�L��ٖf��_��o������ttg��<:�>�� �k�=7S��Q� $Fg0�Q�p�k+z���P��i����1��0b�I�*��Ø��O�x��MG.��x����çh2v��<d�����e���q�Q�zk>��ȩO�`L/��n�\�?7�M^ĕA����w��c��	�J#3^b�b���!?~�ζ��Й�Z�Kߟ)41dz]�M�_�,�E�E�b�bШ�]*�N-j9�"�u�+������)��c� yx�7�=������(3��Y$�l��}��ga���Y��Å����>�-��&�dR��b��cw�g���}�M��*96��B�NK�L��"����:F�T3sj	F�{���B���˩.��V� ���P�e3��m\!.��\�Lڻ�y!��#�BP�����xLG a���M� �R���<y$��ھ&A�|��]R>Ԑ<��*{h�L�� l�h4�UoKU6{]*����_*f*-*/2b�]��@O~���T#���N��6�Y�WB�K�q��4�Fy�<�"�zM*�k��?x.M/� �,`��_�q���sq�"�V���������wH��Ŕt�.%�5���t$	9��5W��٩UC�������֎O��8>�^���-E�p~L�ī�LĮ67El!)/�$���/��4n���[f�x��/��ߖ.��mں3��_�;�g��������po�o:�JK؆���|����#���ڝӶ����Ӷ'�j�hl��an��P��-���vz����5��9mG:	M����83Z`Ƅ����Ō�ؤ��F�;�2�X9�痲�W+G�/o��#�l/K-D'��C�7,Xw��/��B��2�@N�)�U�O9�����2�w�`]���O�uh�n���,bq��8�;�,юV �g�)�`�J1r���Z!t%9���)#it>��:q�����$|�+�V%�]�(`�5����/����Qz�~!{��O>@�r*xy���#�gO���Z	cY۵���G��l��L��/��Ơz�.��z���r�T��Dp,c�rǾmK�cM�c�!_�y�,�~|�'�I:���*��Y�o����k�aeJ*��0��RA6���P����/7 *!�9l"�(,«Th�RFUw6N�4ׂ�H�AN��ҒY��£�bF�ɩ�Lm�F�Kł�[������<x����V�o �g19J�uŹg�Ei�	��+����n�qUf�)��Z�.�*e���sG�4�$Z
+��Wt�9�=��ss�?ʗm陃��v�d��2PQe��,t!eI��jy����\�}��EP˨f���'�-1:4Tl�H�Q�T������ڳƼ���ڼy�c�^����/�t���c3Tƚ��+?�H��/qE�����3��3�6���D�`�F-��p˯�?ŕƧ�\�ݖ�m4����{�WӺ��%N����VU��K�q��8w�mKo��o��6|�f��7�v\�3|�;�AiF��oOW��*zK�ꗖy5Q���;��c�8&c7!�*_~^υ�~�g�g<�m�n^�쓲��8��¾��/�Fػ������u��7_���J�/�*eY��Dq�{�0o���޲��2���K?gI���p#-A�o?e�~��mcB}t���\�
���HCh��3/�)A_̕�H��>WX��<���{� ���/U���ߵ^*`�D����~��!�ٓ��W/������*[�7v���(�OT���qYC=֗�A�DW��G+��x������F;	�*N���2f u�z�c�QY'�:��Kq�Q;d�� ����_��7DY�˚@ۉJ`e�)��-�7#Z��h�����*������O��Ib�`n������U���ǫL�**L���)��YH����[ 
Q8��xvi8*`�X�L��й��c�X$�N�3�;��3gq$y�r��]C��Q����L�w����Qf��xe�2(��9H��xՕ~R���:<,�Qn��􄻆�D)~.�>�(��ț�0p�4�7��%an�O*� ����$�>�<p�M��88ֵȞpn�>
���zw1�D���MDrG*;kp�֍\��'�U�̙Lv���/������g]�8_��&>�/m�v\mиkW���~-�s>�owY���%�ܩl�븛�:}v��eZ��y����o�}�M��|�M���M-�K��y�<5�9��� ���MZ�mB�fr4ߙF��4�5���	lK��r1vM{���Cn��6�l{��`_�$5~��%II���6�2�	μ	%\�%�[&�;-�06�,��� g�}��>�<t�����]�b�U�lPs�펛':\������[�M�/q*\�PfF@Z�/7%N|`"_��R7W��>Hi�ВFC����^�-^��6Qf�a�)_(�QX3���K���A�(_Q��ia��x�z����ųG���z���ol>}�$�!w�ʏ��}_���ZɸC���\�Gt$)��I,q�%��g�r��}�q���]���X��m���.Y[�T�k�,{�`,g:rw�#6�k<~��M��i\�B���`�}$�hP��;H*)�1�}�ͷ�������o���#!�4e�s���l|FH�H�#_���V[=:�][?ף����,�Db%��9������y(gr��l7�'>h�aT�� �O?�!qv����ߜ�����w�����lv*0%i����R�$h�h�sx;!O����l��$S�Џb0Φ�2�;��(s�b��J��╊��$����h�qU�m�� q��4C^��By	HҺ�LB(�4�Y-��ጎ��O�r�����Z<O|���]5��3�MK�	s�G��ʛ L5��J�Ûm��a[��!��4��iE3�)�z��ܭ����]E-y �+S����m�p^	��?�J���gp���7�σ��`n���	f�o~nr�]Ҽ),��}	3穿�[�w�iu�&w��y6�#�L��:}�n�_���+�Ư����u<�z��&�Q�4�ZMu��:(�զ�ަ_��_s�q�c��_�ϲ7�M�^�%��U�y
�Dot-_Y*,�V��f*
���wb{�}V���?�-h+W�� K�k�\�!yѧz��O�:e����/�c4�����/��GXsX��ұ>�������QB��a�� ���U�%F�qb�(�@Yr-��[�:N���Ҕ��h��h$�������%��u���->*���M���9Ψ�9��z�]�v����b>av���ѮJʭ���p�����կ�}�z��d����=�#gT,���$~u�Ǉ�k6/��[����k����{���[Z��Rԍˋ?ye&�2]T\�$*�.zc�m%zqo���B��1������;�'(�*���������
�I��S���М�}t�|닯V/��M���KCE�����R� �ʷ�U�R1:Uq��a�8?�i�X �w�yN����ޱKP���a]��7�(`��8%ex��U�S@#��T�NQ���q�Ï|��~Z���t�����h�.:?s������B�d��-S�60W�E�d��,�����G���I�e�@�T`M�*Ǉ�v��^i�R	��Y#�$,i��m�V5&�0�!��Px��A+���5�J$���e��4�hy �֩<�����CH�P����1[�lf1���n\�o�m˫��#<� {ῢ��7t�Xu���0]��.|��y���T�.���tg��]������G�ߔ���7\�vx����x�7�l�5n�5��<5~ô��s���i7�U�>3ŷ4g:7��fƝ�o�M�*~:��L�^���ND@�<}o�m|-C鄖�`�_�5G۫t�k��%6�h�����eW�L��[�����5y���'±(���L�F�y���;v�����|'�1�����H5�0�v�����0q���t���  I�?RS|�DK&�����/� 'C��h��_�Ex�8���#�
V\d:ю�&���������D\[��\��Z�T�vY��B{-�Z��(���hg�=�7�z����~���%q|w�q�������y�AY;������B���շ�(.���LQ�Y�m�UA+c@�OyW�I�!�M�ˆ;�O^����KS�\r{���a�`����s6 ��pt��Y�H3�T(`���[%��_�)����O���W߮�N8�E��cC��s�Q�.B��Q
���Cu�Y(�����L#E�	��ؾ�V��	��#�>�G���}^Z2�����T�0���|���P̓���ɹ��*{����c{��ˣ�����؛w����g�ʜ���l]%�]B,8�����4����C	�CATo�+���5rQ�V��;��x����h�V���8�l�
`�:�d��e���7���Ɣ���Y�դ�0�ÿ|W!�ꁿX�Hܡ�*NQ���C�/�7���.�b��L�� �m>*o*`>b1�܇�MF�\����l�k�J�iS��I�{�9����S���G����?��)3墜n�Zn���&ZMg~��G��q�/��[��'|��ov�f�k�nNk�vMۤ۾7�m�ٵ��,o�M��f����3����6��Ҥ�����g�r�w�u���[A�#�
_<~ť��D��9G�9t�|M��]��M����}�a�/�<n-�}u�tN9�|���MM�{�4����c/��G�<��������w�kH��/�x��IQj�6��b������?(Z�u�4�!%<�D�u>L�&�����
/�Ƌ�CXY���ʐ�R ����]�F8�6�`�],_A�y_N;~������������귿b��	�HL���]�zr�bR�yǸ��os�c�p�����<ɇc�u��<���t��o��-)D��˘P��!F��m���Z�ę�c�Ӡ���S�������R�1^~���[����ʣG�W�1D�.L��>k�6�2c�m��C���-?���J��	�<��a%Vc�.BwJ*q��#��aD�`��䥩RA�f����[��{#M���'�U�2�,�1���T)B�z��0���1/5�G�~������1��x���|F��/߯��}�E�����H��X�ܮ{NyT
ɣޞ�W	��FyM������O��r��iē&zH��BH^�M�c/�
緼����%���R���+�(^%k&
�`5�z��H��l���]�*i�V$�����m@��6�����-g�-�hvm6�kz�'���R�"��e��Lҿ�?�e�nw����f���?��6:7�w��nÝ�|�
�4f��i�.M ϩ��-��h�����o�k���Қi/�:�eY�psx�mt��D4�L���<i��+e0Sˌc�iO?�ڻ������8	�7����=�W���̌���4r����RrX+0�ӱ�:$�3�П��ZI3W���/4qЯr�ej��,�$R�x����Hބ�rr*� �x�p�cn������+�P���H8��y�wz���8�f�c'<�}����3<B�������~�b������g�OP��/�P/��cB�$�9$�jf��XZ�f(`��&�E�Vo@	Ңy4���X{�wr���7JaG�}�%ew&H�
a꙲�LK��m *��U.�n"B�ӍQ������#{��)a�IW(��<\=�m�S�u��3G'X�($@n`����2�1<9�d�E�|w4���+%EL�f��``�Uk�J.>�]��/����
����Ap�e$5T�� �n��}�hZ�<����:��G�&�>�����o�?��ְ=��:ek�L�N�><~��.����x�G�c�������o�BT������ ��X��%޸���C��3��tr�(�W���<@!8�2O�+�_�W�bb�G$�k:���_�+��7���J�4@FAm�L'A^��7��Y�V.��S˾�<r����?�]��J]�\��������}/y��A��m�t٤��9�;���}�1�LsN���&���7��a��/���?����j 3�/��K�M�������4a�x�_�����?[�&��������~Ɋ6�ê��4��:g��Xm��Ve���.�� �ZV��.f�Nؙ��X}��%2o���:$NX�Q�0`�s��e-���cՇ׳�(�n�S�͹�J^�g���AFR5�D	��KX_�G��WQAN�>��i'�c�p�%��G^��h��5ء�����s��0�2n����MW�o�z��_��W���7����܅B津2W��x�7|{�o�"|����٭�����X�>��J�>;N/ر�������ʘ�=y�h��D]�S\�NA.u��T�K�o ��B��86��b�Gb�?R�;�����o�^q��	e�3=�9��㜳��U��Z��S����`3�|T�s,<����p1��>h��m�Q���<�U,,E #�_��u^	�Њ��0�C�Ρ03��V7ij��qϬ��$�J�"�9WCK�B�"�Q�>a�K\]u�n�W'�a���\]�L9Y[���=���T����6$O�ϛ	<ˏe��\Bm�����W�%�S�MCb�X����+�@xJ������B��A�$P�=�_9t�@�'�|�b��{�L|�Lc�G�5���[�J\Y����6�\�h���A�ީ{��B��b���a��M����Öy��i�-�����ujplKk�/q�~ӘÝ��7�Mn�0}�k����aZ�u�ކ�q3���tt�ٖ�s���]����a��R���Fc�k�K�t�/��L���{��ݔ���z�7!���u�����Q
 ��[r��0k��~��b_#�(��ɮk��'���B�������-��ܛ~���Bq������z�M�d+��j��f�NB�i �R�0���߫c�'J䂸�V���G��A���:?�!Y ��Q�x),(\*���{ʽ��r�#G1���y�l���|����~���w/9bByyd���*��|����Y�"�v��hQ��T����1 �Bm}g,�,~�:��=~�'��-�G�+JP��
Z�[��,�%&l��ײ́�_���<˓�P��������_',�:a&��u��>��^0��(`o�.]� )@ֿω�$��y��ϫ�M�.�F��{$��\ԡpɏI������p�y�!GZɸ���@��0j�&�J�x}��uB�D�1-�&I���2xG�%8�/�1��^� <T��o^���_��Z�o��g�����.�xk�"=̹m�J�3�.9K�I���z���
�ѯ��Z?V� �����Z�X�@;�n�X+�@�7����RdL_ު���m)�
����[��мI
��Ao���U���YGM�V��Um�ځ��z|��A�l����r�{�rv�
ߑǦ�sN]�9n�ߕ>��~��k�wܧ��v?O���M����M|ܔ��K��`缶�����.Ǘ�ܞS�6���w��w�}ҥ��6-�:f���� m����5��I�'xב���=R�k�A�����n�f_�W�	����Z�;0^8�t�!Q�rVf�81"��b
Bѷ2ϱ:�~� �*~��7�3x�1��T▽L��z,O�pc���47n��k��N���$�X����jk_��h�B���uX|��G�yﳹ�S���߮����5�_;*g(1T���=F�'N/p��gϱ&��p�L�1Z^T�2!0�X�X#Jϰ���3֣;E��ͅ��7)��g�b��
�0�'ĵ�d�st�O/�k�d y8���V뛚J�7|���͆O�}B����Q����f�L;2����p"ķ��oY��{�*+`�] ��%����fM��,�R�*WV�&H�,�͞ǵ���l|Z�,A�J�j ��(9�V=��Z��A6 ��th�}��y�apw5~@!s:�>\��b���|���x��C̑�T������=����fJ���:�vw�JA�g�E�����Ѥ��T<��kۓ�~��P����%}��@�7���D؈�R�6�oAD����ð�B
�:Y�UW��M}e�����E�����`%��!���W��]��!��*eʭe�N���aJ��jM��,�hY#��#?m��+׏ddI�@kTÖk����2�T�%|ӹ)�N_��?�n��]i6헟N����g�7�e���&t��j����[�wz�3/K�%O3윶��F{��K�ͻ�k{����a�C�m	����b����L�,H+�}�p�>���z��N��(b�y��p���;�3�i�Dn�2q�2.�U!���^4c(���.\92;)HK�+C������@�?�j$�����:��&��4�ʵ�V�P�>c3�񦔜4��@�T���f��g��4�5�o�z���~���o��Xn|#ى&Ƙ�|���;�8|�{<��{���գ'/��3f``��B�c|�@U�u�Cט���j޲`���1�0�Ü�C>�Z1u�Kx�J�Tr??9:ʺ >��8?-��*�m/��fX�\����揟��a�Q!S�*�?���������n��{r����X|<�Ó�&r�p(`*MS,�f��V�(~�����d��a�$����
p&9��&�"���v�	5a-M��q��N��9��b��%~��]�o8���m�*^0�<@@�]�6hdv��8�o��B);���Y��?q���ܲf��瘬�� Gj�>Ծ�P�-E��dWqi�;����$� ���%D���&&�twd]�ɯb���ͻ<���X�+'(H��r�h'l��0��"P��딮��֑$U�q�~vA�x�L��<<�G�S���Z�C��[�W��BJ�Ed��o��L3��_�ܖ����7ћa�/�m����F��4�Ou�������)����K�1��>�f���|.�m4�r��Kǅ�<�ןX��_���s���zi�ﲯڡ��Ό7<�YB������A�e��uA��6fa�/X��~,b��2����� �����|I��\*`Π�㍙Vf�=�x�lZ�W�q�0��K�V�g5L��@�l-{�*)$.A�O����,��Ͽ�ư1����D�DT�q?+�́�0�b�8���ߡ|�������8��i���h
:Ɵlƣ��(����w_1�?"�Ml�3xN#2��a�L�`9O���r�=p�����S>��O߳����[�5��{�GΊY7��(aZдn��k��	u����ܮEs=�왵9:yGQ�<�A��I�l�����]T�� �k�; \�~��gty��7�>�p�5�yD�����o9=��W ���B��U �N�jX��*I��M! �Øʑ�-Cu��)�=-`jLNj�;F��c��8a��P̀NM:���_��5g�4�+*��iNy�q!>8���~���J?�̶Q������ϧuʻZ��s���9���i��a�?��i����#DH��3Ïh"�,zk7��2�y�������>"E[�P_�QUI!��zl-�U	��%��ж�x�'k$�d�����?J�F�%�i��.���U��t.����F|��潼;�n��a#��:�0�������r�����t��q�_�9��o��3~�M�q�t;��nә�縙�9�&x�ߙ����v���Ļyݖ�����2�S�ҽ���&w?N�{3��-T�����S;��d�)�W(-�����H��h+�j�#{�K��1P�J��5a��al��^�ą�^���0_�sn�*IՐ���"Y!�-%�&���\PH�k8�IE��h�\p#��|G�k����uK��ı�ST�<fB%L�/x�1���W_�|�j���2�Č��F+Q�3V�����3U�9���Z�b3�JP�uz�e`GS�%(�Ld� }������)G]p��3Z�Y�3�\ �4UOu�t(n�^(�փcS�>��e��ܨx����O$ez�dF��P�SIk9V*Gj�^�t��#���hCtz�F4R�yp̹Ǽ	`ir���t����L�_��n12h��4�l�a)5e%G�o (I�������i;�Ҟ0���7�+�>����=#0���J���d�K��7�9�;���,NeQ���O��5w��4;%����P��R9���oX���?oOLAZ�[�,Ѓo�T���*��+>��KO]6t�B�X�&eWiM+A�ǵ1䡵��ߐ�r=T�V\�*�±$8��OvU�Y`�m�rUI�mC$^e�:����D���pU�/8�O�6�-^�g���˳U����Muv3���繡;��:���?�]�0�e�z_�c����߇f�{��`���v�g_����6������a:|�.ޛF�m˷a�m;�t��g�����isz�-a;��K���5����75�P����y��)��`v_�,#o
��ż����5ϼ�1h�ZƯE]ˆF	g/4"$,c���BƵ�W-r�7x���cv�1o*y.����a�4�)  @ IDAT+�� ��L�p��O5�E.���㏑�@�&�A�� 	�q&������	a3W��g>E]�JY��$���W��9˖�Xh�7��[4\�s6��(_���'-���_m�bM�a�]�����p���}�}!���G!M��9�@���X,��$�~>~��q������՛ׯV?��w6r
�m�}{̈���̸����v�SZ���MQf��˴N��*�ʗ�vq��[�V��LYB�y�X`���,�]@�W0j�.���ɠ%s`<8��*I,Tw��뢠E��Z
�5�,��z���ؐ�ő49����w�b�r:�9Y�${���0��z�5
�L�^S�n�W��2'H���9��W����M��Pt�YF�Z�H�mw�LW�������_������ջ�������p-7߳R�$�M|`���!��ʤ�����5�*�^1@懣��ZIn�!m�p���E���rI�[@y�D��u�ҋLu����xD��.!oe6`�+W�#��%?ah5�:_;L���\6h!�NѸjS�_�+/�݄��N����)n��q�Ꮏ��g����wvoʿ�����L��}ݦ{��>�o��o|�Z��F|꿚��7�+߻җ�5����)~�Y�g)Ý�ęÎ�h������<���]�'_���E�����Q�1�q�1C{���	;��8��T�H�xJgi�U�����9g��V�\'��qlYsd�%=�K�Y~b!�kk�6�����B�?h���ˡ��][�q�p�5MrׯM��7 ��Л����A���s�)������4=�;���z��m�d��/J���9��=��9��Ca�|xX�]�#�N��U{p�R�������]�=;����NcUK�0������ӕ��v�?�2��QUho�S��Y�-e�I��L����F]kq�T	bKc�@>,W ��\(����z����9����]p�W��f�f{|+&4i�ry�����7 �������(L|9�+����$x��]_s�W�?��
�X��JAQ�,-��}�pp��nu��`��P��I�9��</�Xl���v�!��X�~��_��G���O�7(�>��er���w��璝_a�D	˜~�
9w���4���0�oԔP�D$2	i�)X��ښ������::���FJ��T�%�x�(<*��7o-�?7X2W���(UC"���=혃X�i����A)"/o/��*��F�q��1?Xy��5����[�t�Vg�_e�G�c++E����G�}a��������}���_?�q���S��a^�.��/�5�v���e��7����<17a_}�����u��U�yl�6�(`��} ��;_��oe��)2-� ܱg�`�ӢE��M�����ٗo�y!���Aޝr;�s<�[������YƦR��;J�cy8g��}��&?p�� v�5��<?I-�L�F���7?���g�^5<�,�1���� � �R­�nD$�Z�e�/��#<y�t��'�2�����ʏ{Q�F�>�K��m�+�8��N+Gf�c��k����l|X�:��x��R8V�`dq#Ż��W�|b
uY+Td��H*��[�)���.��<@9D�rm�
��w�B�8h�BJKW�q�R =\r.W�b3B�="�0b��L#n�RȬ�����*��p�-�Ft���7Mu(?(*W�	K��ątl��F�Dо�-��,�c�֮'O_��`�zĎ��XՌ[�*OG2�#�(��Ï��m��2u�^�b|JBs�4��<0��AR�^��oT�NW�񧿯~|c���y����i�|�b�sv���f�F6>0Up=ӥ��5���#t�֑kOŏ�A�PQ	� m��exs�	6h~H������]N�a��/���p8�j2�Gj�U4m��զyV��|4�P�������Hrr�WxL�x`�c�~�ۄFv�����ĉL(MkN���pnw�is~7�6�m�]8�|~ߴo�o��ӝ�f��������^��k�7��
�p�ϰs|�������iw��0��7�2�����i��y5���af�e�?4&wN��l��%�蟈���c�9f��-�?�f9?�'��%�+X�UKH2� �^��RʜӔ��1�%�����v�Q���@Κ���򐿜�Og���'�q��JX�f6x���JD�Fps��|���B�j#^:�N1䇜�٤x=3gt,�>
���Ϊ�@�������b*��r��ǡ闙ya<f��Ɠ�� +㑿�]_���K�C킍~R�ji�AOPOQ�v	�]
��#E�xDG] 	��j�t!�aJ��y�)�5�FP���ᝮk<O�ƀg��[�d�Ѓ��Lv���O�4�Xu=�a�O��AEX��⒦��4��"8L�;D^a&��e�{��׫G�9������|���9x�фk�-> f&^f�c�T�<n�7!ߝ���;;U��:���(m�A����������L����j��H*�Ʀi�T$�$`j<�oŭy�E�!v�j3.#&<���ʗ7�|@��K����]��x/��v�c(����c�����T�R��3�x�t=��<0Կ[��mp O4�_�\5�q�>�z���2��͙�t�Uz�O��my����N�&��J�	���O��_�7��:��z
R^���)��\��=�%t���h���u��ug���83L�lw[d4�i��w3~��8��9�pw�o�6<���]��O�v\{�<��=ä����Kj}��>�?2�?�)�"��Ͼƾ�����������qo]����q���(�����u׻�=�=F�|�"w�;��/:��2>�3(�!����=�rk���Z�c��A��B���)�)L?*�q��T��-׉U�d%!/�SK:!tH%�������c�L;p5Z`�:d��7_��꫗���r<�ؑ1]��:���,RO<���e�I���xo�a<��O���pU�RfQ�����Z�=�@k�<�g��;��@E�s?UU�X�D�Q�!��m'
�6步-���U���Wl~�@�X~�Y�)W[�$�b��L�v���۰������Z0�^s�æ����Pi��jE�滛���Q9f��L������ �*����{���C���R�J*�<H����U��')�s���=,[Y�E�q��S�W/�����|���k�hLWh�V^6`5s������7u������7m:q�G*��2�fBJ_�뺬X�o|�����T�Ƌ����mJװ����[�bs۩Xq�4���qFZӷ�U�����
�i�����j�vZ���T��YX.%�Ts�`�r�������&L�����B�уŤ�	�v�S��<>b��_6�����U��������������/��G�v|�u�����W��",+yB%�Ս؊�@�.Ü6��Jo�5��p�J_�����N�������tf�ҙo�Z�3�v=�IU���!]-�����鯉���U_��9
�M?�o�f���JC�}[fk|�9��si��sO<g�P����	a#-=�e�:{�b���X7�/�goO9U���(#�\�,�c�����1e�$�S�$ho�k��v�4��N��{$8V$�X��ї��qDP��њB C>>st�����S����o��<��%㹷/�7��PTx!�>ߝ�~�Й��,)_���闕�z�t�}�T�U1Ѕ��ϸ�@�X��WlJ"�㕂�j�E�!k��Y��ta��������Q:^�8��xфF� k�BjL�E]��l��G`���!�u���M�TJ��,�`C��s-���a+�Gフn=U9�ʁ�T�����-��"mBu'�B��G�5m�@�\Hog|���z�������>z�z��������O�����iU�`P�v(3՘���z䒼�Yq��T���1�������c�E��Z�7��bcY��r�7�~��/I����쳁Y+���*�c-��Wot*Hɞ���ھ�<@r��iG�ã5Ե]vnʿ�l���&�]kŴ��3N���V^
��,�.�g^RH��KhN�?�[7�ei#��;�)����p����m�q�M�M�݆�F�a��.��t��my4ܶ4q;�݆��
����os�t�:�3/��]k_�9R>"�y�:��G���,ϜG�Z�݄��o|�N���%͆�������-9�^�`��m�s�窠�ӿ����k�pl�g|��VE���s.$��vۿc󗧧g�/ٞAh�!��Z�.b)cg>]GS���q�?Q�l���C�y���׹�����F�k�_���O?|���(Ͽz���؞���K-}a��Q�8
�G�u���l�'���o���j�b]a3I�4��Д m# ���Q�Tt���_a�N�=}�|��%E�]���Cc��X�U(�0
#o�_��@��#~�L*G.�N����s�NM�k��b�Z�p��Zs�^��|	�Ѯ3r��v&����f��*�
�_È�|B�`��$)��x��8����!��qZу�<�5R��ִ��+\�&�X��x-�.V3����e��W����t�Hr%��m$!n)������<;,���<i�F�ǥ�8��*�Z%��0<��Wo޿��3MT�hh<���k�ۘ�����<�ZF%�Q�m&J-1����#�p�Ԁ3���jY��~W�ThH	pep�*��RB�[t-�m�ۃ[�B�J�V*)�|�7���k��Ǭ�P���E�2�?n[�T���U9 |���ۮe:��1����S}�&~�$D�˧R�jI'�O�Ձ��q�z���� ݊�iw�KZw�oKo�洙�\�f��ۖ�q�l�%�e���m�iu��6\��HX�atU��mt&��7�v�	.��;�/�:���t�;Ә��v���gܤ�v��n�mxsOt�������mC�SD,z4��%΅�XߥU�K�*`.���qg����7���2���brH kYT��IQ���%ї^_4��	]����e_��H�!�G}�r��`���7����;�c��v�� ��^+����W�;��&{.%�'�F$҄�%�����a~R���DA���&O�I�t�ڮǌ�8!~��&fU3S^���#>�S�!G�sU!*ߑA�+��LU	L�k�AF؀���%}-�&Pٱ�����pE������3jN�FqK�
k�Kps%}-��5���kAg;�&G��4n5�:	��+5�6��E�(lh��*K���` �?�-�DZu�Le�t}'��O=��C:�E��ވx�QV����j1{��I�s�[Bͬ*`�i&<��-���K�F���}þL��~ ���0w(p6pc�J��-�Q�]����xRt�-"��+,A�B�\�Y�� eQ��ĩȪ ��&o��*��T��A!$y.��Q!�g9�s�pQ��IЎS���j'��uMގ�,���̃��"Z�(�}�Uu�y�f7���	|܄�to�;�g���2�&:3�O�[��~Ӯ>�&?�7��x˲�|3�n��[���i�v�Jo8ݙ�9^�tִ�9Zě�#���LcM;U�i��FO.OF��/֯y�R�ǒ��i�[Q������ʚ֨�$�wr�����u��u��?�$n�]����y�<�Q��ʊ;#O���e���������iO�U��z�мТ^��HS>ֲE��y�I�r��FD7I8���&nUQŕ�R_A@�j��j�!Xm��B����"�cd�%���^�0��:O#w�K��7���� K����.H���p�$��ԝ� @����5:�Z�MʁR�=��0��[���u�/�M�u����ɒ���*�o`i�&=�@M�i�
�!x40�X�Д�]�� �@r��7ٍ��
��� ��}]��R͉Z�"\ߒ̛
�
��)�����~����i��� ?�z ��P�·�%�_g*�#���m�L��oh��z�
Ȧ^ء4(��MM@�8�.-y6\n��9P�7NI�:���ׄ���zI��חE(���9�����O: ('�[�X�RyN-ad�Н����W�xI��k�D+�%�2\r���5p_�F��g�����-�L[�5�g܎���Dc	{�mi3�O�k�xs^���kwN��NkW���N�0o����5����p<�� ���#�G�7GPn���Y���tc��#����Xe�����E~'����<
ʃG$��E��ٙ����x�Z.��c�s�D�]�;�0^L�+��1O��t�Y菝>T��c�1���)�{Xg\�OF��#�5�,��|�n��?�p��Hz;@R%��+��N�(0	3�����PC��Tj�M��gL�-�����O�d���D��Mb��פg`3�pl�FB�����C��!��YB��T���R�I;�W�ռ�W�6�����p����6m�^lob���a�PU�xu�O+��
$�WV�h\Q�(H&��g#V��i}�O
�@hT�`�	�:T��MaI���Ĥ�\}�_v�Y2a�G��`x�ˊ3���<�ᕩ8�[s��2�$-�FkTU�(I�˟���˭T�WE���m8s�Jl�	5.�E���1�U7�ip�*%�^��o]��u�Rv��E˩E�~Ҫ���7���c�"k귺�R�%�(i�5���#cAl�"]���W��8�0�t��0rW�-����������|n�6��J�inß����83~�iRic�W�?��9��d<���l�׸%�g�����|.y�ex�O�٬��{�f���3�
�Z���E�핅����Ur������	�9��dL�Ū���������0zzҾ�ьvg���x�yS���`�`DduO��<���`f0\� ���w�7Y;����f����+3L<f)�)�Sfr�Iꮊ0nqt�F�Wm܇��+˔�%��ӟ������p��{>:}ʆ�s�H&��?�;[s�Y;#/������f��lG���ӕ��z	l��C3qZK%M���Vz�rKh�#,ĐuI����d?\�ſt�[�.�Z,��Q
,��C���)x�K0������ Ce,�������)Dq&��oyk$�)�z�-G�k�+L��0�+c��;�y)��Ŋt]k��bu|g^��֙"IJ��j��Q@���<HgL����zX@.;Q ՙs�}�Q1v_*k��讑��\>O���s����1�c,=��6#/TN|-3Z>��Lª*r�/���J^#�RQ'������.��-��(���;��S�:�Ȋn:��=�2"��E"YG��2# XN5�gXx��*�x�*����kɪQ��ѻ�
� G�I/�-ݴR�Zө�_�wLZ�/d�M4��.�Mz����x튧��;]�;�-��6q��w�;��D�ӷ{[�M~����M�o�c3�M�7����N�7��7�M��&����9l�ͳi���ܙ�17�	�z��4���x��E����ݗw;���Θ��3"�[�5�\~�ЏW�ν�a�[�J���l�5,`��6���AVF���=�����F���}��I�N�0g�"�j�$i����S҉�`�Br	$`>��zP9^0��X������N�(�B-���Q�D���o������q��د�`e��u�݅g��0f�P��@0���^�&n�����R� ��q'�����'T��Rl�nO!�3E]�����m�5|��
�i��Ke.:U0*ށ�����C�glЅM*Aa,��O�5�����黢[�52�A�e�͚l���SS��'������6��"5i�B�bY�M#�D�e�.���-����2���?ĊS�:Ҵ^KD7H��q�MH��4�U�����ꒋ�\���L��ECUc*K���&�j��J[s;z�����␵�GO�d6-*K�� ��_���:��1D�艔C!�}���V�
ik|ˡ�^��@���~��%�:��.������_��Q��H���s��-��s�ޖ&z�"v�����T�=I��&�[�5��a���[�=���[m�I��3���þ�|�����:�a΀�g��� �/��L�����齫��ۯ]��=v�O�gL1�=xt���̶���Ov���s�8�Mgǜ9���OE��v"_qW��k�iA�O�Pɢ;�򊺆΄��$ޟ@կ7F��<�g	2�ҏ���RWM�BN��X4v�)'��o���[S�T�(��&�t��&w�u�x��!F���d��O���Yڦ�}�`ͳe�O�縂���6�H�$jIG�&�(j���)r6)�e�s�a����3����0�^(�� <�/F�[i�nc���� Ĉ����c$���Ҙg�P]�`}�'G�'�=���U�lě�(���Ě�Ȁ�}��_��&e��uQ�J��^����$�!�嚾��H�ȣt\B��Yϵ���b�i�1ˈ�Lҡ(��u}�W�'{�	'0R�߼ִ6c���0َqj���!d$?k���CW�W��m�f�j�uhs{�4�����6
��8�)�6Z3l�3�o�7�팧��Rc6��ܛ�����\W:�x�47q��7Ý����6���$��bi��uw���H������=p��r'�	��T{�y�Y.�'YglR34"�˜��@�U�ѿ���
��XuWZ�;)���Ғ��˛z����x�p?狹�x��v�2�g�I�d*�2"�[�d�����D�r)��������KL�TT`�S<%�v�f�w,w�q�4%1�Y|�����E�~toC
 �;6M;oҙ�R7\�����1`�m"�V�?dR���L��̼@�x���d����1C�݅͡S&�'`d���m���Ţ���A`%Nm0��-S�f]MK�̔:⥸!m$��$'�x6~6o�.���H��/�{E4�+��Y�,����w�#0.Ȥ4~HW�F�f
��8�o���g�P��&Χ�j4q/z��tE�O��J%
��<*�eD����{gTvR���}r���+
��锈������s�Ζ���֏p��K州(��{�cgH#�)"#�� `�kd���u%�|�N�|uk�=�#��z�>��k�-�MkӝQy�;�QB�yن/�����:/Mw�ݖ~����ߖ�����-�����8��ތ���W�~0�e����6j܌���>ڂwn�ҕ��KE ��G�⌋{P�[�!_7rٮ�g��r��Y0)�-��i�Y���M�65S��Dv6>e�ᣅo�RF��;��'�ߌ�|V�C�3����r�9��9{�N0�N0�NϘA�\7�y������͐0��W2R�$��F�B�0&��4tթ�Ò��11�M�yf�8p����ԧ��sv��\^��r�O&�1�k�(ςt����୙1u�o*9�Lm"����P�`ƮN�� ��45�.�3y�y�B>\��/�������pcW�3��wq�9	5�r��V�
[ީa�ݙ� t��*�tC.�kn����Xo)�N	Vm\��*�N1�дM�b�5���!� �D;*�^z�`���n%�{�Oj�ʮ$mi#�P��e/��JjP�o앢�*�ǙZδ2Gs8�|�)FZA,>�V=zΎ3hf�^���t#D�*��	#?wc���%��R��v���1#%�ѕ筈f`���/uo��:�����LK:McFlX����f���[ަs]��#Μ�4�Ż�Ƶq���Jp-��l}���f>f<)t��յ��N��r7�ux��w��tL�<�N�V5���.e��f{/B7���%�H���0b<����z�E�I:�jDh�d�4�� ��~�r$2��V^$��h:��'];L�I�⾤D�!�!H'�|ϑe����L�Ȝ��e����|�q����+�/�埸�H\rU$ѥ���G�v���BS�1��I���>3{������D}��۱B�e��r�̃��tQV^b��8��B�_���xGV@��ʐ���.Ks�'�*�s�<V��=�s�(`"	H�F�兓%+@�]����R~�E�
.�.h�H�D���Wh�w�T�o�S�D�o�&,S���Z~ڠr�I抄r���n��#z�1v�ia �a��5ӛ�M��*�''|�����t�Xu Fz�Zm�ȎVq���G��Ft�IR����ȸ�h�*^���h�f5�Q񷼸d���I�v�݁�*'�^�4i�9Q/y�<K���s��XFO㌲$�t����v:N��ʯ���k#E���n��۝D�����Δ���d��WwL���|����T���FS�W�s�m�s�m�s����h8������k�����t�\������/�Y5�j+W�NL�7O��&]m�*�T�6��Y�S�j�D���{����9�ڻ�b�P�+ë���/�4.jϫFY��Մ��:�����3Vgi����߆dN����E=-�D#C����ë������R�N�O�q�-�X�3����if��b,�
b��"�<�D����Ȧ����)y�`2��:�D`�{iH�a	c�H?2^ƭ���-�N��#�t:�è��.�[凰\)��l���*��]��cN}�_yS�� s�2�;4�dL����NMi�(%�cV�u���3��ֿ`;�N�k�'^+�n2��Ԓΰ�(0}7���Ӄ
_7��әIVn3(|�v�$��Xߕ+��<�2\���߯���}�n���%����E�o���"��#A�M^:�*�$|��,h��A�A�"(H�8�<G�Y���o\� ��7��>����@��d^�c�5���x��V��Ҳ�4���+�xFOW�� ��0�=��]7i�m���:����׼(Ϣ/�����k�k�+iyrg��t��8���7�mK۰�������6�<����n�w����u��Su���>yJ�yKi�o���۽	�/�m��ſ�n�k;�����	�-m-��\����,�[P6i�1��Y�n�ﭫ�}����gpd���t�C�Uт�Gi�p;�o�^ެ�`�X��R�K���8L�����s��
�1ʣ+<P֙�>ƩN(��te���c��	+7�p����a���U�U��5d�p��L�wܔ��0?\���4�|�ZÊq@6��uȋly8� �d!��~_���c^�PGW����,^�Ƴ�5�?�#ce����R���!��ȓ�[���p�y(f�>rGF�^ͥ͢~�LrWX��j��HUҍ����V~���V0��D����	��۷�F�B�G	|�!p��}�C���֫qLWr���)�*Ț�V�Pq:�|��իܧu�lmļ��Ө|��+DS���3T���,�|6�l$,�:I'm׸BR96_]�6֪`��$V��,`�?���yc���Z9=�Ɗ盐<���hD5u����N��Ȉz@yg�Q\۹˗�pr(�oZzk�*�OLvn���ӧ��N���Яt��?�_%O�TGq=~Ǌ�i�n[za3�ƹ��9r܅�_�~Ձ/+{����s.��y�2ݤ���m�w��y�q����`���]y.�6uOy���&�����ޯ��]`U�e?r�2�!�R���[��+)��_�or��~�ۇE���9S>���(3^.�G%��K�G��ر:gt��#o��n�������5�2�@���g<�����Ȅ��o�X����j�6��:!�Zʭ�~�\&E�����)P��D�q�oӡ7�O0���)�� ������<_�~���K_c2�lO9=&�=�Ya����'�$���[��-��-�H��~�F�kH���sΊNM0�5o3�IS������=���A^9F$x�\����mSSsĴ�WS�5��ւ�����(c��Z8fԌGm���aYgҤWyR)�/�k��aHx�	���>��� X��S�N��v]�rz�����%F�3`�V�KhZ�q�4����i�7c\�)��"�1VyAi�lW�
,E"
Wk"D;3&��!PU;IF* �qI�*t�+�u�y����M{�}\n6�` �U����lP~4���_::��<i�'c=S�n�c�JS��Pћ]?�����X����<�gK��;��iZn�]��v�k�wqg^M�.�g\i5��n�;nN����ޕn�&�%������NwS���["��6�� �?'ox�vX��?��R���U���_+�<�^�_(l)����M��)��_i$����}�{�.�d懲������9���iQ���g�U��Q���o���e5�'/ǲz{\e(��qA�X�����͘�$�B?o� %� .e�$Pr��bL��f��kQM"i'Q�SQ*��A.�TԲ���'����G��F�>lUC�c�<��2�`��<��0������8�����M�R�V�JG�'8y"�9r��g�1/����'���vg��l.t�8�!�p0ؔ�/d�AM|v�W��7��Ur������̬aM�]1b��g�T,k�f�B�;4,f�{�.��$F��r���-�1Vb͢X�m���n#�!2j|�6D��q��g#�//^�~y���T�*���r�Eo�j#���4d�.�f�mH�
(��T���Tl��(p�r]&� �>��$��,re�Q�׭TťhT�7I�]~������ �i�)~���C��Ӡ��P�D�tP\�;;�S��	NC������4��I�:fh�ή�'l¾+7��o�4�D���4�n�e @�NWtg�_׿.�5_a7���7��w��r����Gs�N�m|f�����Ό��:��;�_Jki~�N��M�/�-w`�(�Ն����s�e��7)���-7z��w��P���g�r�R��?���9�u��CσdIM#�fH�G^0�8^�{�~��������%�i�tQ�K�Ϸ!}߇��St�'zJeh>"��9�؝f��l�I��7�&m%�ůt�b��XKe^9�� 1�
jx~�_|��ep���t���_� �:]��Y&tA�g���5&|\�O��c�2F$��Ƹ�jv����	ċ�C
��}�>�MN����,v�v�4���kA:���s.-߬0S72uX�B%�R���G����s�_䂨 ����P�.�5�������u��oţ�����Z������@�X�-G�Kha\�v�D
>ɗ�ؒV�
_#��Nc��8j�����_/^�f�&U����>�}��a�]�Ҳ��,�K����r,�.e4V��օ^M���_�ɒ�2%d��D����Y.����ӳ���Z�P�'a�j����A;o��;�؋3��-��WY�����4?�	X#�f��{� ��..�R��䒏��.f�}�'��Te��]�K��M͟��H��.�o�3��.�q�<;�+�6�����Mw�m�w����4:�����v��a)�Mr4���4�ϴf���N��-<Ӻkڦg���n�im�k�-B wN�|u��a��Ϊ��=�:a?c��%=g�t5\7t#_���0rf��Hb����1$\�$*{�2��`�ާ̴�c`� W&��c?3.#,rH>r��*W�\�o�V�J�̨��Ûd��T0�R���� �%ird��!0�7�A&�a���z->�R�Zz�C���I���=ot2�u���Z~�Z�a\3O3���3��:���ć��7=�7��3i�4:��^l�0��s�x�؉S��&(��fT�v�!A�p����YN�dq+�c���S�d��̾��a�TT�)��1^R��p�\09	� +��5/��G���ge��}��Jt@���V�׺9mˌ'o����|�� �$� Q��6e�-*��q-�1JT�5%�7hҴ� 3oidݚ��|�Tcp��sۘ^�x���痫���{]��b?ܭ�/Q���I)��
�_�V'���΁�Q��!d���*=ĸ�Q�fџ�J9/�ڸ�	1d锥�	�oDn�X�i[�$+��C@ Wю�Ұr"D:0h��T�?��t�߷X��#�g�%����S����QxF&��}ò:2;J4s�GƑ�����Ԑ�t7莼W=�܌���7�f��Y��igՋJ�|fXӺ��Es[�m�g�L��;~3N�f\���L�M�ρ5�v��<��װv���ǩx�V�:����ٕ��m�lK���}m�5\��6ώ�.͌3�ox�M�݆�i��8�-�4�5�n��'�vX
B
�����%u���P��ҍ������0o�����P� ߐ<`,���ߧ�7�w���5�G��}@��/�џ���t�{��ط��e���C^a�1���Y�?�ԑk1��t�^%�Q���qW��_�x���FЀ�{��{�r���2�L3�u�>���h��R�i�þ]s�1J�B�7/�'����d��͇ջ�����s�I�Sq� ql�$c'����<�귫���1���Ea�M�1�*9���X�Ii�~���,w����Ty�l��Tn`�_�6�)g�!�k�s�N	9u?���C��`΄�V�����=��(����5eWn%����K�@����Q�B"���N�[s�
��b/�ae.9	��T,��|@�Ae�[X~k���_��L?��L�R#tf?B�]Qn� tz����X�QVo伤!�/I<yXA߽=^�����~��G�Pq0��k�׫��V ��R�a��~ʏ�p���5*u��f���:#��a\�B���$���!����µiz#uhq��e��C9T�a�G/T�>� ��.�z!�ӱvP6Ro~(�.}r,�&���@CL����a�)Q�6��oy5����z6�ST�ո𒶓+�k�������$����I���e>����&����3ә�)�9�o�9�M'�&L�6��Ͻ�^�7�i�v[�:��N��<�zMw��<tۿo�M&a��F���ь�� gjgx��M��p ��-���וOcJ������c�7?���g�2coכɝ���/�~�>��axI�~����E���{E�-��Ւ�2��W��y��X�s2�����d���(��6�׬��,����3���]�U�ß����(�rS��s$�o�A��u�K����b�Ӌ7����]}��U�@�>��1.���ȃ��K^��S̒�3R΄�&�����X����k<F���{"�k�q�w��{�?�L�����:`|�H	 �����
A�@���n�I�l'g���3j��ᅆ���.IC���^y՗$L�D�Cs
�%�c �>��&��՘U���ˈ��Ǹe�}^S���G��8��"'Z�'���QZ���F��'�>;
�JRr�J ����H�2�y������|�&���O�>.��/_�]��?���?��c��'��YLa3�������ʜFh�Hd�itD�p4�7���Q)?�h��bG�i��]�4���-5Aњ=�j�=B+I:D�8����-������B
Di|����	��k^f�>RG�a�2��2Ux7_*�4k:\i�ҭ%��o�ѧH��u�EDm9M D1Ӕ�
W*��<�n��Mz�(�QnM9�
�ː6��2���#�em�.�v�uG�;|�����4M�����A�B���F�]4[�}u�ɒ�6���B�z�J��!��eq�a�W�O�E��0�<ɾ�F��.u�ظ>hz+���ԧ�;�Ξo�1���35�Y2sr���v��|جqC} �i�򔫼��Ցt�,.�������wet~츊�����o :fJ�)��)���|�O�Y}JɁg��|+�đ(�2���t�G�i����y��o�7=��3�q��/VO=b����&�j��O4��>�q/K�C{�ggǫ�~�3���z�������gϾY��K�5��s�0�SG�d
:�AMX8��yo߾^�z�2{�T��4�V�l�H�bKPGS0JYZmGCXt����!@�-�K��C>1u�c��W�$�X���l����-����Ɉ�ğ%@� |A5��/Yj��r���ŝ;��u]�kP�* ��H#F�*˷T�%���OX�l�SQ�L�l6^�^�	������_�L*�
v��,�  @ IDAT1�W)+��R)�pV�w�W?��b��o\������R�`�Ƙ�>I؆U~5�� 9�FdA��4�aU&��`��P8X��:��ΐ�?3�a.iU#��Lm$���F?U�Ɗ��ǅ�?1�F�P�T~�y3���S�t���<�TH#�&}�w=���g=f}�%^嗘��<�������0�Xx���gH[�s�~��3�b�� ��/<T٧<�q�Q�����o�K��)��ބ�.�ץ7n3ݮ�utfYn�7���.~��w�Ig3<�Sw��[���w�g����_�o��p�owNk��w�v�o�v��f\Z�m�{˕�ejs�rnI��vJ�Dj��:�g��a(�[ʗ���of_�c��Z�A�n�������`�G���X��[�*fAx�wLH�e�e�4R�����G\<�K�cO��o�p}�\�l4��y[�����j�Ҙo��|q�g�8c�F�,5_*(��|(0�Py���Qw�G;�T1W>�+\����U���%R������V_�5[Pp.��6�Fg1$���1
���NL�8~8�e��q���[�\�'�<Ն��(yp��%�z���/~2�q�ٯ�w�?�(�7���S�l�y;�L�	˘�"/m��ĉ3���ʘ�a��chj�s�@wY<�nrbk\�R ��lܔ���̳~3�FPJ�Nap]��Q�Lg?nfĆU�է�m�E"5��l�NEV9?�o߯=�j��o~�zx��Լ��^�X�MbdJ�D�Q����e�:+��rg�Ύ}��8rg��'�>�p��~�e��w?�������|��|���n��"=d*�/أH6+Z������hH+�����@O a�Dԭ~,p	Qm)�C��it]�i�*�t<Q����W��|&Z*�<�k�	�@=��O$ё�0��&쟗��F���5}_J����<�z�hu�xx������M���b�{K��(�u�bc��`>��w�V�+���V�>����)�_�$w���VT��t`*�����N;�Xe�L��q3��;��g]�V>���q�t��e4�nX�\�ކ�L{�m���uE�O� ۽�Ct�M��_��I�3�F����o�~�Ʊ<�ѿ�A_J��}��=A�N�~�5������f���0��s�˙g`4�N;Vc�� �����2`�F��y�Y.� �ư(�#	�+kh:F<`���C���-{�~�����ׯ������f������g�V��11�J����%���c�@�$w�"Y���ǡC(�H,'f�D��ٽ�#D=d�8cl}�!���V����Y=}�r"�_X9=y���}�l������ϛW�˿������50l4�0,�0,]vu�����Yj��x�,���{1��0�B&�7w��?�0� +�+�)�G7���h�(g��Ch���o��_ɥHߪt�r�<D�gϿf�)�GY���%T�R��@�Kݖp�bĒ�u��?	f6&y��F,;��>�����C�R"pыԑ���T�p���0Ϊ��x3�`��ϖ�R�:p�t1Ȇ���Oj���OkY�/	��Ɨ�ﴊ3M)��H���_����W���oY��@�B9Gn���b�>K��(Ӎ���P��U^hfTV�X��V�uխ�,�b�j�m:��%�m�:�5Ӌ�s�'����k��?R��Fp�L�H^�1����^�>}���N:at�<���o����������?���T��I�S��S/\���X�Ƙ�륪a�S�J�W�Ώ�G6�D����ul�y���M�Nn峓�^m��n�gZ>�n���]���x�mt���N���ix���M���m�����G�:�3�M�M~�\����n��J�&��o>�6�M��7�m��
wz��7�·����Vc[B;�^����{Me�d�p�#���7@ '���c��y�vV&34ET�kx�ҕ����������w��o��?�g1�:�%��#����=��3�Ȩ�
'2�M�1��C�a�D��zL̙��s�7�0V.N�0B4FN�����z��S�e$d?c,�8��n�w�C�#���Iƞ����84�?/�1��a�i����|s���nkr�n�	3r��f,��$6�%�G��5(�h�,����-e7�מ�6�������×(|����?�Ѓ�܇Е	2c�_e&5����V7N<5i23
���>aS��������v&��`?b��afP�F����ۯ7	�uQ�2����N�������̀Z��k��y;D�:3�e��AЂ�� ���k�NC����z�R�;����o�z�쫼aPF�J򊰥��b����)Lg�S�4���k��l�3����u�_�]��������?�~y�t��>�9���픧��Q�I�cd�s&�ڛM�ŝ�!�b�3�	�t.�4��H\n�dZU{P˜g�?�k��E�-��9(-��'�r���+��� ����K�
��$�1�к;��\����;6H~�ݏ�o�>^���{�䧴�cf���~�R�)|@�s#�T�lL6<+�O��o�S_��/{�ȣ8>y͗z����K.�ʚ��4��T��Ӂe7��JL���"�.9z�����_"��z�u���h��}l+'1�-�ƿق�݄m�T�v�eM<��}��δ8Xr;�9�u���=>�?`v��5k�8�w�z��)����y��p@����������g儇R�h�Oʽ�Ĺ�O�k��t7P
qɹ�ط�z�	YYr��>���-���1+3h���7t��]Z�=��FV���;�?��!F�C�߳��f�'3G�r�WF�6�� A��"����&F<�E�����s	�q�=F߷?��^o�~�L�(����~�#߃t�pK���򐱀�E�7��C��ua�<F���e@',���|j\>x�^0��$���U^:�cVԱ�B-�]��4�E����1��t�v&������C'��{.s~�3}9���p��y�>3s�%�T��l�������v�wzսO~X���[�����=�=�����[0�@:��}d.9�C���\��Md ?>���Tfx���n��@��l�y,����?�~}���u_�L\j�a�f�Ac6���R߳��ǟ_����q��o^��'�K3�.v��I�<�@՚���
�OB�f}͝Kry�u)$��k���1�)h-GͨiӘ�&%���ӎ�Z�$�?OaNI��S�ӰE3y�7LI.�T��AP%R`/�s�Di$�i�
���}�K�"�>a��N�sK��z��ibg�l�p;��Sv�0^:�d=T�
��븒��,��֞�ݍΒ,J�B u�
d��o�E�S�6o�o��K�f�6��<[����m��n����_�:y7y��Su:�m�i���n�.w�Ϯ�+�����4��6����m������� �ǔΫ���˦
�&c��D�/q�b�A��D�g�oeϖ�%�h�	�V�0�q?$��8!Y�S�@���o;^�����~Y��s+��K��x��D��?�� ���Hv�Y>�;��;�����}Ɖ���2�9��8u#���Y�c�<�=0������p�Eʪn
��$ʐhxG5%��D_���c�:��x#LT_�r�Ͻ_ޭ����8��z��)
�e䛄�G�M��:���c�`䃟v��<�� �PK7�ɤ��	G[i30��-�R�[��⒬<'i�[f��L���g0��"��zfeG��p")F�xh��Hp߳2��'*0`?x�x���!�G�p�;]�����+�֜|<S�wC�;�6�����	-�K�*D�h�̡z��BSl��v#�K8��0��������k��������O"�W_}�:6���go�@��¸���\��O��ur�~"���QI'�g�?�b�����'o=����7�c|1}��{�Q��9�1�M�L3�*G6�{�G�����{�@U�)O�Q1p��5�Ϥ�[BVl��^��=z�1!;�c*!�4��D��_/�?2㪊Օ��P�#�r��F:!	�o����O�޼[��Y���_����W������M{�/h ���ﲭg帿B�ڎ1�QwЭ}��F��y�,�|��$�R��R�����G��Q���2|Rv�]��R������~�X73d]���7�nn:�l��ݒԯ&�̯e���g���t�v�0���J�ўB|l������qH}!w�6m�2#�?ni��s)��z?=盍>t:&y��Nm���z̀�ݏ/YV���V/Y5���{�}0�qeB^�[�đ��S򮫴S3<���rђ7���������5��N@H5�F�7l�q��q�+�p�3%}����c�v�@ ���8VdOu�O���U nW���Z?�btL��r����b�?������j�����_�����,<��<E�մ:�K�4l|�7��M���A�=��G���Y�L9��\b"��A4P�Ϭ�����\ї˰�,]�\̟e�MCK��3VF���p8aV�����,Q�z���߬����s
��3/��f�>8c�R���ʑ�YL�)�G���p��ުu�`�>+V�kh)[1}�[H�$Ҽ��%bc�LQ��4��i<����0�@zs?FՃ���"cΤx�K*�P�)x9$<��l�O�U���=_������Xv���O��ę5ᛎ��%4�1��mg��@�	O?��@��`]�j�n�oeڌ}�:먆W�U��c|i�b�3%{�l�)e�)dJ����Fγǜ�L9�s�Ή�e��T�)������ŭ5}�gJ92UG�T:��G���N���=��~z�
��ϩ��3d���K>����=ʞmc���VD,�Q��ǥ*)3�eh�`���\��N�yn�e��B�tֺ+W�df��`s�.��ț�mKwS�-lv���6�������ٽ��w�m�i_�OU��:<����|6iߕ�M��z��7�6e��p�o��Lwƿ���F�dO4�E��;��A����(��sӳUhC� �Ɵ��q����&���C������w���X6;�o5���A؍�n���-�?b�����+�1t��U���z�L��B�B/f��_c͞��U�F�B�F?\�N��8h���t_Ë�cw%��p8�c��ǌc��
��r��Ҧ��n�k�2T��Yv��6���2+z��D�r�욆��x��:~��p��1�m<����WWO�G����vA,�ԙZ�Ւ#�%���l	�-Ȭ�i�9])��t��X���j�L̏q�*����&���#�9y�?��w�\��//0��`���������'�����3���	�R��Cf��؇��/���S�Q$^�'r9X+�y��I�㚋fɞ4V������O�>�y!OY�w�oй������+���?�`j*��}�O[�;\fҥK׿U��?���-
�㟾[����V��߾]���kf�h<��x��%ȣG�V���=������r�?��͝�B���E��g@ix��+�� QPTZ�kŇ<���#�����9��ݻ7�?���}�yȴ���~�����V��=�S�0�ǩu�e#̆��B�솓
4�\Z0�l�yrH��y%�y�?���7L|KE��J~���5�W:������\�)�S����H���[�H8e/�TV��a* LZw�{���<}�3�N��ȝ�T�s~�Z�TG�J	�2]�[u�q��/�!���.�.���f�&Zwŗ^�i�׶�ۦ݅7˲����T�k1n��%׍	�J��/)���{���2)�ξ�G��-
�{�\i�I.>��g���1`���F���p����IѾ=cG%8���q���M�S(�f0|��5+ ?� �g��nY!�G�ԃ���̋�;�ȓ�U�&��<��8�r��N�_���Fo�ǌ�o��|@�9����+P�!�����|�z������A�����b�i�T/(���t�_�s"�=o��	�C� :�wV���.��L�� ��K���~w��ßF���_^���W������Nz8oǘ�����I
�p�U��sΜ�Q�i�ʵ�Wup�u���R��0}�%�vcrI[Ti� �hb��#�JSeLHz��\ܖ�N4�U��A�~��1A�lY�a��[�9�C�\���- �	` }π��blhCy���^���笌Ɨ�}�Q�H�E�p-���a,d2�Va���Z.*&��bGhqo]���[�'��t���f���=pɩ�c�I�j���~� ���l��3i/9>���9��_1�����'��r�=�c|��bZӷ����(�s�eOy�����-��c.R�/F@5+�Ƨl���~��a	��;=�1���M�t�3̎�q&Ʋo��Q�~�����sR�Z��BG���˪Kx�0~��P	Ё�{�ʺK���D�o���O��g�b =d�ѩ��a~��I��mVV�(ӱQ9ŉQG�牆xه7u(o�ꖀ��֝BG��
��W2JZ���p{Z&W7��;�����m���mK3�Ȁ�Jۆ|G����i�}G��n��]>C�Y'�Ϡs[�6�vgV3��7�m�7�L��~�I�nw��M��]���Qw��A�~��傆�p�I��}������?F�٧x9��_��ho�Z�����>����!�7o^��kεz���W�V�xC�e6gͲ������j_��+H� "0z��4~L@��Y�������7�/�����6?�wq�$�ӧ���X�v~�7�����X����I_�K<��U��l�A)n���#M�ˎ���<�+)����ql��[�.x��Ed��
��#�������C��֨,�*�u��qؙ3�7��o�9����=��_0��%Y�J;˲�=�.iȥ����͈�lt��˔�E�������޴Cb]�x�ю�B�<���|/T�m�������:;��Q��8�	��,����:z�x��4�0p`���G&�9�!͜�IV&�m?3i��j��[1�����>#�������?�&��#�$����iR�(SC�iO+��͆�,��L�3S��ʞ�?��[Z�#�5O2,or���}a�` (�����V�N���~�ɣ�C+��kd7�u�BM�&�.��_���D��x��#�y۳ЀN?T�a�a�|��[_=e���r��㯞�K��=
������;�D�1��ֲ�S0&��H�BK��x��'���JOI�@v��|����fߞ����߯�ӳ`I��Ӡ�۬�x�@��!���apUg,܎S�ζ�������x�����m�Jk-SB�m	n���'�Վ���_�p[��Ͳu��)�f��x�M�㮣�8���~��濂�+U�+4�1�`���4�;nB��;�٤9'���ui��-~��ou��Y�j�k��,/D�l��@z������K�f����X���3���"���F�$�_͊i�<~�$oj��xN_�j���lϡ�sx��/��������w���C�=�	������g{x��l6��gr=�]d�/fD��a���w��-E��(�]���@N�)3Y{���|����s���<�G8�Bĭ"~�H�M�ȝ[����$E�LDq�@&���
n?"A($�20����$ą7L��r���V}����_�a���0�|�����<]��맫o��;��QG�i���:������p��pD�0O�����u˓��A&r�0�X��$NeqG_I��Ё�Du�������e��^����^�x#S��+��H���/~�1��z�Y*����tg9��7*|{�a�ң�Ua�>!�*�)q4��Z�L���K�TiĘ7���!S��*(�9�h��֍�~Ux�-3��Y4T1<�K�����`ǼT��T��~��O1������O�X���M�-v�:�?d�/7��i|%�SQoƸ�h�PǸ��>/�`���j�.͘�9iA�Zajj5S��ݔ�%Jt`��Y*�A�Ȣ��
z��aV$�$����0�1R/��8���X3U%W6"O:<�M}���ᘏ�2���w���i���+������ԕ��jLn�XY-rdr�-S�i\UG���2�\�HJ�<�QG?�o�[''O�4���O�����ϸw����Z���dj�N���v���Ɯ�6�>��Z43���I�3�g'l��m��'�[X�����a�����ɯ���	���&�Lg�~����Ѿ��!l#vօ�Ԫw�M-1�HN*����M�߸�OJ<�Mn��w�A�4�|{���n�y��5�`o������Av�r}�����
���3����,���l�]bS&��U��#=`ZV�����1/�L� �yp�n�ۙ�\~���+�/��B�=C&�����]�t,�����#�x����ĭ(~����Y��91�_��	������w�O(�#����w�w��pN�/?��������yS췿y���^��#�Qu��Vw��u)Ɩ�PRxjp�Ѱ�:�5����<�1�����8t�K�K�Ɠ/�Ƀ��g����i	xff�ȶ�
d>�1V)\���%�`{zZ��̌���牮_Z8��T�~�4��ae�Jcf�7sGH�o3�6�75��I���!?|��y[Ҳ�h�]-�]�_�����G*J�:�Y
��oi4?�x��z߮���G��_2}�c�Y,��mp�ˏ�ȉ6�����GN0{�as�2�<u�#��Ve��+��q!��3].AnC;����fkk�_����4
H|��H6�S���:�㧤KuP����U�ɆKq�L�F$���7O��~��*�v4(;[�o���a�6&�cpJ�=�U��^�f���ﾣ�|�z�>5��pVH��}"S��C9�U/r�qX���:�D�)hj��.����37�\�a[Vu��?�������e�m�o�I���R�M�&���mڦ=㷿�\c|�۴6S���߸��t���&�7�M��~��s�m����ƹ�V�Ko 5ݫi�cj�I7��Ժ�&�&��2_�u����&�M�nJ� �W��MO1j��r�6	c�}���ٻ�̅�}�����@�q;�j�{�J�)�Fn�yZ���%��e�f��?n�EuIW�v��I��8�-+:�ȣ�{ -f�ػ��蒟c��U�}�Ri;&�~�g Nɓ�j�ً�������c��� �C	(rk��[�0�X���7��\��9Ap͓��,Q�1e�b� ��H�
��±V?������Rd�h3�3�]�AO��o\]}S_9�D�NT��xk�x)�?"D���PI*E�h'��䛕�c̽�΁���z�����ηi).E֖�1̷�<i��y"=�¨O�����Ͽ�������C�~�2�rG�#'*Nf�I��4����f<�i�W�PP�K$�����ҁ��c�\�Ǚo�Mg�^�Q2ط�a|y^O.4�*?���{⁥n��Рf�1�u�' *�F�Z��C�
˓Ri�h��KfGY�����D	����#��Sz�<G��;9�E���TLs+��c�g��rNE8����#����#Oa�&�b�Y��2��4�F���FI�R6&-����\&��w��I{N�<;f�'��={�^�|�S�W4 d���Q�
\#V��`���m����{��*\_f��kNqv�m	�Ғ�t��oz�'J5����Ȭ��?.KY�z���� �+R��Eh����;�v>M[*�I�dh�kWD��aa^���[g\���?E��>�U^��ȵL�ց%���Y�&_R/hw�,�<\���z��E
���Z�M�*��BE���)p��-��;�`[9�2�,��߄/Ln��p�o1�殤�g|�kƭ�==����9FFˁ~j�j���%��4�O�,����&�y۽���m�~d�������O�{���߉t`�l�$J���ޘ��T�@��^B�2�֏1��޾#����#F���c+(���8�`Y�7�{ظo��!ޱ]̱${�4����rum̀eLP�6��RO��y`�2�E��1�AU��m4]�/�p_`�j�z���זtO�������W�X��}��Oe����k�U�$�4\K��5�.~r��L8X�x�T��sMC���Y�èRkj�Y���Rj<h���uBI=PF��LX�>� �#�D�8e�ќI2xZa���W�G����������,5~�"�����"���!ӊ�b4�|��Y./��:ϣ�+��jp���P��#\�D�b�/��Z��Y���}B���0�z�[{����BYV�Sf��0ZN�3E=dVɩ�l�����,9jѐ��O��4y0���TP�L�&,�!�:_Aτ�>ň��=��c��=v�?��<���x�9bZ�����>���m�ӌ���t�Ȇ�� u���ș�҄��{�n:&DpfO!�d�����a㴡�`6>On�)��]��<��^+OG>v���'�7vt����G���	{���@֗\T�2�A����)��L��S��s]���i�џ�(?�d/����u�"PF�tQJ�v+�t�"p W~�� 5;�����u��ؕGyBm�ךj:K9��-��Kx�N����	g+��'W�3n˱�D����&����箴��JqE��O����?ߥ���Շ�z*�E���T*[�r�Q��8�(@!w�7�+m��4��$~�\���o��+N�_X4&�Hj�U����ߤg��!K��3j�ͫt�E�:/��s�WP�>Pۯ���v������f�y ��钖ˌ~���0�1Z�9��AF3�g����ݣo��/i�d u�4�Wg��C	˓UX���|��t�T��Fo\���%{],��lJ��^�Kpθ?ȏ|���I���Tngx��s�j�5(k��;b�K�T�*#+y�ڲJ�0/�{��㻳>�X�Ng�å!{έ��q�4U��qО�]flq4PE��\��X�����Fx#1x��85�QxEKK�N�B�* ~�d����~����+
D�s��a.C�c���r����H&�ۇLj=a\�goyNU��<D��#��X����]9�
~OE�x���ā������T�e��T�d��,���'ɒY��%̻��_ �rk�9@ꗶƋ��ƠƗֽ���Q7�b�ҝ�M�F�=,�}�ɭ.xū\�@ϒ(E��q-Rv�*�[丅\9�_7��R�^�;PF�z������G��+|]s@!����4�1 �߳��c:�l �r���Q=�(FN,f�8cMڧ��@��d�!�lfoe� ��',�����h�fF:�6�j������X��Y@e�%��O�~�Q::��§Lk�F�On.A���z�p���R4�G�	�^D�*,��WuDZ�3�z�7Ӽs�����a��Sy�w˶6sh<a�v�o���:n��i:���
��&ߎox�:xJ��g�S�4�W�N� L��7����o�Z`-�zg!��#Ek�4�W����Z�w�[�ft�t�l�!7��J
	q�)ma4<AiV�]#	k����'�Hq�[�R��ۯ��"��PM���C�>��7/�m߭Y�p:�>�ܣ���C�5�.0t<~(39�ul`ȉ
�霣�2� �|�R��x�l�5V�Kåt�x�8)Ғ*ᜩ�����S����@��#�}Jɘ��9����������yl��M��Ն2F��
�b�)��?�\����ffY��O}�F����c�q�9w�!���d=䭺"e�ԍq����B����
�ǀ�Y���&�%��즙.���UFO-t8F�D���_xj$[*�cl#����Ĝ�7~���Þ/z;C�Um �����f��a7�ɛ�TD)�ڵ��M��agXj�@"5U��zG�C��$���d�B.�TF�RZA��:@f(r҇��)�ٸ�m�]M��"��H�.�F�O�5$�@N	�8]rD)N�ė�{�q�>,���f���@�B� "x ��V����Ӛ�(�C��z̷5����(�Y��O�#����O'��p&Z̓�{��44�J�j$i��1�!�[(>��|��CNV\x�z��I�Pz2s�����G�A��2af��BLA0��@}�l��������_���Ȫ����>8���9b�x����S�eC�:�ȿ�z����_�}X�ζ����v����L3��ovx��\�5hlҟ�츆���ۺ�y5�-�����x���4j�]�+H7����t���D<�qWZM����o�����m(=�m�p:m5�9�u�4F�ե��u�n�U��~L����7�}�q��x���$��4,�p�Ρ��v�1q��]�l}ĵ?��(ݞK���_d��*�JP �C��X�<b:���уf����l�bV��8�Ĥ�}Ɔ�O�V����	����k�:�9S?����>�]o�;��'o�3v8C%����F\%�_Ǻ�W_m9�/����O���Ή,��-F�-Y�3Ͻbl�]U��2�|�O�����ҪP�X�h�n��V��J�^é���Qs)h~�W���Ӗ�o�S�o�ܣ�x�G�Ig����'�8V���R���!�uc_�C;��93C�D�2�A���@*�go��:nβ�`�1���A61\��<���L�g�̀��,a�@��ϗI욆�%�&��CcRc�x9ӥ���	G)~&��]ju���aqa�Ti�/țv�ˌ��{��Yt�\H�K*�_ޠ�U_9'K�<G���g�ԕ=u/:�-�g @꿩ۥÑI��>���8��VO#6j�y%-�ԭD���k�#S�72�J�h|���F}r��Ͽ~�z��*+2�!��/a�ͧB��a���_��1{�/۴����V�
��p:O3�]ɢ��&4�܆dxSw?���o-�4��hw�$;^��=�Py�qۿɯ���۸��v��eޅ3��<�p�׮�Y�]�Nk����?�'��0l	\eO��/����*���J�o�ĕ�L�n^Í6Ti|��K��T�3��������l�&Y�`/�
��"]�N��W]e�{xI�P(?��C)�{�4fz�3�S8��r�hl�Ѐ��t����3&^�~�}ǃ%�e�p�LGǌ�s�U$��a�T�3�h�6�՞7��5b�bn�'��)�Y�ꯤ<� {�Q�9`�����I?w���S�'{�9fy9 �/�7�g^E�G&%$O��(R8.8�fS:�p�p拇����烼��T�Yvd֣���*�������~�����o�@�-�Q�^�IU9#y*�昴&&β��O��|�-ѩ�v)��\��ŵC<��ذ��b&��I+�����f�|%�O� �8�zUb|0�#������*<���IQl�Q;�m��{�(K![�b�X��X�g%'C{Ս�LEP�E�*���
נ�p���?
�ؒ����T@-q�	�N@�����1]��(o�Hٔ�J�[�	p�Z��H�؄�y��-e�#�2��z�1�.#�,��ېY�G����+p�m�2&��U�K,pБ{P{Ǹ}��#���<[�'	;e��$��]6��`��B!��=sl�- �"�%�\�|Eq�a�OW���߬���忰om��߳��|{��:��[�1��m���E���ITA�#��n�W򛟰��t��7%6�8�7���Ɨ�����_ח���f\s_q���_:�F���;܀��窬�I��v�����ߕ�62�6g ꆐm���Z�C�W���L�_T>�M�/�
`���)�@�o0��t�/��l��~�\�m���-��[mn�¸�o؂���!���AƠr����m?��~��ҽ���Нx�y��?���C��|�eg��x{�����g�)y�g;wdt=�Y3�N�n*a�2�1Ҩvm��t����A���г���?bqb�����c~��}�.�BXa���S���R
nM0d�*H�E��I]��Ӂ*�8�͎�\�,�U�#�G���[���:7�;F��]C��j/l�ޗ�u����#Wʜ�*ST��k
.:
�<u	��g�+�'��?�M�6]��Kk�s��XKO8Ɨ��;c���XM��I��0�0��� ;�v#�)X�(����|�7*X�4]��Qo�2P>x.��,��aФ��ޞ�V�]����d �J�(z�������l�&��'ЊՀ2^Yn�������C�9G�+9\�U�N�FC�7\>e�,Ђ���#s�I��@H	3����<iА����9�dn�a��kaۈ�G�FX�ܺ}k�A>ƗYM��F��Ty����a+^8QS�l�'�x8o|8u�ۿ�����{:^�~�G�KC�'T����u%/x�.~�G��Xί�+߾״K/���e��toN��ӵ���k�Ǿ�Y�u��g:k�¼�t�&5?E�*n�ʹ�⧿��]����R*H��K�7ݻʵ.���Kq4A]�O+r�y	�HnM�P��Zc��ߪ��pb��W�.���M!�Z�v�隝N�+�P����"�$�5�STr�&��Ce���Kt�3�R�<���w����ܖ�>�� |��c�!��ru��F�3J������������VzUyC��7�x뒲w��ƒ�iJ����"ٳ�;d���g������4�O�{�^a����B���Z_�K�o�=g�|�
�I���S�J=�.��*�� �"����6�N����e��zB��
~�wq�T���m���=���ҩ�p�B�)���T��,��JmA�����?б�3��,N@����#>�L?{��c {X�~�2����ۀZ�g�Xм-x����f���S`�bX��=����X��W2�c��B����,zETH�S�� +( |�wW��C�����'�TX�p��ۊm��y��쬗�Ɨ�3o��(C!��B�J]�/�� �/W*Sy�C���ڿ�Ul�sw[�i�"	";^g�
_�,�2�ke�,�aV���_�Ȣ����<�����!����#qsj(+��B�N����%�z}ySF��8��p9;rf�`��S��={_�S�X����Y-�g�?���Oq�#�Ur���G��r���nA7{~s�z����V��a��2Tm^�S���s��1��v������M���m��
��y]�m2^�]���r��Ls����:Ӻ��pgZ�\��:�l��	��6Z��C�%Ө/i�����S�nݜ�p�����vB�l�m�;��;����H�._�J�%����>}�̥��#�B�i�l�S�����㍷U(�H������O�!�@E����T�9�'�����A��Xg䞲�������u����wƉ}V���� �##?G���cޖGnި�KhLx��Z�����l�rt�2+�"��Vς�ґo�2�jt�"�>��E��?�)ˠ*�+� �c9DB�]"'�5*>u�H*��U%	'�|��P��ː�J�����w��r.�h{�1iͧV=�	�Ӕ��<t���o���d0_,��ݵ�k���u*4S��v��/(x_�ͭ������Y{��#�[!�� ixE	d�Uc����Q!��E�B��t�Y@�>��RpI3(���yk��Y.���6T*���g��-���U<��-M�#-i
��4U�J*eڠa�Ium����J]�w�OM,�b��A�Dg�2��W~y�+�Ɯ�piV$K�>�AU�P���y�!k��I8т�K�:O��&b4�����#>�O\��F�'��ͮ�xSTO�������2� �
��j!
�Y�;I�/uz�a7d��S2��o���CP�o���m����3k��J���Ob�f��%nU�x������o����tQ�M	;���f���W���voC�:�]rv��g��:�u���ܙ�:��o��k۲�kL�;��@`a�7�l	�����ę��a�C��It�����m^���#���̑}�oc���!��9X�~�P�a����9��[+���)�]p�	��~8�*}d��_>x���r�/&=ee�G��	���b��JU~A�c�Hz���4`L2��r^h�1ά�(��K����|Ԙ��]v<d�1U�����[C��������iR�D  @ IDAT1j�%�/�e���5D���O��Oڊ4�o��㌭���q{�-�
����rL�+�����pm ��#_۵p���z4����}�c챘D�.X�T4�0ϰ�dɎ2:��b��>3bΎ��ռ5��%�B�T9�Qt&I�(��*L �gTT3��@�C7 �
m�&�����x�{�+ˠ^�IP��
RiCq�ͺ�/�Ũٸ����R�l!��սS��MO�BS�ʔ�j,@`��L^F�՟i�܄HNQ�Q�F��}��AC�W�1��ܕFV�F��nt"]j���������d[��Q��e��cģ�L������i������Nx�<滕��9{�r�����̻K>Z��s�7�K��g�n҅O��m���H}%r[�����ի��N����)���&9;ޤ�67�����w��rlW2s���_ͫ�,�Ͻ6�ޤk~;��6�f��\y�5����8ו��Rxǵ�6û��%\y6o���f���mmꖬ���9Y�W)@}m���'�	�.R�ikC˭*>@��V?L�A�#ު��":'zNư� ��`�eT�)�Q���u�L< �����|�O��"'�c���#�����3[Ύ�f�j���ٟ��d������=���L�h4��=�vbgpTQd��ȭ����ai���]1q�K�|��?�
Ӄ:.��D������1�ˏ�\C�ѵD�1�Kz#����4�<�mؒ�ud�b$&M�3z�(t��X�-S�Yv�������u��U�2Ts�FM$��Ơ��ʓ��c�{����3��W�����uwiL$p��>%\)Z�ΎY�%�P^����O[�/\3�Q� ]!�
R;������SL�tq#�J9Tʪ_���ZL�|Q3�T��O�%@�*��M�A)l��p�/�¼˸*Y!���F	��o�a8z\C/=f�e�1,�z�B���d;=t�0��:F2�/On��Rn�pEFX�N3�ױ�9	t?jk���6�t-���kz:o7��h�<�q����cđNͭK�d�E�H�б����ϗ���
��X�(��~g��4f>)�PY��$�r(m�^I}m`�14-��&���U�6��&�U�w	uym������x%jZ-�a�m�7�6w�&lN�<w��*iw�������ێ79^o����w��t��B)�j�?�WP��I Ɛ7������_��g��f�tP����7N��w&��+��i�Ϲ` �����K����!p�����ޤ�O4.��%��eU:�ٷ��B�K��}Y~d[���g�<i�V��E|8��
�$9�Hj�o�`�w,Ѽ�������n��4�x.�p2/�oꎕW\p��<��rM&��J����l2�z�d҈�McZ�k�+u ��x�B�k��.��p�d�a�Z�%5�#_�&D��N�{��.g��g�6\��bV*���B�|ο\:���Y%1���'�=D"4dJ����i�~t���V1���p]kƣoCM�Fb8@�a%/h��7?$p��k��E(oˍk�"f^,� �Tq.āo�ʙы�2�ruJEo`���Լ��"����7�:4(�Dξ/�!G�8��a������W��TZ���p�D��$�O:��4X���W�����.8|�#$>|��G��xNǥ!u�&>mV�3ʱ�f�"���:�g�B>�*�(	 �9��m���Ʃۿ���7��){����n�x]|����E�6iM�E�:���7iu�u�g�/�l&�?��앆��V���DfY�g�����涸m���I�ƢHc�J�4�	�	�i!&����D�NN �#��g��� ���ޚ_��������N�C�8ߣ<�T��>to��P���������lR:M�M!>h�W䓡��t�-}2�� �\����#�Dאcȹ��ՇwoW�|S�!�H���}Ȳ�����V�������+{�����g��fwO�8i�#�oD:�U�����Kȝ�5���h�8G��Qhr�c	n&WF��[4���V��;�wJ�o�w_嗳���j�PA+~Ď�7���6SD/�|V(�7��7���̹�\��r��@GELy�� �������3���a|a�G���T��?{�V��dZ7��̺ ��;�1�~�^S-k�o@y����I�$��"�e&�	��m4���2c�d���&0��ʰ�B._W���]�5V�������x�k��q�x�l,�
���G�K|B��2IE��82�U.�ֲ�k�xĄFW^>ѩk/u[���o��(ס��|����Jӕ�6O� �ҽ2�7�H	�i1�sY����6�NCꤓvdF�ڈOx�Y�<��ͰJ��čdݒ�ZWׁ]�Z��_�QSy�/�+r�w���w�����XJ3��i'(N��[�DBC�T6�6�x�i	iz���_�uS�O�x��s��_��%�]�e)]��O�Z���Q�,���:W�V��4o[܌w���XWӛ���v�z�Q�.��(�9w��Z����Յ��[��_��˒Is�rg�U����9:g�����?�nuumd��d��y��#�\��_����f���;��C�4m�������1��'W����Y�|�[6�sSBڽ��o��9ﺅ'en�>�m�e[m�O�C�'�m���a;m{���
��޹�ը��n]<�>��I�}��������y�7�"֯�K����]c,����Rv��Q`xdC��'צID�Co��6�T���$�	���d Gܵ��vˮo]�V�pP\��׋}W�;r�F� �����A~P�����iN??��+�hួ�+F��
����I��(tÃ;_��(%�#�x�m�s���2i1�ێ~?IgZ����P�����Y::�}��&���kB�A:��r�t�����bRͪ)�,OJ�唁�._-�Q�XB��Ck��7m�A1��2�)�u�RM7�.��?���$��J�AN9�Pˡ���^%�_�Q6et�B��i@�%N��X�sXo��)��,}3�4����{f�iBo���є��t�q�[��i���&L�/l�U�5X�u�\���,W�r��=�}��H���C�\s'�W�=b��ay�皰��>���e�3��W�&��1Ѵ]��\Kl+��#��l$����c���9���l�G��u�Y!�-�#	n����b�d/�,��p�"v�������%h�^~P,���Ĺ?�_���8����y��=�n'Q��s�S\�.��K�	D�ӏQ���?���Wm�mW^<i���8��睆s��+�^2���9��p)�NP[َ#i�s�<���?�����|>9t�Xy��U{���}�,�k�-A�+oi��瓧��_/�f�v>u�}� _���ۼ��l�Ok˵W2�Y(#��8�$(�{ε���ß.A��B�+q�L`A�S���.���@5��s9��̜��r8�s2��a�WR`&aÖ7p��ɴ~7�����)\�A��b�>�\�vU�Tq�'Ek\�W!��Qy�m`�Cq�F���O;�����!��N�؝��+|�e`�����*N�<�j�`�b�Ze���2��SU��yA��G���`n��K���8~ D�6�}?��p�<�H��w�X��X�N\lN1�a�#��h��S������GS�9��465��Lv��+4�J��̐��*<�=�/�"x�����}c�c���H�辛B3]�U��Q\�X�u�2c2��tH3�4|ut�ʺ�\o󳄲o�y+�R���F"��}\[7��UvN|�]��������Cx�&Ǒ�#����kt(��i\'����lm�	g�>������[.�o+ߙ~~(ˍ�7�W�w������o�Ү�E0;Kϛ��=��w)��F�F>Ǒ�No�;��:�p�T���M��;}ɿm/�m��f&��H�,+����ú�+m���ڰi+ɻ9��ӗ%b"��9�:oRb�l'��[.�L��	�U�ߎ���_��1��2��$˒��7i۽z�:Z�?3�M;:���^�m�au!D�c�ğ�@�^��V��ke�4�-йYY��!�]���<C����}��Q�'WϹl�8��ĀAo����IU/:A޲z��xWBq���L�����΄��&���12Y�.�\ք7�=o�L����	c��(�g��ͬ�G��[�"�PF�\+4�k:Z�7�x�'�$W,0M8N�y�o�CPC;��
���/���axdB��P���"�g|�S�Q�h|[q��ı��E+�'?$3K��s����워~�|u�k9Qf�ЭC���7f
=K���4$���6_����Y��#�����fɹ���v+S�$6'��c�����J�񊮕�E$Ϟ{�֓��/8��ɒ����í2�$�y�����:�zF¿&�h�T������kq��v�>��O��6\3~v�>�K�?��A~����`��U���M�\����M��e���y`�;V(��#����*������\��1����Nwڍcyq�gk�O�V����⅓ч��l��=�0��I�~�O�hOU�θ��b�eh�6r-�R��i3}���H�*cu��(Q�i��^�/�f��F,���d�8�ꔆ�2�C�(Ӗ�-B�LN�+X����ͼ��y���/�K�����$e�3�����W�}����H!��EHNC�v�M�ƃq��}�L��y�w�����Ȭ�/�C�M��J/�C��3l�dTq��)�Ц�������:�L&]B�)�;��u����S'�������J����t��Q@�4�ߵ�3,p.�(��&�<�
vJ���#�)?�i����u�"�λb�䘣��(�ؠ�B�3
Y�{�ר�s��S�����M��Ph�s�&*��GPq�tQ�CQ�%�(�b�ƀ�7��K�,��8_o�����Զ�<�/��}�e��aHo�bT�{l�O�DV��.�m\�,))�X��*��9���um!���ș�s�k1,��H�)w�.��\IG��
���8w��9���Y����N�����R���[g�ü2�0��y	���ؑ4OY�:`#{�I�d(��t&N�ù��4��/w4w�c���N������W8ʭ���.^6^����`�0�ʆ%�w��x���r�߸��uitۺ���.���an�&��ؼ\�K���W~B��4�?`/s5�p��פ���!�͏������)r'�8��uIۖ�H�p��c�
{��#�ծ��p���	�:si�,�)��^�r'��Eo����G|���i=��mI�Y��Z����m~g��✖�]k^QP,��϶��x��$��$'V�LIBg�z�ov�܆�t�i�40-l��0e.ٖ�m;�!XM�8��8)U/�l��L�6>��?i�2�~e���L���:zJ����,.����{���&YlIj��/:'��Y�]޲.	A���+�%˪����?���Zʑ�R-�a/BgkbEK��$�:�Mܰ0�����M�9����7B'���Iᗲ_'Zg��~~
)�����}(�6�DP�ebq�\W>�sΜ<�&�u�e�Dϛ8Oo�G�m��|��Mitio���0��)��l�\�<o|�X�Q��R�RTz�cu�ɹ���}ʒ<�H�	|j��.��Z�X�:7z3�����F쫏2������' �NeS�M=@O�ʯ�����Ք\ٕq�0�ǿ�AvZ#=W�a�@�m��~��D­H�9��ێ=��[��i�,?���Ç����kfB��!��9�c�Ap.��Z��_�v?�Ȳ�m8�G�WÆ9��x}�?�Vv����}�g����S�w��?o^�9�t�K?º�y���v�6�;<�J�Mw:�U�<�9�o�k^�8Or�c��4`�#�ƻy8�7?��T�����uv[�`k?s���k��l:��g ���γ�	��؋�&�Mf��]݃�/V]��+?���&�~�����7%Sߦ���݉��M�I����_���]���Q�,}�.��ŘO����R9;�E�����"J����I�l�sS&��i��a�2�M�\M�-?���N�,�J�c���'1���='�͔#[t���.�v��d��r�lܐOi�Y�h�l�4ke��������O>�sxazQ�)SW#��lr���\<a�Ld�Xz�+���jz/��0=&�X���.G��xyrc��	������F�'!H�DGq��#��ܽ.(ᝢ�x��%���}-�t]��%��jy���\�v)�x9��dVs\�\�|�w`ϕȊ�� !����4b�scٰ3_��XGl�^�?Nt��,�u�}�|��ӫV�g���4&�~(�k����	-HӤ��R|�����x��ۉ�(�c�ǹ��]4��(�8j'������u�:�DB��!��#�g�UXr�d��v����wxU�����}�?��9+�*��b��%8ALT�c95�#x�!;�>�����gS<:���f�sw�:\r�e�!m_�MU�0nʸ��}70sw]ن��e�\>����\�<?H�#6��g����ϫq;�γ��pt�SR_��ӗ3Gz�ҽl���$�	�G~��M�q��4��!S���a]7P-;X
g[w�vn��S�i�}>�����ݕ�]�ߜ�[��)���aџv��0�D4��RWF�z�(t��ȫ�uI�&у��o��<�ȄSگ�"B�ʠ��Ɲ����;����qw]�'~���mIK��̭�궖�u���fnz�o���x�kv2����]͆�8^��Ioy��cG��'��2�f.a��5:)J�p?� =�;����<��`~Ź������޵�ɔa�PD*E`��:�TF���r�����Ջ!��
~Xcx6^wCY��C�j ���̤��o-W>$��({_�S�TK�w�"�p[ `���v�)OR`��$Rs�/�w���O>
��A2�\on�i)5s�N~e\�ٌ�O	�	5���0\B�9�̙?���j�`9_�q�������:��������s�QfDl�ǣ�ѥF�Y�{�n�Ƽ�Q�k(i��f��ৱƫ�E_����+���c�x��;t����]|��W_�5�=��ؒ�J�!s�#P�e���7yjӵ'6�6O��[Y�P�R���vY��↿=�#�2_^VzI�`ܼ#T����+�{y9M`t�:���n�~�.��LB[g�׿�5����ѹ�dM�p�'{ �Y���.��s#�s*g��i��'G�v����;���Ҏq��c������M���`�-y�4��>Cq�|�8����CfT�=?��n�ɬ]��#���-N�@_��OI�V�&��g��ݣ���7>���	��S�x�v\m3��;����:=_]�v��`:%^C����/���S��[G�gv]�tc=q=��P�WdB6u��l�F���H������_���>�Z��Y�'����ԏ������H�T|I�^�Y���͡=����T��>�J�\\�s��&���	)su�4z�CbN2t[���W�#2{�"��ӑ.�J�������'?�sd
�����y��AR\�'�S|�3��ɕ�]#�ε��	�5�AФċ��?�X3����������P�u�v��}8��m�6�G L���u��}~Z��ˍ����e��o2 ��ΎW���H[�-z�b&�8�� ����^���ރ���/�%��1��͹�*�(;9�s����φ?����5#�����"=G�&��o���k}����׫4�Η�x&E�1�~�{T��2����c�ѓ�/�������Z�Paa	:�e�4�ŕsK�mhS��9�7cn����[g�@y���>�]�S�w���e^ǮӺ#C�*�i�8с\��v����c��¶�U�.���S��+Y�s�o��#��y�6YV@o�T�W�ɏ�e&�ɓ'�7�Γl9cxT���<\k$w��E���3����l�X��Ύc��yΫ�#/�m\"�ח�Vڦ�>���]�7���w���ߕ���g�]�F�;l^�,t��[�2�ԃ3(�Z�������ygS����̱�����L~4_v�a���+�pˣ�[�����2�͆� ��|�?:�c�i�
���*�.��ֽ\����B���� +�gz���"�U�ݖ��>�w�rh����Vgm�?i��n�(�8}���.98G��Ik�Ń�趲[��"���e����;����4�&^?��ɳ�<0���:�9�`���9=)��t�a*e�p�_���:a}�}&e���w�C��8G����1����;���rTx�E��Ch�0�r�܉-��f_�7��f٘'~�2ҺE(e����Xkѕ=��+M�9a�E]����}SC�4�Ix��o�@�*&���P�03�Sη���B9�h"�a+CJsɽ�S�t�D~1^)�>�4��a����Da���]��=�ԐXa_,��
&L�w�v�!]�B�+mh��D+W�T�7it9N��bϗ�|;@֞Ub3`f�|��̑�O6���<��O����q��w*W4�ʥ���ֽ��}�z�Ru�4D9аLȨ�d(�.yC����3p*G��t4�;��F�ƃ�X_����⼟��(��<�Kd}I�����!d=���!TN�u$'�P��s���Y��E��B�nG�������_��)~ݎ�y������s��>�4��q�+3'dE���2s�\�/�k�:�P�~6o[ߛ?��YIj���gq�����c8޻F�w�=^oؖȏ�����	pHذ�����<գՀHW����!}�L�5��Mf��.࡛��dG̾�?gFS~��>/�8gz}�1�[��/�{�����,Og�C��h��.܉�1���~'MO����|'�2nY���^���I�*�)�M_֥�1�u���2��˔�6ѵ��SlU���;���h���e��>�����U��~�O }�ݷ=y�<��o:U�Q���y�x���w��c5� �Њ���kQQ,<�w	ga�����6d�}��e�t\̌��-���e�r�<�dc�����!��|�2���ɞ&N��7�w��!/�F�|�%��
-7ע3C�[���t�r_��徶#v��-G�3�Œ�]�+��Y���y;ƭ�3�EK����#�w��=\S��鴾�:&1GbV�l�a�GX
�)M��"Dos��kJ$Х��h�	�� �u�?�;ﱂ`	�}>�MD~�ʑ�
~�'��q6?U[�͜�Kt>��6?5�u�*���P@6�C��9�œؤWo�o:q�q�Ӈ��|3r�|��͛�m\Өj�5�^��;V�c�=_�>�"tZIC+Pߒ/_��}��A��MÎM|o��,�u���:晊f`�2m?��e/y��5��q�����k(�l�s�Dg����!�J�D�*���NBUܪؓ.G V�fcst��'.��0������SG�~��.K�_��iogɬ
G�aT)^#I��}N���/�uv����C/�w�S^�g��|�gqG}J��a㺚�]�W�}�^��w�]�����}����1����U��x��Q�����Oթ߮�<mݰ3^��ߊ~��/R�b'tF�!0�����Y���d�7oN;}�;�������o���8g�G��N��F�s9H�-�ˉ��;��t�ctUy��
["e�Nq��#�7�f�Fߩ�i�y���ɫ;�,�zۅv6ב\�@0?m�zS�������OA哥NXy�7��m��/�DМ����z�MM���6z�e��U�X��[i����]����P~q'庝� �jJ���"D:��39J��q�
@��+糌�T��`&����3���X�`.��C��/#�\�P�j�;&=mh��o���_�5�^��u�~l�O�
IBc�Xc���ܯ�ҹ��,N �$`>����D�۹?�,�/�1��]9�z�1* 6#8��z%���&� ��X�W�	g%x��{ 'x�9�i�ྖ���^w��T���2�4��g�W:�T��������1���r��	�ǵU�k����O�����Y�������1�����Y�R�V�% ��Xq��+1ndY��_?�,Mj�|R���ދ'����S�-�ܥ����Q�:w-M�%��g�� Oc�����nj'|�?|�\�~h��.��s �1\u�����XVz�%'K��`�):��ѣ�Lmy8f�g���O㰙5���?����/���g��"�v���)������=C����KS��Ӧ��_!���@�i���v)�vqf������#͍e����:�Fe�seq��<��ę�j�k�S��Y?^�]�mf�̀n�Cǃ̊�ϊѭ��o�⟎�	�k��z���r��?��s��^����O��g�ο���9��Z��A�8�6�[���`�>���BYiO����8o�U3@�Wf��
rLt���O<�G�V�G{궚������vOG�ͻrLY�,�8�m�u�;�De�k�n
?�{��S���Ry�	WK��	�Xg͡����q¼�n����af��"[��
H����>�4�t�J�尟Hb�\��5~Rf�o8e��c(�"����R��	�o�0��ѕ��m�<WS9O�����1[��J�ī�œ<�9\e��봜�:`��-J�2t�!�H�t�7�B�X��ɹ��r>ċ0g�$�����+���q�(��A�p�ٸSld:W@͆�[z~O��m��W:e�!&В�!� ��8`f�,9��e�Wark�E9���8O3�d�+���9��4���࠳^i<4ڦ�u��7�Q���tkߨ�F�6Z���A@�{��x�l]۱���질v6�+0��o=[�2�'c�b;3xS٤�ބ�L4�B���O$��3���ލ�u\�$ ]#3�+��V��J^��(�ɑ:��Ƀ#���YlgG���v�"��I�[�dy���<	�$�}��GշG�͈�s��q�rtI{9V�����Gw�SY�ȶ���X*�{©�f���1�x�щ;����G�����u������]H6�;�n�<�nKbwDd��Yӏ@��};���W]�/N��~}�"���>ӿ}�s�ef�9o~�a>ҜWS$ݞK36]v��4x�8����l���S�����/x��5Z�w����sbq]�[����{u�-�z���K.�c٢����SF〩�S�G�*�p�l���C�r9i�.B��j�����H��u#�q���Mq�-���!����[�LT⦤z��8�LH�呈� H�"�(���vbTYf�e���9}F�8ja{9�~��Y#k�+M�2(�x!�Ŋ*T�� Sg���N � 7y�pqK#s��rU��~��T��A���T����θ��I&uvy���u؍_"��2e����x�)Q������,3тh��9��?��u#�exYd�9w����A�:��(b����f`.5[�ɻi�#���U�\e:q�6�Kc�ҿ�"��h
\��rT�|E��Wt��m�'����j�5�/��k?���~�3΍�`_U��s7O�P���U�gy}D��L#ޙ��e-�;]��J2g2�\��Og��,�H��C:����q�$��O67Ri����̃ �|����N�L�H�G�K��';?rrb*�庍z.��L�R0��%���Ύ�2������R����_|��'�Nu�:i��C��8�p�������l�o>��{���bf�����ݎ��t��������a��~Ü��������~z�w<�\��ԪC��ݪO���8�/��t�)�ѕzȱ�.�%d:���_;�50����L%�Cv�~�d����������q�?�۝�~��Sk8�c��{9������Zw��ۥhmX2W����L�^a���"�#53�ث��!�=ɤ�8�;���-�8n�,�?��<	Im�d�C��\z�U�mAS��m��0�X�7��M{g�b���f�)9�B�$:x�w�P>1'ۉ�N�
#�({QF*?h�}��]�ks�`��'�  ��1x�fd��[C.<��.͹��yL�8ǁ�a�T/$�_ډ9�B:��Ȧ���˴n��SxI��2e��m������<��&`Uj}v��̖e��p^���	}�V�i��~���=#3�ʛ[�y�G�ljV�0!�
��4v5I.{{���NE���?B�.�\��>�bp�~���ꔩ%4�8�O'�}1���n:cA28����m��}0�1̼Ӕ��4���i(v�d�|-'�3q����#�8@����{O:*T�1�O̬��!I�ȯ�⬽���}���2;�
y⚡���8���B-Ox1Z�k���Y��>��j����
��|��3�p"�����,� F��\�~yX*X�\x�IL��Fd�[g�I��jE��K<' ��"7�i8r�t�!3Ac.���!���;뜝���t��٣���!`#�����c�V�%y���ml�����6�����tl�!p-y`��9�ʹ�N?��k�A7�xwލK�w-��Dq\;�8һ���켭��S�CE���֌'G�ao���x��M��{����7閬����%[��W����M~2N6���>�b��=���?W�ym.��Kq't���}�	�W����A�wc�]Ռ��~��R���,f�,�}�'�c���?�E�e��>�M"B��k�]�y,L���𖹦vi#�=����1�� P�:��2}�8K͍����A��>p� @��(�%�����W�MJ���ƑO�>�*����+�Xe���t�J #����1�gɫ)��'��EB�O_>�Y��z@��g�#���e�ϳ����6vɎS> �+�"�ٵ_�C�����bsY]�'3;�I�I�b.��p��:wk�I��(�Q���;9g���L��
RO���ܫ��*K<+~�r;��\*������o�+��(x��q�|�А�@r����!,�N�1
!dNE�Y>�	�u�a�7�Mg�W!�3(��b�� �Ćh�)�X���i/�!<�s��g�מ�>�۴:���'�o����mt�3tt��d�Oi��:l�9OY݌As�9EFX��Z�SiG�\�vKW�:K_:��� 3p��D['��>�B���jf��ڈ��q�!���d���oǶ���Σ�S���:�;0ԥ��4��vΔZ À`kw��� �SdD���|�8�|ѥ�������¢+�r�s�S��S��u�e)��>�ْ�{O��A�3���M`qw���l��Qρ��kXU��Qb�?%��;ߎ���[�O4*���Ni W���;�����I��c�ő99�)�׽�9ظY//�5�ũ��/��(��9�kx�^-5ҝx�!1������w3`hxY�'�̐�u�Q�<<�����U����OT����ٯ�S��)�� �RR̓N����g3��ًT�bg�s6�������)N;���O����u`�	�6�I��G8K�?G��2g�C�ٶ0�mk1�8<zrSC�Yx��h��/��2j+_�?z}�:]���Wۓv�x�5`�E���z<�;���fk��hG�ąF��������y�^[?�8�کH�2����7���ak�K�\��v��+X`��gK���;�ٶ�=�/S@K㬅Hjc��i�8Pv�����Jl�ȼ��}�̃/�2G��=� 7�$	�ZM(�*&/�K\ğ��2L���T��[ل���ފ���P�㒫s,��uf]T�M;� ���+�Nw���5{�d�c�.6���k�G�k�����ZHz��t$2�F���l4be�z pu��2�dU�Ы�%Ƚ#�'��r��b$���vG�i ����ϫ��2��e����	ё޹�s*���q�T���t/;�-XlG.�"$&�l�:Ȕ��1��Cy�;�]1[��3��|�M��XC�V�Z5,]`A�wj��'�Od�tgZ����Y�i��)�9n�S7�9�횼���O��α��sGF^E �k4͔tC��Ҁ����I��c���|=|�0���|�i;�>�g�Hn�A�p/L�le���=u�l`��i��0x��S�֝3<�����C7�P=�v{ٴ�Y�} =]�3�\�����m��9�7����-GJ _N���X8�\��h��q�u��/x��3��
��?����m[Alɒ#�{a_�,��F:��+��\)�ǲ�s��ܛ������q����w�3��p�_r����_�T��mn�����8zspj�n��嶛7m��\G���тs��y���r�̒�kn;m|�u�͢��S�I+��j<	p$�ղ��w{��
?9�d ƚ���/ѝoM0�?%)t~��z�Yo���`|��j���漷��J��5��ewx�T�՝�9�)�p��9l�D���:@z�	d�W\�]y[���h��MqL>���e�Sܶs�Ŷ�͓-��F�ڙ��4�r܈cާ��7yO��4om�GG���QV�W��;��i�<��32V��!MF�<}qq73_w�|���ٚd�����w"04E9�C!�V�|荗)���k�S���$�	s=i=�R7w�'�'x�RC�g���l�6�3�c��e���8I�������5$���;^]��Gj��TұA�E�l�yp��7s�"Η���Ɩ��y]A��w��v��Q	�43ż�t�u�s����(WC�ǖ[ɿ�^��}-�e��*߷�f�xF���e�w�á<��g��A��x���x�As_�&/��[Ѕ��7I�/	g�a�a�9���Mj�E_�r�D�3�#yd�6+����sK�'�Ζ����	#8����t/]|yi<���
����4���Fq�4�,f��>�A�ݿ��<���ȷ�.�D�N�x�N��"NgM�95A�O
G�Ȱ�ﳸ���5���v�ը�4�i���z?�\��&����#��nw����AtCǖ�����p��(3��>�&���Dm�l�~KNu���~�T[��<����µM��ˋ_�����|K����O̔g���*��Q�3���J]%�����h�b�����/2�t�����_p�e4���Y+q:l��.0]h�K�i��[��q�:;�oߐ����e��܉o�ST���|���1-yE	�IJ�^ۑ�Q�������O^�R)����U���6���U]dqn��A4~j;���贅�#�,NB�5�?�l[;�D����>p���w>�SY� ����U�[��]����·�;��U�dK���$��2�����*��?�l�g<�tx�L�;��G�횝���d՝LVE-���/��دr~mO�I.��k[�L�"���i�0��A�q��F��3x����EF^7�I���������)�a��Y;��f�x����b��������*��ؼ����L����HH����g��'��E��1�P�1�vD�k�B�X�33�q��C05b�l�����|�A�\#��cFp��f�r���H�iDƉ!�n�\��3�u'N��M�Sw�%��5s��u�K9(}�XY��0L;�2Ҡ�4��K�Kw�Nا}�2m�O�����Fֈ�
��FH�m@������I?��U<����6��
DP�Bx�����������L�ͅSchK<Ǭ�xYi���,����⎼:z6�J��v�<�ݲ߲.��-}0�Y<���c��p����39�E9�k�_�s������JO>mtג_�ؒ]��H��W��O����r��1z7K�0N=��O:.z��.���������ga4�ʃ<�ų��^h_�X���+�;�4��vv�ĕ�9*|�e�6�s������#�Ϲ>�+̥��0�0�[���|��@~rV�JG�R����߾�>/!O��wa�Ӂseꀭ��7{d�����4���s��罗��n"9b�������!*�s�9��YL�]d�$��n��L�R~^�a{��U��Y�Qʕ�<��F�'L�#Ƙ#`�A�F�*v��}�I
�sVQb���gu,��䧯��x|d�L%N�C̆ ~K�=�5�����	 ����S�o�\d��|;/��ܾ*i;N  @ IDAT"�I`�gr��n�É��\�w��}�0�Ўo{;K�9��KXۯ�a N��W���<�l��(731QM:�xdϭ�U
�u�Lw��F�)�'�4����p6ř�0�r���z���b�G[ [���;@�9A���\�� �ч�fjU&��TH�/��s�R�Ǥ�F�g��ta�ܦڂ?aʘ��SDS�"d��:�'[�&x�q��Xs�:��8|�Q���s�*�h���R�v ��\p�	��|�������Ҍ@=�DGk�?���,c�D�E��Jv3F�qx�ݓ|BGc�B:�s���.O�T�7��c�����@N!N|���<�^����M�ܨߍT��*���6T�D��9������� V�}�¿X?��:b97%��!E�82���lǛӎ]~�����	�4�ޚ�O��O�4��D'(~ʋ2_��������S�!������������;~�w|y�79_JI�Op�C�#??�!��K9�>rr�6��XO'8iM��R��ѫ��kw�%/<����]NS�M�:S����#��.:�s.t>f���i۹��y��,?ŵ��S)8˟S����c�xt��l<�K~��X���ʺ�X?�v�2�~F�`����m��6��޿�)�{��?����Vӑ:fyi�ޖ}�s,NRt7�ם8]��J3}'��t��|%=yqG�w҃߉��EOR�9`�?�$�e�L|���#�f��r��d�T�;q���g�,����]y#˨���e��v��a�x�<�<��k*�&��x����^��|���{ك~��^�>kg��e�t��S1�S�3�`(x��O�3���g�r��f&2>Hց��,��q�sU��s2�r�>dlG[����>M�l��wp�v*'���𢟾�}��i/ji13`7nev���0�x�����D؛��R&��L��Kט¼�SAG0 ����s6S߿s�8�tz��̼N�/��>{܎|����9�x���Z�]8��,�N�uO�(a�;��E�*Qg& �ϠriIП�7��w�&��F��z��m�K�7�T*F�,��ݓ���鋋�2���v��~S��ռ����eX�W��7���}8�G7�F�f���1�t��)�<5�QK��'/��WE��!;O)Z���r���=���>�T�:}i���H��X�2�hh�u��9n�U��=]�4��o�Tƙ���`�cp�Zd��f3r��}^�N��:a#r�:P�� �a�b�N�x*����2Nc3v\����9L�d�b=2}���e;��7���\��I}zS؛yiH�.6`?�ӧޠoS��,IY���%ɇɗ�X�n�b8b�x��V�^\i&���~4����3�	�HG��A�cڎ�
{���B}�s�����.�.�>aF��6S?cS�=\r�k�"Y���瀙��*�D�2;|�ƻ�9:��9� �[g�����O�'�k�?��3��2���V@+�n[�U^��Y��[o��9�1�e���1�T���Nf�SO�����>�׷��m,j���ы>����'�VE%�㹨^�O[j�#���r��Y��]D2T��X03_�|�5�[�up��`c�e��o�Y�쾳����+l04���Bb��m�w�EeI5�3L��v�<�h�36�>����y�s�F�5�-Hi�k}i���䛸�K3#�6-�|���3xO��A{n�C�i��#N�8��o��������pރ��P���8��op�>M�+���4��ѿ���y(|,(��M?�0��d�ގפ?k&�
�XxT�<��o>��|�T?I��s����z�<�_�6_2�J|�2��m�����O��/��w�'#E�B��9�#)�(SD���=�`Uw�6����p�?��gU��'4b*����N_���M��T���=T0&O�r?��/ܫdU�R��L�~�Z���.�6��s��w�_��������|�o��ŋ�"��� *���&|&�mglR�/�i�@��E�����G#|7{�셲��Gǃ���=_k�Q#�!K�c���b3(Μ0�S&F��:�o�P�#�T�-����F�i���Hǡ�fê�H�C�ɡR��I��u:�i1¿}�����wOG�@�H�iD7�k,��L��!��1��V��Y�?�T�hA*+���ٿhhb oF��G�Ȣ����]��oy�='�}�#���s��멃�LX�q�!�x���m�tJ�6���?�ۻ��;��~�l��R�������6P��rAi�s�FMѯ|��'^g0MY�hي
������r9ߎ�rt��8_Ż���m��c��o����AMIic�S��!��g����'CeZ^Y�WT��K��6��	�w$��f:�^���^u~��xt�O�-�E�r� �a�ێJ���z=!��ؔ�����C���%HŇ28���p�4:������3+Em������̭v���řѲ�6��nhh��O=O�<��7e���^��-Z�x��k��Dʽ/����O�[����TԹsN�Y0����ׯ����7__<����$=�>|E��c�|�~�A�,��Ǜ�e6�F��V�0�&�2)v��Ù~̲ܴ���м��j�$��H�a�F�:Q.o=�Yތ��,�?�d���{Y����x��oE_4j�1mQ��RL��B����Vێ�����O�"�Pye��kS��8%mX��v鷂8��Y:v��e�(����0U�)�8�Ȟ��~f�o��Z�8���A�k��)����)��nmUk�����>jߗ���m�C�f��ܽ�NA�a�j_z�-�K�����=���v���.����8{6��Թ�e���`\�G'!�E�6�z;���NGoi��GH�V�`������'��ghۯ�ܙ��L+�'���U�
��Y,IakHK����I���\��OY�2ŋb�lob|��I^X����B�?�%�1 �Ǽ�4PB?g��!eo�5
f�,�հ'g2�2(Fg��a�_���vI99_�g����2$�v�L�s�� m��_,��W���F;xS��^�寔�ѽLE#�:zF1�W��K��.��H����ͣ�]&�����<�G�il�Hfj�Ȅ""*O�Ȧp��Y��U���f.�d��K�����SVN�5�?ԩ��-�O#v	~:W���O�ڭ�����1	0��X�	�� ��!�v�xu�%��5hߤ�~���F��Ӽ�����<ݻ���O�A�B�̦Y����8ʭ^%�r�&�M�z:��x���]��
��{�N�����,�wd�A�����@���χ����)B�O+�W��*�U��`��Q����5��7S����F%lk�J��L��_��]����0p�?�r�q�2%r3��;@��5���o�GgŖ���`��p��c�u��RY�И���N��'��Γj�N��F��%<�ym����=�:�k��Y��KY���T����n��J�t�Ϟ���>��櫋'�[􋖈��M�������y����m���*A�D9�.b0�ԙ~3��~)w�0�dc�WY_�NL�.�\��+>8���
�t/�$/��A��~>u7myz��5���s��d���iy�~�ѽ|�>S����p��J�8_zQ?�G>Q���hsS�\f�\?}ε�Wʡ?bϟ��J�����}�>�,�0��7��O�{1͎z�Ӛ٧�>�lR����;6������o2c:��6�Caܼ�ͧ�.�����O>��vy�!�L8�� >�gO'ɱ��w�%pD��o_�~�	���7�C��a���<ѥ��y���qN��M �������ƋG{��k*�)s��"�(�,�$=Gx�3g���D�ah��w�y��fA&8*܁c�PE��)��sY��Zzt�f\�S~3F���e�x�,%̚���ց��'v"'�b���2�c��|�,`�^��|yGG�4#?��|�S?y�K*<��4��9fϑ	�D���58׈(rz�ɇ}_�g�}��(6c���޴oie���ENl"�4�T�S��t����G���ME�>r�b��:6��.pt�,H5n����NwYvyڡF7H�C�A$_���/�@�a +�׿����AM���C�&z��ieOq��Ch�Wd4��ۥ:�붎�|�V=-��һB�vH�z�l��Dwq��� ���'e
����^�"�����t����t�?Q�!���6n���Ҿ����KG�����!%�q�����?ǎ#��3ѥ��d����y�YUѝmf�~%.B@��zW<;Ϝ�^^�Bj7_�:嘜?�h� ��X�[UT}����Hv/���r�O���"Ψ����1����-��U�q�]�#^w�Ky"����L�ʾ*ؽ������vl�|�ٯ�9^dp�](�;��lfĴ��^d�*��M�zcw!��=�d�'q��8=��-+�����\�)��֘i;jt�MN|�����G�y73y��L�꯬�hr�q��U%V���PV~i�?ͫs����ŗ��E�q����'�ҧ��<^�䄙�>���GбJD���2��>g��0��^V�>�Caw��
��&�J>�ٓ���� �X'�8���K�#/u�U�eR�|yR���G���������3���v�N�ۖ��˚�!�Wq���` ���of�;���{����W�@��Ŝ��ü>�������F��Fu��	�Lu�ي�=S�~4����T�'�a�Řb�(jw�";y���8�aR��p���tN1���8״�த�9<t`gdUK���e�sV7C)Y93��C��|�8Gn����=[q>�p��2�5�6ۛ�����a�1���>�U8IT��/3j��=wf��i�r'�=2�>5/�1o˥㸵����܈��zx6#Ff���a��.'*t8l�95�۰�F������azv��J߭�����0�#�
Z�'\��Yi���=���͸a��%u4�W:�<��A~)+���b�;���2��E�W�k&ћ�=��U:3`^G�&�t��'��k�������q�Y�U�t^l���Y=b�Fj�S����[��� �Ki#��)�������ܛ�>_��_�v�c1Gj	)٤ԣ��Ҫ�z��{�wP?[�V{GG�3p��b�W���;��!��g�%�Xڦ6�8����i1(��+:��A*��T,��A�mKx�q͏��K�d<�����̩X��'�鱬pॏl'�^�� Q�t����W;���c��LN���&��i����C{��W����Gt�-#�SgFl����_�UO/��`�:����̢{�roB��qW��.�Q�A�����������D���"(�P�;�����_ۄ�+��v�%�J�oV�\g��*@p��J]�Wn�?����O.�鷟\����8`y�(�<w���Mui<�gf�M���rı���t�}�Ed�g�l��j����0�Z���Yq�>������{�O��(:�(��տ�8_�og����w0�s
�=O{��S?����>�'�6q2>�~�V}�+C"�e�3���8O�l�nQ�B� #�*j�'�
�2F��x,Ř~��{�1ƣl&8kbS	�	nΆ+����п���QJ�`*�[���Ѐ�����<r��h4$^~��S�䍷�������n#�YBӣ�Q���K$g�j6b�xsq��	2�T'��Wh�4����a:S#�*50��i�9Op�ֻ�Z���o9P�Y�%��2�A����w��긥�ǚS�	3�|����� z��n���؇��%P��N�8��e�������8�����R�>ϋC?���:at_�G?�m��y�̢��LYɿ�6_�������K�L��t�#X����nG��I�ڔ2�~c�ǩ�����yǡ���u�Lٽe�q��-�Uf����G��˿d���[�[�w>��u�k7�ہ�C}R8|��\#��<[6��̬}W���Y
��u,0hO��	�ڑ}����K;������Nݤǆd�Ym��l����۸����]��è�Х>�����ɹmjx�֒����7�K�)��Wy�V]듑ɡ��ml�N����#@<F��+x:�p]�}�mI&�JC�&�����>V��e���n���E��}��ş��ʊ�ۃB9N:� 4����<{� �p��E�<:�+8����I�M&�q�Î�*�S�/�tq/ލYϛ7���J�8R�2�|43�]\�A�}���KL�E��n 	=��f�K]~9'
����O��	�)�6>N��+����2� ��kvW��1�q$#�L�$�~2[�n�q�s��ŗ�}t����_����&�X� �gV0��"��Wy�Bd|+�����)o�,��)��raz�$��%st���K��P,3^��n�	/t��~�(rL�����`�i{�xh�Q=|�ty_�.�3U0z� v����|������=rOZ����R��I��`,8�#��䜃�!��Uح����#�3�+�ۉO����H���( ��V#��SR�$%����(L#���s�iV����N�5����Wi�gf��L^�8�3��=�K�VR)�Õ/�m��Rډ�}��d���qh�z0�Q��!k�u�]�Ll#��xq���ց�ݡs����u�v����1
1�e֌��@W=
͌�ѻ���5���S�ޮ�63�>�N7^�L ������#/��"C�o�k���ër�D�w�Z�|p���	{�b���:|�9?ut�����V2-�W��^m^۰���]��e3�l�͒�ۙ2���p��f߰�9�8lh@*������r-/�u�+2��ڬ� sU�'9y�9��H�ԝ���4�mX����!ï��mCR�T���M���\���v�u����/�:\o�/�G[�� ��Z���۶nXj�U7K�O�>�c�?���<��Q:�s����V���WY����N�>�tٶ|�j�����-&�;6Z���-�]>�;�m�WܩlB9�'�t�-�k�L���؟u*
#ee]��丐gDg��1�)n� �Y{�'�u�{~�������
D�:`A�-���i��vE��'��Q�6zī���&?o�E�,����"�v� <�{�2����s>�0@t߲��R�7|�F�� ���s@q$-z�cǁ��w���*:ŔILh����������g���x�-���a5��Y��q�f��gg��Ͽ���������uں�����)�%{��q7N�+���!Y*Ƨ�FV�VXN����Ir���^�U�Dt�+}'٫3���8�`���'Dnҭ0X9��ǕJI}����e���Ë/ℽ2H���ؙ=}tڷylfL�S�k@����C����<
HQ
���7sߤ��j�wzh̲a��y�?��L�/�,�I�!$/��`�#�8�p��owk�p�rD%�7+��Ԡ��!�+#˕k�ҕ�W=ӎ�SEo*�j����i�(�z��ud"�"b|w��K�3��(��a�8��ˎ���z7X��>�4m4�PK|tm���Uf��m�Ӏ3Z#�����%�«|Yz</W�O�N�:Zr�����|���˔ϻ�5윯N�ǀ+?2
mNF+M���M &m`�Ľ�	���N�+��<���}�]��M9��u�Pw6â'��N�L|�O�6⥏�t�F'9����f>8�:K3)�`8��������䝇(̎=���вL�D� r��ڙr���А�/��͎h̮��G`v��a���n��G~.��"l-���P����8��2vB/�t�2�5N�Y|���%��T�e
N�;��|ʣ�E���{�:v�]Q��'i��_�z�XN:[��7�G��6����c˼��O�������KM��ՑN0� �O��fW0���������_�7/Ǻ-/��Z�1��\?�&�i�ok>I]��Y�s�U��|���\��spH�J��ϫܼ���q0��q1���~���yf��8��3����㊁}��^շtE����r�ɹ<!�x�ع�^΄�2�y���-s� !6R��&,���	RV���̆=�&�w�^��0yl�׿|y�����G3���=]�'U��c�ͦ"��#^� iC\S_V�|�O��t�)y�H?m���9\K��ڱ�P	*e�L_�[dNӮ� ;1Y���%ԗ��f�Hz��Chw�>����,>���?�1us�T9[m�$K�i�S�=��1�x0�v�DK,�MQ��9W��)7SL�\�	L�	�ŏ�\Yvpj0-vA�ntH�=�I��w:b�
����Pܹ���q(A|�P�Q@�tDȹ����A^��G~{��3%�aO61&�%%Ξ�Y�َ��ˍiԽ��g�jd^5�
g�J~�w:���I�#<w��x�%���rڔQ�.M�Bw<�h:��/B��ӏ�d�V��a�IP6��_G���&�,��`�*��Q�%k�aVp:��Xy� ��
�Q��N�_�'[��T<'��MnN9`O����S��3T��z�N��>�G��32f+�>��LmgIC�-x��I"�U|{�v�J���w#��{�4�˹���e���#�Ǒ�<E�*�ǩ��8���Y��]iW�[�Vf�?J�*����:���j�1~_�pE�Z�v�`:K]���~�����]��a�@�Ouغ��>�:_���a]u3q��p�Վ:�{{�6"���.������|�m�9�v�ey��gt=��|�T|ͼ~�pUN��}}��\��>��	x��ٵo��5��m*��ex�L2��{��=^����x�S|�'�=e��y��t��)�>��`&}��n�j�*���Wq���]P������g��T��=�Wʤm6��<��M�궽JO�Ϟ%�r3���{�%�Sw��]���_i]���rnf�Ѹ9�ໍ*󕧲��I���sF1-_��T߭}k�M�t�3~f�U�%NU^$�e���_���>����䡿Ŀ�}�QM�f�tB%���%%�W��t�lZ�:+���3z�L�I�P�g���;�gsx���mj}
�1�ȓS�ʥ?�?�4�����{�J�6k��So��HFJ�хv��f�<�~�߄���x�F�����1�TP�J*8D�3u�b 9��u�@<Y�b��H`p�9V}��!c��uނ�:[�q c��1`B@�A
`h��k_��)��Pz��]��
s�6h�����ip�0g��8P�Hz4ϙ�F�M��ڐ�)7�Cw���|Y��x�����=��x*�0oŏ�
���'��蟆V�ˉ
m�V��l��!�q��%�e|1��I>�>��"�)p�!���q�n�qߘ`*����s��̍w�(<�8 �3�
��ˌ;�_ȑk~�Ce�7��������i��?Ө������<+����/��F���	t���Ȅ��,r�Fe�=��?�hf9ʩ{:l3�ˉb�#_�2��|ٰ�����#߮/���(�#y/l�.� �@��w��Jo\����,�rӛ�^韧�C�ü��cw*DF���D����t&�:���#�}}Νv%���nYt]�FV��U�:�Z�&G3�_}�u��70m�z��}�O}����t�o��zi+l[0�q7�%�t��}t�}6@v�?m��ֹ?����5��ffI��5p�����8z��3�`�ߴ��;.�Xf����ĩ�w���s�e��~����b���cu7��2rT��]�:t���!�(��2�ǯ/���w�He@�&�C���I����A�2��z�����y�~��>����\mJ��O>�4�샋�?���Qwo�m���߾�.:��(�>��̓��si ��E{�_�9\N�w������4�>�-n�8!I��y��B�\��%!��7b��t����K�<řٮ�����*/��s{#�E��у����_^��?',O��-o_��a�'�1O��A�ض��3c?߷��$F�jR:�^�s(ƴI�˃�q~�>��y9�����s�V[�(M��S5��~��2y)��ڼ����V.�A坾��ޢ��yf4��׊DH������|FΌ��kNA��}F�N�{��z���7���#�P�lu�5�2�2D�4�s�r%�5G8a���<��b�I|`�Qz�YAT� bX��T-������2��'5>����<uQ�!����	a�a!t���f�kʖ_��;�Oy��(�{�8_�u�Z��á��b��ũ�d�dۆ7��Y�q�x�k�2�{�t���[Y�|[�G�Y�,	ϼo�p�.��v�ng�{�1�%�N��O�hu���\e�}[Ꜫ�J1��2|F]�H~��>a���g�^�a[��`�:�ɧ�hٝ�"M�ɳ�r7<]���n��,-*�\�@�v��,ܟ7��`:%O�h0Tt�r����y3`f���lҥ7��T�
;{Cj/��N���ԑ�f�إrK��e���˟���u���t�̒�t�����Q�4;�uP<)@�6Tk�S�������{��9�׻:�����S�l}^ͳ�8��m��N�0����dO^X3'��W����ƠI��0x�X}���,Iϒ2=Z[a/�o�h�Ƕ�P��X�yaV&4;�;�����j��9`x`Wcm��t��a��4�z���:�_<`�h�k�`�����~.|#��K�s��闆e�+��o���8`�iHE�٢+����;"ʹ�n��M��q�;'���J�ڞ��|���Rg�fC�ۗ�p�#��q>ݓ6�r�e�:�)'���,y~�͓�ϴ�}�~����:8�F�엺[�!� !��+G�[�>'~���)�r�Qp�@>*פ�m
�b����y��ճ�yp�����S^O�(�M��x���+�b�^=�V����*3_ڧg��L.��|�� ��TN����*v����'gv��r˝���^��)h�ͤ�������9�c���5C6���N~�7�{�Q;��s3w?{v3��G{V���\gdn�e��GG?����O?�,k��\�K%5��;s�܋�`�����[�JHZ��᪊R�d ���n���4���@�Q��L8�z�Y:�g��y��&|ީ7�Z^��a�NO<BCd*!��$M���*����,j��$���%U���ix������Ѓ�e
/��V�+�0��s0��oGh;_��`)��lc��+�;Y*���u ��2��̉�+��I��,���h���7�fd�}b�g�`i���#�n�n|�<��4�-�	�5f<e�@��Ca���T��dx�b��Î>VE�꡴Л~|��}ya��&no�\�N�y��M�-{q���?�3#a/:οq����L[�}�4O����:���|��l�9���t��� ��U����������K_��aqt��'��/N�Q��f��$i:j������Bl�j8��jگvE�t%��~/�K+����CN3Y��42�P�8u�Y=�ky�Jq�9�����0O♅q���Mޱ���Y������i�8{�r��N2n	�&]��'��r �ֶ)xw�k��N��rs�u�X� ����Ŷ҈���'�W��ˊ6$�.:ʓ��M���Z�"�v�h��ul�|x���a�f0��D>���rJ�;	���	�xn�g�&=�Ef|�}�i2��K=����t���B�b �M��<��сu����{ʥ��,Lp�|-c���B]j+���/]��-CK���#�rŜ#�ȳ3W3��}��Ye� �A�i�?�{�O_�6ˏ��|�ͳ�?�`�5������뮺��>�Y�=M��ׯ�D}�q��݋O2K�]�p���P�ք#g۩��9�O��0g�����s�[��L͵���z��{	iR��?���T���$��9X����I�Y���u;���7������r�q$3�_�-��򷿫�z?�#��0����M�Wq\�v�����k֬�֯3��t�<�r�@yU�岀����j\9s���W�;�ǀ�E�݄��mg��Fy���B������ۍ�*<!Oc�-�p���=���^��I7{��=)�l*_�'�2�T�_�Q�U�U�d�#Q�L9��w����Y�t|�1�tuJ�M���	���Nˎ���`cْ�u����:Q)E����2�-G]i\�7�{i:B���!K�:E�Yy�24g�E^(�ı�m�`2���L*����FR#�|�6���q�W;Uz�4]��C�E�q�2P�2�|s:��w㎻��!�����0:`�M�)}|���d�o���܏�7�t�:�N�/�UZG6�8��峜e���M� �[�=	�t�6qGG��hΗ�IGMh�t��B�}�Jw,k�6��Վ;����{�{��wY�Ws��O�W�p��i��]��'v�����9�W3VVt����A�K�
�a�=�S�l��A�܎�z�An� ���t7�\m�^��מ�A�o�yL[�c�_�拋�>��MbS��\��.����҆�n�q%.�^���C:9��Y=?�>6��vɣ����{�0|�^��Y�һ}��_F����g��� ֕�Ի:�-Ɣ�D��
�G�|���䎃aiў)v`���{L&��!�R��'9
��
O��.����u��R��o��搻�p�t?g�O�h��gI��-[�>�V��M�p�Kv��G��R���J�7ݿ���fo���sL_�m6̧o>��sNp���lU�苲�^���dk��<9��@�4�_�&�铼Fǫt���>P�h}��H>X?�� @�r����L�}@� ���0�
>�|չJ������ڜm�4�	/h�UD?���?���+��}`_�N��=����4ϳ���EF�q�ǽ��ӭJ�2��X;∑��*��:Z���wt�|*;�0���Mc�ͷ�z����C�{?4P�f�`����Sa��NP��'��hp����:�g�D�f*	�:f��̎�E˗��?�j��/�ٞ_<]���xEv�{�3ViT;���Tz����g*eN'9F3�՘ݪ����a��	�:|�3ˎ���5�/"_�m���[��y9l��:_1��K�1^#k��g��M�O0Z����^r7�/^<��I�<��n��sݸ�I�9�� ���$㉯�^_�dQ��ϭ�_7D�+�э<�i�lc�2�y��bw��@M#�F�������){ʟ�:b3R-���80:c�ᠹ���M�4���������Q�#�.t��-��1'��8`���i������?��b?/��K�.����ӏч|�lI�2t���m����h���<�м���\;ǻ�G���a
h�*��_c���:���`OL��)��gK���m����Ճ�'H�Yv�=~k�LGpH3�����g���l�)�U�9����ko��g3���l\���XBx�.g8����!\�tw���Cn(�{�����Wآ#un�)K~�A��jñr���9���/u;m����˽�Lf��ª��_���ʝ�θ��8�`��@�n9�y���^!��ʋ�e�.�m��
2{n��^ۻq�����2�F#���<)�0�s���;1�s��]$$'K�D��`����&I8����H��u
f���+��۷�|}v��o>�3�>�Y�-��Q7�d�)��Ϩ\�׫#^��f�,���v;�q��_f[�Gu^���_�f��;2!�i�"��a>d�4'���<Ӧ>�O�Y��5��M+X�hh;M �BŖ��Ix�k~��Υm�Yq��x�en���aZ��q;�9\����yAv���7}�����_�.����w��M�>t;Sj���)��=� �rL�8F���Q��J�:�tNJ��ˍ�$3Y��iu�s�����z���:j�Co6:� f�f��qL&S���W�9>y��,EYF���Aa$�goxO���R�����H6�D�>3��#�#�0�����t3/������,]�K�q�Ҙ���iЃW���S�FOf��H��d��:{1@��}$Ň)y_�3k�G�sO�!Y~m���˦��ԍ�1p����;��C��=j/` �Ù1����L�o��O�iW.��1�D:�tB:r؁\v �_8�+��-a��a“��'\��]I�Cp�˶���v�v�V���L���.���e��������5Ӯry��}��$9�����%kkdƍ,g��	 ��[��g��)�9]�i�u��h��W�]����y���ZD�Q�q���,k����Y��+�2�f�M^g���ی� �s;���A^H>�͏Sď�8�=^q������#";Ӎ�M���#��<���ʋ'#a�~?��{ΰ��>~�vrC��ě��	.'��}0Ȃ̻WUʀ�}�)#eF7�c-��\�ɳu�B�v|7���
i�����Ik��_�5ó� �c���+~�O��T�?5e�%�x�%���G�v ���~����Ƀ��O��L�>���9e��W
|/�
˹=@�ѱ��3�a����1����7^�K&�S]���
/��{{%�h��9f;u�S��N�����S%l7�З� ni�׹(	(��|pȁ{������ذ<���Y���)���R=�%����bc
fKX�:<x����|��nɑN1��B9�C�e;ۍ��Yi�3Gڏ~-9����q;633����ɞݮ_�<H�o~�NT�����Ŕ�7-�vsF��le�+;*�g	.�����\fu>E��D����|����!�����1�8"�j9
S��N�k/��uG�ą�>�)S%J*�z͐<�w������md��Ouq�I�!u�+ |���26F��W{�I��z�X�g���vㄨ���2r<�EҰnG�� ���Wa�1��=�hOr�5��������Hr((�uU`�I�/��Y�w�F�i�F��|�Nl�8m���L��i�A�頽mQ���(�L;��5ó�=GѦ��Y���Gܔ����wq 8_�jh ciN�1���,0%����󀑼�S<g�N�#;��C����QO^ף*�����)�G]l��Bm�'�dFp4�#���'���1�#�iK��z��ڞ<ms�,��	��$K#�<>����1[�O�8�=�_x�3|�n#$0p6m�����^��p�@u��=���%;C�+�@˦	>`���C��:���ԭ���_�`0��[2�����[�fژ��E�+���z��Z,�f�(r�S�d���޽쐾��F�7��>��r��뽽��qO�Ŀik�W��8�\`�g���Ln�8q,5��
1��*ӄ��yy�{��@{UZRZ�؍=<�џ�=7�_�.B�a�9��u�lol5�z1�k���(�����Jo?T�\�d�Bρ� �{������3��M閈�������3���� ���}QN��'�0�q�%�q��;P��'�܇�R�ރ�r�G�2/O��,հ�W����}��>g�톿J�����׼�����/��R'{�S���+Ӫ�^σ¥Y��y����ϩ�D��J'���g�~��V��U�q�.yIq����#,_���y+�3���.ʾ�eVA��m��V�����\�{�E��^�q�+��s�2A���~$=�)ծ�\F����vF8t�UD��-���0;`Ѽ�g{�:y���� 
���9�Ð�&�2��VP'�Mj�;gĐ��;���m0^ˆ�6��gy?�x�"�0:���9��&������8
�I%�h�>e',��m>����>�L�П����/��DÙQ$����yjZS�i�uvR�F6#�\OȻs�G�tx5��3�>Dt�W�3��C�iG| ��i~:���h�7�%��O���E��p��:u]�z�޷�8|q��:3����~�7��4��x o�ϐt���	��)���W��[ж+�u�0��`X�|b;��n��ե��;���H?�O��3.fh�1�Ei�
�t��F+.���r�#�dCGA}m��5#�����3�\u��$�T�㌠X|/ߦ�턎�ǂ�is���z�����z�t}�<����r������C��~�9�'l�����:ӆ39��Ȃe툇Kx/�0e  @ IDAT*�[�� �@�w�s�)G�3fa�z���/�{ε�G#h�Vց�Wv(I>������,w�c�'��(L�w8Û�;��U]��%��чh�*��uaĠ�Y�[(h�]��>��0�̚%N����|Y\�?1P����f�!O����elp��=ߒ���;V�k��O�v^d�l�#���ŉ��((�X��C�Y ��WH;�w���zW���\
�S8�:��"��FO��p�D'.������EU��M��1es����&L����һ��mM��t�Ύ�e
k�"e��ND��:W�����l��������N��?��
918�x?|�7S�q�o��F�q��ć���L}r����X��2ypԁų�G�Q�ɳ2�K\����^&Gq��7/����S��r� QO�Uɀ䤘/MB�dI�.ӎO2��u֢�r�B�̇*G�=#_Y|7�AFe��پ?%��<��h,���������?��!�-	ˣQ^�m��>�{�(E&�ѧ�ԭ�i���K�o��N��`C��յ�k�)�־k��4e�`cl5�>�v:|�d��2���!k<�;�*On1�]/��5Ζu[����Yh|�7��=����8)� __
0ږ:���������7Ů}��rOn}z�{h��,8z$߆�tk�Ǚڡ��ݓ�i�"��O�/�OPq�9�q*7����0����G]��9~�|��?Ǵ�ܫ
�u��!�O�{��=3�i�n�`
����J�Xy�M0�f�dk;�菩�FG�9D������ږ_�cj�������Jt~�-ݵ���ܮ�y_����7ҏ8���#��q�;v�}��|;����]��;��{:�q�[�$'i���<��,��o*�意�}�h��S�:ɍ#ű2R������ȥ4�/�l�[��c*���Hv;�CÙ��w8� �
�_�'^��[�]Z���/s�p ����um������~�1}H�Ŵ���5����z�W<�:��J��N.davᮭ�[�#�C&F$�z�&E�����T��#xo�N��E�i���O�׉M���8#3�`���Fdf���HN�	k��z�\?[��K����٥7�=��)��^q"�Ӕ��)&�0{���!��rl����z�@b��ᡟ�т��pM;^z{�.�+۲d�:_F��-��{�]m�W���K<ϣwIS�)���^^��#�/>ϺK/�\�i{��7�2�&���U�(�9{q/-�������w�ۑ��H��h��ʐ��u�َ7M�v��y(kJ�١� {�2��[j���{�a����������^J5�֌8�8������Н��G����(��)��1pQ�0C��F�_ޅg>�b4&oZ����'�Ԗ�A��������0*�F@�mI|*�R����D�E�s��m�y��h��5҅�il�������t��cu�i�{��Њ7��n+�����͝x�5�y1�6',0x�`s0��G�/�X/Η�����)S���s�𑣠>���u��}�
��?�C�FGT~:u+�S�	
F��*�b�� a�O:�x�$�ˁWgW��:0ZX�v��1�9ׅ/��yε��wR˟�+N�4�³�m'm�!g��{|g荂p�t������.���x�LS$��-��\yFP��|�����(���i:�Pz\.�7���&iKnh��M���}~U�cھް�y��N��ϯ�{��p�q7�7���x�Xp��|�:�An��y�
<��)�'3��(�;�k�����q��*C������;���k�6xG���o��(���7�v��'͸~ڞ���'I��Fw�oXIl�3���{��5Ӧ�up2���qb6��N���(�C��%j�o����:`�������\�<{��L���d��~�k�����9�"s�Xץ>1����e�´V�����v�K=��)��g<Alr��Y��X�q��We|�,˫@���܇�\���~{�`��ѝ�\8U6�q�L���87�q�ne2��;Փ�	ۘ��r��HjZ19���C�W9<�l����~�Ӂ%�C>C�^�_�܉=�cưs�~�oB6q�ȿ<:�uuM�GGN���S7��2O��3쳨0�*R�Hrm�Χ:���qΫ�jg��
�P^5�J@�߀��{/�4��N7Ơ��|���
ܪ�pT8Gи0�Y1
g�k�V���>��X�1Ĕc�ꌸPs�:*���)^��O�^h�F��wV;�i�F|(�~�p?�����u�}�n�f�(��r��2��E���a4\�S�〙wƘn�g훼E�\#aDȨ:�tuc�l-bt���bx�ѡ>oH*7_H��?��r0w���?��P/�Wx���yrI��{v��+u2�F�f �(�-L.N��gČ����h?���搸3��3�A`w@�<9�]ñdq�w0Qn�x�+����34�|��^+�z)��x!n�w_��aǸ+��6�x~A=p�� �.��CǮg�٦c�*�ny�?��z�F�����+������sԏ��g�=���:7M��Z1εP~x!ω�I�z�x�={�6�=g��@����y�=kmp�婭�,i;AWǰ��(���6ޮ7�M�οӑ�䖕�6t�.�c��8*^���H�wRF��� ¥�%���<��!&m��8v6��S�ScE1rbS��vK����y�:X���d��F}�����Ǆ�%Ǜ�਋��a�o��p�������x��sf��/m��yIn�˼��p>ɡ���/r����#��� ����S��K��X���9��������P^�x�YF�7�t�)=�[Y[�<��p�|��XC�v����������|����d-쯞f�w�F>�Y��{�5�Q|�=b�}VkK�Q�t�w���-{Zr��}��s�T��m������	�M�1��te�>Fw|��]�_f��
�;Z�'�
��B���it$FD��^<�{�-��Z�x���,�
�#�|Stӛ��<�.8��퍐-NJ
�P ���>��s�]��(�$g`�,R6��@u,�m`ΎbU��zƀs��[��؞:M=�F���(Tg��N�_eb@l�0#_Q���<]��QBOG�q�`�/�iǎ��N��SL���f0O1�(��(Ɔ�\?���g7��O�ث�?4ލ�D���I�p�x`tk�F/9��$yr(�;�q��5W��h��O܏'=\����ɜq�{�IK�͠D�x�G~�)#�)=͏4�1�	}�
okTS�<��|d�G�+e�Y>�xH>:O�tK<^��Ȭ�� �W;ȣN�my4��?9�D�x=mHҎ��CsO�����v�ew�/�����:o\���ew��+���w9�tCa��@v�>k�s2�I[�u�su������溒��E�����t��94�s�%a��!Ѯ��G|���o����zk��ɻÑG;n�[Ϫo����	�jltzwhl�:�Ռ�ϴ�$#�<�K_ /��������W�4��;��!���ș4��VT6-5NG�e��{�sۨ~��2 8S��S�9��J���O��!p]d�r��5�on
̳nB*Jz3��B��]y��lp:�"]\�Y2��8$ax�����K�'���%��pqh:��5UF��4�����������G��������
o���1��7_f����뷂Gڂ�m�@G$�v�T�D[�e�#Ӓ^��b|2
�2�L�t�7�w�\��cv��f�ݸ���6W��GEMI���,89'�C?�-�)"����U)��w��&� ���eq�!�"�(���b�y�nϧ!��E��S��r�v�V��=�&p3ϨR�!/ǘ"�w����:���<]t��mR��֨)C��/��X#<�)k���2y%���煌|Y��9�W����o��Z��9�v��9��k�R.�e��1����>[M�Cq|#��'����{A����ٻ�Ww<��B�)w���{���x��m�8kஞ~=y�3����B�pz`�����ROC�PvB�>B�\�;߷Fc��Pm���St"%����7����5���Ϩ���r�͔UG��7��Κ�z��O��$�4����i[0q܊,��b���栁Wg>�&�����Ai�
�lG>C�'��x�[�4�~��w��u�h��(��8���YǾ�~֡��+����LB���Z�ҩ
�⚎��u��L}�]����
q �9 (�
ꀓ��#�h��8Ϛf����!NBGs���]Z�sή�n']9�o�.�Y���5��mz��k�	^,�M�|�~R4� un��ނ��]o���S^�O�ܼ~���fT���Yô��Yե�^�N&�aJ��KB?�/�1��kKsƧ�����X�o9��TY���y����쏵e��H������E���*��H[�>����o�:e\���G�NY�،�lGݾz��fXS��]f�'+�٪���w3`]�α�Y��Q%��?08��=���ڞ�<~�͔3Rj���H�>�y�M������Ŵˎԍ_bz4�>�4В��>��>�u��A>�v��f�>K\��|�/��Y@�UW3���[���	1�3�gX���v�ٰ*�"ú��k������m�IΔ�q�?�����7���`��s�������W�z5u1E�+�K�8d���12C'0�NnGc0��4#�젷�^Q��;��r�5_��C��xS����`��	c4Jޑ�������X2�pG��`�PS�����5j�9��R֔���.�W_��:|��gH=J�����¡�5w���gX��j� �;���(�N�����Ȅx�8�T^������[��H�ҍ���|
I듬����8Ɨ\�����Cu�۱[^����t1��i�{A+'�������쮳4����ˆɟv26^�`Wr��q��q ʋ ���-�����?;���=�Q��>��x���y*��n����fǃ{���s�cG�4�=�Ӛ�|��������'uj/vD����	�uH���i����#�xe�ץ ����7Kow����CI�:��ϴ��+���'�=�5�F���J,�ǌ�"?����Z�m5w��;��!�.�^����6��Ɇ�utrIm�(Ԗ����4b�w�4�S�sr�7��5�RǞ<m4p�?G�So���Oe��`Ft9Ȓ�6�i{^��4��82�]kQ�V19��j�'��͹�!�	�v*��}=�A�����l���t�َft���/��Sq�N�^tY��
�O(��틜Uь~N�W�8�%���^��>N_�$r�kX
�vU�E���:�u��~;�C������DV���SQ��r>��w|�Q�X8��8:���惣Ϟb��A��c����U����x�Z����#BC C�l�7�|��I>C�P L`(�W}M��3bƛ���ə҈t�9��E(��eTz�=
�3h$5�=SZ���~�Ӕ����h\���#e6��"sh8A�c�<�<)�I�p{򝶋P��]8q�|F���v����C��s�4F�Ǭm�3a���,�ψٳ,�����H!ǡ�5>pCK��yk���=�t^͞��!x�X�<��'�.:?駰��ܚ~'��h�;���٤��X\4���7p�嫯|��~kx�w9.t�0Z��G�|ByY�/Jy�8`���#��@�1���h��S��ĽC�W�fgr����Fit:W��%k���@+���Nu���ӎ�yn����?7�z�9^o�G�]�1��_�i6(F�#��,�3��ʒ/�h#���J��&$e�D0�����櫼�`_�S�7���A�B��*/}e8��H��1vT�=�n���p��:y�C���-���G�)x�OYO��ݑ¿��U�O��v���U��&c�!��Z�t�n�����+�$��[ƒ�J1��(4��t���ct!�|`��é��s����G~������IHOٗ�Ъ�jCg�)݀~4wK%1k@^�5,����7��M�"�3�`m��>���G�RRW׊�.O�L����ؚw�ogW��tN����A�G͸�&�>�f=����a�ӸԼ�9η�
z{J7jS��غw��Һ�_}NMT�n^�o'�]�Kj���:P�C$�slV���0q�����c^�hf���8S��Me�D'��*l�7���k\��J���5�����k��=�A��4�3��S؂�4�~[-s@���@�9O,V��v
2'|�ä����،<;mi
���$�4��|=`>/4�x-��zE�btխ�.����֬���|lHg�pOY:�����Q�9�#���(��uڂ��Q+L:�i�I�|-oe:�?9����9/��֍��� �+_�FQ9_�?���7eu0��}>ƕ��s#C��Yy���8�=��%>e��n�;�c��S�1��wdQG1|�V��rq�#�I��a�\���1�ҳv��{�t�h᪫��<~��ޝ��O.�K?�+���_u^��TǈW\o<v]�w�Ӏ)ltOh���OؼضCq������*��'m�4�7���7;�~m٧���l�:�zI�,�ulR=�0���!bu�dJ�[tB>8?xx����m�2�*��B���cт����Z���?z�ȟ��';��nx��>���O<���'���t��\N��)|����8<�G��w�-^�0~W�O����:p9��6�X��Oۜ�{y[�A�/�@���/,�8a��-�ɕ��>�?=�~4AvH��
����Z<�S��������q��@y5������=~�/ �P�GmJ���Cg�Q �>�S��|�{~7��Kr������2�K~|�S��ח_��7�ɒG��G9_m���	�y�N~�\�;�#���,j;���?��X���|��o=EA�7��9�p��N�!��O�܏z��Y� �*��ޯ�M�,;}��MAJbZ�15��]�ȸr��)x�ΏFt���0mI>G��V��aל�`�'9Bk%��޶a���>5���O���ȗ�y��W��͏w}Z�������Q쎔�i����~w7��B>�dq*S	�3��h�5f6�����^�=z���4���D\<���_��7G�!�rZ�wmR��7e&೎��R�5�?۸k<�Dh��)YA�۸t�zU��59����ۣ��h٩^�	7��}��e_��T�;�w���<OҌ���)�^��U^��y���H�}�c�7^��_��<���Z���A:j�
��y  }��y9�����t3��;����Nۑ��C�Q�)��-���G���Yr?�!X���{gC竂�:�} 	?��q/�Vp�`���l�C�M�ɔ̻��TC.�z������ U�g�2�ӟt�EQ'ǩ�E���۽��<�ҵ�A�>���K�NC�(�-I;L�)�t��wM����u-��IO,����H�ж�t�!��i��j��?!$��W3�<�$���uq)��sm�D�������ef?#��+򕘌�$}` �O~|�)A[�p;�w��F�Ka���ns��xsZW+��o?x�oKf�(osߗ��/�)������09=���r;z��nx8�|nZ�w��P�k�S���'!f�6B�K7�N5�D-� �Y�����=���9��Bc�L:�r۫S�.]����ԝ$M� �	�).ْ)o�8�?ⵗ�2���r��i��>u)q�o�n�n���!�8!?ُ��,��S�ĆS	��/��T�$xi �j��|�i:%��(���&lU2�+��:U�v�IZ;b�0��:�36����"��Ι��Ԩ�W/��#!Z~bV���&n8�Wc��'�P�{e�1��m(�q�;��@�<J"�Z����T�F��2��m���MCe�9�,;嘧_g�*[6u��e���BϞrMc�Y}�'12�bX�li����R��7�Т��к=ρ�3wW�������)b�����u�~J@���4� 4���[��t+c{?0��X)��D5���$�"�@�� m�[k�A�(|�c��ҋLn\���ŵ��|��}L�ѣ�Ѝ�C�lp��)���������KHj�;��x��N��S��c�y_>2H�qǼ;�xV�[y���k< ?\�r�U�!k/w�7��oX=/zY��|����`�Aw8^x��bTkF6��C���%��L�$r452O�ڍ���4�QHf�<�i�Ns�YӍ��@�ΰs�W�.��#`�>�Q[?��u$�Q�8i:Wu�����--�<6���v
:�@������OiɅ3�'(��ė�i�{�8y�z�|�ܤ�ױ�ޒ3[�\��Q�nօq��X���3�:��t�isj�e��Ls�{��>f�o�	��,ݡ��M��:{��\��,+�3����� ?��ٺu�*��];���Y�d���T!Wm{��s���O?E.��C�-�B�����u�l.'Ӫ���_�}@gh�ӏ;ߜ��58,�eA��Q*�	�a���Q(Z�6O�����8u��pgd�@&ԥ
���J���s�9q���i ��(���ĳt�_��_e��|r�;��  ��2R(��|~&��;�sķ��g�^R,���3cQU��� �h)?�JF�V5���m�	��QS�.�Nk�6R���Vu�\�h�f�c�l�i]G��>�b8m��E���o����׉2��!Vʵ;
�a�]ǯ� �:��!���@R�Q:so;Z;&��H�1$v��"��3
�1"�K��?�q�L�u�M��eߑ�����T\Z��y��mF�v����pxS�Nb�۟*"x��\,����W��Ό���2E�{�����܍����S32���Om	�X�g{�_�h�������߆��#�|�ie�==����֛��F6��7TW�ꇋ�qsV��F<�VF�����k<��>:�]�yO��O�ٴ�,������㦭��/�y��u�x�#�q��l���g�(__�Ƀ���a�&���c���SQWyi�}��j]��ퟌm�褏l�;ps���gu�4������}��e鍺��6H�`�W�>�|�2�Xp�O��I�|��N�����%�~& �9�v���w�L��uYH�D<6����>ɗ%��sC���'��A5{\���c-�Q��%^X��%�������$���3<���sk<�������\���C�|ʷo;]�K�=�D�}�*�1��E��V��P��E�J&]�S��,�Ğ��Y��H�)_ +�$o|�������ک�pa SY����m������qVϘ�
�It8��Y��4���<@N�&C���;�^��r�O��m�u&O_��?�s�x����ޑG@����+H]�W\�!�Ð�@�'}��f%����ӻƝ���������]u���;z�:�S6w����He�ȵ|M��S�Ry�K%��C�ܹ�i�M.P���)��J��]k,A�@R��Q��-���Mu�88:��������R�VʈםL9�<�7��8O����y!�J8�Q~��ӝ1��<���A�ӗz}�k,#'׃Y����E��~J�C�&��!.�����*�|.����3^��#�=��Ӕ�����:�J��N�$��Ƒ��N���{_H@~��8��z뭷�XO����0M!�Gg	�Q�����qz�V��8_�:pt���,8�H�����{�A|ׁ��W:ONB(oY�
[�K#�,�����G��(��M�u��˽C��>q�c�%���\���Q~��5���g��1톣�:w��T`�V.qm���硦Ve�c���ۗ_~��/)�)D�!Agч��U�U��.]QW��\�C<�����$*�t�c��^e�){ݑ/.<�=�8�o��mf���{�kx��tL]��{DvZ;�K��mJ�<ǲN�YYv��x���T�H�y0��b�^>%#�=y��A&�f��yF�/M��Vzp����n��4��w|�0��}G|򆤼Bf7������դ�Q�D(h��,�q~ӝ��R��rr��=�O�N.\o&����%��z��+�+�$
�cSl�SN. u$��w�F��jiHҧ�yh��o��L�,���l~�ʭ�I�	�{r5k~Nu%5�l}���*|$�x��/o�Q�^�39�e��/�{��u�G�w�]��\F�>��ݖӘ�?i�c,�[�u��_��=!n���7�I���F��2���� X�sS�v|P�^��8��#s�W>*�{�Pjͪ�bl�=�X�"*9 R�����Q9,:4�a���N��t�����z	�XG�0:�@Tr~�~�N��1�4��=��8g	���RF\g��[7)3�z�k�v�Ҕe�@�C�Sq�G�Ft">=����ӡ7[�Y"J#٢u��<����3q�"<]���ȹ�H�!�[�b knv�˘�t���9�ɓ�|�����裏:U�٩I~���:K<�V�m٩8?5��py��5�ѯ1���'�t|��2S&�Ƃ��u�FF#���F�QM��CF$`u�����o~�?���q���Q�DD�_Z�3<;n�/�E�z�H�2Ń�v��Y0�r�����5~����0�Ty&?'���?�{�O:�d,���9ә=Jp��Ѥ8��|ڣ{r�s��v��>\:�=+�h���;Oҵ=#��9`']��"g��+:
����'����{�^����_�7o%�qqG���c�;�:,�@OqL�Yg�c�HM��+V�s:uݶ�I�2��5#_\�`�I6M����;yX��}6�e]�Sm0��ϡK����W���Y�4dG����oϛ���K�?ض�Y�c$�M��Nf��1�GeC����G
�=U��К�8�aq�J��5:�����10-���ɭ ��n)���M��������t�uI*��7���M���3W�6�@��Z+ܙPz�V=�$]I��u�t���tl�݃��uΎPU���n��;[����T��]��������집U���T �Ċ�������,���WK�������9D�7r�}uRbS�����K��hƩ�(Q��R�Y��}���k{̃�*���D���I�W�:F�87��_�)�'hG�o���	� �(pj�nؔ�!ݝ��g�*#0�,�)G��rCeaj@���Y�_	�4X����uf�)�dj��~��!��4O���Q|�O]�d��:��:��?� Y���N��vI��5ge&2��g�Tx�����/n��>�T�G}x��?����޿������?��ԉ�_N�>��S��Փʛޠ�1V�j rnǹ�C��J�Ξ���^0ZxR�hH>tTFɫSy�Mt����(���`p������m:�X:�:�x���lHyp�/l:w�}����;�N_5%:W�F��~T8�#�� ]��>���N�U��\�d�!wz���߿��?���oq�?����Y�2y?~=�K{�T���@�#7�������|ۆt�K�z@ޜ�EX`��Г�Sf�\M/;o�Bwi����`�#{m��(ٗ��&�w��]GǺ��ތ�n���k�v]nÿ?�Ŗb�m�:��������y���|�u��VG>�ӎF��^�!-{�W �"��=SX� ��}��w���@�^�{�2���<{4)@�G�+�\�\�g:3�=7/�)˽N��;�Q��m�I��%I�N>���i)۠�]F�Sy��u��<�΁k[�������o�Q${��5�]N_����Ë�6����CC�:g���=a^H�=�i/2����&-1�k	X����'O��Ĩa�_|:���=Ǹ��*7��r,����{�皀��q!I[WU.B������Эx��<}2�2D�;P%nC��S5�z�l�z�s=�J\0��i8���D�2R�N)V�z*��Q��kR*p����^�8%եZ��L��&e����ڝ2�����,e��اӕ��G�=��Gt������R��5���b{4�3J##g:Y��O���z}�~��w�E԰�����6x~�Qa��g�~��Q���A�~ey�)��>��|m���a�*��"���M�&��u�@���x�ì��:�G!H�:տ�������ſ��u�>����pX�k=�p?#�m��Sˤ���3|��9�C��}���|�f�ӑ��_��%�N��;�߻���[h��e�e��������H2��3��۬z����6M�������Ag��o;��ʣ�S-?M�~��q���'�$�V�I�3{*O�4��?��]�ۿ���_���zb��3Z���<��h;��tO{"{Gm_tH{�m�A'�{-]б���9R@kY��+xq����+��s7u½ԣY\���S0�}���8�q`��a�����������������Q��v�H9	F�s-t�k���������QU"��	�m��(z��{��A�E���P��T��]7�5MW��˼�o
ӄBJά���"ǭ��¦��#�O^9�c��-����<ᇩ�\&��c���ά�5��W���{Q#ˤ�;0f���5���E�RHz�`��������J���c/�%����`z���RF<;4���3�N'�>�C��-w��������3�i�@�s�?�|����r�������6�����K�#0B�8����g{
��6�^�/{�2/_D'T
]9�;��f�;5�f��	��\:Nq;�F� F!��bCG����0uD,  @߿���VS���UEN�u�sr�S�]�ĥ:C�	x�P���J젼���"e��s���<͜4��3"[��4��hR��Q��L��nS�I��~jܦ�^{��Ń��M8��/�LaX\MqV�%�4P·dOs2�Q^#^������'�-RШJר��;��k�q��y{���Q\��.I�������NY�3���	�\�`B��}��rw�>g��a�~���?���/�����_����T��Q��_Ж����,F�u`��[f�v2��u���װ����S2L�5]�d�@V5Ќ�w:/��S�z4�/0l9��;owd����]�C����V��*� �%�̄�I;�U���隶9�~j����?�m�V���s�o�=��'p,�M#�ĕu�s[�-����"�}�)G/FpN��?�t�q���LC��f��t�)}0�:�mé��n����:� �G���թ�c����t������Yu��J�@�SP.�+6ƈ��L�Nm�S� �ئ����>S��TL����5�dh����K/��ב�Yk�:� ���Ǝ�[$��y�g��O�2[��Sm�ߝ�/�0~�V÷d�ݼj_�?O3�s��ցs�B7G�N^r��Q�pb�<N_�ixe:�/���F�+W��\|��#Eܤm�ֈ['_%_i�#N9b�|�k�D�N�c�}2�M��95v�S�[���:>�⫋O?��❷��{e�j��)�����S@��
6�(������w/ߊB�И��*���k��ɽ'�=�K#v��yx�5z�-���0��2�]���m4�Z��:T�E|�\��$5d�t����f[y�Ch��������!��\�`f���멪��ʨ��t����_�eD�A���	�~J`8������J^0f��s��ɖ\�I[�dg!�$��R�-u2�;�����UXғ�`s��̓�!�.9Nj^\��z��,U7���k�2����F+�)��V�^�$���I��|eģNT�y����~Q�o����'F��G���16bv��|�Ȉ%���ѣϾ�����/>}�u#�.�y�q���E�FW�͈�ehg�Lk0|wb�.�P�~�W�C�G}�] 1j ��Iu�0.w�L�p>��N7�ǿ��⃿��{��qZy�)Y�����`�Ǟ��v����u��S�����B���mKCt��'����6:�驎��\�U��xi5����#�F�5l?����������㴙*�MO:�:r�6:�����ӝ˥���_�
�a�t����9'��L !g�s�'v�R&a���|�E/���G�X�v�H��!m;_F�����}����y��ì�"S�`�e��W�,Srlc?N99.x`n=��<\#���OoM���$��>��.�*���Ot%�7�7��ĳ��8y^�{Wi#O2��������i�8b���[���״��6���Գ[�I�s�ݿgyO���87�9��^=�*tO��S9�����ؿ�|חX҆]߻���<#��{��j�U~צ�l� �"����8���l�t��2�݋M���ڎ�ZS����Z��;m)�[����]m<��N>}c���8{��<d4���K�c�Dԍ�c˺��p�e�)8нjy���mf��?h��Ma�����D2�#ۤ��ᣯ�|�ٗ~����~�OQW���^{����/�]�yĻ
���N�_f}vz����$c�{�?c<���oB�+�H:ސx}��}���i.��ef�!��w��#�d���ׯ�dd�et��Uh�Ы���F6��a���`N6�]Z .���7���A�3�v䋀/�����S�ܭ
Ie-��?���0:�;q�t�M)7=��;	Ҏac)n�u����)|cNj��9��㠄�U�Q ����l
�F�w(YD��F.�������7�}%Sr��ƶу��17���n��K���)���1p�}FO�Z9�����-I; �#��b�(��a���P��	P���NÞD�[��[��5��,�Y��|������&����1���t��U*�Kٙ����T��t��<�v��(N�+��3P
- ��ҶTG�lG%��RS����q�>OB[������	���3����U�{��ܖ��s��I�1۝^ <�IX`�*��ܹ+�|-�|^m��C)?�h���'w�?� yЛ�֬q�U�r�4��������N�s�S�J'=3mP�8	���F�xxl�v���AԄ�D�cˡ��g0\�w�y��,�;�u��`���依��m�y���'�&"��`r7F�t4Ǥ���G�6���[��R��-���-u�)�Q��F��c�S��ƫ���<ٶ��}�w�d����ёl#;�U���o�ӟ�',[Ud��6�a�dW���D���> &G	C�:mb�?�	�|�r���L[m�i�ͽ�����=�[�����W�+��/�/)FB�6:4c/�l�����kϪP_�f�l���t�8�pi���9&h�7K�� ���7<�����Q�|��R>x�f�s�0|f-��PV�Hv�t$m�����Dg�_�m煐$<Ljt]�:`y��*e�ِ�*gg��G��<�.��>�D��[Y�o*O�=��K2�瘇����,n �naG���Lt"��$����?F���\=�ґ�޹���>�R��|�vh�8X��E�ė�s\�n�I,s���Q
��Hm��9�� ,)J2q)&�>i�JX����Q�Y�	>
T��J �0���b�N�N�0�=��>OJ3�W���粼-��L�ɵ)f~v�;Q��Q�����d�l,^Ȳ��@V�<�>�'fX��U�g��F΅��`��� ��Ay�5|��4��Ėc���y�}�z^9�F!e:j峯�����W��i��MS���N����z��?����2rf.�v��.F'�G���?5����5�6�𾎫���*HE��/0tÓ��αr7r+O�2F�TT#u�d|���,<�<�2�K�N��0:r��e]���O~N����8X.xӺ�邴�k���f�S��+�fT=Фy%l��N(�+o+P��Mw�=�)�hB�����{�M�K{����7�a��F�ΰS�^��k�&Ӿo9�
��s�l�����Xd�\E�u¿Ail�	��]h�r�8ތ#�Ck~�i������zX2z�'���)j�}��;�xGlÆ�7�?z�&ɬ���5N+Ӈ�\��~T,���lآ�U����垚 �^:0�S��Lޢ�]��  @ IDAT��/e����������|�_�O#�t�z8ve;�3��F?�w!z�����M�h��'���(v��㭝���A�i�����|=�rz<|~�5K��AwD�K�[��hb�2L"� �y�I����Y]�˹��d��^����wF9j�vG=jS"HS�1�}��|酵����{�3*l�IF�8A/2r�%\�1ps�eU/7��
v:��%�cF�9;�TήoŁn=Cu�n��tU���6*tD
;����?�:G�D���2��u�)�8\)\~�{�%4f��J��|��ڇ�_(o�[��Ŏ���w���&����W�:�ʠĕ��8`̽����ҥ:pਕK�S�{r(q¢}i/y����چQ�Pj�ڎZ|����9�(���HTT~��g���%��k��u�&~:ò;Q�pPP��C��<�p����4q��v/����n�Oʠ��
agm����]�r#7�(�8_�5~	r�0��f��^~�ϮDL�z�~����xW~�*��������'jȣI� ���`�1[�Jx�7��D��'��+�3��5_i�/�9��	�kj!�=�|y�.�]�K����������-=�1�޺�>x��A?ʎ�U�8Kz��1T�$�8��gy\����[��0��@vF/b4�d�r�SU�H��}����BVv�k��r��jt���p����&�u�^�g�(>:7��*4���$�8���3��(�Z'X��.���^�s�+��MJ�/|��{~v�fمs�a���o��S�C�f��^U����u�"�~�=xE�ʩ�īv��1��)������sHb������#.){�X�k���փ#�rd�~2��t��Y�@B��g��iI���G.�~�nw{$EY����������R�C�9�c��Qܻy#r?����5����n�&���pr��x�з��x���)�����ƜF�3���)�ϳ�̗��FƝr��8Y3�2�
/��{n�.#aY+�^�w}�O�����J\���y����ŵ�|��O�|Z��/u{>�`PÁq�S~s����۵]�3�S�r��r��+5: x���D'/�C��\ӝ�ϲV�y��ϲ��LC~��W�gj>6����,��Wܾ�89^f���Og�^F^�h��N��x@�>'���a��䘶a=t����`��9�>ӆ��~,���u��rAEs��n�.SI��+�G��"��,<s��:�F>��t�d/ )JCd�$�,C�dotSs՜���LSpJ���?'or<ʑ\�6L�������y��(�Ґ2[ǰp9!���]�,�q�h�͹�)�hŰاu�7��谿L���HM9ۿe�b�O��`��Ο��sA��WZr���>_��`L�IQVc��OV��x>Ot���t���3�>y�"�<�Ũ�r�^�c�C�q�f�~F��Y'�j2b��QdS�O�<ɓc�zq;OY�0Ӕ��i  ���R�P��r�=6���Ou�<h��촟r.�O�}�?:᭗hgG�>�t�Q0<�?G�h��/.C$�w�����v��4�v���7��0�¿3l�t����)�O����I���2p22&����xR&��ӱ0����o���CΡ�1,�UW>�c�F���p�N�I��bo��;�6�Fߓy;$[����)>�u��f�`�m�׻��jt��In�;���|�j���XѤ^��h�gz�����E$Y��z��_�X�*�rt ����ܣ#tlx$~�v��w{�x����t�5Z�_ֱ^�S2�oD�eFO���)�����m��S�p�v��kDY������.��d��,� }ֶ���o.��_�5{���m~���D�����������mr��J��њ	��+|���'Y?��7@_�n���'����	�(��(�};`/>�w�`{g���Y3+��2�E��B�,��FD�J�������{N�,�&lGj
�~�l~���z"��7����Web?_��3#������Ͽ���W��]�����k��_�.gшS�c�J�B�7��ӏ�~q7N�[��6�O֓�:n?1]�B�ɬ�� r���F���E8zO�f}�矶�G����M�,��]%O7�U�r8����Q�KtE Y^����{�!5}q�( 0�Y�h�P4{ULd�n�&��ޝ2&R<X���a���9�<E�]�5���ZZ����yu��y�)�Rj �	q�b���bQD\�#��o�O���.�.��|�z��9���^Q9�a=���<�hR�m���h��Ʒq�)��ҫ��7�����0������>1OpF�,ַ�"{o;r.�l�(���u�J���/�,2�\���13d�,��ߎ���a�ɰ%?����9�v�
o�Qpr�8ё��?��c���~Թu��u"x�Z^P�_��3�od�ǹթn��M�U�tj��\�Vz�r��Q|�_EO�g%L��[��Í�\κ�q����"?�Ӓ	��3���i��[�2FF6=�l�6~�Ӿ��_��Pc��g�8�.Y��U�W�|�0��^�瀢���en��eV� 9F<�[�#��p<�;=:�"�F�N#^-7Q_;�Նw�`�c`L�#�ԫW�p�v��\a`�>$n�*L}S��]�)��?������-U�؍ڑt���1^p����m7�#O��� �s�`�+����zC��a��Z�EP�w��Ǐ.��w�����zf��(��	����kI�����Y���z#�[�<���8'W�m]l~����7i���`�)uHs~!_�,���m��)=�h�#6Y�}�ȽrHEv����sv��@����,b�.�&Mƽ�XR�l�K�Fh<����L�X�d�(CVB�?���I���7/.�3SՏ߿x��7z��0�^�ʧ�23�e�JKa2���3ڵZ�5ݦ�"ٔ�xk0sD	�9�q=�̌����'O�������<��s~���h3B����I"G��GR4>L`�;����f��e���*��n�rP��F���qf�ʸsO�ƨ�݄�s_#�7��k,���"E������T"��Sb6��'�p�n�4�%X��F���w�
a�c��d�a����{8�7��9��,թ��D�D�7�+cQ�Q��U�l��	�F��}�)eZ뷫�:�S�m�R���Ea5|o(=��y�[_|e�U����#8�t�mw���'�N+4C�)�k�F�����5�?��Ȩ�7X5O���>��#C��:q���Q4��'�d
����j�������e�78	ŧW<�ڻf���a*^��=��"7�=�t�p]h�����v��{U8�N�kt��	�7�@��Dt����ؓd���w���t!�f���t�#=7����q�>NJ�#-�
��<<��~x�1t7�{ �ί���4=|*�r�H��.۬4�����v�J��Ψ��%PǞ�������m;��~ח��S~ip���ְh��o��rژ�9��4�̬UH�C�>T%��r�~�ܦ����xa�ۛ����=O=퓗V��Ӻf�D�_�K�$�|�x�Է���Nf���!�h����w㠽�5o�\�-_:�ӟ�v���-��������..�aF��V>u�#e���u�Az�L�y�3��<Sr�;j�ujF���.s�^����z��OQ�I�z7}��x���Ds_f���v����] O������[xXW���$2:aQ�Y":�W����!���\}���v��ރ�B�U��� ��ܹ����6X�	&V9 ������ٶ%t�����_^���?e��ϲ���޼''�Q3��~]��O��Fw=_�8�>���� Γ�=��f�L�3�v�%���ʙM<q�7�a�`�/���=����C˭8��,�G���� p!���tw���k��IC]G��G�8_��;����\��+��W��T��o���|�[�� ����"@�).(9X#C��J�A�ٯE�l|ñ�ϐ伲!�Q;�}���Z�F�=��5 .�Kq�N�tYUx��]�V�� )=�z��̹0Ro�Qk@e�6�S1i(iI�`��j>S�.:
ߑ�E��ڬ1�����`٢�8_i4ޜ�T�{��Z�ȇB�лV$X�`���Ŕ1Leн�Yg6O�ɦ�{��L�[j#����8��;-z��:��
�t^�!���#_C��_Ӧ�9ԭ��gS�~����o�T��m��ħ��rux��Q����=�z��N��=����fo�I� �N�+~�D&���\��A}pT����@gs��V�������Ĕ�aӲ��Ǵ�_p���T�!�f��K�8�����j�g�a!���Q(�m��5�������3��9��S���-#}D7rf?+�f�n�v[�z�e4����0�`ôY�N��4b��զ����&��n�' u�l�o������6�N�h�/]�ɥ�����=ȈG��ü�ə��������z9��qz��}��;9��Q�����˼%�W�֛����}2�x;o
�U��8ai��f�i�u�r��>��rџ���D4.JiP$}.��a��#�e���s��k̛�m�$�@L��DF�C�A��:��i��|���	{?k$�\��Ѱ�{���}׼�e*Vlz����2oRr^-�����Ҩ�.}Pf�Hf]���'Y&�7�=��l���;J����Хy�u-��Dآq�1�vt��Y���F�=_>�[����~"���T�:����$G+�h��04F��E0F�۷
�
g4�g�Z=� ���e
T�$�ty��4ǭ˯/��_~����.d��`ӊ�g8Iz�YѭC��;4�*A�D7�a��ly��I-Ը�M�O��Eo�m��&~�"'b��*�	R(�:z�<I�(��ki�\�'0��,ͅ6�8sfg������se���o��q�J���o��b}o�
}�ROF�(�'�����ʓR戾�)þa}*<�]〧���xANx�S�NG�۹�̟0����?�w��4#}��<dX�C�cw`�£�Q%��,N�|n��quBo`�6S~vǻ�J�7�S��z�8r���X\:����!TfF��9�W�54��zܨ6
_؋G�	j��E���q�Ǥ|�U�[}������v~e8�ih�b���x��ڱ�x�#=�V�OYF���O恴�,W}�O~4�R��+������%�����ND��5x�9�[I*8��6*N�~	M���tj�̱��~i��u�v�rMfmG�Ǒ��t�.j?�g����ͥzspv��Œ��ٜ�(ESW��K�A�VF��y7��d  �R��t�����+�T����=��׿��S�V׃}�Q�`P���H;�>lJ��	��`3���G���I3��sB��<�T����E�!��S����QK�rΨun�ƦOI��H����/m�'##g�W2������F'�G���j�C��b8�Gsd�oz�ؑ̈|���ſ��O����_���e���\�%�4����^�ּ��Y�'y��i����Çu���z��܏�LI�4{���,�w��mT�=���u�3?����D��G$ʋ�B��I���:����s���g���<뤽�f�����|�m|�C �o�����G �M��a>ӌ�����ax�F��|��ē���tu,�h=��Iw�{�0�<�Y$�(���R�>D΁�t��9�W�H�A��1�t���:RS���#\CK1��!xU08����(nι��u�
�O����3/N0С���"�gW0�U��WJP#�띮*�JiD{�]���<�o�v���l��'={�yU�����dq�b�~0_�w��Ȟ@o����?����f��}��G�w}�	'�C�`�N!t�%-=ç��)�Ϻ�p�Q��Q�۸��F�ǉ9�1<^���E����o�L�?4O]��=�/�;~�<��7��W�q�б�Lma@���A��X�-���k�w2N�qq.:;� }*�*�3H�=lb��ĕ��W�HS��)���-7%���~�p�w���h���;�=F�*����u���nTc��y����M&�at��^0�w.����X%��#����+��	N��F;i6! ��۹W�� �ڣ��]t��Eg:�/"�l���ld~�yh�ū;
o�̶�H��[�e܋(�H���g�z/���c`�	{n�P�H� �4ޏm{�q7����O�,�ľ��^_��������3&��ޑNU&���K#>�?����1������R����5������32/>�	|ݪ��]���ճ���.y8����o���p�g&���F�嫾.��e^�J��>M��8"O�V�/�08߾x3ts�^�+���
d�a*��܋<�?�ڭgYs��g�׬�đ2X�/����Tf,y�e7�����^��^��?�a�ѽؗ;tM��K��']��z�;�MF���&e^f��g�e����C;b�Y�<����yx�t��"��T%���l���d��*o.�D~e��uT�
��UB���(�X©֍��
q���ޛػ�7}���k�3��V7��ŊaO�	�Ʃ�BF�9��<�pҌ̍Sh7w��0#�"����8���|�/)M�H��'�:F�*�j��9�/n��7o�ڱ����sC<��ꘞkJW�Z:8�;�<O7S?��V�l)�I��'2ß(��,�k�'DJ={��'̚1�v��Ȃzڢ#��l���.��w�����u4���������=�y��~yk�柞�q�18{w�x�#���̐����h:�1%x�wn��B��-��@e�m�
+���o�����OƦ�x�8v8ֱ���[V�}�@���K��t��s�*�;S:�Cyj2�����=����5u�͠�+���$�H|[���u������@z��|
�i�=H�"��*�&���<�3���X?�P)��hΡ^���C�\����|g�O�鐧��tX�����G�ʷj���i�p������o� �����8X�d(	��s~V�?��q���<L�8g_�;�r�,1�a��VΔ��p,�[�{������C������G����&�n2��摮O��U`y{�v�⻛��f~�e	[�/��0t��3�S��[�gf�2�54��,���6"r�C��Q�m�3��.�0������#�s$�ȩ��U>wxW]���ڧ��HVw1H��2�vյp�U��gq�>��\��D�����w�u�7��m������w��:�|Y�s��eJ�Y����)����:/�����[o��-Eg` �J�|�ʙ����J*Y��҇yH?�ud�~s�,ui��3�I��e��^gWW�!�f��|�q*��yPz�񯺾��66��Q�;��(kC�PZr=��W�څjl'XΌ2�j1���)5.#�~C	q!�	H�l��!�n�MÏ�؍@�$m�'��}���ҩs
,��p>�)h�LM	��_�@"L��c��R-�uq`
�|����9!�u B��-UTI��4��< �������G�.<&O����I;=�:���غ�\���N��}�R�	:�r�`�&�kG��o���g�[�O1:]�ris�3*�d:��T�#�,����/i8ofh6�~�A�c���)Z����a�Kˀ:�Wi
4�.vď>/rW�ᕛ�a'������I��t4g>�|���;�&I�<�|���]���,Ƥ� (\p�����Ld�'�m��A��VA�jxhc�v�5&1 ?85�z��ħ�(t#܌9gi�]d�A)��נ\��v��n+��������|��EۖN���H�h�;�;-�	H��:�F��,���*�J� Z��m΂�Һ�ˣ��,�s�2y�a����3� ��V�S���s�AT�`����9��<:Be'ǔ����[O謋-�qд�Rw
���u��d��3��P�][:8W�{{�j���t����O2�����ST`����I�1�]�E��O��>�#�d^q������-R9�����N{�f��ζ/n��h�R��f�݇}q6�����N��Wߖ��0�l ��T�w5�0W�"�3o#Zp�e��`������8F��}N|��?���� ����^������9(�����O�e&̧�F��HK�y��ip�V�#>菼�p?;��k/d�:�:�G�}}�1Nm�638}DGO�fׂ��������ٝ\3�R#��3�`��y>�n��<�|�Q��x�_�y�6���L�3�ڑ�L7N���.l�;ľ|AQ(O�GN�2ea.BN��+��3m�e1(Q�P���|B����~��G������)�7�x#��ݝ�}0�s�)����O���@�t}�ӮQ;8�X��rKD!�E� 8�d�A�C����C�PB�=;^��A�JYno�*}��ʿ2��;Z�:��H��܀$~%R&�$0 =ڑ���7tL18OP��'�4�QM�4�=���9o��b���Z�F��=��� C��7���_~�����կ�u��`�� @c��sN�]{����$A�i+g��SNp��	�����).���t���j\2�,��t�I�v͡�Y���G��gM����nN�8��T;Q�L�TY���iZ�o�u�T5ͻ���x5? �Pn��f-�|�o�0񓇼�7��i;� �'��N��RC����J�!r�}��Z��Z����J|Ćp��RǴ��4r�V�=��O����L��L]K8�3tcd��@��D��f�L�lT9W�[:��lG��,u��"�f����o����#èҤ;%lu�p�}ۇ�+�ؐ�k��m��g_&�I�n>#j��bg�z;(ڰ�I��M�m���G����e��L�Q�$����sxZC���)�M��w�~��]�6��L���ë֯M��y��2S-Y�U{Z� @:LWw���m"��}�z.���-���J����K�����^'O�����r���lu�۬�%��k2���V����%N<�T�f��͹�&lS�?�����\MC~����߹�(�f-��z?�j��#�����?����ʖy������g�<�(���ٳ7�C�)Ǭ�|�&���~�%}"��=�|�6C�J\��n<ڴN�����pw'���d�Lq��w��q��`������}!���j#�?T�2�z�Iv��X�e�I޽)��X�,���G ���<����%�۠o��d�~R��� ���w���3|���WiE���s���p�p�4Nس���,V�#z�.�(ګlְA�SANP��Vo+�$r�(��#�k�0䚋�*��������a�z�z^�&fb���9I���qf�%]�a�� Î��� c��9����-�F�'��ů^�p��e�����|�9{o����p��m��� M�N*�q�����h�?9l�l������<��Ae��i���c܆!M��ͷ�6��WB�Q�zh9a�7G��Ox�.���2T��5B���[C 4X��On�dRS�TD%�a���
f`4@����ʜ����? �֭��c�]���|
���˟_q�}��R����\��z�����o7(�Tg`��sT�ڱ�m��EA�ϒ����S*i�����#w-�]�t�V�h��MDB��#�յ�2�x�훗�B���OQ�����c���Z���3|�x	�@N	ڸ9K3U�롬�ѫ*�����7k���t7�L��і��T]��y�����u�S��%k�L&�$�}�+bg�r����؁ ք`� �7���Bnt������@��w�j��<�qf�7���q�K]y�z�A9����jOyD�x����Q�;e�����Y{���Xu�<��zs3M�M]��0@��bI����"�֏�j��	�լ��p��U�y
6��Jzf`}<�ƳWN�6�6�n�A׺�!�S��x��!N�7���>���t�p~�m(�/�N����6��u�ì��f<�m�;��G�G���ҏrI[���S<4�px6?�y�=>��#J�T~��e��̵w��,z���"�u�$.�y�Xx�r(c:�^�偓3�0`��у������Kf�@�x}N	)������L:G�8��=��(���/����cY͑rK���ǡeP�S�{|��@����{΂�:|�ퟣx+a%ﮮ�����ӕN7�-��Өå33B��W���:u%dD^{muG�Y�8��y-#���f�0Y{c1�0©�;��6�A�)"��l��G�B�m���Aޡ�3%�z�2�5��ԟ��tpt���~=l���I%�����w�ܢ�|x��ï�#���x³�G�.}gɾ�@>�u�06q�x��w�yg�c$3�/M��C�Gϱ��/���:��y���-ؼ���c�=M�ε���wc�nڤ'y�Z�m��V�uD=䦨w|Ұ����ki8KZ[��՝��)�qi�vL�+����O��0j~k�#(�8<�H>���G�]S�~����蔇����m�7/��"y0����٦�L�_T��}����i��m[�����l<�u,��z�C�?(�2�u�!WN�Mz7�\������ʪ|���pE��o�v��5���ϐ���F�E����ђS�^��q#<��t�r�-��8��y�=O]�5� ��qo¬��,�6(����+fk���������(�!;�?d1�Kgo�:�
��2�8�.������34�}�����%�٭,�љ���E�AY태���P���;	a}��϶*�oP�;�2}��>���)	:���I���G�Q��3#D�����5}f}�� �	c��~�݄�	$W�=�r��C�Z��sV���������&���Bw9��6��__2�s�Sq6���)�<�<���)������Dk������f;l��/Z���(r-��+ɣ�<��}���t����	��|���F=�G����n�������q��=��z��T"rr����takyr������CPJ*[�7�R8-^I����RM���D9~N1��нqz3���E��<�[�٠�ׁ\E�4\SUv���6S�.�s��΢�_�}{�i�����r����@���Ό�g�t~��i�^FP���y��z
��U�9��oc���dJIo���^Sre��[E�^u���L��aڈ�e�Ԉ�d{h~N���Ǉ_�q�7bݨ�7C|�V�ũ�\���>lF�$h�o������?4�"E
�4��R��(]�tg��>l䭙�U��鵿���S�*�R�!�È��!Mu��Շw�_X�#)��p�86����X�g�a�a�h�%�Eۆ3gމ�i_���Cg�8����
��2CJ%��&��ѫ8�bX��9����˔��Ԇ�wL�mrg��q�FHsா��'��I���P{1f��+y5�6�,gz�J{d{Ýt-�_[��:�Xu��4�7���(�П�F���b񏮶�T�+�\��8}�O�?�\�s��OC벽Ug�l�\+|t�vi[�f^�E'�o}�ȵ���S�ԧ���-ƫ���c<t��wyLv���OX8�8�-e,��1��?�㖪B�X��q���̎I/�AqT�[mƒ��ugc� ��7����uތ�:�����	��9�Dv�A�I
��W���Ti����j�[�y���E(*���%�H�0����*m��	���%�O�DУ8��p�\����mf���ɧ�⌹�H5�g���)�|"��q�Ёl����`���]�d"#��CRj3�8��e ��88y§�pA�"T��Pྊܶ�|?���?�t?c�;��K=����,�>ᵫ��ub�
�o�nʵ<7�"s �N�j>�/��H���`���@HP�0͹�{�(���V^o�A���
��>W��[y�>�k��c9g!�N�3-��� "�LT��%�鐤Q�4?`���$�ɫ�4 �������q����S�6p�g&���_���h� \� �<��2�Y�+l.����)X�8�T:��3���=�D-#vi��bf��Q=w� F~줣%�nSG�~�!�DH�A���t�_�g$ﰖ�֭;AG�� �E_R�����:Au�\m'.�jz�a����Ri��!E����˸:M����k���xl0�FS��l:M�Ou�Ntt,�έ�κ�QGgtYS���-2oB����π/~;�7��t��,];m��>6 �����a��3�|p/|	'��s�Sft��t0H#z0��7Ǆ��\�9�s�gaB�����or`R��[�N�9O�AP��O��>d��6�3A��t�SN�zX�p���jQ?�ˑ�<�9>ֱ6Xl�'*��7�3�a�J=Ԇ��M�k�f5p�����Aڑ��V�֝�k�ħ]j;-rL����r��Z����#���L�_�JE!�_q�%]���8@WnW�����ik^{�?ǻ�쐧M��gϨ˫/���ۙ��M$�t~�?�n�b\�-ۮop��x�;�n��G���l8�-|h��^Y�\��_`G���M8A�n>���(��K �d].��xRAd��D����¯�\~�ۖ��Y̯� ��x�Ro.;2�O��*X(��9��@xI��2ͯ=��|�1��i���rˉ�;��c��K=#�y{���޻�xK�ç��vF>��=�u�%���މ��l#���&ބ��\��"�>:�"<[��Ҁi�\��{ׁ$X��k��V2v�n�y����߼J�tv�kt} @�r�6V��B�=ci��u��3� �.O|T�W��]�����w�����%��2�4�Vx�CgR�Yz�hO+��휼��Yu�"*�穾!�J�$��Y�%��<^o֚$��䣕#.	ֈMo�Ζ�Ge5BR7x���)i�g���!ce�0+?�,e}��ʴ��d,�XTB�����d_�Vq&��� c`�d�q�Zt�aCz��ܺ&��>�������H�v�3_��}N�ϒ:v�n��':/��?;6_A���S,i(ύ�ϑ/��O��X4$;����FO����Q����hG���k��(�1}f�L7-�KO����il��s�uѳX��A�Gu��M;B���x'��k�֙N���o.�7����|9�����{�n�u,m���]��#��^�G�R�)�i���S�as���e"d'/G�q?K�Ε%MC�V�8F���8��E�%���:�~����{���be�QW�� �q�j{�p��~���p��:�欅�4��=ge<L6�M��z��O�=�t�3xs`|����_a�s��l8����2��d\H�s�L:����/�7�!��q�����V>�s;���eE�q����T"5���0T�6��d=�� =KxBG�u#� �0���B}�c^���VG�βe,*�൚���{ۛm��>u�}���>6�TF��/hr�0��>�k97���m:`�<�r`��v#�7޶ooU�6������g,�ȓ��?�M�G,;z�}��s��>��y���M啚��m�I�V0-�ڣl�CPG����W�,�̳�5��g=T�E���n����\(;/�y�ح[g,�������������݌֗/Ə8y�ۆ����2��^��*S�p�޻�>�ɇL�2s���������4�j	�`�0j�El(�)�eԘT��Q�јe�� R�2lu�0�i��a:y�<{8i���s�JU9H�����a݄r�0OJ����z���f�N���IH��|p� ��=�{��̑I�M"A�Gv�w~ԣ�9��| �!�������T�z%��g�qa���X�Ǻ�w���������l'��
�c�|o�ׅ�w��u,'�R����af����QB�����L��_<)�ԧ����nt�Ȱ�g����es�ý�<�6ȣ0�G���>v��Ӥ��+ڃ��n�`�n���4f�j�t�t��e��P�d�61��w�����][�D�E����u�����χ���e�|���yW�lK./�G�(S�UgFbqs��r�b��_ʞ��E{F�Z�לA}����<��q�$�Y�.�pSH�<ܻw�ْ燯����i��&�t�]]O9���	�H2�{{����8?��k��~�uVy��؜70�U�hp����=v&�4Ü��ô�Lӆǎ�3�l:�Q�L���L�����<B`���7�$���=�x��|�#7|���q|��p�o�8�6�����g�ܔ�;��p4��N�*3O��:��P��[ P�i��,�g!�]vȿ��@� ���[:b�f�c���OU�c8�ӎ��2��'��?�̓.3�뼍x�/U�g���-�9��zl��!�y|h)��[\[�7�3���<�ki�KG�(��U_q�ر� �>�ͷIw�/i:�%��`!_�9׿����|���?��e}���oI�������2�����6�65�w��^ԩB��0f���8)���j�C��g�k����c�K����<�\~p������g�lOq�I's\ʄ�'/^>g��c�@y��'���	�O!*ɯ�sV�z�*X��OB2�)a<#g���[���8`P�����JS95#|i�`Gh"%��YVTV�{
]n�[x�����|�L9��k;6�l��P�ȍI�����ҘCP�"�")�|S�ⷼ�1��᠉�CKr��R���a��sL�8�P6����)��z���3���GL�x�ݻ�w���ǐ�y��9U���<��,�R�w�͵i=c:񡯋�z�|Ķ|�%�q�-.?�A���P�/��P�7RϝI��{�g(��X˷�F^�n�'���Hn��t��:�/_�y�1Ë�tm��L����i�>JQ���)S����x��)�x�W�Y8̣�;�x��~��߲���<J�4NETP��U��꿶6�������C۰G�c�n	�a��z�%��q�㴷�[�ɚ2�'��2$Skǌ���Y7~��Y�O?�$��3�/G�M�{Y/m?�[��<-�E�u.���ޙKg�W:~�1�p�*5�4����]G�Lz�8�ceW��_�kjt{���&���mz-]�o0�����̐
&���B��Ńr�YA_� �����W>�8�1@;���-D��ѯg�.� �=.-�l�W�Y���~��Q�M�����]?���6��ط�x���o�2�`S�1��1YZ:h���<�@���~�uz]v��ԟ�����[TV�ύ�r��_}1 O	%�����`�IW�*����,�V/��k�U�*����k�	��o�4[���~���]e�Ы��:oA��I��˒��q��zй�U��4jPT�Љ.I��؂�M�J#lm"6|�=)����9����>��q�E�8�\h����:�)�Q��H�qC���|��xM#{���Z~6�)׼��q轻�:��6.��ܟ	+n�T�C���1΅	[���t��AG���*fM�\��1sI
�m7�S*X+ Nn���_����`��.��k�;Tx+�����2��7�@p#H�d-�+٣ׂ� 3�=+�0�t��^ZP�+�$�Q��ja˳87���Q��6����	b`�y&��?x��>�Oِ�5��q���}��8�Bt�5a�vj�ε�(�J��X�>�	�ԥ��#�o��!��]�4d������|��G��������������`�Ҧ��+u�3���V��=+��nrp{�x2��\�S�P��-O�v����Ӱ��l��Yx?�6���G>��ׇO>�$����Hshϔ���^8��z�n�"c�V�1?�)N���	�
�I�����g$���3�o�/�#��W>�\_(����U�`���/�����o����\Bmw��k(F��}��e�Fq�r�y|�N�\ϭs��Eg�o��(WU�Oq:���zm����vb���ҷo�	�g5|�k�yNY��0�_�n`��ʚ���X�%�h�=�1��h�4ۮ��2���j��y�㭒��P  @ IDAT�����I6�7��n���u��mm_�α/ҝ���߾"4� /��ֶ��T��c�6@�O{��b�?e�&̸(�g 3�vpB�?S )PoҴj���/���}Q^ӷ܄nlM9"omKn�%���7{n���5k���Ҩ�۸��Ӣ/���^ab�ang�`;�!QmQa�q&��l��Ϝ����̣v��׊^�<�G��f�AR��Е����ȅ2�GC���#4�-�'������!�K�Q9�/��W�����ㄳ��q���ܺ��u�=t�:��ߚ�9����1_����bA=~��D%ZEc\Y$3��ICO�7(u%�	b+�
-�`��0J%kx�VA�T��Ma�e	�\�m sH߸?���IVi�>aL�R<���8'�i��Ż��ꭋ�c%���re7��� d^���lL!$���ƽ�!8�=�rL����+n���|raRx0g�+�o��޻���¼�C����;��N���y$���pq85k'"�`���� �r���O��.p&����'�o8/ݮ���1��;���[>�[�:c֑��\$�8a{#/��7���q������"g�|�1x�0�u��(#�����"���)N���)_��Q���_�������?&�]f;z�.?�=zϛ�Ge���-MT>�)@lh%����;��ܜ�;���.Ǖ�c�/����z��'�m`�3�s���8�9z��q��}�0�%�	C�L�O]�1�I�jC��q#�s�E�L�<�He��� �3�=��̆*��z����Gf���t���-bj)�pxZ�ʅ#0�B�~�e����,�#M��n�c�)�}�y��:q�^�?���nm��R�)�p�q����Wg�[/��a�@k�<{�_$��X�i7��28�Tn���V��8�i���%��A���T�[u������a-��-��tĳ�&}�mZ�gtNy���͜3^�1M�o�Dd��џê�Յx��tg���V���Dq0���u_��\���t0g8k��6c?�s��tV��a4���׈�:�"�g�r��ǿ��O]�\��j�fX���]�NX�^��Bgӗ'�^��C��p�|zQ[��@�b�xe�e�;�6��?���ᔯ��U�"Ry��O�sp������T���
0FC46 4�a�
Cǀ2�bd)��5��_��� ����s��U&DQ���3���[����-}�	�yF���y_��<���0Mwt�۪���s�]�*rly+�`�)-�9Q�*nu3�+\qu �=oC|\�0�B�-�B΂A*4�;^c��A��Ct����������-7b��F>�z����W�~���᫯����'���p�ǖ�q�p��`���#��5-ߋN�z�P��b�y����\)x���aQ�fFƲ��wԖ�0�vP�7�#�ݦ��`n����'�|Y��V��ϵq;Yub[p���k��7"��b���>&��ީ;s�az�°O�ޑ����]s���}�^�{mG-o3��g�([eT�K}��	���/�<����<ps-��͛���|ӧ�:�$���n��&� ��4���֡U����o���f�ěP>ȵ�����{��s.L�\��c�<���/i�_��|�Jz�*�8�K;�7�����a,y�s䷌�γ����d�I�d �F�'Oq�����Ų�[~��E�B��Aޕ_@�P���P����f�:̪[�qr���cZ�2�L�_Ñ�3Ao� ���_���7e��m�D��o�?�ǉ���b%aG记�?�x"��C���P�q6���ڙ�yq��8��J�K�3_:�]��)�N~�m�:�,�é���:�R��T-cb�����ܭ��Z���O�"�n)�Q쬑S���o��}�N��?'L�8ۧ�㞓R��L1�x�ڽؖ����$`�76'��=�W�F^�Lڈ�����זKE�άg_
t�=��+�(���T~�5n�����љS��wx��+7S�8�܁q_���H�%^��+±ǳ׼�pv���*��|���JL�쟇i�=+�*�EXQ6���|���D�1����8t�����i��Ŭ�~4�K�x�)�9�(�z�������ef��������6�{�N�(0�)Ж�ܦ91x��<$q��?������x��Փ86g`Bv�]�;��L�"4�.��B�x`���p%��xg��wx\u�&F��6�<�wMQV�1K� ����[�=�����g��a%���o�a]NǉY<[O]�_�6Q���`j�:���>\��T�����W|��q;@V�aO��7?��� �4�3��m���=�t�)�~�Oq���\q�\�P�Kg�N���V�:b��e�g���4�!�W-$:1^�W4��S��p�%u����I��سe��a�
�����]�[����A����?g�'�<{h�UU����q�qv��������Y�lz�}g�t����5�~q$N�g�3޾�Ŏg<�t��Z2��}��G���yMg��a���s�:Q��ZGi�M�GƑ]�yk{(L�<ˎ.,�	+k�ؖ�4.��<�n��*����F���7��.��B~�E	�mz� �X]�#yU�֥m���.3˼�J�{�c�0��:�=�)�Z'�q��RfJ<e��g:��	�����
r8��Y�їU���7�ӵ�ȱg&_��}�/6E/8������C�N��W�0g�ɩ��-����f- )h;�Dw�/Q'�t���|lӗ~^�C�:��R���ͺ1�#��̡L��I>�IR��r196�CDx��e����t�1ُ���_����_�|�Q���������+W��ZN��5�Nt��39L4spEA9������C;x��+��:���\:`����}��z�	9�~�ʿ?BxL@T.5�N�����A�&5�j�u����J��*~�����Х�-1ς����[G$.�@}7|�K�
�֯#���,�ؓ�N�rG�qpęCs��a����Q�L�|EHTY�q��K��9.d�|ĕ�bs ?�g|,��e�=�<��/�ĩ��Wg_�&���Ň~��A���C��`p���9w�?��C��o��1k�>��Ǉ�>�����Xxh���8��"�'%p@0h�(^���C���v���p�������s��+o��[��H��O�%@ʌ�e}px'���<�Ϊ>m���N�b�.�7]�#�>"tV˻Xm��]�s�����@�S;Ӂog=�X��~�̘��W���y�3� �9���:��H��2��*�Jޤ��y[��os�t�_Ə3������GE�M`u�Mj+�COå��d}�ݻ�^��>�����⠟~{�9����2K����?yL����=������r��f� �cs=�+ӴI��nϡ��ڵ*0�X>�v�+W�GK'�ʜ�~g��8�#���b�Gۢ�9�}f�D��f>�[J��@?��?�9�v�]tnuh;�����k�7;'�~��3ĎO����$T`o��u�{���/S��<Z������ҳ\�Ⱥ��u���V䱣��Hx��>6�m~+���ˬ�7Tk��`�e�N׋�]Kg�={�G��	"Oe�+r��]�2&-��y2k�\�V'�W�g�'��p�L�)����Hj�b�z�s��U9;���=��6��?t8�wd�s�(�o|۔�Ӵ�5��ȶ�D����3He�^/��8H]>�{J���R����J�/���sT��&��Y��RB���|͋<ts�o�5Sc0�uN�??��0��?b�a�N�3`�=B�4��Ҕ�2�UsN�Cj�Q�NeY	�VQ�
�K��Q�]^ P	��#�,eEKz*�
���N��W�U�L׸u�;8���B7��S�3�q�5p�<z<cF�����iEj��� o5r"W�B��Hi�cA���9�m?V��܎���5�����Eo.�����δ$��sj�+t���՟���G>��C7E|��-O���.�n߽s��7�~������߳��]�G��zgSB!R�R�������ˀ�Wǎm�4Ǻw퍶7Nձޭ������F�YXU�,r���&��g���v�YG ����������Q�g�����D�P�~�>A���Ka�L���l�x�&i3;�P��J��0{`r&A�od�^������pE
/�]��0h�9ח�r-����P�M������ȑi=�� b�<{�r��F��+i���3��93�,�k��9{���͟y���;lw�[	ݿ��ٜGy�)��g��^�^�oB����5��r:��:e|7�Nd�W�w��4yW'K!�!J䞏�����T+4F�#�N���}v#����ÿ�ۿ���o�dy�f��-��̟����+R�e���mHK]M��@&��r�b�R[����m���!+3^�"�U0��#>��o���پ�4i8�pʆ�փ�%k?ḙA�q��о/�d�|����e�	K�2dH9S	��,���3+n�y�X���i��S_��+޺��57��9�W��Wo�h�'�����N����^��1=����>���-�~sL3h����`�Q1�A��Ox,����S���ig'����wϰ�>y�㵗|��)1��_�̒�B�|u���؇��S=��po"�mI^�?GI`&��0	���Jk6��ԫU7�u���ʷ@��]���L��2̌n��/��x�7>	Q:�ũUY���Ȥ��\	r·[�,bJ	 g�^��V/:������R%L�xrM6���H/4)���y�ɔ��<[V���R���Ka��y�u��ԏ� ��^�ؔ
>�J��ⴽ�-����0�����������7iy��}6����6�{�V��{������g6矾��|���@�������]��O>v��_�#^ �ȘH�t����c��s$��[����W'�Mz��}��|;Y;��A���4�������?�?��Yԭ��Nܖ1_�mx��1��i���9��������s�H�C�!�J$a`s�s�8�,^V7�2��c��ƃy���&���oΣ�c��\C{p�YΣ7�S/�8e�1Ή��e;ܞ��6��U2��������K߲��������{�?��۝�^�ہ��w���9jE�wm�<���t��zDfP|Tg}�
�3����<����Ď�'��9w`�Ko]�K>2ˇ�MG�	�W_}u���t�����9�˷~}ܯ�O���m�y�Zw��a�s8O�v�����	�ܙm����>@%m�,, �k>�DIw�Y:��x%jK����c�|�/�W�C�|L?ԾQY���A���t�`�\��.(�WYR�[����'eem���[�����H�[�!��
�^dw- ���cf��Ι]�T�0��IfWW�5Z��U��[�[���ȑ�c?4�3 �0_X/}�ٴ��9ߟL8�S!�V���~NXRsͧ�;�S��L�Nx^ �.�'g�kzl�f拵_��p���p��^(��t�ho�^8U���&��)V2�qy�I�TO���	���
��Z##�DԎHw�R1��G�VaxP��R�b�B�d�I�ʑ�<ŋE�yuZ�8Q\�/-#MԄ� 6_�鶱��PX�z���`_Ε����gx�Q�+��������
��y8�	�1���q���.<�����w��h$t�4fMY��;��g�3`������`�����Q����8�1wV���e�n�툟�)�aT�Q=oˮ�9kࠛ
�v^�C�;��A����0lgl�K����ڐ=�E��}����/�<|�/�,;�B��~&�m��mS�78�s�w���z�J��.\�>Z�4���#C`�M�����3i�i��a�nb)o`���1��8Ѩւ�8`�oy�9��#�);:�y4[�)3�N��V7ܼ��.70�eې_��S6��sp�1���l>���q���<�$�n�Y��}̻�c���l]\3�0���o9�-�J��7"0g�\�ԓ6r�N�Q=\3�
���?e�뫯���cJ�c���u	�o��̷m�Y�萦�踓���9rJit���8F�W�c8�A� ��e4D3�d��+�2��tm�qn՟8թ�g�:yC���4xR���g�q�/��I7�aa�3c�{s���q
*NE�M�z�x�
�r�2���*��+3nQ�T������yD(2��Ϝ��ku�Y���o��u.$c���UoRr����elK��.w�?�łlT��Sfq��\�Θ���u��»�-56�����Щk�^���.V���"D
�d��8!.�{'g��8���oՕAz�5�QrR*�
�`0b�mH�����H�C�Y���� �q̛	N�(7���"�FG�S |<o��4��Hݼ1"�&�j��/���NM�����S�1�r7�)��M���`C�|�]��q��tޗ���
T�0C'�ix�2��뺇��گ[�PLg��u¼Sw�ųg�tq�)ww���_���w�?�1z��GJ���ю%W1�D�FQN��߱�����kو.���
��� �ݙ)��{�,�>�#FM����w:
��ۘ��}�A��×_~�-"�#�����L�� ��C�p�n���T�҂��r�ϔ�2��}��Cvً��ݥ|FGp���Ƕ<�~�5�9��3�"��1t����e��~ʚv!ε�9V�6a��d�)gm��
��+f<�㬊��K�p6须���Z��|��=6��=�}U����ܸ���Z�o���w���!�_ۓF7�ç���g�)��l�m�7��B|LW��F�2r������^DY>D�����=k��g����q�=z�����W����<o����g�P�m�5���r������Bnf�ݞ��������/f<�D�20�aݰuk�X��������]�P?�d��RęQ%w�N�;�&�{-jw�C�p�'IY{$���vm�>NX� o�6�F��eʻ|dV�'H��^�ؔ��-1Y7LiY�	�:R�Z�t9�&h�3�E�)Y�M\���y�^	H�(�8u�vgLR��)�5ȟa�w����`�b1h����)}8|��&iT��R
�8�:�ڃP���K%ع�b=��r`���㉿F����K�f_�F�����/�۱QT�+P֊��6$.=�P8Qd�y��7ĵ}3�R��r�?���@��PA��~	��V�� �)m���&�UD͗B�ϻ�ʻfdY��;�$e�/�ē+e��=
K��2F��1���.��~�N6�e"	�Bs �Ӽo�(��̎o��ܺ�������b_�CCk�}�G*/��� �����y��8���|:s�#(�p �ϛ�&q����r�MN�h˶�d]�,���u�ة;~��h�e�����@�ؙ�B�2�2�l|��9�(�GP*޿�+a��6P��_c���܆����$�iW^'��((|/�ٽN[#~��ƾR��!����M��R�4���|���$�����Y(Z�`�n�ƒ�ʥ L{B�/��Ke6H1�v�ޙ��3��|��o�g�Q։���5b�%�Jx�ik��S>�6��di_֝zqP������ ����2�H�&>z~�yiϤ.�b��\x��.ס������,��:�G�:`:bqb�$y�Z+wp*C؀��r7� \��N��eYK�ü\q-!�u�+*c�g��o)������o�2�D��(��8v;b���qѵ ���b���Ϙ�#�m)`����=a�0�����#�٨c�c����-k��#5�,��Fo [,��1|^�f��|1��&�?J�Q�)�b�h˗��C�-49���W�4V8�)_�c�.mj��H)~�y�$��E�n��_
|�E�L�����k��0��*w�����Ys׉��V����p)����yj �%3&��Y��\��lg��靇�k�>�s�z�
��=:YK��4�DR�y����ifFLz��B�J��0�T�p�h��K�ˡI�i����bh�R2`� �4+Պ��1�A`���--%�=S�����{x����`�������~�=���[�l����:r6�9�}��{�~?��)�{�ſ<"�3w����}<��G�Jd�n�̧�8���S:����e����M.���?�k'���PV��ؖ�c��Z/y����֗w�s8+�Z+m�@�����/9�`=�kO����沎��?�JJ�#�	��_J+��U�Ƨ�֞d�?
,�����H:/��|�s�f.iڄ9֋T�L�E�[:���s	X<֮'L��+��nfb�O{�mz�0��.Z�^�Ͱ����A�o����9��Z|�jfS���^.L���wY#��_����w�e��k.o�X̋F��m(�OE�b�q}� I	s�}[�CՁ�pY��8�Y�o�����s��d�p1�:��>WoϯN��E�;��c��!Y�ۣ�G��� �ێ~��5;���]�)>ew�C�-I��Cs^99>�SI�h����5s��3�ɡ`� QX�(�"m<��#.�-:]�/θq{�i^���?�f�F���Y1�+C����X.��Q�J�:�Є�����?c���Zt t>�F��d�!�c1ْ��O��ϛ��(��Y��
���A+G�H�������ZZՇz ��LX��"]ݏc<�,yy���ͶktO�{��ѫ8�=PȦ�P>��Z�‸�;��Uևq�#��>�7�}�3������XQ�(���y^�JJ��P����J�Z��(	��C~�!.>��tt�r��8b��j<�F1�)�!2�*�E�^�}�pô&���S7S2�)��^Y�C�%\���3Q��e#����t��n(OdF/���0�c�թ�	��s����ŝ�FJ^,� K��Db�p��\}��:��u6$��$����)�|��`;�ʋ����!��)�a��k>�k�!�P�p���5+������X	~���`ig+�77�;g;���w`�3��<��f��QQ�;m�Ψw������w�v�􄍈aø����Y����V��g�U7۵�{q���I����\��_�^hɶ�>l$�k����GG������_����gC�ڝ1�nr����aO	�lI���3?�m=���V@m�;%�/Ka��W�
v:��W���I�58�QW_�[������{8�e�6�I1~�������c����ދ�ԑ��E^j��p9G�Y�7��#��+]mRr��<�t@�m@�K'�k�,����U������O9p����M��6-�_
[����ChQ��|�f�_^m��3�4� �u���	sK"7Xu����̏p�'���r���fف�c��K^N=>���������r-��7��F�8e�_7�n�W8i��!��%Gd� ޑ��:�L�-ˁ� 6a�]\*J��/b#���Bn;�V�w��؞�R�k��B_<գԕ�<��POg�'�B�3ѷ��79���:�MH�dK*��(&%��7�Ȇ=�p>O��M���Z��t�Y�Q2��±p��� ��0��ٿ�c��̙��B��֤4I�
��39�*6)��L�����Z?:�҉��;���&����*]��,7q�[n)@���/�y2�3FI��}�2� �*���3���{�ICK×B�P��J�cnh�-�o:8�	G��������d��hE�(��(�8.�j�-6 �p=�S���|��-���;*t��d�A`t��2Õ;!v)��%S�o�\�6w�l���q���軛��8��O��0�xlխ���:4[���}OY)[g�A�A��X�A= '�~5����N�g�v�k&�A�N���lԦn{*0.�Zc�e1���.���FK�|g�|��������g.|�,�ڡIe�� ��#�D�vp�J/Y?���+U�l�H���?�{l����!�Eb���zȀ�n�9`S/�,�җT'�u��N�yCl��,f�,i�g�-e=gy�~g �`q��m�3>��L|1)~�Sԇr���l��;��-�ډ^��t^j���t�R�a��I�|��Aߘ�s�!�ļ�1����9@���㠉X�q���Z xsl/�=����?�ȷCя���F��goPҏ����?�W�
 ��#�kN.��t�^���K�k���ޭw�r9�؇��Nx����k�G�:a~�'���m���w��K��v��){�a�ru�7�иz�y�����	4	�Vv�9�$۷}�	�t����$ �O��ge��bH2iR&�}��dϲE/�O�X.�9�؅�ik���^q)�J��������"P�T�E �d��9�;/?���ų.Oɷ�Š��J�0y~�Ȥ�I�Py+�)#�m³h�M/s	�L�(��椎�/n�����B!��v�j��������O]��L�<�I�,A�I�N0P�����'�N���L��Ѹ�&�&�����tО<�,�	��cB����C�ˠP� �IY.bh��HE�Nq*����‚`�p�9��K�jي���ꀫ;�	d��A�ǲ[��$+n?jtA��|a����4��b
k�R���MZ�FL�4��67��m���ಓ�0� �t����e���우n����8�~VC��/3 �#��dߙ
�Db� �`���aY��/[B����^�뿢l�&ƙr�5wC�>~�p�|��5��y���{a)�f;Q���GK!���Y[��1���f��(Hc���5������O|�=����ҎH3{�����1ܠͶ<)�Ϫ;� S6P��>�҂E;ԁg�q6���lp	å��W����!�A3�z-δ��u��A�4$�����.��oB2S?�ɾ�E���k[k�V$��W��2>��4H�T�i��>�2:�.����(����em����i���2|�~��I|��A�5����m�˦��}|���;vMz���U.\���P=�U��CY�~�Y�bG�'ۘ��ޜ��gMf_2pf�7V�~�Ń�q��މë��f$�b�CG�#���NX1� S6,�b�/c"���b^i8�ȼ	>�-[�ͮW�\8�sa,��Ƕ�I\eq �D68S�W�6��I��WP��6ol,9cv'�=gVu�,*}�(]/m����0����R����J�Z]�c�,�� i�o�	�$��ϖa���)m��/h���vr��N=!3����N������C �ڀC<,k���� �d@(��i��^�E.�4%��N�L:@%�zA����Q�*B�h���Lҡ��t�dF4����	�)��ҹy�;�|k��f����V�:��w���R�����d���3:Qu��kg!�t��SÉ$>��#<}��;K�_��jc�VR��P[�g�4���-X�7!����gK�s)�ث�Y�7~�
#sJ��w��m,��x���$�vL�bg/��xg�\��E�OIQ�w��i�L'0���v[S�j�N�6�=,=D��%�/�T�u��\�T���gb^d�i˛~����[V]Ic�:7(��0`�#��j�3����W�~4��_�«� 8ğ|x���H����`7��L��S�:��؅�Cv�m�b5dk{�y�mM��A�x�5:�x�0#��x��b׎|�.������\\z�<���#�}�v��Çm]D�w�����nYA��8����ڥ�u@䑣�7�-�·ȥ mî�^_�u���bv�d��)��猃334��V�a`�9I�#���. 6o�U�u(�O�x�`h�틶�)���;vcf�rg����ue����*���h{�϶��S,|�T
�}l��C�gL���|�#Ã%|�/�:���M���`1~ޜ�yp�=Y� ��'�m�����>�|�K��.���c��Z�����se��o����N�5k����H=�W��|9��G�ڼ2���g����3p�K��y^H)i]�S��	����z_f�7�۬���7��o��]��!����N�`4��-��ߑSR����40��~�,���ƽ��`�� �z`{n��C�mt�W/�!��~��Ǿܪ�OJ�D�f���~��(�

����w�����\\I�H��
�7(����웽�F�V�����RN�Ȝ��K�7ٞ�sh�7߼�3��?��2�MTU�v$
.���e2�c8}ίY(�b�7��|Z�)1�S?��3u���ΩX��Sc*i�Kr&LJt������x�q䘸ס����m��ffpGS�D�![8��G�`�]t�2o�HW�k<>����̋t0:R��� �#F�����:
dC�鈩#g�<���٦,��:,Y�U"�V͘�,�zՄ8i�`�69KQ~�Wd\���r�%����\ѷ�Kw�K�>�:��deQ���'�d��җf;��S7�`G1�R�h�'sc�Z2'�)�Ǎ�IL��7es����@��P20� ߼�"�9�8PCg��>�����j̤bU����G��"7��%�_�����݋Y\���ul;t�A��Fs��c<r�ԅB]���|���1=?�^��>s`sn��V����D��{C�x�����:�)�H\ݨ���f���y@�� ��<W�C�	e��j�۹�i�XDSTKǥ�����-��)$]�o�ҷ�V��S����/\�5���co:��P�^�s�x#{��=ov���x����� @翾L��A3,�y���bFw.���P�l��b
�����3�*�g�DE?A^���E�NZ�� w9�_>?���~>�������������Q}��N_*m���52�6����o�æ4q�`DM����݌�d�Z9�R�.�@���?��a��82c�����aCNmK�A�'�>iMhܫ43`
��&��nH�g̦�O�|��k'e���,��A .è�%�"��Bb)c�Y����AފNq�Hґ��kkqŅ�qy'��<^;S��MP>�ێ��>D�gL=_=��Ɔ��䇥���#,�s�G�WYl�
<Wf��0�9w=���i�:���M�=)rZxd�<�tx��vG�lz��#�x;�{�:`}@�Y��4&f�Y>8�����]|�7@P�y�����+6�t������#:g����,j�GG�����8u�q�V/u�,K������/�I� ��@�K�=o��A�࢏��cUy�SvmH�WNgn�(��)�n�~�sn}����iZ�q83w�Y�A�x3X-�#h�6���؞��o��<�a��%4�����a(�8�ɓ'hIr��H[�	A�OxH���� !^y��Gy�\���Q��sfG[o<�eF�q9x��#%~Ë:��L�WhQƺ��6�_�pXGY#&������h�رz!OՕ\��xyJ�&����y��L�M�dL=�r�	&"�ʠ2*����֟mM#c��ҵ�N���S���E"��&�����CX�k��Aqv�'�%@�<ۏ!���kt.�I=�m�KC3AF�3k�F�x8��(;�P6ۤ�R�C~��)��S���c�
��h��\���W�$.#����~���lZ����L��$�"��[�΂������CC0"s�"JNӑ���t,����(7ٌ��2�W����ؒ6����~���6�_�W��X����E�L�ܼu����_~�����O�p�p�l�+���P���K~����Ѭ��7$�+��PO�.:2�e����Y�^�M�M�$�o�w r=B� �2���H��KFδ�7?��.�����|� ɹ���_�u�
�ۥ���tua&m)�bRT�::�:�����#�.׋��S|K3]xC�Z3I9���;�B ����ɳ,g���6�{[ ���E�D��fu�8`7X ��ͳ���O���x���� �.�;7�G����[��\릴6 }]�������W�V�3GM[�s�Z ��L[�iӹN���<������妎�Ƭԕ*��]7a���;@?`��t��7�:���8��YY�P�I�؏�>�E~����������%٢�2�$�ɕˆ9�Jcv���ͧ8d>2�?:��	J�c�Y�v)��%M��K��A�O�?e44�����2�����~�+�m�@��M���d�n`�Յ�b��q��������̓D˺S�j�,�.�
N�`���n�g���A�:D���s�s��8�jI���'Ù�:��Ua�����VL{&]>�1��Rf6�O����w�;P_BJ���S�&�_�B��~t����W�������'������ɡ�j>2��=���,%C�	c��s��)%�l���=I�)��33��*>�r�}�%�� K��ף�ԑyV����\��n �`Be���;7^�o�sh6!4l��`˳�Zo���ؕ�`��Db\ǁS?�
�g��K��Tedi���#i0צ������Ζe@wً��"���F�D�E��)�E��o�-�����l:�wz��L���+�xs�٣���?���]�#͖~R�۷W>�o<�����������/|,�Gݶ'e�E9��L���V�z��^��L9��ə+���Na�[����JY��Ӎ����Riٳ��d�~�� �(h$��9Օi�oҸ^dNl8H���"�B��R��U�!�2r�'W�Q�"FJ�I67q��%Q&�a\{b��OS-HG,e���T}�vz�u6z�O�ΞsW�������ͩ�x�����m�P�z���d�r͎�q`C��ކ����4�����H���\tY}�ӽ�������MSV.r��	o�!x��B���U���xY�nU8 ݼ�: 71d��ǂ�ܺv��'���}���s�0 �`�k��w���:��pϞ������F�ɧ���ֳ�e}ˈ����.6��?yn`�M�bGrl�N��y��������n��<��ڈҐ(��->���}�`h����"��d _�<ʵs3]����]NI6����`�&g���q�㺬�ȥ��un��e�~H���c��6̶��z��\Ϛ��+}�0�6����:�I/3�y>ϲ�������L���v��=Ǽ�!��h�؅�����"]��kSOxp���,�8�`��Ƶ�Y��r�dX�������8 7��s�δ��T�m^��Ȯ<��	7���NҚ��m4n��Χۗ���O��.4��˭z�9q�{���^^@�������U�[�ʢ#f����X�hfܮ����)p�3zQa� (�ۂ�j�꨺�V����<����/��r ��ҭ9�]:io��ggˮ�G��5u�p��b=�~gh�
��b��oM>c�i]�kL�6���&���ԃ2T��kje�.K7���]�����N\\�ؔ���l?^6�}vdkJ~8P���,��v���3�gO1q�:�#߰����g�?���������ɏ[���x^'��6D�>:�67`K)�k�X������F�^�W�㠎�s�G�\U��8.s�N�lR�(�`V�Mk��0��hzq��&�����q�5��� o_�a�71"R&��6{Ӭ��� f�E��P���Kz`V|2|�/�3�r�w��$m3��f���s7KcC(�Γ�8�v�v���J�K�t�������8��Ι��(1y�6�*z��vh�˸��0 ��4����G���QEqZiBj�r1�Va�\�W���"��{L���U1V�3��5v�X*w�:d�8q=a����e��q �	;=.�:^tHG���=���_� �8�ΕyK/al�,/�jx�e2׫�	tʯ�%��S]��G)��@��a����U[�ƕ���g8�>�2^;��<�t�����e1�&�sJ@i*ƒ�H�M�^�ҖhY��k�I��:��� �۟��XgE䜭t�֑.~�V�2���>B�6��G]؆��ѻ3��k#փ׶E呾(�.��<�^�`�-^���+|�Iy��7�Oe  @ IDATKH��O��=�MZƁ���u0��-	�tA�5���_s�lx�m:npq�˂V��s6�#Ŗ_[}�8q˫ϩ7�����_"+n���^���+ޘ��@���z���z��Z���=�K':��� ���la��r+?l-��!σ#mEFV�vbq�݈��#y`��`e,m��[&��כ�o����m��<���ZZ�!)�vHy�l���^�t������n'���"��Y#e�բi���^TEo!�D�c.���!N��� �%2�V�+�ӊp�Z��'m��M��l�ΗjV�f?��%Kt�Q�%���G�.yκ��l�q��s�M_�0��4���D!C}-�v�#�Z[����<7M������I�@�T�V����`1u�A9לc����zT�)z$���Q�i���Wq��zIm�x���N�Џ^�$A��Rs��ĔN���+0gIF8�Ij�#��"'�Yڞ!���{JKǴ�Pǥl��*��?�&��g'b䴜��q��S���<>���3�}x��	`Z��]�qGͷ��&�0�XB�:�`�M������������_x�����W	�6T�u���7���Պ�S��,��t<ʻ�	i�;�IZ�\��W>ۧS�qꄹ��t]+28���m,��Ou$�/���>wJ_��{����W�����������������"o����B�^|J��Gf����9�|��qބt�;o�:=��R�VG�����|�t8;��<���V����������[��khM�^=(/i:LFv�ڂ�
@��*�b����ё>|���=;[������-i;����3Ŭ�)��)A�:;�Km�}�[S؆6�D"=�x���MN⬳ g���m �fw�:���3i�זT0��_ꛙ.w�w_��ˁ�MM��Vo.tƲ9��]���@�y�>n�3��P�I�7�Օ��?����Y��絭u�_x�Yp��o��_u.M��I�5b������/]�q*y�eFl���ۤ�(���K���:�@�9Rq��L8��l/���>C<��Fз���3�R\��&x�
q"��M�^̯;�6z(�֍3���S������ 4�>����_m�҉�Qg��DG�8<,z�D�g]��-m N�W�h(O��x��ԣ��O��N�e�C��k����1����!���-/��(���I�F��ͪ�qX'8گ�K�2�A\;3d�Jǘ�ޥ2��?��ҧ�_	Çk�r��9:e�5��U��좑��2�A��I��[�Fw��ң����U��J�<G��_@q�]Y������́wz��o�rx��7�W�6�%9?*ܜ�`aS�)$�SZ<-�7�`�m�dv^b��R� ���
����H	ҁ�N e����g�;^��gi���Q�H+.�%����:�e�-�ܓ�Ev y�x�pa�Ȼ��0��
����#�gv$SO���Z`���M2�9�s��}�wAu�(�u�����%uLtR.�"GZb;v׀��?�#�	>5���%0�FC϶�ڦ��_�Wiʒ�NK�l}K��������t��Y���ɓ�0�����R5Ц��[Ɉat5���^~jai�3�Wa3�&���O29x���1����9�B��"V+�J�8I�u�%|����z2=w�8�q28��D���ȑ4P;#�3*v0��������#N�t�_�k+�2�A0rxm~����ЁM'�lp���c���`��,�i�F�s�b������ ��Sl�N\i^�!�ͩ	x�^�Mn0t�����7���\6 ��(_m�#�����t��uq��M7p�@��G�gڿil~I��/:֏Υ�l��E���u)Q�8t��3.a��r.��N��O�=�V���}�]�3N��r�֟~���ipHK�t����)Q�I����9.�ީ��M=��B�3j�m�߹i��r�����������gO��Q�}DE����:9�[���EQ�L���!3���3�9x��<��WҶ]sK(p�ك:+���^
�;�ltC1�^�3'-Cx%-�s�6vL42؞�;�2Ox�z����-^\�1�Kĵ�����x���1�H��+�Ll��;6=�Z���ʣ#�����k~���)�`��?�I�e���g�/%T��z�G��va]DLsl/m�B��/Qt���d�Ʊ�N_�U~ㄈYa8��o	#A=&\��M�r�h���\b��6�p������>:$<#�P��:�g̺<}Ƴl��_���Ѭ�����|Ϟ�I��v�K�Ȳ�ǝ����Vx��;|����+��K^/�b�Мs؋o�)�%P eHPf�
gH�8�-7�&�W�|��8](}����3:��w��͎�N���N�خ��Y�Iځ�E��fG���髯��+>o�5��,e�6uAߝF�A W�|��������3�'��f p�2����h�e�p�Q8@<|���q��58k�@����?2�?>�Wr�R�ʑ��{�4/��A�I�Ǵ5ڨ3j�vʣV�t8~��'f}�T��K7iu�꺖l|K�5����
�_R:(ʣy�*��A�A��r?~�8����}�n>�.���f�|�n�g����L^���R�<��>�P���I������=���:b[֑�층�8� G�d�pD�ri�LxFW�϶w�|�8�IS&٫G?�H98e���U�΁?�����h��ufT�p��ҙ�?�@�յ���uQ�u�t:�Ǵ�i��P�׏o���v^Zxg�Q�.|~��{�g�����>�C�$��i�Ge�>u0�N�vM�m�����<�PX����|�M�'ߙ'm9����f���yS�����e8^ڠv���Gan�&}�H�mX�8>n�X^���+xpv]y�'1�&���k�t�eՏfA����shi��8��ڐd��Ԡ'C�όy���m(����Pʐ�s�0��V ^���{qm���a;TJ]��d⸜qeg(4���/�C�~���.�<^CW��TK��[��û�><���Ǉ�|�֧�g���o{���	����򥍶�"i�uZvxaH�9U��©3���n���i���C�1���Sٓ�}�&��z����h�� J\>{��˜�QZ����E)��)Q�b����B�T�f�O;:_K@΂�t�))�+��rp칀�n��LD Ӌ/�a
(R�����?jW��R�I��x��]Rlh`�\_Ҡ��,F��0�gl$���H�Q^CHc����0���)�\B����G+{ׇ�Bֳ-�}��§�X�̽�S�C�?^�)7�*�������ttg~�㌎�d� [�t���*�#�z.6,ꂼ8k�k��p|4�w޻������D���^8�Y���a:��S6t;�'���ٲ�u:?��L�w�>Z{��a`=��)�G�ʠsؙ��@�o�e�J'$�C�����Ϫ�ʯ������_�5Y���t��k��R���(��P^�����[��a=� ݳ�8p�<f6�	3u :h}��'|����|P1�$��TWq�ѣ<YWʖoÑ�#iu�� F���G�D��~���K:����άWʋ�e�;a���?GIiPf�<b�Д�)�/u�@��dp��;i�5�Gu��Y\�mKzg?N�e�w�R���	4�Sg����L{v+�3fUK�Θ~	��֣���Ξu;�~uP]ȗ����L���m8��bsevS�kמq��V��� lCeEK��f.������c������d�f�>��?��UW:�����_o���_�EEˏ|*�Ε2(��m�nH�9�|݌S&��@X֙@kHGT�@�q��wXGj���?��L�6(`�q�ӎ;���]Rβ:�:�XEu&qB��$-y:[X���But53:�}/]WA�:X���t�ϯ�j?�A�m�`M��`�4[���>�!�qPgB*�m�o@����e���|�Kl8�q���{�f��9��3�Ln��ީ_}*o�˃�Y
mס�z]�Zec�h�ò]r$c)<
;u#ދ�2I�7@^YX�GaGP^W���缲3c��NHx��#}��!��8N��6m?Ѷmy6m� �MO}����:f�S����~�<���G�F#��F�Lʜ��iK��\�$Pű�.&ӎ���u���1��E8�;l��!e����؛��g��}��)����n���od��G̀�P��*Z��/i)ĥpl��W8H�rz�1]�͆Jx�{�c�:b\��6ڲ�AI�oG,��~�lZ��9ʁe�]����<^������U�V;��`݂с��W)�����A�x�*¶#��ӟ�g���޽���ϞqgN9�4J��ѻP\�汘@'��&�	{G�]�5ζ�:$��la���@��Hӌ�1��;:�릿��h��%p�H��N߁M'n������{�+N��"��<|��?��� <�A������V��fЗO۱�Ԗԗ���̀a�g�L��.v�y��7�����?�����~��@ԏ�N�Lי���:z��}m��̀A���u� �/|g	�[�B;�g���\G�N��q�ԣ�U�C��m��R���R x�{i/'=8��!��ĩ3(�::S�:Vu|+�ft���8�2�p��Hǻ]�G8\_1��5N�31�EzB?��3+������[β2����<�T�^c�f�U?��5[~P{��8_�H��Rq��u��l��ڴ�T���اN��9��)/�"���>�4ۙ��G�>ű��=�	�]����(a�Oi�8���8h�W�8GN,,g�i��4��%�����}v�,��o ��f0=I��=G/v����%�Z-)�����/�撒���)�&\FDFfem��hvt� �~F{m���"���A:��(fz��m���Foj���3Ffx'S?#��� ���O��v�:��i9o3��)C3�E�eYN\��뤭��l)�B���#��_}r2�s��g�{0X�����X��z�QǏ��v*�C)��/��x%ou�����w?:�[��v�+�����y��&�������{����nt�P-ݗ��[�.ȣ��<pt{񾂦}����b@^���_��o�_؎�̧�9��?՜κP=��?���ʛ]y[���ۢ}9-g����g0���2Q"�a�t�ņ�ʭ�c_��pX��
�`;���[?9�L~��+F=�$p��̠I�iL"5K�M2�'�<+�2J�h�9�p"]ϛ�)�&�_K�]��L�}�'�c���~�G,�*|�C�`;��Q��l���x��D{��2��1t�EhˊS"����m��g��<�y��sJs��ޜ��r\��Oחu)P�G�s\��� ����FN���ͥ���j��R�7�.�]R�ZR�*��U�L���{�U��ʗ��M�'B�rs��sF(?+�����u{����F��,|�
�:Q���+R0�'���Y9tR��|�����w8O��>ʷ2�`9�w����'��d��OM�&��mxc��p2�D��N������mc�NF~���D������d���^?|X9og�w�}ג-��<��R��L4�\�6WO)xQ��:�L���p�m����d���>c"ޑ���S��'��=�B�]g�l�rF&�<�=��5��7�wp�h#3�7���-���²�=Ï�>����/�����ar2ϩ ?z�@��w�o>���Aw��a����`=6���\�&�[�:�,�,��W&<f���������6�i2����6\{�խ#4���LO�	\i�&�r��9��1��QZm�>p��q���Κs2��=T���V�p�v1�Y���ڼ����v��9�C���9��|tpOF��g�m�����M;�&_���e�^8�������Hg�)/�:���<[\�v��~�IxY����� �9��9�t��)�>?]8�	b�oZ��6"D��H5�G��v�VC������*��n`w9��l�Ǟr�J�r�-
l�ODɵ�{S��Ũ�-�Gn��O��y�$����)�������%�'呞Ͱ�;/�gB��$��L�Û��[�������E�$6��l;��)Y]m-U�!é�����=��6�V!�;{2�O�έ�ȿ���J��x�3���<��e�FlJ����%'[z7�빡�y0�6wo�'()�v%O}}�JYB�h�5��]�l"f�q<��Pqd�I�{5u{��^��ͳq1S8wS�m˘�9����\��L���ѐ���a��\�I��nJp��\��P���գG�__��[��c��n��˼����*SuOyҔ�ף���JC	s���j�3Qo�ޮ,����--8F��"Cx�}�	�+Ļq���t",��������;x���1��A3T}�2-�� �s�Z�LDa".kp���"5������k���0�;�#�;�!���	|SPp��gC��/ؤ�{6����}e�6�����>�]Q/N�톻uF��"�|����n������J$�s+jԭ)�B>Ng`����ʕl�Jv��8� ����Z��GM�\��S�u��3����&���Ýn��g��$괃Ky�1 �0�ǽ q5G����'�d��G�|=��h&�n�x9r8�0A`(�W��C�a�=tQg�6�����s�ށ~db�/󧆷��xȥ��ku�在MeL;��"`��3�8֜-��8i��z�c���Qv�|�jqޡV�L�2t�5�.������mc�10/ܞ��~u�Et�m�C���Y�LzU�hd+����	ǫ��>��Ƌ8Nt��a�$�t��<�,h�E�*�u_���D�k��:d����J�orV�j^ys��E��'�Q���]��h�t �� v*[Y�e-K��m�������S�9�*s_uD������yr�>}Hwb��q�����柾�S.���<��ih������޾��]�c�8ŵ�Y=(�4����>�XR��n;�΃���������|���rʹ��S�캫�ɲ�Mn^���{Zw����9���oj_��b-�L�q�EH�	�kDLYY���C
<�S# H�	�a�K��>�DeM�w�*{���06�����ฉ�
a�Qc<��|�P��L��'���t@��P_N�(����qע� ,�(z����t+�m���ӵB<������LJ�J�e����^w��q����[�^e+N��4D��ئ̄_��Ba��@�ݬ�>J������N��pJ��޽��^3]�ۇ�v�.��J?�2���$���;��7���\!̽CY`f �Ygo눃���'>2�� YCwy@�z"�]��iu2���艷)_y�eX���s/�FV*#H�Y����~�����)se��3�KAh�RL@��08W�D�u`*h6t��s���{ �2�Lz,���|o��ۄj�/,�h*�÷ Չh"-�]����޼�!cpr��y;mi�IІW��Ņ�V����@U��+b����1s��Iˊ�9c�.�Zc����Wy�av�Á�,�c\)�M�u����G԰�O 1��#)���Aq/�]�,!��30ڻ+�����!;� 6�<�z:*dryʹ��C�x��:VF�z��{�7t���Y��î�'��e����Kt��wW�|��:��U�8'�h�9���I��+]�)��F9�����W�6Hn�Q݆`�e֤:�74�ިƔ���2W�S���o0�W��&� MVNWւrҩ�<Ss]��������0N��}�y�������I��l{G��'`���M�Ϊn�K���%����͍��-l�m�)�j����p��~��Ndo�ؔQh��O8W��yJo�yS-�#_�"�#<z�=zC%�dƮm�g�qy��9r���S���M3�/�{������#��NSnmcҡ��N@��}���*\������D��q�u�,��-v����w��x�����<��Ϳy�8�ӛeo�AR�|?x��Y�S ��vv���x]�I��v^)�YO�"e�w�׸�K���2��j���NgE�0��!y\�W��-
-��Ex�!����Ԙ4�u4ի�`�p����)���� ��%���`���2�d��5�� ��y��Pfs�iW���.'ϡ�?��R��3&Ӏ��=6ʁ�ĕ�s �~�ݾf�?L��3$p3<P�����{�C�p����Q�e���*^m�|��y�*�9h�P�#ogu	��.h��yP/3p?�6������$yJ7xE���,(�z47����p)W4H��zg"�3�	o�0�&/�Q�h��
��J0��۲�e�7�D���C�����j��P�>p����2���q��x���)ˎ��1�~(|������\�0�����9W����xU7gTڇ��y����!G.[��I�������0�����E"��A��ʌ�LsD���s�3���	�#�H���ۡ�}�r���r8�_~��ٽ�F�2����r��@�"����޸yT𦗔�9����ȿE%u��K��C�$�����<�CYd�~o�I�PkoNN����[�����Y�w�����L��D�f�TV��V6�q8��fC�)��Ks C��6�l+/+Wh2��t��q�Or���&���Kq(��u�+�U��h�s�4�9�O4��G�ϣ�F��Ng���6�)=�&C�jI�Lw�(m��C��V^�I�2P��Qg�G���rk���җ������M��Ћ�=h(ג[z�� ^_��'}0�V�ib0eL��]~:�j��6���������7ڿ?4qow�R~mڿ2��z�t?z��[�d�������u��!���-{��%��>���*�#���rXhG��o=���m�ՠ]��ÿ!��9:�/��*y�F�iڒ��?&J��I�l'��.Z�p�u}+���~6�v�����-}[{���lcb��������+UP��\tbǔ/"a�V)���'Q���2#�!!�dу���H\x\�g
b���>%�q�߇��(�m���xR�<ʷ��g���k��cY}����)_��JY}~�l��4�'��I��UcW��x0���̈́�
��a�8ty�<�_l=fn�C8��vB|��IQK�K����ʳ_n��6Gt���T��'M��hM@����I��l|�M
����Go��&b=��/�q�����}�kp׌��XG��g/�TJ���ޓ��}��z�x���'���}Jv��`�)X
��%J�`��y�AГ� -�+zb��|*)�����Ѓ�rE��[83�b�����|Cw��7Q=|u�����И���j�jh?xu4�f�F�.ۏ�9�$Ouv���Wẃ��q-�m�s|����f��$pN�1��ҡ=tNg��Exą��7V�+R�Qo��m��}y���0L;O�2�臏��p�{Z����菣}����ѫv�{�/9>7�k
=x02����|eAǆO"�/?�y��`�*�|��P���!��Zq6�r��Pܾ\P���;'�W]qd�m��h@�(~�?~!�����P�#M�cp����f4A���C��+g��� ��	Ku+�����.�:#ڈz[��j"�,
�>彗9��svxW�D���<�59�pG6����L��%Jf�q��i�lea��S�:����6d�:�)�ȧ=�?��!i����(0���?�ަ���-��x�'��Շ�ô#�Z�u�<Sd%��y�ew�����e2�sѯ�:�rʺz�\t��Ώ��|���~�������s������%ޓ){@��?@Z��#�Sf6{�oY.��s\'k��N�`���]�/��e��,t;Աv7σil�{48l����F��q��8�m�3�%�W'˰tM4��Ar5�;2$W�r]���^5�h�R��"a�����ɯ6)_�hv��a��8�Yt����_7Q}ވL������֗��G��l:�D� �>���qv
�ƏQ�LV��<>'rD�(d�>uy<J�@&�ܜ�� �R�qQ���:轰�ߊ�ӻ�x��O��_}�i�]g�A�$8d�.mW��)��\Ob>�AQ��N�=��b�Id�hy.��S�<a�J�~��.���� $��qS�bf?U����d��,C`�o�9?ǇǤN��V0��D$�"~��^}�*����0֚z�ZI�͗��z�.�$��n����5�􆍋���M*{nQ�����{=yܼ��H���� ](�M���>�bP� k�l����p��f�+���%�p9s��rr{�I��s�Z]��3;8Ѐ��?Y�.p��Bw.9�(w�d|7��8`�ȩcxV^΂ȃ#��}�^>�yx;�ɰ�C�>��:W>�6�`�P�1�W�9P��2�����d� ǲ,���>�e�4	�P��sB�=�������
<�׮�q����b�:�qN��O�7r��5�?[G��06�m{��Q���C�Uڡ3�����V���yz�=7?�F���Jx��3�<�-fY�H����Ï�>z0N)�R������qhԻ��&�d�.�ǉ#C6�Ï��2¼ >�)_Y��f��螣�9\<���<�������|���h�`�(eyLR�|x�����s�A���Ǫ���+��藼(�N�u8�iW'�� �e�~�&jR����0��W���T|�9b���n�ڂ]������s��}!Eg���4Q�r������� 8��r_=��۶,��N�2>ܨ|d:�r<�[.N4��͓�yW6w��b.3����:�K��?��t�Q{�uFֶx�_���&Zz	�����F�0��G�L~��q�|p��X�J����O���O�ZK��])�6.��ֽ��O%v�u�;��'�K�
 |go9�GFK1_�,A��~lKz�쀚d�h9� �izV���eao��w}��j�I�$��^O��_m�A��o:�zc�4�j��%b4d��E=�[�)E�&�z�o�>&U�4.@�H{`���3	�U��W�GAx����;6�4?9Dذ���8$x����12�0WLt��]���T�cyq��6`"��m8s/�Ml�=���u���I�<�B3�(z�H�'��:���3�繚�p�=��6������GE���ޗ������u�}�k0c�S��烲��àS��0������u(�%#��,��`���Q搘�!�l,�ZK|Xպ\�'��_�[�w�#G�3�9�/s��p����cu<`?�7B�F9���ax�������a'�p�^���e2k���3�1dw�B]�@"'�n�<o�Dv�%-?ů�:Q�� ��G��Q�F�����E��Mɩm/�8-�w�g��y4�F�a�Z?��E��1��vԵq�����5k��=��k��6�	��ce;���qU?�Aٳy��yiֹL.N�M���5������V������៞)k&�:�N��b��yy$�df���(!l%�IW��h��Y�l�S>�O��9ǆ�M���_���FVї�ٖ������򹴜���.���z��9_�ݵ}�
G�pz�q��Kx�7yT�-\K�u�+��;���:|��]���8��N<��+�Q[�V�胡+��|�]���6��Z�)c����J��l��j�����d�G=��s�]m'���2B��/��KD�vKܻ{{�fa�_��)d��0���"������$m���K���I�,��cCͥ��N�vXn�D�f�zoz��}2���Q�>�t?-~Xw*N����ɁL�\OP@ڞozݹ��l1|��v��)˴K��|5y"K����t����pq�D��4�^��q�r�+�0�!����r�z������;�  ����Q��{�[���b"�Ic�C!��h��u�=;�Cm�g>�7��ܵ���[�&� ���7º��H�*�_/s9�oH�"RJ�xC��U賔~�<Oi��F
�F�#�
��^$��C�٫<:�3ys��t�n��Pw�7Ŝ�= h���>߾2~�
���Y�G�Ƽ�x��"*��ޖ�J�h���L+�X�uM�~���1Qgp7h^�)���h��l~�`T�)oO&�e�贡������������x��Q��Y_�yea���.���M�	'O����aJ��}�{je_1uV�{���6$��!»7[?��7�r�i=�IC�?&G�`��&,��bk��P2d(}�8.&�Ǹ��Vÿ_d&Z����}����9<����f|�e��p�=��B��\���U�)�W=~�������	��oÙ�l/�1��:A&�2z"C"!�΋�yp5�u���d��`�o�E���V�o��&}.�����p2�r+Z�j/�3�`���h:/��h�%��T�)��}q���(�)Z��A ��ge��1����Ũ�uJt�N��u4�v�-��a4Y�������-�2{�=��%)�wEW9����hZ8�g�R��'c�q� �$�E|G����B�"~d���Yю�Gr�>���P�.��ݔ���|�DR_�i(^���N�􌬨�'��L�C-�y�I��G)���=�E����hk��ޙr�>=����q�[�n�G�s�u���R5�E�'ꘗj��wm�X1z}�[y�����D�7�ܡ)��o��ڔ��Ik�:{��v��)Q�[M#0��b�ى��ʡ�oyQ�ց��hM��ء������%�k��lD�m#��m�:hbj�bj�l������ӟs�t�n�#z����!�D����>�4y�����1���?|�\�sz�FY�
^���$�� @��_;#���n��lI����[e�<���'�o��e(�m�>n��ۍ��g�Y�����ҋx�Ͷ���4�a>.>j�����:`�	�=�r�����6���u�vPVd(��XVv8`�)�j:��<�#�ZPa���Q��7�fnqC�/_�;ܼ�p��Y����6Gc�ׯ>��b�SQg7���o�9�5���U��晞8�Ps�Bg!�FĜeXy���0H��Ӊu�._�Ŝ�@ϡֹ�{��h�`GP�H�r��/Q����fu*�=��m
���c��I��˫�D�E�͋�`��U�:D]�����6��?J�8~������8���.��%��p��pN���ֻ�M�Z�dv*��$���t��.��w�j���	��;}:$����Wg�[��W,�+?/�kHw�3fE�.��-�{~#':g(0�����nM�����`������;�U?��X���:Q,��V�qn��F!F{�u���4�g�0*��q��Á/�2�xC^i�;}�C�o�Cfʂ���w�y���L�&�Qd��f��9�O}����~���Hcr��B�A�Ƨh�t��[c
�d��FK�5�C��s�h?�����t�%<�ˋ��˹Q�:Jǐx�g��q����� U�D�)����s&"`g!M����5�˸��7�ՁLNԳ�<�|��#<�H�LG[�P��2�!�����g�F�"Rp��K<NGN98p��с�.C�Ƀ�O��r8_+�Y�xB��&�{;�o\���x�i��b��v�=������5�9s�DWC��I����4y~��V`�h��J�����δ�ڃv���Ĉi��~�{�k���:_�/m�ypv=x�f�Ʉg�كaҜ��6�=s�Oх�"���- ����FH�Ó���#[�v���#�`���������#|Js:tq�97�D{t��l���t�܂�H��t;��5.~h��������/n$.���&9B�m'#��B���z]`�u����`�M5�V�Ew�=Y�a��+9k���]�4�*8�p��w���)�������N@Y����Љ.sl���@ҕ�L��{�Ϸ�O!�u���P�k�c���e�YM�9Y9b��_�ݺN���"�n���-�� ȳ�-��2h�U�{}� p�jOڹ�z��Ę�Lр��-C��������)��2z:o��R^�ۺ#Zмє�g��d�s^����l���*b��z�"��O�lb5g,<>3��
�9`���Qi�����tv�p-���x@�c�X��ܵ�����nҾO���q�G����sBs�8��A��Z�S�O����i��9F�C����R��g][C�i��R��s*�_����ݩ�xc��g��(�W9f�_���&�?M������r��S��1�dً�����1|Rj��/���r-�BK�Q�u�6���折ph�4wG���qnX�a��\�:'��۹<��3Fֈ�v�m�[h����%_�W޼�9i�N�<;Y��^pp���X�E��7��uLk�v8��3�ql��9�9�)Y��9�|�Z�Y�̺Ϙe+o΃	�=?�c�N�1�qN���(>h�`H�f�+V�EA3u�sv���պ1���S&��=��_����1�2+��c,�7���s8]�y������.�A���9d�3�l�O/i�������;.��I�?UЦ�q�å��$=��2�(��*zzF�Я�9�`��{��F�~�Ӈ���s�JcV���1�i;Y�cz�����Zt�o���Жn�&ڵ�Ec�H����w��������c�g�\�=�����|d*�楌��|��휨�iy�m�ո�q
}&��IX��z؍:{�:�r�$}�������Y�R�N�%�㵶#�	(�E����"��Vﴖ�^�ww�?��r�=�����t�.���l�����b��n�s�S�@գy�g���'l��[��`�\�=<����[r��9�?���Yit�ޞݿ�����.*�0]�$!�k#t�K�NN�͢Lw�3�O:��?�Wϴ���9�=�<�l��Ej��n����8��i�C�噴v���(��N��$C��ȗ���Y.�e�r"9��z	���^R�By9`74��P�v�(�ʾ6� ��Y#�@��i�[�F�sVXVQQd6>zR�'��gz�]?O�'��9����	��#������B"v�!`�b��&��ޕ�y�Hf>����v�<�'<�]��XN��9L��}�l���+w�7I繟a���UC�j��u�I��?�+�(�89�"\�&(x���2���#��aQ��?����oI?}*�HG��PSL7n��`�6%-\�p��u�fo��z���B�9'�VU��5,�X�/?�?�a+�؜ ����_�S��⍆�^�[
b3�'��Ə�R5���ɹ�ξ���r�s�4�CbN�O� |��+�3�S���nh��fX�DQ����%����S�=���$({zG��
Wa�M�qt (uF]7�Ӽ�g�i�r�Gy7K4{p���FGǄ���D�z6Cik�]��#��c���w?�}������m+�������8*w����B�!���h{�o�P~���2������z;��K����׵��pi/��?�ē�3T\��r�_��h#C�tr(��I���}��S��?���w�3���5N�DU5F��[p�0 �J�8u�,�P�T��![�m�;����s�:R�'���F쒍�{>ϯE[Ώ�f�5s���.U����q��C�`VwP�5�k�>��FL{�1�{�
8���1ȼ�!�
���8IJ�,��_S��`�R;�ސ�;���'/~|�ݷ����}�hUY�um��}�15
d���ކTشAskƚ��w5��q��cs�*y��� z+[�ﶣ�=~X���);t�>4���a�]�3�M�O�~8���$>�9�/�V��65��>����F2#�����iLd�	Ll
5�6s�))����PY���Z����m$Y�Ar��Ұ۶���t��m�S�(��M;H��d	�Ny�w#�����f��&W�Xx�c/�5���~ε!�"��;����<&�%}E����;>�Yf#l�P�o��[�E�0���ח�7��|���8�<CX���iT�Q]ڙ��)�`l���6S�33Ɵ8&?���V�s�P������u�+;��嵉��]��W~��U�՜�����  @ IDAT��Nl��S�A�z8�B������Rα/^��+�C���sG���֐�ǽ=4�>%��r	��-�ǥ?	�<��|���'���:Gı���S���{�ƕ�s���%^��������D4sw|z�~�=jk)Q�o5\�~5|k|<�w� ޾}�t�6zѵ�{�n��uѣ�gNKÂ��6���L�7"���K�u�c�q"S�׻7x�?�W���(�բ #ot�v���2��Eo�p(g����Y�N���+G���m�*���@���z�M�Ws�D�,|�n��{���w�s�z�c���F����([/y�}J
#��8c)O8Ý=��^E ���s��G9ʭ��.-���:�F֪���K�gm�����h!SC9���u
�#C�Q�S��l�f�M�8� ʃGV�甾�Ō�.R�G�<v�N��ǝtO�&�,>�MoH��a�i/�f�Cϧ��R��grUzUЧl�"'$��X�	���8/��h�7怽(�l!S�'������r�b���"�z���Q�ᄑOt�7Ä��u�)-��cH��c$ċ�ꞁ���䏳��!�=,� �U��<h3��G.ё3Ɖ��壥ǁL>�9��]��L�Q�Q�k��彙a�������ϝE'��f���ž݉N����_$�����=�[����FE��]-[��%A#Wp��[���6wO�C�9g��Ǔ��e�����8|*���qN��~���pL�Iw�xr*a"�� ��������&>�N+������z��D�p�mO��xM{nakÐ�9dVf�����5?����'}w՜���5���>�����Ë�g<�d��q���A2b׎�{�����o*��<ӯ,&��75}�P�<�+�%�l�E6�ν��g����t����a��U�����sB(�T��w5�z����o7�'�y�ׯ�N�4tԫ�z���#4<J�*�0R)��T��<��]kP��8�qy����{ރ-{�(0���+O9�>_rSL����6�"T�;dcZ�6Gћ�:�n��_�Nn$�ބ t[�9��N1
���K�4*�Ώ*d��T}Y�$b��;��S�[��M�����8������ˬr����Z9����L���j��k���s7���j��g�aB==���խ.*��1:)G�eDE�n5�}=���Wz�6��ys�!��j0�2�<�Eq���1Ǡ���S��ٕ��d�E��|NIR�S�hSȃ�Ը?�z�Ѕ�W�J+b��~�߽����	��A8��Y�Ac,����oNFV]�%r5�P�&��%#d�2���T���c��9d�l�AVC��:%����N�=m�mtQ� �d��#5茾�~�}���2	��h��kD�1V�*;�6��0_��lGHp.C�~�8��u���R׮��(ی"�u�O���K&�;Q��h�J,�Y8���X"E
�e;��ܳ��t�� ��ÊL��<�]bc�eZ��>��=�:l�\���C�Y�I���,�"��~KgK��#��y���u��L�h9�1�5����пg�uD��a`ڍ�NٖtC���.����Mrv�r�"����u���G�B���`�ۮ7ixU���-��]J��d�0G)�M�>�P4�q�_�nsS�&�x9�7�2C�t�a��E�p��o2���ZtGZ0>$/�k:!'Y���߶+�!�i���>8Y��}������}(��Ϗ?��/? �֝O27W���ͥ$�wt\dX����N�=/,^v\��c��%_��׈Ń�s����?j1�O?~8Nף^f���C�H+�H�q��8�5����@%���o'�Cz���!���l=��oo-�?m���&ғ?����c�Y��޾�`��O�~=��i���KW�J����/��5��������a޼��>.C��m_�M����X;��U|���z��)RX�ۄN�l{K����4.�<�ʤ�V��{Y�)�(��E���K��u��?~w��^bs��䐉�\��T� �k�l��O�p�QhW���I�T���%[��ݷ/΃��4�=�z���Y	6o�`"o��e9_�;EJ|ڎ4.	�e��(=4�ri �ˋ����3^}�=�{�oP�jރ|B�aW��jg$�@o$���L�]C@�}��E�B=n1�]i��j4�)b��o���B���9�M��1qX62�k���E<	<y"��D���Ãw� �S�w�~�2�:y�A���Ǿ��0<�n��Wg?��2��k�W�7���"v��=��k�E���~O
nhJѿnAc��ɨ�(0�8h�,�T�-:��d�ܡ����99{p"�]Q9��1��U*�3���=�.J�=On�W�4��nN��[��W�p~}�m�+`��6bg��n��8���}��i�����Fn��ݝz����<pAC�)g����{9��i+��8ݫ@�t�+��u2�h�v�:�;a�߶�>ޠ�]��t��ϟ���F�N��4z�ͽYI�^���`�i�E�o����%?8�>�3�u�L,b4��/O?��F���n�I��&m|�S�a��[�HT���>�|K���u�.��K�f�e2��E�`<�otI;m�Nz����Dέ�-G<lj3��dG0>���,m1��y��Em�z���.�z޲��MG{ܬ��Q�OϿ|�ض�Z��y���z0�*��r���F�~#"��E�`淉�q�gfu1���]���땇�� 8ҕ�6��&D����y�5�bf]9[y�n�'����'��vJ:G�D{7I��ӽ?;��?{�Y����E��I����z�M��q�>���n���限���E��'^��^�p5��ș�՞Y��]���|�h��G�n���_������>���"^�;u���R3t[
���t҈qSM�Q�.3p/�\��s����1(HS������_I�Fǣ��.8ꚕ` �Y|����2�L�����y�ȇZ]5`W6�b��rHrhė	!�飏�}���X_��@p���n�Xe8�d[~��J��9�&&�Oh�:���h��C�Z�%c�8��ϥ�=���������o������<�Ue}�	!Ŗ�(����&d���<�O�_r�/?'=��-K�S�|��qh�?9�O8gG�{��A
�Pb��� � ��sLhJ�/�����4�=�����%��FJ�s�y(�����{w����04�����)��s��7| ｔ�����Uܘ�͜�+A�h���W����6)����5��s�@�Ͷ�K"U�gȀ?�����5����b��t1IinD+G.y"G��R�Lp��H����{b���(�y۰^3#"����\2'���u$Dc(�o�&8���[��)��@����.vi0�C	.����v`�<�b����{r!��0N�ln�<ʸW����]��P.Ga�Zp1����
b|�ƕC��uNt��4+Wy��e8?�!~]tϹ�:>��Q4Zgk�6�2����l��zNH�|:��S)ҩ����Q���1�
��1,�@�x!b#�EJ��ң�#Cݰɳ� ��g��K���O��	݄����`�9��E{4�i|��Efh�O0*4�:�I~��@=��X���m�v�P�/r(�����u^e�C�0iC����g:�܌��H|�q�VK��^CGg�^L�G������qoC}����_h�m_t~/��D�t�Qz��ah+'��_{�ro�������K~�_�4�@���l�<`��˗�1��{�g<����2��XtQ5�A۱I*�b��\��I�i4f=��x~���A3ul1�O��Ǔ��>���e)�_�Ա��6����qY�<8�t�!�y�'8T��> I?ʾ�k�60�YzX�L�����v`½ѵ�+�)����y��ݳ/?}t������W9`��v�?����^��铱GS�����Hnkꙍ~�t�{���16�Z�!�L�����9z&��1�����yy
l�ʈ>��׭���E��iO�A2Z���S�.8�&FipJNQ
�e��ۅ �=<{�ɗg�~�e�z'�dGaa���A�Dp�4��s�=_7�6��)Ă�"�X���WlB�⨡�7�4�A�SHh��'��������������������χ:����+�
eV�fCY	���~p����8R���X8i��I;`0vsJԶ����N=V���a���S=G�#�q�Hɉ�P�"e"L:����QJL�Ҕ���K�G�;���s4z�O��ɡ����J�I��3��b�5~���������L�gر�������18?J��e��l��5����8t!�p9������}ߞ���������'��O>9����>���q�D�^�f�F}nM�|��w�O�QU?��9�+?�EX�>}�c����V=��������^����>�t�B�ް���:83z��E>R�=���@�#��K�u�@g�e�9��ܟȎ��i#���o�iC�g�������4�>*�/?¤���I��`$["$Ώ7���NA[�5�F�����/�8����2��|���׿���5�B2r��Sx>�ᇳ����S&)2y��K�I��vJ�/Y��J�!���"�����i+�'�@��P���O?;�կ~}������EF����7<o߾������M:f#B耏ګu�8�'s��r��ߚ��Q�o�m�#���hN���/�蔈�>n��u��{T`�h���μ��7�?B�`XE�$�� ͗8������+ހ�<�q����u��볯�����n0���Z����������O>^p\|�C��ǙB^D����/|9;��e���5MgI�W�9�����Z}�0����q��}��N���ݨSdI���u�D�՚���E$�\~w�=:k�9�W���1�d����3_r�NNE�K2;�2��_���l΃�����y��%�����I~*�}!�g��v������y�(�)��=�O����O����3v�x�lBr�i9����E�q��LtW�2E��L��uŋX�Z3�����������_�����u/]`��vo��������)>`�{p�aL��i&� �a��,��R`Gϗ.����.��?�ȅ�~��.�A�x��V�l���*�m��]�����	ܦ��ӝ��xe/��xY�^]	���~v�������8B�y��PA� �!� C��(FI��?=�(�<o=.^�(�� ����y-SsoHuY~h���T�(��P�5��x�����Ĭn�۔���E��t�&f�e+OJ��p�[�Tc��NB�����g�<�����8���%~�<N%��-����K"�:[�1���Σ� ��Mù���]1��s��H;pN��ky�a���%��1�R1�Tdd��D@
̸��z�7kq>Sc8q��Ew���S�>�}��[����N��'2`��`�ې��*>���ǌ��H��N��N¯��<�x�7*9s/�{�ق��݉�޳���b����_~9J��o�=���4F�3�N��>({���|��W�W�3'L��!�z��X��q1�(����RD ����'��p�z���Y�ȝ{���C�ߖ~#_��ȳ�+��g1����Q\�~������o��)���E��Ӝ�/��b��I�]�fpiN���+��:aw2ğ�af��I�/N&�<�MFÎ����w[<����_V��qL��t��V�����������I����6�u&nO��}���+=���1�?�������}��ZF�`a��LG��`�����q�S�h��_L����������"*D �:|��I���RGF��3/��Α=�!�1�L�92|�!�o:n�s-8D��?��_%��P��S�����Gvr�M��A�Vt8�gqe���@�+Jut��	r�,����/~�n����_Oѻ:��.}������EF���گ~��������F.8a��)��W)��,���\����
7�[dK��K�4�7�8��3���;��s�]��U˔!2ף��݃�][;du
��db"2�KɊ��&
��іe�gsg�u����9�*\��g't��4���{tڶ����-d��se.4�gs�U��K�t�M��J�"�`r��o9�9�&�����$h6�X��t��}��ٯ��ٿ��_�}��'�ю�����g �����-*P�r�\��%7��td��o�&c��S��ڶA�6���\�DrW��h��r霉rI��;��O��w�i��Fv��j����.��.N&�)��!�	�W�o6Y�ν���|=x�i4��J_����N�C��g{\�� � ~��S�p0���b�C��S1V"� ��-u�ڹ� �O��S�`��n'Ȅ�?i�n=������5��o�p��?w�O���컔��(���ء�,�6�9Pf��V�zT�
�\�{=7��gh���t���*)��gwI�u�w���Qc��H��h��z�Ɓ�$h`R7o�xО�v�u~���Uz�++`�Y��n�����91E*�Z�$J�� M����zs���Ӭ�2ТC�9�����ǟ}>s/��	��>����2P�;ǣ.So[2o��y��II3��r|(cƒ����}����)��+2.5d�����O'n�#g&�-g�V�ɼN��9?���Z����G���٭����%+cDAL��=� �◿��~^��U�����k�3gB0C�`�CԁA��,O8�w7C��g���|#壿��a�>	�{9��Z()�N�!�?f�8/�%Y����f�/���������?l��@�:����a��@s���O>������~�_��g�~�M�М�:Aͻ1��� �#02�%��-%�ތ�/X�J�JT��黌�s����m�p���)�_��Wg����Da���όy�	pbo��}���~��h�w����g��u��x�,�,�rK���	�M�`�~����~��O���&�c^���4w%�|�՗��������k�6S�O�C�T)��xm�>P���~���7�u��E]��?�<��i�/F���W�o���%o㿉?x��}��D%�A�j��K�Ca����`#�t��!�I�բ�����"F�H���v��׿N�>�#����}z�漱+*e�6��?���¢��V�_�w?4�r�,YMN3^כj�.�G�/k@�\Ӭ���oG�u9Ü5C���f�L���ݹr�s�s�Q-�B�@7�>�F���(36O[���'��i��I�v��Gk��F{��y�6�wo�*еݿ�rh��=�����tՁ�I�����& �ёf��9r��d���x�w��=�)��0b) 2�+&^�zYG�Y���k�^�M��o�<)�{�������~��gg������~��/���ky3�*JQE<}Y4�~[{�צ��� �n�v����)/8��]���a������K�r�"�U�w�EA/��Wa�頋0�Ff�1�#�p#�z�~�65|If_�y>o�<nޛhу�'�[w�����>�=��5�f{���JG�	��b�ט��}��Y|{���L=��WĀ�H�y��D�_:ib�:��`��Fn��ī�7S�E̱�����o���3�ꢏd§⊎�J�]I9pt�{S�a\G��|������x:�]�&ᘧp��n+�����9�_�Ç�e�\۷�ᩮr<�<����9���y(��q����?i&�I�Q��gpfBoRѯw����2|K-]V9<7.�?gl�)ո8��� ���9u=2.oW_��ܺe9�]�N�#��/���`�`�r�[!���?�sT�g�P�"F�Sad���9s������� �y%�>o[Q�z����нh\4���{9����c!
fΖO�<�>�`�	����"��"Q����̓�/����ƿ���g7l��q��ȡ[C�����,�HqB10�k���Ù;>�n�nX}�y��&��9Y9�&rO�'�e&)�2�^8r9��g�Y���8&�?8�( G�%�q&܇��'z9��&gۮ�q��EtŇ�Mju�u
��&2�hΝ!�u(o���YT����9<g�
�t����E�}���r�Oo���Gz]wM�xC�DW/g�ss?ܟ����1�����|_� 3W���8s
8^�~b4z�κ7|�^���<c�M�o�ߪC�����3R�=�WG���p>zԔ��iO�|׽�@>sf$��1}�� ��3dkr<�j�P�i�
�>N�y2|-Z�=��O���>��Z���n���D7�d��aC�M_��?�^:�.!'cg���9^}Dn���5��!?��s�r���sD��F�pt�O������g�U�0�9Js/-��_���Z|��O� oO�q�^q�c�&E9Z��+|[��[��[����	��x���p��d;���P��Q6��>|e��>��?�O�u~��>�f������S��^�ͷ����괉�x�����������g����_���/�~}���E�M琦�ym����͝ҁ����|�hC��-gk�
���Z�<pvz�OÞ�0/M��)�.�AJ�G$�'����}u�q���?EP�ᖿ�F�'NC����Y���(��	k&�=��ӳϾ�|� (o�1���z=���ezql���n����,8j43l!��i����\�E�z=��o�6��<��@!�#����"39X%���1E�w+����+	��X�_��OS|_�[��������E�L��Twy�՝�^P{&��U��4����A�ۘ���qX7i�n͛A����Ois�FOQ�/&�=i��ќ��I�0|��g%�������qp>�&]��O�p��.�4V�3�w�4�~���jm/���
�_og�.�I���<T|�ڪ��BbO���lz�z���,P����zoj4d@C�Ƙsu�����9%�9pu�k��<���K[���?ʡ�q襐���f�{2��1B^<�r��[M����1yT��uQzW��dWQe^�,i��;^�G|
�2)3I]��:�y��L�|8N��{���ON�N �Q��4Z|�6T��Hn��M*���ȯ�Q��6���9���[�@�I���6�Ȕ�m�ء_D�V���lݞ�\M���R��Λ�z���ۅ�Z0�[?^��}��zo����i�$ZP��>Z�YgI4��Fvϗ?�KE������8��қy�pT�zބ4��$'Ut�|>]?��&���k����g4|�<𖎓�_���+|�)�O�]��C�����,�<gٰ�g�=**�}4n��v��ӈε��l(:�.w�S��7o&���/[l��F{�<�N���9L�����ȶֻ�D8W�1��aB:��	'�[N���?�P���H���e���|��h	-i�����5G��7t�n�.$�t1�E/��nQ8m�ZpsT�����
��viM;�/i�X��u�S�Zx�r��i�����݋��[)/D�9D�oDb�N|	MGEW6�Ч륃#G2��鏣��Ғ?��{�>9��Ϋ����P�z����h#Hc�=����mrC��z���*��xn8q�N��Z����Ȍ.��8�䴲,\��:ٟ���.O�F���zrhU����O���5�x���M������=���/_�lCo;޻s��_=:�?�ӿ;��������(=�Ճ��J�A�$�iW��\�j��^b:�C��q��gT���t��^ė8~:���F��[�ME�v[+�>㼟�H�L`�Ғ֚|ފ�˛	��"�7h����qC��:W�JL����G1�x�O
S���q�sB&=�#%�* I�,�����Y�o�G �8B�ƞw�g�7HR��Lp(e���kK��,��<m��a�b�e�6C�~�-�		�0˸{��F����(�xϜ�g��_��ξ}RO��մؚ�%L�JQ�2�o��S���	��R۱��k�0=�Թ���Hb�p�#�%_��i�2�=E=�n*q6�jN�-׃��=�-ᨓ8j�Q*�L�m
�k7��1���J�b��d���-%�yF�v�vk�C|�ϝ�c~��C|-�^�E=J��x�;2f&苐m�0��O�H
����|k�y��>u�,��q���*��xl/��=2�(�6�:#�z\c(��FAq@�x���9�=��(�qL���a�4�#4.re�vf���n.�����h@yVa��71E�nN�b�|`H|E_�O���i'�n��#��`�	���կ�Jg^�|&*�R^�p�``g��ߙ���5�1�<d{'[{	 ؃CĉsThx��#��h�-Z����ٗ3���#�[�k��4wM(�YJ .ё��6&t��~��E ��[ta�_�>J�#Θ���Σs��J�����]�'�����-��FہZ<��V]�je����E��9C5x$dFv�e���Z��tԹబ�ך_3���F�9G�X"-9�"�����~F����{?�!�h��F'�h�3���� m$�����������h� {KU�O{��$�Y�#�Eg��=p9ǗW��f�N�g#z���:mڣ�X�G��<�u���pXէ]��[jQ{��nў�OP�8m\=�{�e�����32�|*K辗؞��ʣ�fd���9؉d���f������VѠ�o��_����TR�ROa#q��t[l��i��q�'��O�L�szY,Y��ݞ6~�+�>���i=u��4����b�ת<��<�5�z��}Ut����g��_�}�������tt"^�0���t�n��SD����8`�~8�s|Lux��B�-7�&�Y������0Y\�����שg�믊�����n�ػ�!�բ�wr�+�4������Q]�J������7���Wф�5�F�~�y$
W3r����H�3� ��Y�|#.	`���ar�\S�~/`Or<�z܇W�o?%�E?~|j�t!w�a�\�mX�y75�K�gh��h���`��sτ��i�d�f���W�L�����o6�T�����5Ú֛|�o?J��R� ClWR���p��~��p�?~��{��%�D�L6��u�'�4N�Z�M:�N�a�_i�Z�BWW��<u�z��?�5~FO��Z\]bΊ��[�sy�fѺ���p��k��1�{w�7ѷ�e�8)R6v־�ߖ����5T���e���9h��s�9$;�����YixV���IN���q�iH����Q(��;'��"�����ab�㐬f*�,�=��%?E4�G���,w]zx�A�i�?�~l�u)z�[v}�ޚk�r���:F�AJq����̻2��X�L���.�G�]TCop=�1�n6��y7�*Qd��+Co΄��ڕ菨���)?g��u����>g��
6�\�7�u�A���>/�P`�A&��F���'H��<?6mE~�3೔@����{��=G��v(m�|"��24O(�o�yݛ \��GCs��2����8ɯz1�� _u����]Ɩ�Ckm��6�_��o��@{ZA����E��ư���g��[�#E�n�T���I��^�KyL���Q����z  ����}.�!��C{�GNѕ��fDI�������W�O��(�j	o��t��T�*������!�[p�N{e%�c�������-"oT�E��#�C�����,FOΦΌv�C_�0�
��X�H�q$��5j�L����Q��ˆ�,�9�B���`�;f���gEC���3�0W�t��}���=�P�'�`��^��ىn�l��L`��D[G.y�YaFχޮ�$=��K?�y�V��n�v=�!צ � �ҫu9�`�[�䵨,&�Z pm"�����6���ߜ����y���e�^;O�MM �r�=n��|�hU�̭��#���<x�o>��M��ݨ;z~�v�C��ؔ`V>ٳ�\��8���Cs������B|O�F����{7S�}��Ă���n�D���c�؍������O#�<�e��tzcD�y�*3��p砌SC@8R�_�znAMóvB32�h��v�14�,�:aۜ��a�7j�͸�(o��ZA[a�5J��{�Í��y>`@��1��E�(���D�?~��4�����[~9n�b��*¼�.��NP�>�t�m��tu:����e��JWC���?/����V�ݖ�mI��ß1����\�p��U��G��QC޽�����ϰ~��㳏?j(�~=n���]�[mm�w�D/��C���Z��S�b�5��ӹ�����S»-�e2#��a�W�jHֶQL�bPQ%��g];o4�������S#M`H�t	�vz�d�C��瀀ݜ����kN���G�D��Ic���T �&��g�KVEc<��YP7'k��u���ehT�h��_�����j+�9�򦏟�L2��ރ�z��HQ�x�1�zd��<�%^�����]�[��A"��+>����s�x�f3�#��a����
��&Sh�I�HnJ�4�T���:��4ʾ�<����4z�uR�u����oD���$�k��22���q��g��^���Z�`��E��6�@q4���(j��c�:h�(�Ы��q%����8n�OĲkN�ۘ����|�ax��(��#m�T���>����u�u���Ύ.B��0�'j{��}���ñ�h6�� e~�\2�*�W�[Gr������џ��Eq�n�T�L���Z��'
8�=9�+CuӲ�?<����A@>�m�wz��\9, !@޿�`VB0��D˕C�ꑝtfOx���m%��tb���f?X.o�/ˮ��?m~�O�X�`�֣\*�GUѠ�T�~K���܀��؜�Pu<ݗ�+��J��Bm:�L}{��(�n��iv2\="����騜N��g�;�l�z���go�����iώx�6�qq�q+�ů�<���������ޛ����=N)i������Q��:�H�Q��'�X��<�bl�躝n~����%U���E.a�)�t�eՍ�����@0��L:V/����(���۽�o�H/���㰭���/C����{�8P�f��#ST��Ϭ�"�d�b4a.=�R�CEY���M���t��Q%zN���^�����˔����7�p��XBfz$4"W����^y�wS���]���A
=Xâ�y�y��?����ѿy��w?6����|*᪐e�D��u�	�-O���H>2(o��\��.��>.��~\�C��3��Y���{'���c�PN�fy=�$���q�].�U�>���'�RXv��~�%��|�� O��U||^�������՞�ij�������$��h������;F{�6�ss���eab���g���yסz�l�p��?����V�7�Ѻ_��vN) ��~�e�2���` փVY�{���X8��\�i6�s܃��'��4?�eъ��C���E�z�LE#�h�h0�V�MaS��0/�aõ�:xp�-#qk���8�ᵢw��>hy	�yOS�/Ç&D�����[����>m�;�P_9�Q�r/̝Ӟz����.R7�Yޮ�v�^����z���Ѳ�:��-�Lz��zy�P�B��|�C����T2��	�T��v���;����iX�#C�&be�YF�0���(�/��ҞeJ�����L�����6���MV8�3$X����W}��ǾH��w|�(Z�����ڟU�E�-�a��͛t^��0Ò)t)��c��I�([oD��&��*��2�� ϰi��7j��D*��c������Vu8:z���~p�{cњn��G������嵎Zt�Ρo-�2߾�q�V�J>��K	���Iۍ:�s�u��ə�;������d�gMa���^����	��_��DߨH߈��k�7���[w��Κ]�_D~� �dI9of����Bw���ͼ�>��:���� ��:��̓�QeyP�{��j�t�h�D�z��Y�g�t��x�V���\.KM�!t�!k��=ن�|ܜ�'�ܵ��)�|ie������
o���a?{���d�H��ޟ��W!	�I�C�Jd�Զ5:��@S�����u䀥�;���TZ�/�)g~Y?��� [ͱ"�3:���oI[&��O����볿��>Z*��X�ˇ� 9$3��~pv�/��Ȯ�&�C�>���Ӷw�F�Z��-=OA�=��ߌ~eVƣ��4��a2��I�ڀ6a7� ���/����љ���6竓!�Ute�i:*����sc(��h�5�$,=Fm��Ÿ�8M�:��Q~�G";e =�EVAv��z By�R}�����<xԐ��1�H2�FƉ"�U��/����}�:'�U_[����� W���(*�́���o�[M�|�_楃+���f2���>�lX�X���K�
��u�ypW��_����/��r��ӱ2*Ly(�����W���4un�Jxʨ�mMS���Z�qZNһY�53��|:^u�F��L���W�oQ��c���M ����Y�e�5��l�nz	Ex# \� p�M�t΅��m|ܫ����^A�!�@��=�M�"� ?�f4E����gWf�z�7m^Z���h2���9>]�7r�s�S� i�Pu�{�ΐ�9��fF��a�i�㈝�((GKdITEٳu<zj�?Z�&��޺6�[l"`^�6T<�}�!"K����|�ܞ�� ex���Z���-��x�9V�3ê�qf^�{Ν�s�8ʥT�_����Wԃ�W�@w��4��y�[�����U�I��HY&�+�u���RP��8}"BO1�m�̲�:';�GGu��u�:���tVa��'��"݊N���Lɔ�����4D8M�F�JY�un�����	Oy�[��t"�^h�&��&W���tV�e���e�h-���Ot��Pg�u*�n��ӡFtYG��v���!�~�[=��n*�v��SF)� v;Y��Jr��^�I��0�ED�s�j3���}'%=_��W��z�V�ݢ���7x���m��T��';W���|�(Ie-��jy�Ǽ�UzQ�ig�R��Y�t�9^�hdl�����NP0��K�C�'���t�˜����|b_N�8�*���?g���KQ��X�����^�v׶9tzy��12F΂odgj@C5mmG�Qxȧ�U[m9�򼏱-�.1�O���	�ϛ�!2f�#�/�o��l��~���_��g9�ә����e,O�H�a�߼u�����UJW���3`�u��ls6�p���nt�bGr�w���sp��
`���<l2��=Nmt9��3s��sL�zQg��:,�P"���ypݓd� $h�@����CcRD� k�,���$��Ǒ%n�O5z6^vh��,$�Q�����:�SJ��c�^����;�R�6�`=+�6�`kbG����Q(G���y?|x��֮���>��AϷoV]4Y��ư9`��F�-�W��҇�(��=�]�� �89�zB�E�i��sh3e��CUp�����pH���x6��?ʎ��M�SG	��G����kR�g��� r���<���}|����)���0���h�^�ă�,�SN��`�0�����m�����o�r�ZC�w�^<�[YOϾ����V��7Zj ������%c+Z����0�����"8�<�0,K��-�	L�1^R����\Z9�<]䠉�[5���4�G����D!��c��p��{�ބ��$�J�x��ψφ ���%i�Ό��놟r���쥑�2Oi���z��������\�Z�w���@>,���1\'x�"E �]���L:��dg#)��66K#D��&�W��h.K�Ȱ��k%�
_����.8qp�� �@'��s; 8;�0�x�W<��9�߶�yս1�'�&/'�[�޾�X���y�����96��11�����L�m�Ζ<�Dƴ8��^S(B�!H�>#�E�EB�W�����n������ϓ[9�3C/��B롵4é]�չ����ɟ��  @ IDAT��^�6��,+k��^��<Ap�9e�-њ���p��� J@ε�aFx�M�s�9�"j��x�3���r�C+�Z��h1pG���{��9�	DN_v_���nB0�����{���Y���h����� 6d!�[������;E��s<;�c�C��=�萷R����7�*f�6Њf�7c^{(�e,�N���=����屷}�nu�+_=�1��?��G�$I����M������]A�
������ f�g��N����C�c�d����y�anfnfn~�g�j$���ԯ_�qqW�����A�^�O���{��2	��D��w���8A� ����#��ǢѠ"�l���k .��';YPz����5>}>�W_�:���􇶜��õ�:�z�k�:	�Z�3��wb�,��C����nc酒����Z������ݑl��$~|��t��T(��;��e�n��ZSf�l�3��5�]FeGG�d'm�w�;K����N��D|�tA�A1�"��.�����#��ł��z�s�,��َ<��h1/��g)��BQ#��R���JBb5"n�Ր._鸌\y&�fZ�%�[a�X� �/J�ҽyª��y�	x*=��u��ef�ʷm�ix��˟bj�77��*���2�P�a �����;��?�V��^�l�b�'��_�]�/Z|���,��MDTZ)��{�y�VN?�ڲ.�ɽ�£Z�zn`��5�)�dK ��J'��ӂN��������ڼ�2~B��zgM��'(�wm-���h[O`��	13gx���N��0
� {��6d5�Ќ���iB�8s�A�W5k4���x�����}'�4G�ׄv�N���j���kT+/���t�2){Q�_1��{K�1v̯�bszD�����G��Z��w��g2kq�(�9s,�zZ��E��x��54�}�%�dm��.<��VT�_=Os�V[�ZHp�3����FX���KQ���v#~��7�:�[����8Q���,ϑ) �H�|<�M^^���<��ӻV����S�
*��R_��)	�.ց\mG�H�a9g���$�exQ�y�FP �����c)84A��P�ҫ�������I�f�;1��<Ac��N|F�i�D��R�#�2����H��)L\�<�K�\2�1��C�2�!!:&O������fէ�����E�O!�X�hĨ�ghx���{M�^eAqxx���9yCc�����m�����#^ETN|�G�=�7<i�bm'd�4[J<l~�.�w��Ug�V{Ӟ-Р/"~�s:k�i)T�[�������O]�`�ho���_m�7�SO�+K�g2T�	 ��{�bgT���ͺˣ��� PBمoB�{_W����g�7�|��ʣ��}�;yη�wrj�3�:[�.\��z����c���<+�x��G�5�&�x���-T��g���t^���u�S��l6Y���d��0�tʴ}��g�,�ŏ!c�ą�{�֧?�v�xK�bL�O!�V���
�:�Z������|��i7�uc�F�$J�z��A�?�^�x~[��
}�<��.9zL9����<�����F����Ȫ�]��L���FeJ���K�V0_m�dz�В�tv-0*l��x��l�:�y���\x5��lVS�U��P*��VzUJ�3 T6�I��U��P�D3�y���}L��7_α?�x����t������Oy�k�]v�aN����7h���\�a`�q���w�w�Ň�����)���_be��č�����)h�!n8���J���u/��u�Z	�����U��KGq�{��p�ޓv�1�{��z_�zn����M0����q��͏p��x$��m��"O�w΀�i����u�fy4~�/QC���7��^�Q�Ѷ���
KN��Ǽ��\x'��h��-��+����2�����@�f:
�b�[���s<�Ќ푧ō+:!�7?kݗy�:�2!B���+������k�=X��'�׏rc��(OЛD��!ו��eg��E{F�.�V��� w�̽��ڟ��	��X}P�4��Jӓ�Ѱ)�i�*������0��+m�P�/��Ã� �3���8�ȁ!��1�)�%���M�����N�[�����hI�}����!��!��[x��?�e^����k��7��������6��:���B�ߌ4=&�xA>�#���e�^7?�<��b+�4�ʩ�+��l��զK��^����Ɉ�_n8��6#?2�^gH?k���m��&,��Ho�adz��V<��56�n<O���Z8Ѧ�я�����^��!%ޮn�g�Ԓ���*�Bu6H?���𢎐���>��d97�}N��0s.�{v��� �c8���t���G����G��)cW��������9^O�����o���r���=ѳW�{�C_�2�+q�xuV���C�<|�Hm�߆�d�����'/�t�����I*m"��N��D�����_��`��ޒOp5����ʂf��}�=���H�yߥ���ˤt���L�H[uB�E������ޯɣ`�N޹�G&k99�f�Էhޕ&�w�7�"љ��'��a2�wL_
 �Hg�~��U;/�;g���C���1���]�s���G�O�W$r�θP�xEM�޵1�M]�v���O\��i8�;�Y:�%鰂O��p��I���SvQ��i۲Z25��. �|��0���xCI>�>��z��'
/��y+u+�4*�	�z�,I^���c�oQWs18�����:,���\6 83�4D�����*�u.%�2��M�7��R��u���k�ƕ}1O@�[B������)�+��w�j�[C)ܷ�}�~�}/⊽j��~o�M��ß~O&[���F��ӈ�bxV�e��Z��G��r4ʓ�����;��N=����c\ɃuTc�R��7�8�'�|�Ĺ�����w��øФFs �߼��e��u����ѕ@��xb�"�b�sՃ�Bߵ���+I8(]Q 9��M�5�̀H\N����h2����΂��y{��܅��d��� �in��k9z�e�QW����%q	��kl�*�nQ]>��˳�0��z�j���y{7���D�U��V���v �i5�V��-/�7cD�nF�eD@2^���!�s���a��z��SN���
�c8�]˵||�o�]�Μ���c6Ǥ��c5G����x�{Μ�����@�P�����(���xo�@[���;?���g�c�xt��K��lm�0B�T�<�y�̝��Ë�f�}�W¥�ܵo�X��t;���~ojWd�H220��b��c�(�*g��c��ǈ7A~Vf���4Z��w�?�]P3��)�թ�!��jH9X�"�_Õ:�+�V����	|[��Q�� �c�.�F/
u���szA�^��9E9q}�~h���+dw�w�"��Ŀk�B�|��n��x�Sd�+��x�,�`��,�(��z�6kc�~zky�*���Q�o2`����p���Ãǭ�{À�A�Ne-e`���<�A�̏ӧ_���������~��	<��/�e�ֳm�!��)ܮ�KfU��+�����y-���_%�W1�^�V��\��1��j�/>������@?��Ȏ���Ad{�7��36��36@�v	A�:S��VH`b�c�P�~I��&�2�[�������jm��E�.��K�W�a!�Ȟ:�`Ql�g��:�7��y
��'XJ;�ɴ��a�?���UhU��� D��u%��a�&���f�z6������m�P|�V�`V!: �x�4B�4@y]�A��>�n��8�/�-�K�&��F��Q3�C��UXz��;J�F;G_L�R0\���E$K�OF%�g�UwVme�d�,j�8��o8��8�R����8D�)]�^B_~[�[�)bBחbo�x���:���}/Ҽ��z�������׽�	��쇖�$+�X�̷�}�x��iݵçp˼���I��M��k���&7�h����I��sa<�8�4�I���%����Zz��|��sTCC)\�}��U��^�<����x.��P=_T���$��O_gZ ��E
�|G�<Q�l�ק��7M�Vx��R<.Ao��z�<m��ö�{iur�2����üJ[��>.�g$�)�w��-��b�lg���г+�'~^�E�()CL�a�0*	E��->зP�2vxƀ�K`��[��� �Uq��a�
FؘOh���l��Uo�����
��;�'�frl�]��%�gy{��#N��r���E����P�A���jOC\WF{?Q��I6Pf#�F�E����o�SEVxt.�~̍�H��R��72.z[�o5���>�4 �Mm�Cr�s�v.���<�kÃHA�m<�&��y��x���%+gn�]q=�W�{|ul�3j�9s�2L�
W���*e1@f[O^:iyx����;���䩍��Ld���R}̵�O���W�5K�q�>hd����\���䐡ig�)�M8�r*��^^ v��n�Q�A�ۥ�b|�
���)4�=�G?ٗ�ܷtT]��s;��@Fgx$���P�E��7�,�ox�q^�n?8���٭��*�9O˛d��M:�Y�f�&lA˺�7�(gj������ޣ/<�@�6��xK�ש.���<��\�G�<��V?Ӟ�1;�J���-��ׁ!�^�^u}\~d�O���2���F�����7����� �`*�ksgh^O�[)��;. ��7׎������q~|m?��e�����x;���cB��7�L���O�c��#�1��xI�~@0�a��P��:����`��>�u}ؐ�Z�CU*@y��
76D	D0œ�e����fxk!	�f�3�"sDqg5מ
�(HW� ؉20ŗ��J4��<�I�����`E߮�5�����璶���D�Q�ϒ���`�I�A�[��j+����V��ޗP/��)gpN�*�=�U�8����>��"�y(o}[q�e�R���2W�{+��X$�{\��g�b�5�A�l�۷�'�nd���"E�&zk�]���w�uƃ�<�6�x�|���N� ��y�l
��EO��4$%�<�q�WWS����_�=��7tL/�������L���:��׹��})��e���<EB��Q��م�|(��"����\�#^R�=]A�rm8)��6��Y�L��f�h�!�1�\Hi�� {gD�0��g�˟��<�_��͓�m����b`�l��A��X���-�HI��ݓ��_y��ז���(���1��#H���I�'�[g��ڳi~����W���]��p-|?iޖ�<��Ù��63pj�hB��/ʋ�����%���w��-�BS���m �������w�ٳ��1\Z�_�I��ޙsX��Y��^A�����:x�)�	�z����慰*/9��f�:6��l�ݾ����ɳU�Q��HNC�nXr�-R^V����9���9�E[�]�0��wsT��x��_+���{7�։��^�b�=+��摙�V�ħ�Fs��2F��Q~��1S𧍑)��o�Ca�l#�;Җ�����9�M����e8k����U����͋�_�3�~����hʘ�|F�w��S���)ޫ}ŧE��^:�{.�uR����x���vټ�?�#�S;�A������Ow���ۇ��x��7��8�����UO�(b�`xD�X���C�%l��9�y���NN�\��������Ԇ��f�kE���Kw����L�H�Fp./���*h����V�t���x%Fm9r�Jp�|�K���y���kUi��!X���N�NnΑɤ<�ujME�*nu�/ؘ�������6���ܿ�!�cq���,Ю�a�2=�g���,�3�+���(��,��ˢŔ���E��/�Z}I_�~�V�&`|�
yj�{F��>U�ӌ�WD.9BT�î���wē�c`��A6$��h��n����	��+33�f~ΪYq���ZM9�B��l�c_az]'5\ʑ������8'rV��8c)`�L�[���U{u\�ڟ�q��K��V�ar/����j�t�k1�^��@���CC�LJT]��BJ+��=�?�NˉW�`����ؤX�ŧ����S�D2����㏷����_}��j裭NN��.�s�{�-�Ye��L���J��#4{��{�����P}���Y�w�{���=,�t ����|v�j�d}>�D^m�����9~?��c{i=������z��@ƌ^��<�-F��~���׿�]��5~�
�V�)@��Ue���e�i��o_7��j��O3L�?��~���z�D�c�S��f��k��*M�;�!�{�r�$��6���������?����(�*҆�R��mg�{�fxВ�j;t�	�G������߷BCg�����/sk�i;�	?&�7�+��!W���)�~������b)��)E�=��w�e`f8�P����6ߵ�퓩3#�I�ڽ-�ǎ�2�'���n��s4�o���f*c�.�9G�"�W�����9V�08���iRF����;C�o����w�E%/Ç#�D���țt����<6VD�흧�y�<o���&��
��e��筤���أ�my�}��E�yfv'�H�7<�������mx�zy����B�{<�C�~�i��dT��}z��{��$=��ɻ�!�cLY�y=~c(�/��~�Z���B�<=p:�rr#��gm�J�����9������w�NtȠo; �۵�Y�	+��Q֫�(��f����ܶ0�����V"���M�'Ω�}���7���s�v���މ��0*�C]{:�3�6#ۥ�`Y�B�%GJ�{�0 �ē������χ?g������m���c�2�t����ɺ?�U�^�	���í�uo��9QN�H�⋷ޅ�k�-8��eF0�tL���%��"pG�`� ?�MV�iGu��jҕ�'�iǳM���G����d7C�Q˩�Fu���|0�M������YH5�#ˠ��'z�P��+\�-���9HҐ��Ļ�G[�-���s�P���f�9������wt#�bM�4�6�]��s�pyzu�A�e����;E��oE.�=��4��{�D���(l�|��
�j>�1M��oҕC���+�Lo*��p����M#��oemW���>��1�W��Wq(��6P�K��o��ozP��p@���2��\����+������ك�g	��<��wS�-Ζ��W٫�J�w��ޟU�d��-l|x�7����Y����!���d`���/!5�_)�1�-SQ~5�R�%�s���Ǜw��^M�\JA22�6�T�K�0� �X/��I�XM�}�&���S�}u�ex�J�%?�5�<|Qv�#��he�`���v^jX��6����5;u���83��҉G��mx~�Ԭ �Y�Bz���+D~Y=6�4ρ��a��U�vg 1��c��K��yBx�8*�p	�I�SJ�v���>3��W��Qy���e"�''�I�L�4�4ˢK?£ZF�c���3����疥��C<�.xO�X]��覃��eI6ޛ�-ђG�B^;Ì%\
��a;�!�<��;*��C>V&/
o8��.��[%{�4xxn�>��7�-p0��5��i����~�$eP�o��#N��$.��r6q�v<�hx��k���V����`x;|�a���./��J�;��x�gZT��qlm�W~5H���0Ʋ#X�e��u�W����L=������$�\Lǹ2��ByP9�3�ѡI�CF��s-�����]ۧ�!#>�ε�r[μ���]���R^0k'��,�H>�K�2nyH������7|�D�xh��ŋy�����ԯ���W�c�f�>���:��jx(t>iԳ��
����fϱx�1������u<[�׽��M��yo��7��׵�۝��׿�t���;� �Y[�	OxY��a�.�.5W��_ř�+(�W���;��?\�>r8x�k|:����&r!Y����ԯ��ɞ���X�2��҈3S,��� �|7�M��d��"���Ck�Ͽ�)�1�Vf�ώ����<�q�{醮U����\��V���7����{a��ӵlx�J	H|���Ц�4�_e���@�qζ�U�s�'X?\A�!p{� X��X�`����]��� P�!�����2����5.B<�ӅA�`���+��ʚ��kr��+�<G���)x�=�A��/�BH��G���i��(����b����3_|����w�U�)T���ɫ[����<�oo��g���U������`�21���t�'���-���D�/�֕e�r=½�2Z����}����ˋ���A��;F�T���������ӝ�?��L��w���Z�p�ua�}�؞:6�#��l��x�U|�Ý�^<&Hʽ!筽Ϛ`��$�(!��Ủޏ�͠����������F���o4l������~>=�;w��4Îs�]ϵ�kQW�vi�&~����ܔ�L�vϐM8[��>�!SHW�^1c�U���rܕ�����%=��'�>����#�"C�j�"Y��C��eh��Eo����7�>o���+�ŷ�Z
�u�|�~��K��E�0^�g�0�w�W_{���~s����!O�����k͍���v|�T��4�EL��}�`�R،�o���o~����[yj(<�pb�Q�����շ�b��+̍�y�f��>������N1*�4��i|e(��<O��H��4dF�������~7Jo��<�w#Jo�q���]n��z��.��#g�v!?����ۯ��Ms�6S��FY=7�
:0����d 0��ǻ�	#7o}M��[t�Ϣ����K����=k8H'&�ؘ��]����&Z���?3�l��M�2<l_�'(>ô%4�i�m� �����:�S7�����V;6��I��Z���s-(��/D���S�5�j�.�����Ra�-��a�K�����ڃ������Ό��!�U^o_:^�}�
��e�p�9U��ny>��L�1u�f�i�1��xI��(}�90�]��]���q|Ҋ�/��nqAs%���@��#{�#��BrR�	��{��of����^�3�+��^��M�0��CF~6ɴ�����HK6��"����4<8�ON�p������
y��[�ʧ�����k����"V��O\s"�v6�ɍ��ȧ:A�:�`��x́=#\��~�F��l]���/��!�x�cz zM��w�0*��� ��b�������Υ������ս_C�2�ɘ����n({�ҏ#f��s��#�Zϧ~�&���Õ7A�����	�*��� h����s�6�������DM�+��S @B�5����7���?����?-h>K�ǚ��Ϫ�n�*���dl-�)	X�1�;A:+~@o;�w�I�!���Ut�F)� �w���뇬l{��s���Ğ��{�G�ʒ���4``p�����u�^CW|I?�7��|���znUF��`6L�������xϥx꽫��f�@*p�߯V�S����?�%�����KkWl��z�?w�L�1�������r����?�l�'�ߧ�ϧD�g�S�`Ћ�yi�K<<��z�wv��;��n�H��D!�(Ey��63�+�6,��C^��;��V�A~�dpJ�Rb��1 _ۘP��"9�d�I|���C8a�\���d�G:��x�ΜyNy����G�:��/[J�i��;jCLx�UB��͍��9�sv#q�ޝ�&��M'��fq����> ��'� �I��p�����ލ�T���f�x��JJ���'.�����m�t�4�.^g�5���_���^G��&�P���^Z�MஶC��g;���1y��7� �Y	�A�ޟ\}>�a\�� 7�����>�]�D���MSD׮��aa�o���ݟ9j��u�9�NU0'�AH��)JI�dZԭ��7&U^}�^��	�xFԅ�0������;v%�7<cҾ��-U�]o���Gᆗμ:^Q�M�
�e-�[u�#���=�x�LX��E��!�:�U�����F�{����?���ڷ��f�P�'�6i���m<ys�E��=;��s��̳ʧ�6�ng�����l<���C�(s��:"�����C�V���[y��
��H汛��#���<%I���%�%�3���'Ɍ���7�#��K���/o��$;���|1�|��K��g���lq�t?l���r�0�ǘ�ǩ�HE�?9��T�ʛ�����*��$�.�v�W�.8.�<&����?��p�g��)\�BIƑ�m��쮹���_�o�E)�9J�d��2�&��a���f���Cs�^��1��|�0>�0�2��Wz���	}]�1���N��&���~vMpOI\�0+�������(���J|�QVЄK J꩝�e�peo�"�����וh����+����l���VО�������v9���y+ă�c�A�'4	�a�_�1���ꇏȹ_B�~Z�Ɣ�q����q� o&�����γq\>&RJO�hY�1ô'�C=@C���E�@�θ�>��|�>�޿a	*cp!W�D0�R�zb^�C��+�|g$	�>p��46��"�a1B����3��쁭�%��!B���I��6�$����|&���[N��l��_ꁚ�b~уxԆ|��3/'�5p��}�^���S&.��<�����/��<��U��Kך�������< ��G��XX�f������oY�l	��1�_�s�>��N�6��4c��a��`h�
�z݆�����b�瓳;��Lަ��;gS qԖ?�^�R+�:כ�c�N�^3eD�~���V�~C<J�2<U`�6�i*�9`�U���8�6Ό~��l^BJjm��Q^)ꇏ^����$Y�-)��ӳg&�;K_0p-Bh�H�����,g�Y��|V�w<D���DXaz�cG��/g+�dU��9���Fk7A�#�Æ&��# �-��g�(�����e0���D�1���Eyu5��P%��(|������A�Z���?�T��1:laJ�1K;��Û�e���ɐ���Da���h��+�v7ĩ7֜�汼oU�q|{��w��Y�_Ƹ��e�0^�k���^^�7!���2,a&�?��v	�ߥV�k��g�?�n*6�J�ǉ�`p�L��q�9T��h%�qv�ŌC���fn/��k����ps1��A����ʄ�`	N��.�Nش�i\Յ��������W���e> ��]�;�H�-��]�oa�Aɣ���a���<c�*�3@ߍ�+����o������G�����2�r�u�z��R���<~F=�f�=�-���6�Q���N^u�1w-^w��g���P<�o�
���!L;&g�=���c���P��������2a�B���2B�;����i�7Ų�I~��P�l^jۻ�<!���
�$K|n�s����'#���0�u�b�i�>�|�w���V�����AA3��G�&�w��������y�*��߃o���ˏ���?���nzG/zr:��NK�۞�d`��{���6�
��춰�������MN�d�ߑ�އ�
�,cK?�����)tKq� ��|Zf�.�-_1ֵ�#$�Y�C؛kCؘ�U��\��F=	��ԓ�] ���������@�J��]��r�)�
?�懀y�aqda�b5x���A�-:X%İrI;�))��)��+Y1jx6��)�V6u^�&cU�Ty<ӘT�b��(r[Jo�ͤc����2ؾ��{��|�\�Z�7+��V4=z���׆~��u���I�z��~�kۄK��[���u�#��X�Fy[�d�5�ey���j>u-�x�9!W��o
������s�@j�E�>�£�H������GyF�,Q��)-��̩���^5\v-��$}��Y1��!���<@5!4Z�2�'�=Gʾ�fqy�ְ�{󄪚2��mW�ks�MBg����=+����,� ��6a�m�Q�������&�S��x�R��1���C#��x����f����91Lz���kQB�����$8T�Rp8�_U_[�G��+�~�R�,F�;U�Af5��6���Wn`d�^�i���Ņkˌ�h�������5�z�}���!���?�<c7�Z�hq�󼓭3,�M��ܚ�3�I�ʱ����`��Az#��	�ku�"(/#U��!�����O�嫃!�M�J{b��G*C˰����Ð���~�kTz���w�뷠nʋ�6��[��[C���=�2*��k����=�?��Q0�[�Cn�L%���̼P~�4-�t�o������u�����������Xp5���\<�:ZX8�$/����b�B�(���N�p|n4�t'��E=����DTv��W��[Rt�`��Xi��:\sE+'�����xD�d )aڬ���)����쟑|V�����I	�Z�Zt&?ƺ� -����o�	���-������z�>lמ�ϕ��e=�<'���E(��m�i!W`+\y�U�e�y�������h��?z��OPVY2Z��}����2�8�L?����[u��@�aƈe'�
��}z� �e����G�N�_Fa�0b�"a�.d8%"�oK�#(�w�F�;�E��}u��������{wA��X��6	���\
>P��5��,�JF5��ܼ �FR2�U���os��H��D�XI��5� ���L��;%�{ќ��9A�? @���o�~scN�Z��z��Um����H_4��O�f��_����M�=���8sC�T`�ں�in��7/�f�����"��L�~<��QG���p8�c���x�n�.䵹�H��N)0�Ëvd^��jd�tp:C��~"
���qsK�Ѥp�xM�O@���ke�^�#
��8�[�����9d��<_���7�nc��X���p�R��vګ�UV[�`�]o8n�}��<�S��O]�
���E���AQS��?1򚉇�	v�̞Z)9i����oP�+�Z�F�/���ۤ�7��e��RF���e�	#;�(lt��/[Ug���{Wu�)�Z��fֿ�Y=�����ĵ�2m5q��᨝�y���2\��_���.ϵo��}5F��Vr8Ԝ�������;=ó�#���I���i+]o�|x�駻�.�1�A�3L͝�O�L�/Ɣk�-�7��u��(��N��|�0㓌����kf���-��p.��ʖ�j-�,lH4�M�z�ǛW�J�ex���.�L���;���D����#��ms��'��=4��$s�{��0��b ����̘74��a�ވ���Ml�a�|�Oqд�7/3��<oq��餕��q�_u�᛹�y�f��ȟ������MB2n$�/���W �_y�!܎���v�wE�U��w�Lɭ`��x��R��:�:�:s�9gr��?����.��7������#�pm��LZ��`H�����}�iY-�d�90�I�*����M#0W K�q�*�f6��L����I>L����+
N�dCi���S\O�g#80 ��x�?L�e
~L���&��ׯ���9���i�2����c�l��Q�Ӡ�_d~����|܏n��D�N�/�"��J�IT|��r���F���J:E�])D蚈E]Pm��/���?��Ϫ��>l4�bKm��>����C~�/�<��ą9��M�g5�E� �:��<1����{�tVL!�ɿ�<�l���3Ê��L��T�]�d	�����)�+w�K��e�i��oF�wF�,��q)�dl�S��EԨ�4��E�B��|��{�Ќ�]�yl{	Wsq|��|�Ȁṡ-��]�@�95^�ʲ*	%(q�;�Ȩ&���N38o觞-Ϛ93c�Fυ)U�p�̶9�d�[U� ��c��U7�D�gy���ҠN���ee-(s��o�q�:K�y<�rsI;�/���!���N޹���޷��f��(�6+F|C1.#h�}��3Ų�!Zu���l<yS���o��ق��Z��ɰ�#ޭ9ʩ!D���^Z��Kby��������W�����`��Х��3B��t4O�� E�%E"����~f�Fu���(�?�����p�^c�Wf �]��b��;S���2_��fd��<�3h�~��.�˨��y�W<�S$�ȃ�`��Þ�W����i�y��Lɔ.�����%ڍq[9㙭��1�o�s_��A�'��	��D��.��ⓩ����J�S��w�om��?�a�%���E�������^� �B�p6X��ys�35y�|[r'�U��jk��v�x(�	�c�4��lƾ����lh+[=��g^p[�h�-��1�P%AS[���ؕ1d0Ad����Y�8���n��l�O:��GpT��KC1~��P��&M�������J~Ƨ�#SV�jɮ��vO'���.�y�\�)�~�=_g��&?�`hV�}����5�0Obq/d�Y�1���ˁ G�Qm �,�\��?��
	�����y���T�����g�߾�I���O�F ���\�����Zoc�H|����?b��Z�3{qV�������äH�TA���p=���I0:�{��"��/�\��*�/�b��
	���y��%Pc�>(v-}7/�j���#4�<s�j�V +z/}Z#B����UӍa+��K�4�°����&�7\��'�w�션p9�5��oa�g�&j�Y��ө�r^�9�_��S6�Qc��佰WR�n��4�}�k���\���G��������í�Әδ���%�1-��A=�W���J^1��,�[뵇�E'd�&�ϒ���bk��[0[�z�r���;�|���M��U�Zu�gk	�i(M�ڤоQ\��I����I��ma�2��R�'g�UIl��_ɺM��H��7��׭�C"��|C
�E����eH0�g����r������I݊�H88�`c�0�>i�͍�t�<�s����GL9G���#h��@�����E��r#�Ϛ�4�#8G��=���_�Qw��C��s��qr\G�W��j6{}Q�c���#��1�^�Ng!�j�x���O[qw�{N���nJ�E�xQP<0��U7D>=wHV�`���q���s2<W�V̳���x�v#��x['��(����҃y��۶����8��9�8m����;�Y�g�6�2�ު=m�s�W�0R/e�80�u�����~\�/�DB�{�U�9�Ӻ�/��?W�g:�����#�G�)g�����ly�����+�����Ջ����GT>ꏖ�(�e�Gm*���v}��^��ݜ/��[Da��U�,�w�ܔMo|yƦr�+�/�x��L:h9���a�Q^��˃ʘ$�H����!�h�w��U��rF-�9�[�.2�bF���<���H�����&ry��,�7�+���5���e�KY˸݌�`���{�-U9nu��/ނ�<�a�>��h�ۗqj_ܳ��e͛]xW{(��+���Wߙ�Ϟ� ��d��!v^*}`4E�+�П��m��>�w�}|��ζ��`�������e3Y�Y��P��i�[&��d=�^ͷ[GJ!�0J�\�#����kC�G����^["��z�4=��p�=1L�Y�P��Qp�8���b�ʑ�8�1����o���k����h ޶Ɠ�#p��qj�0w���a��O�1{Z�Z�m�ߪoY��/��K޻��SxZx|la�S��obcɤ�.8��e6{z������߆ f��zt�P�9]#D�r4<����{q�a�}t6�'Ah�c�Rfزx����	xn�ni,���=׼�+�&���lN��>�������8� @�ӈO��ፁ0��
#��fDY5�NaX�͞-*�7�<q`�X�a�s�0,��ſꈾ�n�<�,[����}��"tF��-�M��=��$a�R  @ IDAT�_cޅ`@�)C9n�%����yG�N*��S�|m����q1C�0#z�$���G%���{��2y�h���x<�alS�VZi�P�	���MΛ�e�G�f� �c��ͳ��l�S8I�2*��V{�_��V��.�iU"޵ b:q��8���WM�~�����Ma^]� ���JgsU��7p������S'����� ���M]��[yɑvVV�Z�c�+����@���GTJ�܇mF���&^�%�����CC��1�Ѽ��ţ�l<��d2.�?T���&��g�C8@+</�?H`���eU����^]K���s��;���f�yã�ۣ�o���L��V�c�&�M�W�`Hn��vA��k&;O�[�~3C�+_�U*ru\}������Y�r�/��v뽰Ֆ�6Ym��+���5e�D~k���n��YL�JJ�5,�W�7�C_��q_#+��
ڢMR]���I�޿�QlSzAᩚ�� xq�k<0�/5�<'�d��y�E7�l���!憺Ѹ+����(�,�۫��x�<(��I�w����2��c	�F�4E��c:�S��&��-��G% ��[�3�tr&T�/�Z�^q�U�)�C`Q��0�" �D���~/�	(�n�V\�>q�|D$U�H�FV�iS��+������ߏ�!L`]7�����}�p)~O��~ ���uK����a�*=_+k�^'1/\1�M|��f$xV����r�-f�>B\�$��f�t�[$p1�{P6�O�3�T�Lx���B�������{p��ҙW��LMN�w��9�p(+��\
<a�o����0M�=j���hEҕ��V�o��#3W^�O�k�	��?���ʌ���oc�sdÁ��QC<)��wU����*���}Dw�;\���I ͽ��EWl݋��U~��ad
������6�C�Ջ�&� ��[9�C�8����VVpZ��τ����.����>��Ő/f�C�G��eU��^�d��l��0�z�^0@f�#>���O��9�O9hG��#����5���_F�yN�TY���(��]��
T4~���k�#~�e�R(�0d�I<j�ޖ��k�S��+�V�1���Rγ"�����y^t�(�̚�9xg�>�(���o2�.v��P��y�3wz��8�Pg~	���v�^:�~.��w�A��PD�1��-���!��z����ˑ^e6��Q�i���D\�C��x��&�@8��Ъ��sV�GF�<��<V�pf8W��?��O�ou�xt��-��;�D�i��\��<s4YS�í���ކN�,����k2h�2]}7�d����p�Р�:�.��v�߰^ւ=ǘ�.C�>����M���o()O���b��=�_����
�䌰1�õm�f89|��!��ph�̳���U���[鵗�����嫁�:^��c��<�Y�٪}m���v���ןZ�scd���M-9x��Qe�G[�+�gi���ڊ�Ņw��5�E���"�ic��W��x9�'L�\<�-�x����N̳-T�����>���
]�����&�� L����3�1���@ܘP�ex�M�1l�i�3��U~��L�	+��W>{;����-�4��y\�5ď �+�A�w5(�oo�v�i<ðꭞJ\���q-�3����c����S�� -m�!�(4R��ַȫ��l�W��#en�O�_g�'z�SL�7^�`ã<�V���o8��E���� ����z���F7����`l0x <�Xј�f����R�I���j|gg!|�����^.��������zz�o�be�EИF�hT݃ѡ]r�
�'�\��)���C5��Ă����������;�̺�m��1^�Fp3��g��	WZ6��7+.���"XU\�z��4��߅�Q��� �f��j��M�U�~�V ����<c�׏�t������ =���4���!��c'�݉9x�al�+�aZo��憡k�6��ӌ��k�[����2�X[�8��I[Q8wr&q��US�:�i�r�|(�u���e�y����a�Ճ|��ɐ[xE��6��FUmA�M�I�s�R�0�l���*�W]����#��e���e4�&nҤ�[�,�����sc���ʼzIG�R*��~3�.�"�S��W�!��Ⱦ>T^���]l�A��k�I�3�%���j>��%8ۍn�:0�m���7�?߾�a������#�ȴ�d��y��V���<]xj~gh��8_�#��{.ޛ�D[��z஢@�t�K��w ��d�7Ͻ���Q>�.|��|� ����C뤐�0�p&�����Vi5����&���6�ڡ"�<�C��Ԟ�:qMy�/`.�xCA��
�Ư�vI_�n8>��o�S�Q~�����n]�|���[�� ��N^�_�e5�0����o�����(����W�_�9�� l� ���뚰�`���w6Gʪ�e����W?�c�V��xp�=���}���S@�@N2� �*܇U@�%M���Uˠ�䀛��bUr���n V�&��Y��#���TᩘJL~I�l-�F ̷���v��WeW�����
-AR�N`C0%cxƒc;��yg��d��e���^fL37���X���#x��ۄ�I��?��p��exDH|&��Ũ�ͪ�a�a�J^������&S�OQ=|x�E�����v��Iw��[,b(h��|�H<��ʺ��g���}��Wd n���)3X	Gƅݡ_�yդ�<Mx�d����K���(e���aE��Ro��z�v���m)����r�*1�q���(=�ҏ�� *S�v��>BCۏ3�Q���Y��3�΅B��>@I��}ql@J� Xs�ɚ�jΐ����?i����r��������ad������V����,NP�7��ᖓY����4s�+Ah����Q~�;SV��^�m��r�9�U�8����=��(&��տ��/s��I�~t�~�k��+=u�&��Q�!���<=�R[4_�UH�u����D����1f.���u���mrv�'�����Cu}`pP�#u̅9:�)��2�q{6yZh04�H�ov�Ϡ���[3lE�W^h�]��7�<�$��*���l�	��8�c�(en����C����Am��ݟ�~�V����v�/��*S�z�\����9R~m��)�o�|oy񬙿����8�P��=m��ޙ�)�<�a<kn�=�tb��-�x�!y�l�f�U�Y����ⴸ2�
sÁ�6`������>��{<y��ɉ!gx���S`_<���y�ċګ3@��7��2�ZN���y�c�]�(���k�j�ڒ�sqV��#cc:k�q���Qyx��p���ND9Ó2���4��zNǰ4�y,���)���wt������3�Pپ�7�m��>�}#c��x�LO�Vɏ��2L'����e���C���p�VVMw�1��DXO�ڂ�`n`Cї��cu0�4���{��\����7`�Z�~���w���0)���h�����+\�N��ۅW@�v��	�O�0(��&��+�n��%Z�뽽�HR��EQ�\�.V��e�>XFjQg�a}�o �� �߹X<+���;I��:���TjU��;��GC"�R<H˲�v��d=����'g� ��OC��K H6�>/��fR��}�F���&`m��@rv^�vSZ�3XL[RF�0�zM#(�4� +;`�a@�f��MRWw�;C]�cǌo�owq�/���s7&�*��]_k=}ܳFA�NV�(�R�5���0)j�S�Ձ���Wi0չ��f&�fl�:SC#V�0�Czx]��Κ�Q��%ǯ�����	�iV=�����'�"�W�T�`��5�f�Kp��8壥���P�c���p�K�-�V��^��}ޯ�橝m6�8g��� ;�I���	�%��Z�S6�/�}3��eCo�A|�D/s�B��,�:���cz�ቐeTU��SF��<O�iM>��/�]��mk��a��D���V�YY:^��;�`�盔#C�Uۅ8��ӷ;��i���?��l�j%ky0�JB��]��xB����g`��pR��~�+/���ˎT���;y>����1F�8���S�r�	.��qlR?�+�3���86�myh�'��fT��%\�ϻ6��`�$��7�L[�8��ד���'��6�_�5";8�V/��߫�Ig�^j_��ŵ�Au#��L�htZģ���Se�<�棝��ͻ�a�Ҕ��!�;׹���ރ��)|�p>k5��^s��N�!�Ȉ�0�� o�?h�������`��em�?}������Iuy��F��c.��Vޏm�q�J�[m�yۭP�:8:vp<��ܻ����Q�ԭ���NNE3؛mr�[��]�μQ�i����(OÏ� 5�Qp.��;�N�8|�7��paq�!.ʊ'���qp	�_���!(f�X�� ��>
]��Li�훜�j�.�BV���CX��/�����Dളj�x�k�}�[�B�����mF�㚎⡣���p�@}�ꍇ��Z�΢t[%{�V�`7R�Y'^�AuK{�T��F�㦖<:yy��^����V� |vK{j�H�9Y�<�a�g�J�3�O�1@ՓA�3�$��W�Ch@�_�u.��X�w��/��ͻ�na�F�.��;��3�L矼nĩ�ƨ塁��>�����o�J��s!N�){����$b�>��_o��<++Bv'��;_�FyƘ�qp�����ӗx��'�"��C<��ư`I��Az��짓v���ެy�l�\J�87#��+ɪ��p�����,%;+���}.O �Ѓ���H��'U\�����a����s���
�B�d�,Ǩ����LumJqy[L�;g>�	��5���>z�V�8w�Q0��6�8/�_��dpF��VB}�I{:��yզ�&�;O�j�b�JK(eRq3�ohT]��@!j�[E� -  ��
�J/e0��G:x���&��+��W�k��^\���*�m��Ac�(nH�Ǔ)x�"���=ǣ]�#��-�8<:��ðx�9�N��*IJ�י3ap���x]�n{8��0B"ާXxg��PJ�+c���^#��m�A�IY)Ș�&Gۡ�<�;B����g܆y�|����Z���s��<��`��L���rx������g�kM�]pO��@�3W��sy2њ��?<F�2��=XxZ�Q��/�<
�U������.��qË�3�e����7�Q8D-F�jgG)� ��=s����@����f�1�=|��aw���A���?7�z���W�O��Eeڪ`:Ax1D�iX�����V���O���
�s�ٓy��xgN�n�G���o�;�������������W���2�앵V'��ɢ�f�08�����g�Qt�8�6��Ȁ{w������)\4��ƣc�iw����_|m+�Ių`�_���<����9x�Ź��+����ߙ�����=��Y�V�V���,�c8ۇ̖(��r2�l���ŻV��ꐑQ:2��x�j\oE/�������Z��?G�#	�٪��K\�=�Ye��*�f�N��H"�|&���R���q�Ù��X8�R��ӡOX2��I;T��a�|`��8 ��f��I#|� �cr"���:�y��,���Y���}��P�m N��~Sx�;鸫3��L�Nָ���%��xa�@M�˃,�(SH����`%���v����`��vʨ|_�~R[�w��	7���&�M�Ya�n��A0(s<V�;�lFC�3ln��
��Y��.�B�~��f���&Έ%'�)�f��a�٩,+uD�U`�.#�9�M{�����yn΍�f�v���Ӕ�絧����"V�Ll[^��(�n���jcZDص�`��Ǣli�޻���8%���w8`���w!e~C������B`�C�8``�{ �H�=yL8RRӗ�	���1�i	��R��|��x��%4De�W�}�#��ؓ���-F�,��8yn�O!�Nr�ХX����L1՛����^\W���3��t�F~U�: �� ?��;Ct��s�!9{a:F%�dX<��x�(xcܓ�k��HN��>��3��w��	��C�,��DuIÁ�s���0�#! ��7�ݳ�.�<a�$� ��s&̇����4\p�}Y�3�z�V�w��7���f��X�rÝ<�y���*�����#J��.vfc=1�5�y�7���z8�v�e=�۝�w��z�t���&
�#С��g��c֑A��@UC�^���1p����aޓ���)aXo����m=����Ė�p����`�3�O;��U��r�V	�������d ��{����	#�$�����CG�u�]r�թ(� �;��B�k��ŕJǚ���$�}�C�`s�2H���d^��1��}��5Ͱ����e��&��~��Qg��6�sŇ��F]�V˙Ћ攂�wO���/��]q:���>�iX9�Vg����ރth�"9�x���:����7�����a^�R��^�=�͠��?}w����_F��?wΡ�������_�҅�x��<��0������ǳu�~�B�$x�m�Ì�����EVw�"�90���<�����:�~vk����9Fx@�KC����ɃmA���<����{yETo�����9T}�y�
�k���v���y��im�J��3�x��Z(�`��6*�|t�eE�塋������iC�d����Vg�8~2l��dc�ka)^l�0JF�Ƨ�b\�7/'��Q[�K
�%�hC��Z��.F��1�x�\Gz=���&9�/� ��ѵ��P򰕮07� :]<����l5bQyKV�������RƓ���F��4�ɳ��5�/������4_��@��n��'O��h�mΛ�u<U��� O+�*t�t�y��n���_�(�z�������W���r#,�~�S����`[�n%���пg�9���]��a���?)��.s&Ե��V��Βkt�+*'�����r������)q��Y~�Q�4���1I����۵Q���5��`�o�5-vJ�w�����X�5����zm��ł�A\ ���K��،G��=��Զ��\{Q��
��wU����V�sE¹>FZ@)�G�1�*���;���=��e5�R�w�\1Yu���~G�Z��W�s�N�1tb���ڜaV�����]��,?ƐF��m�A��GhHl/�b��O�LO-��;��2`��w���v&�p�ZOo��3�7B����I_U����]�N��1�9,G����R}�m��ͫgE訝�:z�6D}gC�!����R�J5u�A���N�u\/�ms���m{��M�KP�����j� #��:e��e�k��ɣ���������,��$)�c��	isg�C��M8@�(Z�IA0�܆�����ǟ�{����LǠT�����KCg�?y���ğ�!�hz�/�����,Bo���M)QTv��c��t��u�����u5ԗ�<������/�GJ��
�|6��2�x��)�'S��g�x��v������?�ג�}��qm�x����/\̓��+f�o�[a�mt��dL����?����N9h���� �c�"E�'���w���<D"��i�Ӌ�?��Ct~ю�&�������x��M%�E����I8sn�������.ϑ^s�5|�����3��}k�z*������a�xJ�᭤T���N_�#
~&�G�z9���?'K�-ԾO��\����+�N�v�*O��"�$3(>^V��z�a�������[y�aJ� �RȁW�V�2�O�Itʬj�Q��3�_�s����_������Ǩ$�̳�W�b	^/�ypֲ%#�0��E��9���0�d��J�x<��a�[�qt�-f�3x>�xߡ�ڙ�w�vN�}�:sת����/�jg�.C�-�B��-
1�x���霨�|��x�I������yen޼ֳ��Q
^�� ɫ�%��������*#h�0���$Z���?n�<ğ�����Q����_�x7:�rc�������:/�//��`�I��9��xb��Z#_�i�y�2jZP�AgA�N,��~��[��M���@��v�c?�s�߻tx=#������NظV���P������'��׺׋��=�J�<�H�5}}^flөo�[Dўn��՗�������Z,|�y�HJ��%z/����Z��y�W��w� b�kq����K^t
��_:�u���
)��>���=��c�zD�i����ŝь���z����^���!��%�퇧OkLh}�����w/��  R�ǋ�KE^�e�$D������{x�cƛ��x.F������ԛk�0�����GQV�=b0F��(�<���s�}d�d��w�C�T}�M��!8%� \0��+0��b��a�a��L�|RO��a���9F#���j�����S��)��5��v̇10/����we,aY���ʾ�6i��)��>���s�9�6���xk���&����#����ߴ��8o�5���J��7N�Shp� ��4���v#��F�ӋN�jDϞ��3Z(^C[3UA���)�S��3G��*��ye�3�`�a�p��0{�)=�,��s���7������o�����Iyx#v|�PVC6��f���xk�,5`��^��{TK�	�5��ջ{�0֓<`�_!�#�鄗���<L�_�ȓ�~�Q�9Lw���ؼ�c��d]3K��2��^�g^�1tM�f�y��z��V�o�B�:̀"�\�)�^�Q0�������ȶՔ���+Ζ���g�k� ?s�lҍg:E8|�9F`=m��Q�o7T�iإ��4�㵟W��yxG4�H�X��z:�g~C��a�(�_b�p����i�-��l\[>�@*b��`�駟�"�x-ym�Qi��4��P�36[f��GU���s�]^�}��e����M�� i[���	'|@�֡k���ю���3���8|L�a�����HgԽK6��0�t�&��ˊR6J/���\^�♠���qbB���I�a������1�l;Q4��;�W�$��u|`K
s�n�">/�<}pK�V��jD��=�� µ�	v��R!����*<3���74��DNk����/�v+O�'y��������u��)"���� {ӆ�OoGg�a�t�δ�S��+͋��3q��E睂6ʕ�b�3B����(���1&�7��ܥ��<<�IΜK6�<�
���>ׯ~����?�ָ>Ɨp��{���asܞ�Ԗn��=n>��臟��~-�į���1f�3�n�7}3^<�)�npYA3hg�C)����;���O�n:D�%��mp:����������et�x�=�E�NL�"�6��΃���p�N��<m�=`��������4�����|�h��ݐ��gkV�3|�頶�`��)[�X��v�ǫ2�"�'�W�MZ�<hӗ*�Kf��Vfk8�a��7�Z�[2���`̪�`�UyΆ����,���k�Ȅ��gR�a����$������gc�ػ3 �GI���?j�B͐�����	�i�ƒs8��~%@!��џ�8�ז1�)�OH� �$iQ{n�|z�zZ�{���?��_jx�ECG�0���8W�g�|5� ���"�3�J�	�k	�o���b?�'1��ë��_e�������HYt�Nޖ�������z�Je��N�?�ɻ*F�,᠁}1�r����<��6�4��W�����z6W���@�0���a����p����a�*���9&RG0j8�~"t���@�D��\z�@�u���/+�ۯ뙵�9/܋����d�a=�HHR��z㇆;��K�e������`�����!x��3���O�#T�?yb�6���=��O<�}�x����Çk�	AM��[�:���#���s����gZ%@�F��� K��PD��\�e���R���2�j�g�.e$i��/ف�%��[Ou;j�B����E�g�[Z*��<l���>������o���!ބg)|#g���z��Z�-|�h=���P����Q^Ǫ6��3�Qkj ��>L�p�̄�_�k��Go���O4���A�R��Hs`x�i<�1�ͪOi�s�_�M��xg����j��c�_�d �#�e<�z�R��;���핇�$%�.�U�jS�J�}�b6�.��t��nB��z�t(�Rqz��+ZP����	��57��� ���e'`�/�kx���,�����$���6��<�U�C��R��9|�K]�P^�S�o2��?�#W����e��	��6������w����w����婋ǂ����#�upՅG�z1,�B`�Wu��[F]َ�.�au8���P��r�H�����_|�U�-��lE�-(Wϙ����������O3��������y�~�|��o��;唈F
"��4#8�a��8�(]��<+o��`��O�1X�̄�4�>�}r��EF�W_\?|����j�-Hk7d��-<]�\yw�y-ou�Q��!�ۇy�yJG���OM����yӚ�۰kgK'��`���ߢӒ{=�����-��4����YtC����'����پ�3�.pW��鉅��,-F�i�`F~�y�;ɣ�oSL=�H����o����_^�U;\����*.�pm�ޜM;����+�?i5��ں�3�\���)�Q�F���R�u�_Se�:��=\�Dj�:�%�TF���M�㞎��}��aJ�,/Xu ��w�y��.WV��Y=^�ȅ�<���T��U�l6��k�<����k0�XɐŚ�� cx���Q��8CΜ��[�St�I_˗�V4�6/���k	P��I�$O�+�Ă���^D���b���Z����:����$��|�����/w��95=VOL��UK�QP{��?Dd.�M���r�Z��Pn��~�Ⓦ���)T.PFf�4�f�J�
�Ư�~T��F��G���Ë����=C0E<e��6VyвyT̞57�?�㷇���ׇ���j0���>��Û���Gw1��ά>��w⠿���	��ux�16��N���9\�~�Q�����_��W��S�����0�W��\��h����VG�4�khm������?����1�MC�S��Rb���u��9���Q_^�W���޿ύ�p��z�:��z^�a�h<9����ϊ�ݍ	���,!i�Xi��P�*?)v�r�9��9Ƥ��hB�<m��(/&}ʃG��T�G���2g��6Q���f�Pj�[�~�Nջ'��
Oʐ�(�Ÿd�D��Fy�0���m:��f#�#ȫ8�/�jAJtJ��ˣ��ڠ�w��� ̓!p��F����1x7z�2��F[��kU�s�޻0[6��H5Ln�%��x��N�a�s���S[�5��wʂb��y1�B�ԪE�{��ߓ!x��c8�0V�R�%,�.�L	�W��S���e~*�#��>����Jo�r��LoJ	q��(�RT�%��\~�,��T���(�1��i?��򰽌A����c|�dl�#8�\%ڗ�|T��:L�ꘌ�W�p�R{<������e0��F;C�z�e�j���*���+ۿ��T�D�ܓ��|�e�FCV�}V�� p*���M��>��{���[�g�@�z���-l0�M�+Y[&����Ƶ+#/$ �����'��8F��;\Ew��L^���C��n�Nk���ͻ����_�ld�R�Tx����n���|Ĺ�&��|zsr#y�eżm.Փ���z�O��k�!#I�s���V��?�_Gf�4���e��s�>�Ҫ���U�� e�;r���l�^��Y��� 7چ�)�~`ڳ����6��ps���U��}���͛Cɫ�^�QAFgho�����\Y�r̃�|�����%�\�7��:��_����u����I{�E����.����u�mv�F�ߓ�L�I&����J-��t?��o���Ҟ���uK*��Y�������J���<�lX�@ ��t�|��$�n��6���
;@l0o�Ie�Ϛ����@��>�4d��h���'���Qjs(���\I�TxT�lX6� ����Y�@#�P�5�ISCV�M1\;���Qؠ�=��_��*2�Ϟs9"���u҇i�<�R&�	�!�]jGSQFɦ���g�=�Uny]ܸ��εl`�&����"�`¸CZ�sW�:��2�d�8S���0#Ap��5�/.4�����\��Ձ�R��r۰��TZ�Y�Z����c|��ѣ��v�Vӣ6�n5�	xX���v%eG��1^�Q��.�x����;���?�|�%��p�fʩ|�%�x�`��+gw��������[���]����FC#F���b �d�)zw"fsв�g�nyi���mi]�9��B6L�"�A���/��3��N��>����ci����5�l�rӥ_6Z�|>�L�����cVUv�����=Pe�e<�w9�?6z|�_�%!0��YL�Si�:k/�·�XK�&+����LL�������t>�c9�5C�9ʿI�0��_Z[�(�ot���Yc<�$0�.�l�b�� ��Y�����}S��(ax�<hZ�[�QĀҁ�62"xVK������F�7i�;8ux��Q�q���+MߧAOG'�t���� @￻ �U���L�"�Fc�3���։��"|���i;/�k�:�m��O�ڹ~�f����Ӧ��~i*K=�e�C	s1�Ki����gS�e���xGm���q��jP�����6�f������$�U8� ��  �U���yVoè�>��.� ��w�V1r�Sao�f:b/W�`��[ً�	���ê�M�BF��M���{��@��5(�=�<t�s��L����MD�q�_!JO���@(��<Je�:?�����-�x�,��'��r��O�J�ӌﯳ�w�n^�o��g.�|���x�M�5P���l��;Sc��*=�7e@�4�l0u����|3�[-���s���*�A�1�>�a �ĳ�N)N�T:}��`%�y/���]���%i;�����/���Jq+ �JʣN�	���� ��ɞF�����Bm����w�~��A��ʧ��X?F�l5�c[Y��1O>3@�<@VY�-�SV��]g�j�
�Cs�:���G�6�N���f�Xm���l�	�>uh-��]������������G�n�����)W)�l��ƴ�c�gpՠ�eZ�'�Z����ԅ�F;W��*S3!	_������i̎7�}�=�~��1�\}I�Q�pT]�Qc#��%��%�/���V�i�%g#�'�=����f�L��cND�3���=Z��d�&�U@�R�e��fj�" ��X��:	LoT��S���3�Z���ڡ���/	ۈ�}ڙW1X�G*�eSf	u@o�yɍ��5ݢ�� Q�9g%fB�G�n\�TЄA\����ʄ��?���,m^�aJ)GX%��U	:G��4���Lix�bGi���{��	`g��\��>IW���5:�h*���N���jvO�=x|a�.�fz��:����~Ъ��*�C1�\�9�뇯�w��O��.�B�����f6�3���� ��6U��lNF����ب�紀�y OH�-�S#ރ�_Jp;S���^�����.���9ˤ9���hOK�1�o�����[8�����݄�i<LK�%3��8ш�_%c�۵�Z.�����k:�p
y��ם+���6��$�j~���8���i�OUZ��n�$;'�_m|�Z�}tI1,4T?��L%�<ED�C/���:��pn�	�]0#Qt#<��{������h�ה���-|�xԀ
8�O�^�v5�'ώ�.P�r��\7l�I~~T�a["�o�O�<����6�R�^F{��LNeSpB�wiL��ݜ9]}�)mЦ�0��� {����|�l]�������4"?����w�bLm�龎��)~�,Q��GG�Ҷ��D�Z�A��{�u*�l?u
;�)����/h:�;��$z��[xٹx�8�(�fR�7ә{��G挗@1�#	=����c��Y��+l'�q��	�KAP�-
,�2 �ϵw#l�Zy�4�gj��jN|�t�7[�p=l��ꘁR0�Th�Á�]i�i�W60�35�&PZb�=� �|��";�Ӆ]-B:���j��1��.����r+�^�2���o��W�"^�&dt1���d&��S<ji���\�At�V��O�.W5�a)�T�UG�۱oĻ�u�g�����ի�,D�ٷ~l1�����fh��~قi;+]��ЩË	&m���"3�L9v	`�RR�Ş!|iQ,:,^X�1OӢNW�5����
e�r���|�J]6��';].G��T+./�k��l{g�:���Bu'!Ơ�v�y�'������3Hk�^݈���/2�xwpIѢ1]�_�w�`��Y�R?+<.��]WU��E>%��n�78e�JK�р��XL�K��۶IZ\p�;esuh	z��b'#�9��sL��>*�'Z�^���ؐ-0�ʧ���X3Vy �w	�?h���\LV����5��U0��,U�l�Z�z�w�1�o���b���fC� �&T��p�{/��H-PY�"�W��G�K�FUAl�rP���rZ�xdC��0���9Æ��
����aK� ���Ǽ~��?�y�F>y>d#����#���>5gӏ#��^e������Lg*"٭J���Ng{��`��*���Yu_���;����~v�^�����O�����LO��rr�p�F~����~����1~�h�B��d���)%�Y���b���t���N�������*�o�=t}��������W�h�@Y��}u%���2Ҽ83̓|h�V��N�GP�%�/�;�Z��￞��\��/�P�q���ۊ�F�m.�ߴBm�;h�B(��!��*�ɉ�~"Z����u�B�<�z������':���	5�Mm��`^�*���M'񹁅09�m���q��	�)h��e5L�t��0cC�L�rP���X
 3���|�f���S�W�� ��>��d�W*+DW0-PzWľ���>�;��׫��n���wGLa�MX0�?ϦT��T�Ѽ�;t�:{J�����ի�ow�O3�t�3�V��t��4���xXgV��h�-)����^��6��*��~�a��������a.�@e�E�Ԫ[~�*�h̷Lws,�����Nb����֦M�:e	��Xo���х��]ո�\���*��sC����V�@-4��z��7���
����J7�y`m�t�Z:a���<�Щl~^���tt%d��}���������l���7��G�����#�>��\�l������>h/�����`7`dJ{!�V�_�Iy�>��5�i3x]W�6n����n�Wz:^�e�bP"<~�p�I� �&gw7�"ŋ�0�~����D.��)%Nv	_��ն.�#�cw�b�7	M|�X��	S��w]	u���E�x�_��ٻ��X�t&A�D���7R�iY�x]Gc���Hd�F����u�q�[6�K(5�c�v����q�CL�3�TX�_6K�m�
��ݟgPs����cZrn�����XX�{����j�f�w��+�Y���f3C��ޖ~�N����M��?�<�����w;_\:?$ԧ���b��=v��<zz�p�3��iNN@]# �C�W���:��D�:�/�0�5�����1��v�+��-G��u>������c����e�R�%WD����!�W�3�3{נּbWa9��9!Bb���)GZ�#�-l��&�O��lx�a��(�sU�VC�)�4Tu|9���7B��i�A'�*`g�DH�T5��~�%Y2�`	  @ IDATG�3�b>��:z$#���������is��P�ٔX��3��p�ڹ�HFɻ��1���
A���yԺ�_)V+g���Tu	U��aà���jg5�O�Ί0a�}�N����_2�nD�o�<��}��ȉ��;�5���4W�̖ĸaWҵ�n1���k��)|�N�1�n�1��:�{5>ӷ����U�L�^h_/�J|�����#,lG�5xZ�2�� WL�<�_���&���NN+��Q�������J���w~�ۉa"{i��PcD'c�����$И�~���E=��W��:��hnl�*Bd4�����v�*��A��h�b���sq,����ro�SYU�T�Jw��� �i�e���|��ʠÜ)jyX���uӁ�ny�+7h#���b��B��	��ٽP���:/V��[��1��܋�	&� ��	�	�\:�AøR���si���������<¸-Q�g��;�{��7!��ө'��H�ګݍ�އ�=���~���~?+�,vy� q��ɫ����;Nn�0`K�O@�?7�z���G�h�����J�g��-WaSH�?!����Vp��?��\��3�����[_��ߕv��>��^���jx�<�i��_[��Gޛ�	��4����*��K���7S`�1���{2�!e��-��K8����	�B~@P��`#�	��+̮��Z�u��A2���րu\ϟ?m��q�r"��vT`z� v:���ף��gi1���bh���v���2�:�����T�|���s|%�:���o�� ��Ȇg����_~��Yn:�a�l�L����)Be����˟����L�i���w;GС��&F��U��럋o`��ַm��w���M�?�������.����A�\Op���yB,�/����ϩ��������v����,>��ۭ���������Y<x��Mmw�A�&�?�������e��1M؇�A�Ư�kE���}��,p����ޟ)F}[���������X�&�xQ� �� 4|!�p>���>��ۣ���ܼ�2�����-�hD_�͆SZ��G�ٞ>��L��w�͓�X޶���˧C�|�h4V��}*�T��x�ƏGG�9[l��@�P��<��
�l��պ�,|�r_�N�Fǚ�;�q�nԊ8Fh(���C+�F3��h)�f��њ��u�wǈ�[~#�:��Oٹv�N�*۔�g�d��u6UN�Ҧ��!c#8�*��T3�[��/ә�ޔ���%}�a�₥x���j���6B�Ճ�[Eh)6����ۯ��t�<n+�೭	�8�h�x�\m��K�	{5���͠�H��a=j�F�l�F�id�0=��HC65J�f��MS����Ay����
��u��Νi
3�Ry�T���:��M�p�@�����Vc^�tq�g�m_���p*[-+n8U�<�����7fԂaq�������������{
�Ջ\=��}������q{NZ5�u��[Z�nk���Q���׼���1�:�A3�d�o�/�E�C�ѫ���D��{��-Oc߄��>��y�����\q�D\��E�2XYIw������{)H�3 `8MD���	��*��)��>c���wbn�'���o3P담�M�c'�m�R�⋳;?������|�ݗ���6^_�u��^'���k�fE/�Ȭ�*�N���m��ۯ�����;?|�M�������=�����wj?�+F{'�	LhD8"�����:����ˏ�w����#nV��IPVp�)���4|�9`g�+,U��S�M��U�v�����$��n	VEݼ[�����S�кI[^:<�� SCa4@H`�Kc0�.滄
����k=�}#�07�O��N.<���j7KPR��,����h�}�����GP�q�Έ������<�Y���S��5����0�Ե�7�y�H���!]Ǖ�_윻ry�d�z��T{i@�&��H3Ek�o8�,ñ4���6z�����^��{/����'6�G_f?�ӷ�?3Q�;�B`�޻�.�5�x�yƹ�g����H���X��g?�<#���F�\�|�/.e��ޕfpRv��M�r�4�8�|�5�	�S����R}� �qvR?�5�	�K��`?\����W�뷕˂�<���2�p��}D�V��N��M9�1|�ݼy#eƵ�6{(�W�ph�L>$7�,0�>>:���KΠ_�:���ә'\>��3W9ljC0}D3�b��ﶨ��	�~��>Á��˓�v�ku0S�=���&p�7G��=
�x�+�O-ebsfZ5�n�x<�3��E���޻��_|�ua�9��z�r��4a�9`l^�}�|s7bŸ�o5>��ƀ�� q��� @@g�ݖk"6�W�	V��@��D5�D!U��)��x��g��\ID���nL9Ґ,�%�H��xi�H�4_w�n�K�|��c���F�Uc��f/5_D��o�a����r."Zࣈ-Ù� dʶa��W=sbD:$���P*tZ��7o�6�c�p��+���e��q��v��sIʗ/���ND��a�hSq��:�H�
eF%�ƙ*�;�ߺy���="�q�p���
Ĵ���D��lڇo��h^5�b���\v^�Z1dz�8A�a��uz�����⨾��4b����F��#8Q#z���`4�{o��wpN6�x0LI��ߣ�Wƈ���?j{�)߽wo租~ڱX�h�u�����Mǰ�a�����$I�B�bsj�/�-C4;g�����f��
�1�sD�Ι�3\�m;H�#-j�V��8[���zY[�H�x�Y������P�z?0N�%��@������J�WY�rbn����b��i���W����6������������Mi����ڵ4֫uc�1��i������e?F��vr9zb:ap`
�=�v��o5�B'_�Mi��(�D��g�[�>zӿߔ��p:�i�1A����r9֯��/}����� {1w���!�I������6���ͷ��w�]��cr�~� =��9&��7��h�>��k^�}�8M�]u��� �����\k��o�����h������hz�S��d~q,��?��^���K�� ���6�:?q��7 &�}'�GsSƣ��w�El���)���=S|�N 4Y�_�!Դ##�f�X�R�/Gۈ��tpe����1�.c��`@^��*�6<������ʬ����X�i�P9=΁����}O�Z�e�[]l5�
V�祍O���ζ:����p�]�4wf3N�:��<H����O���
W?�[��m5S�G�����tcD'DOp}�ԧ&8��r����vfsi��D-�� �V�a���i_�"^T�qU\��.���t3/�
�f�i"��>�Az��[آw��V�v* ���,�r?����������LsZ?��Mmk�2:T���M޻�>��y}�iaS�x화,�,C�{����C��ۣ=1� xǏ]�5�KJ�����g$V�26�z  ��:�Ü4��W{��a�X�Y\T�Ujs��(�0Ԑa>�_CCl�}��,�8�iy�\K�?��H_�؛�V׵�n����?5�� ��;�ײl���6j�|x�Mʻ��N}w�I�K�^D$��k��]�ʯw�{R�!��fJiI��+\�V�����������{�_��9FigZaȎf�	ד�bT��b2�*ۗ�$��h����n��Ȩ���Pr����������`3�!���o��������11�'}Yg�6�Z�O��U���qNL��޲������?��~0�E�&������:���v4:Pj���/�?6[4r��6L��WÌ��,^4M��b���V%8ژ� ?+�̈́ys~�j��q�ss�jkug��&e6+n�y�Jݏq���jF��(��^�"��C��C��u��D�FR�u�Cǋ>���d	�q�c/Zل���Es��O1Ͻ�D�" Aw�KhLٴ�(�fǫi0ݬ�R��_�.�V;[�+<�]�ϝ.[ 6�_o����]O�{��M{K��k w:���V�����a-��kV$���3� G<����Y���G>�g`6�gҞ�6;�
���v|�f��s�r�`�HY硬`7��0�9���㳰'�� ��/�u�8l��\�QG�sDU��ZB�op D��o�I��N�m����mh��7a�_��Vz��}�	����{%���6����浟���Ү�%yhO�s����j�S����o#�L[��W	�)w4"m�Msϐ�������)�^��^��N5m���E�}tZ�<����xYխ���h��0��D�N��M��ղU�5e�>A�b���b4]�-|��R|^����|cw�Y�fE�*f��ޱ�M�3:�q뗴Ji���o����n�h�Qz��>6cc��|+O�)�x�b�3�-ڷ˳�=��3���ۥ�]C����l�.��c�����x��W��6'��}���i��A��<�N9IM���\�>�qgS�k���cS>��}�Ϩ� f@���� ���w��'�|����ϔ7�N��|U��A��^�׃[�_2�g��ܾ����v�=�j|�u�as>{&m�a���b"��"�b �}���[5�L���<��RE�
d3�@�P��}��t����d��VA������Uϴ%4��.Y���g�I�[0�`!�N��=~x7�ފ7ը3Y��û�Uf��:G�Z Z��1�*V\�g��o�2a�A.s��w���<�esn���O�� 6�!��tB�%}��7�?j�"��~�Tm��<g��k7Z�~g�Y��h+MG��QK"��Ikr�%�G��a�T�h2bF��"z0-�B,_�����8�����2��<H-�$���D�T�ĕߐ���E���T��ۘ���t���~�JǯZ9�������5����ꏝ��lec4��8d@]6��SuH'��ўe�`NB��ly]�|�w�	�	`��ch�N�p-{������~���i��r{���|gf
�1o��j4x�¥�gM�4���6{�J�$������:X�0
��h�T	��Y��xϰ:K�#$��V�F��J��C �b����0�����(�>a�2Ѭ:��5��Φ��m����3z�����7-��`�AID1�6�M�/yT6���z��D��p��n&�Ҝ{��w.�Ϧ�{��o����I����~��WN^e��� ���ò���$0Y��e~�8}�r��c�Qg�KGѴ�.��7����;=��Suj�הR6/����Ɨݟis�`���5�h����g���M��0�NA�a+�zvx(��#���F��Y(������܈�M�`�n^���n�������M���d�Uz�/S/�u}r���o�r�l ���*��ʰ�:�.���h����|���mt:�;�⩇"�L�|�qS��Yx���'�����f)����믾M;uzh�R��*���9����>�hV?�e�±��p����L�Yl` ��~��,����V�%X�|+^�/	�[�p�?#���E|��~+��O,����&�q�"w�V;�fϟ��X�Q"���Iv@	���L�^ܿo��>ŀU�M��ϣ��@���j��/K���?l��æ��rf����Ë�A�)���p���Ƨ�Dm*�ju��ؚ�pLW��ev�������1�ov��ӌ����q�a��u�O�z��]��}^Z�l���>�_�6j���6}&����l������� -�[���9FcE �����@�g�7w�����:e4�EP���������e���B;.�x�·sBڅ��R5�r��ٌ:鍣Ó�	[+!��g�VÞ��W^xb� ��Av)_d���扡in�,��)�t=�9ioa��Y0H7*a��n��al\��mI��;�G�7JyB��6h���rN⬗�:OF�{������� P����(b1T����ʅ@�RL�~�4Tv���*�Q�E�je�7ߵ�D�J��}��w�\/ʹi�0�4cȟn~�v�rܙ�4B�����;����Lit��k�׮g�����G�?�+뱏i�R'�ީm켬\w]������$r�ժ��GX�5
<�=×	jV�]�>���1�$i�~��O3����D!vY6
\�[2��)�{��6~7;3K��;
�ə���]�ʉ�O1�h��C.D^���F�{���l�!F���ojT���y�R�#{'�^xR�ǞH�_7�BK����:3�҃����u7����:�����dEh�w�\��O��йЄΨ%��������y�w��z���i���\���v)�~j�`s�z-oG�Ն6�����;�K�e��G��)M����[�+�M�A9y��t��u�c�����9���/��(��w;.�i���c�O�|��k�\݆��D�I��
�A���4� N '�+��г��k gtm۱�1y�0���L�_��N�U+~�$֧�to�<����8@f}٠k�zئ=�C_�O���Jc���^�n�l��GHp�����-\�g�tJ>�s�6Sg���+�?�Ia��2�ZXW��/~��V¨r�g�����iJ]��j(ӹ�,ad�IҌ���;��Qt�V����r���� `z@k�$�s��@|�4"�Q�>����[7wn^���K��Ƀ_���}i�u�^G`� �)'���v�5	�)/��h����_���gM����߼9Ҡ��h�][�d�{�d�6S�f��=A���
.���.������f�{?w�Z%��@���F�y|���vR����U��N�,
���Z�%d��	��i����L��zV�Ő&��?'̔�����fgw�N�C��.DՆkߥ/��~�xh]�􁤰�@n�42:�7C��	�w�k�J����K�?1����7��[��*_t4t8�
0�B��
�貹�C��ϭԫ2Ȋ��f��&�n�xo�w ���@>G���RC�tE�˗�Gچ5�~����T�E��x$H*!�6'�t��#.�����n���m۩�0j!)��vx�b����aR��z,���(A3�4bp>Ik�K�Y�޻�6�a�r[!$��an����F���Hm7���~�I
m�!�A(�*��؎�*XujN���v1 �N����5���w.\j�˹6WM;t���1�T^�?h�����{M�Y1�nfKc:��y8G(:"�'���{�&��Უy��y����Tx#�������T�@�d�����+o���8�p!��O]���8�e���Ʉ�4f�u�c �l�iM#���ރ���)mis���x)�NO�(zo��Jт%Z�Ͷb7!n7��U����~W�Sڎ���*7}<-۫�0n�!J��#$�H�ȆA-�nm(�s^֍j+�M��&�F?�}�T����chc�y�p{��
�ʀ��A��&������M���a���w�I�pe�t�v�yґ��K�`o���<�pé��ę�&s���0�Kwr[�8C�ݬ�{�����H�nJ��׉㵍kX$��0:�&���|��!:�̴�ae��r��7i�մg �N��#|-:l!G6Bgj:)u@ ���RXf�Z�;�0f	M�3eP��.lJ��G�/%V詿.p��_q����O�p���D�jK��}���&�IK�+�I��gy8�����۳��\��=�֠���`il��w����k= q�����]���j�@��f�	|)�c�o�J���K�]�?-�𮎼z��ES7pO;�]�~��l�:����pA�/�U4!�ai�6�~�Mխ��;���цt�(3�`�s�, smtS������a�so����>�Z,�H�w<Og�s���N� ?�?�,B3����iȇ��n�	KxPO&`�:�*g׹d8�O�F���-t���ǲ�f|O���~�g�����i_�XG��A�oe0�޻m��av�(�h�R���}�f$�lgɄ���hE?I6�<gO�ʳ�㪻�4}���"��w�߁�	����8�����҂��.mhϣ�g�cA l��వ��c���_�Z���j�w�'�A����?�8����,��yl�l��r���	�4��	}�Au1n���	` ��>*�΀�HF��?}R'V%%��Ϧ�*?91�"��`d�iu෍��*5h#�m�o(D}��k�g}"S�`Sy�Y�S<?���j#_[���������i_��j>�m{�}P�	����W\ڏ3g/��tٔd��W�<}��"L�!6���0�ʭ���o�~# {��R��|h������e�w<50��=ΌD����ō�˃G{�= FC�t����$?3��Q/c�TV*#��Uje�	V� �2޽�g!A�������0�b��!��MlOB˅4��[@P�o�K��-ݒ�Y`#���ҶkQ���l�O��FNP��`�:�J�Xb1X�^nG�����E���)4u�i���-:��m������Jsy�\6g�n��S��]���������� ���}��{��'�c�8vu�ix�����iQ�s��C�`�d6�E�0>Π��-HWG(�>�/��Tw�y��1�i���"!U�W�z*�X j��(���6��.6rў��l��g�S��&g�@���<W�I*"�!������������4�	����
`�~�����7�S�قa\��.M{�-!�L�9D��o�����3��t��LrQ�-͙V�i:s8^x�ױ��42U��N���'#)�n��p:��)�7=��Ʉ��+rG�Gא48���)�<����M��uՁ�����|~�/S�^�4���/��?�<��0:�-��$z����K糍c�����2��hB%�O�@�=I���(|��j��5P��*슧��&�Frux+�+�vPf��#�����$n%����>����-b�=��9���G�v�Uo�Ԭ�.N��T���c͚��F�A�ޱl��o��~���xR[ɽx~>|}Q�ga
�Vf%��-��1L@Uek:� v�.0M�޼q{�f3�:�*�T��5%Jp�f@ؚ�Ǔ�ّ*�@�@�P<���1ڝc�������efO�_a���)}�j�&!����E�(?h��/A��&}.�SC��U�h	�pG�6-#V�TKIȫw��Y_H�8�g�����i�����k�]�W��O&rτ�iw1L�����ë�sn7�>��E��޻�Vm/�g��-��cv��^�E�7�'G�i�~�g�����~<��4�+�����9�Ka��F�-���H!AjN��*vz�
�w;��:(i�Lt�	C�:�I0�����1#�*	n��'���Kg`")��U��H�
��c?��_�u��	�H�|S��^�PB3�7�>��4buڴ'�J%H���0$|�c% ���]�A5�L��֢D8U�/��8C�Q�NGLД�"N:�i� &A3�g��ҡ0i�2�69�~Z��|�T�54+����Gb�F�X	RK竱�Q��(���d+��8�-���V�,�,�W���iN>�,�H��k�g��M�L���0�xS�`e�@p�0fd�pZ˄gLdh����#iP��>>|�t�Ǵ��L+��mg��T�Z�Vs��0?���c҅O��2[����C����m뒐Ӓ^S�GL�(5����U�V����su:��tl.s3���2՜o:��0��(�Ց��rR����\��Z��h�Ы��Žr.��P�e�'wtf���oS��W�3� ��%�?�k��4�^�[g)=��Y���9k4�?ڍ��)HD:�s˨A�X���*�L�Kug�d�)��O��1h�Ľ��H�ޢ�TZP�U{�U��s)\�Vt2u7n�8�RzG8 ;&ļ�<λ�ҁ�A�
?��yBO��(_o���<������hN��1q�̣�����9]�Q�]i�����1	o�yx]1�QX�K~���-�� ��sï�3�m��~�����&��Za���T�f�A��=m�lk���p"���=&7��p}���E���V�s�
z�$�ؔA�6��ުw��؉����h��]1�W)�a��2�Mϲ�z��Ar��n�6�WM�Zɼ��!���������{�}ӳ��/�ș����:��4�϶ߛ��˴�w�Z��&��&�#x���γ�l�6x�;�i�7���� ��K8y�]��In�����k)���W�7�+�����ߡ���uёv�	��錿���p�"�A��.�v�TB(1�+�B�I��w+^w�� �DM�W��j�x]���И|JV�J _����8>ÿ�ˋy�� ���d'�y��IդШ���6A|���n���ϻ�#��O�&X}�[BX�(zL �	m�HB�������vyo����_������*�y��WI���A;#��%/��$��5��;�8���`����?�-��XL�maU>��R�e�$��Ժ	W�����u��zg���PB�~+#Z�Ƹ<Th#�ʮ3\+:4�:�vT
re�B���f��O�PA7�R޶�?����j{	�#�����MF"���7��8���-�vh�U�� ��B��-<�����7o�mJH:�&��%Α��j i�j�'�d��+{x�dS�y�B]�3e׽�݊X;<� �C?[Z���X	0�X��*S�L��
ɧ�A>�NԘǐ�fo��2�+C�4i	OʯA/�ji�d-��ԉμSex��<�_��	�G:W���~��˝��t�����ѧ�H���Ma��b��f��o2����Ke������^}�0��� �o�	��&�
1���c��}C[��Q��1�Aw�!,�W�5q���,�^o�.���ɣ;�`��oÐ|�@���-x:����T�D�b$XK�6`1 �+4F��0_�y�υ�c���1�@+�[�����p����TL�7��ͪ=�����SAp���R(#�R��$系�e}�_�
;�S��p��h�ķx*�|0�.��w|�+�,�Ƽ���s,���^ln~}[
�+%��-��Ӟ'����>)t (�6K�n��s�0k5X�~f�c�9��[͡�Uq11���a�����8'�@HYn�����^ �X|H���)���~�?����%���Q���b?ݼ�Y�ݝ_�("[�?���H\��c�H`��9S��ie�A�ì�[]1b���݂�k��n��,Pnxʟ�^�f8�����`����΃��G���[�t���rkмg��N?�������vUV�g�xxzع��--w6wvXoʞ�ӟ��!��2�TU�m?���a�R���  v�َ�5������{�~� �"�_��O	a��{�>��v����_KQp<���4UA[)o}%�������"|�o�����a�-��Q�b���EA�{4x��^�E.x�6����T]�c��P����Nh���`�Ǽ~�����
8���J�CݎMп���;iKc��
��L�F�fm�ך�`��T}�~6w����|i�H"1ɐb���>�MSh�i�Qų4F�&��H�(&	9Ң�Qw�ro� 
������.��<��gyҷ��%�Sy �JK�����k��q*�gP$B��B��g5#fQS��vQl��6�����ӏttVe�{����d�<�X�����j%-�n��Uք��v��Kc-`XZ��y��(�Nf���ǝF�����U2?Z_����#^����3	,�tF	��ͪȃ: ���Mc��1�0�X�X�{	D8�u�u\n�Tބ�$�7��1�+?�tyo���T[��Ȅ�#C�(*<�2Dm��K~�!xWNb9Te�c�:�Q�/#cZ����+�c�q��ݘ�tZ���h��?:�0VYb�hT��!�~l��˦��Sy�j�X�)4��Fe���^сŸ6
�v4##�(��b hr����L�1��f�Y���c%T#|�;d�7@���ʡJ,IV������J�2n�����T>�m�6�aj�K���3�F���~�����N��)�z���1�5�O�4z緕{�48��f�ތ��}ۖ�6��t���=-�3�~?���*�A�*�a*�A �6���򊫣7�����$C��
���rlL�+�����kp5�T�jk!�\����:����=/A��[�w����E;��M���\]���g#�o�)��(���sIi,!��u?�ػʊo����jM[V��v���c�?��i�P����oW���n	��V�rL�����7��6.���`�ƅ�43�Z�n��iWOgq�T��a�up�jũ�lꌫ�᫽�ҐNŞ�[��_e#�􄖹�x�֌�����|;�A"\�� �7��7��R.���F�'ꔣ�<��=���I�ʧ���"�6�x�v���f>e�F?�L��[x6��7�jÃ��QWd5��d+v;M� ڴ��MH�!����d������w��<��!���Gئ�U�<)
V儴�pGr<O{Y��c�-��t���B��c^�4D%�E����_0���^Ӧ���d�h������c�-9tl���!��m�D�i���� [��w��߇1@y��)��i2.�Gx�brJM��);���Kx$��1N=-�G�LR��"�̩2p\���jۜn���,���Iz׷�0w���` �\*�`�2N�u��c[Pįt�QwﻂT����$�y��t|�� r��"�*�@ND7D|��h��Z�b�T�� ^��X�����	�Fy#|i�:�)��������V�ݏFM�%��eK^-�ՠ�;�%���P��~��V�u�KN]ms���h[��u,+����`����Ν�wG�Y��������F_~̗ @�=�M �ަuZ{+v���9L���βy�Vd��W>u�,�4ϳ��j�J���ҕ7A�Ȇ �!
1I�fvh���œ��%�Y:|�p���?���ow�]�$M�}c�ې�ہ��n��mb{x�Wf�mgBRW�@��2�����<l��O��٭N���|Vbz�D	bc����!��v��SCAh��1z�y'�����RJG��Nis���T:��(0i�I������}�\�(�@��y"����s���E�	a�G��&vDF"�pg����u�\
(%N�|~�\���t=��k���>�W�x�(�U�C>}�Uoоr"?�U;+l+q��pEXmz1)g��t�X�5�B�lu�ޅ۷����v�q�Sg{�-���hk�`��Y�>j��vh+8+�.A�o�q�Q�%�S��*���u3p��\]
�Q瀵ŋ�s�eL$�昗�M�yF'�T6s
2��n����^��^&�~&̦Kۼ[q�����wHS*�{�����}��ø�w����T�9�W�n��% ���I<l���Ē��~�vU��A�F�zݔ{ם�=+��֑����m����i�W�s��lk�\�X]]/�U~��S��3}�6m=��D/�0RE�P�0����r�*���W֧o�
#�� �}�� ���.�*��yϜ�����F_>ˠ>��[� ܾqs\�}��;w�e�hh��ԥx���x��/�N�6%9B�2�7�9�+݋�B�����]�{�T�&�}�F����´Š>l���������hO{10_x*��e2��ģŏM;ÓB����Y�D��re?����0��i�= �;��'V[���ɘ�L�W�O���)�Տm(���F>q�����X���zlh�;�]qz���I?��@P�5DM��Kё�fZ��y���W��,M��$��"��&/�q)�f	�[-Cʛ���|]�%?�Pa�HB�t\@ \�:�������2�y^`NX��>kth��
�K������&�`���ԬP*c5`�{0!��So$��{��<�F%=9k�-���_F�j�&�ɻd�`'ܬ���e7�Ԃљ��4s�J��˦1����ɹ'��--���+JN����C�|�Ҩ����|�����	k	F~�%	{�U^lc�ˍ-���K��/L�hA���b�E3E0Tƀ
���ᙽ���4�W�q�t�X��8�LS:�~JKjd�d0u�X��z�mx�E�6/���!*�0�Am��$�I�3����@��1w�!���w�Bd����p6O {����.ėo̪�ܫ��Uxp�V�I��k��I�v��*��Թ�j���d��������+��j�=���`ŷ��P��v7�Տ+��	U�G�F��:w��o"L&���
^yv�N��{�ƅ�A��`�,$��g 1�K#�y7Hܼ����v�� rNٺ_�i���휐,���P|hi�څ�1�<{W�Isn�J;W6�e �5w��a�6bT��x-��)���+xfLx�1�h��}�hw��`!����d��6���{^�PV�%lՖ����h�=U��--�݂m�3����v{l���p&�@x�����s_;��n
��
?����e���@�
������Ww�}4{��X�SQdW��yL�5��,7pz�X�+�2��W�%�O��M�V	��G�S��'��ЋF�<�����%h�ʛɃN�EuG z�U�" YLt��/m�sz�����/�ն���A�Ӧ��J�c[N�8x/:lڈP�/7:����^�ҙ�ŀ�EQ~����h*�_�	%��D��[����̆ܯ�ՠ�]����:\a�e;)0��B�Bi�n����HX��	��G�Zy�v*�S����J���h��ާ5��*[;��?~�R�n��絳 �#ͮ|���+|��v� I��^����nЈ�<��غ�y^*n@��-L��w)������!Ѧ�!����A���sS:�mN�Gh-�L�N8t�(YYA3�P)ы9�<,�V5�f�Ѫ=�+�#I� YE%A�&�Z�3�%�}h��۷��fd�r
TƟ] �lr��|��nS��l������+l�v��A\�$h�B'N���K����L��4j�����y�F3� �P:n3�L����De[��ѫ�z�Mm�[9�IgK�� Q�U~<������_5zޔ���CR����_e�~�e�g��*ɀ`��MUf��&a�Aڢ[7n&@͍Å��iر���J��_���ӡ��K�������z{�ȹ��E��
0�y4����4��&��-:#�aJ��Ӝ�n�������U��tmM=�;�߹p6��i8!��!���
�G9�u2�F���d��P���]��W��E�Hɇ]���	�ƎWc�)<Y���,m���LY*�����}B�G�v�ک��M��B2k�^̕���#���"t/na��bK�`'��eE�
ӹI��ţݐYK9�LkU��Y������-&`�����,�{���ʤ��AJ@��+h�%>�.�m���^>�����/�#�Iv5�����B����p�ǁ�ɫo&��Ul!ד7ّyQ4 ��\z�[�b��7j��i�����2�=���g�ܺZ������x�C�O���ν+700��|?Զ�C�X���1��Y�[���}tԱp:���
�d�����y���w}�؍)5�)$,���X�M�lk:S��Y�#<S�C������~|�<E��Ei|�P���C�8|���W������8�����S:R5h!�׾�N�;����g� ��^���^ƙev��[EN��<�X�N�vu���3�h��ڵ]3��?�S�l���/;w~��z9J��%̃	�Y���d�<��˶c{�t����Z)� >y�kOږz��;�t�C�� �s���|�����^�y��t��j{����K>@CS��PC��
1H�>�w{�Y�[x$�3��ڴ|l�Z+_}��x����?�?bL�[�iqʱ��?5}z,;63 O�6e.���H�g�E{{�:���f0�T����B�Sx�J�*���9�!=�,%�`C��q�o�8���/�T��\®�j��H��c�-	5��k�Y�E�¯tѮ۰�#�ΙI��������t����5�)�Q����2���6��1��!�J�C[g��^��(~�  @ IDAT���1�؛��f�MF�l�c^EQ�a�!v�>�|��u{������n�o�m�M�Ib�����t��9�0�:�����aY�ƽ �F����0��
V��+�c.�ދ������?x ��4�i�� ֱ���~U�gc�"x.��FK�n]�`�-œ<�-;�>�?~Z�D@'�T}�����򬃯��6
S֓	jW.�����ۑ_.�e�#	�u`���\U�.��߹�s���ݲ����r[_|5��r>�5RZ�wo�%�gs����w��m�]�\�;S3}X�@�5n?�W�����t��y���KPv���*-���WL߽Eh8?�m��[�=�ȿ09TG=?ݬ�j��B��Z=����#��ٟт|l}�6RŚ��7�����6�%F=ږ!�o|d�aϔ@�ݭ�Kq�bĐ$lð�E/�!���t:f�Ѭp��R�4W^��W<��/1��Z�}L�ۥ�`�Fˤ`��E�'��Ar|oZ�*a���L&'
���>�i�3�?�z�W��`VÓ$�W9�y4��ٰ�a���&��_Rak�C�fp�IO���{e5}�o�UvN��ʄ��@�'<�����6�\�ݴ�nDƄA~c#�7X���$�c� ��u���e�'��,	�K���z���2��C����i�-V��'ZU����&�M"�o��I/MO%,�+��6��lwu��A2���	ϥ1�"_P�8$�0SK�v���Yp±ic҄neh�g�������!�������9-�Ր|#��	k_����|����K�ÃF�T�S�)�lڿ���WJ��h���t�@;\|��(������a�c���y�o˴�<�#�K��o�O�H�~uu�)U4z1���39�R4i�f��>��u��*��;ȩ�ү�lP|��s�b�-x��{��0�T�T�� i��)��/������}�N�45�\�=r�d��.�$��p�M��|T���������@�m&��M�@	��N9zv��iCu}BG΋��g~��]q�n�A�����+����M��0�Hc�q��=ϓ�o����>��]Oa�'�Fx���`"��d�f�V��LF"NX��U���n4c�H�ӡi�f�Q���:�*p5M�4�򎢭��ƾ�>A�R�����/� b!pPX�L-����4�ӈ�F �༼)�(-�\��|��1P��|����m�%eG���Z%J3Z�cA�JfF�!�{i1e�pp�T	K��e�D�Sv�Gt��F�4L�4@��$�����L63�]�����m���P��4J���bS;���H���K5Գ	{���<9ƫ4`�5�o��M�C��.b�i.|�$���
^�NƸ�#��WmC�����\meLG� _�2u���˂׍�^�H	|[��a�U|�l��ѾH�v�d������k�H��܎�OOXe�!�4ziҢ�cuF����Y�D�:~Z��]a��*�A燶H������1��641xC�����d�NS�� �������B�F "Pkcq�a�*�uL�ݙNc�j�I7�2� \��3�� ��V}Gyc���P/�|���u\dtu?�PWr����޴�n��j����j�PD�|�P���kK�A��bD:Zԓ�ulj��8��᧲aMxFiL��OV��͟o�Iv��'~���ay�6@`�=�a�T���+_�;ФU_���^:��n�-M8�>�l,~ <]x;�=�LVYGP�݇�h��W"SmS�����E�:�i�7�ɛ b,�NBx ��{�Β�u�+Ak�V�����'��*nZo�ڛ��Yܱ:a�>.��>�d@
���>Ԗ��J��:`Z��70�����q�Z���i+(ў2(�U�V����M��i�-��eN���!�������fl�h����fPQ��|���eM�+/%��|��#��p6Bw��̀wiS[y�"�\6�W�^7GcV"�
��u���4J 4c`���2g�n(^��҇����4Wf[��#��?�5:�=�ybC�4�g0��;�^Nş��mS!����W[	j� �گҌ $�ةhV���h�7��>y�:�yww��b?��8*OI/C��H��{!�˧h�vPQ�3���ʷ���"���c�=���^Y�[D�������C�����G�S�h����%z�M����������{��X���\��捼�-����]�SQ���uoX|��o�Ń� ��/]!��9ܯSE���"�Fw�x�rM>갚�������!�AT�<W���4����^'~��|�{^׉?� V���0��4��v��pݜ����|[��d:l!_ׁi��_��x`�c�V��r� 8>¯�0:�)X��=�a���~3�0��c���K����o/�����7�U��Cƀ^gdo�ȇMc^I(��U��6f��������)[]��:E��j �S��^n������9k����Γܹ���#4�?���i�.�m#�a�W�T��{���mB+cD_~���-&�	��IM���e[���T��c�5r�U�Z�򯢳Z8��� uP�^J �*\�a�	21�]�����	'xp�@ͫB1��d+�)�B���9*d�p,�J��3��}Ls��O��3Z������`)�_��� 7x)F�:�Jm�G�uC�b�	�G{���H��T�����w�B1:��7�it����X{��+��.sH��j�`�f��W�>����y7>-,w�~�v��箃���
�KQ�x����(�f�g��c�2j3����C�3`��19�4�iw�{G�0ڏ��Yv_ ��L4`��NxY]�&����>iDs$��C�W=�r��n�^��$4y�f�o���]ؖ��^ډAu��������`1$�yoJ��~�����2(^��yu������&<��G�@W�ܭs�@S�_z�-�x��%[/��Y)����n���e�=+hk`Gڥ#�9,2m\?P�h���{���MW�y�٪�4����aB:A���V�h�N4%y���v��8��M�+��{ �er� �"��?s�\8�6��*ky���J񱃓�G����q~������r�r�v>�NfӸ����m���Nf@�Z�h������'�
?��Ƴq~�:0@50�����w�~2[a����c8�ߘ T��](á��%~� ��M��Wn_r��5��3���T//r��$W�Z4`��W�w�ڂ3�8_�dA_�gr�vr�ԾTξ��Iy]k��Q���AȄq��և­W�n�����ލo�G�~_����M�ɠw�y=�z&0���z?e�5��{��U͵v���JpOCQ�a���L��B��z��J�轕WT�=��o2p��{�cd:��4�p���1O�S�~�WzFϛw¬�Fw��=f�i��o��w]��U�y.	�)��J�4�0`��z9�V�[����C�}�X���sȯ�kt���)<�f��0}r��d�O���w����RM9L��T�т��i�����|���i3��z�1��������{��ǐ8�a��������i9��2��	��x� �������ۍ�Ĭާ���~�����_��bf�N�^bVX�߫	[6J�5.�o�f'�i<�SL ���\޵�ӝ��O;?�n!B�V{r�&}d�QayXi365ڱ��Y�j��2��V�SG���ʹ���;z#���5vn����B���6�t����G5	'Fs����(�]�Fi'���ZaT�3�%\� NpM��Ү�#�����t*T�~g �8�A�r�7�ǎ����~S˳z-���f���?45*_]Y�η)���;��縥I���b�L#���F���Fb����ws]8�.X(�ɵ�6�r�Xm|�O�Z�1�e��.Z~�7u���ђ0��~&�b�����Q}�z�����|w����%�KS5m잆�/l�@Q�2�|�B�<ǖ���5���&m���n�A��4�Wi2�8GU���3��^�[���T�M��Y� �ޣ3����BP �Qف��O8Z�W�������+[�	
;S�-N�H�W�՛[�
��V�|�Y�8	���:WS�Z��*��!`�Yko5���Y>��J~���K��om�p{	vc�|��=~<�f����{��(@n�$(F(�'���	`K����
�޲�i�{��Fc��I�e��A 4�|���rSq��stL<��Ks�����"�L�|2>f.�/��
9�?�=��M�Z�ʂ�C��vi��wA�~8��m��Ғ�l�ӽ{/v�����u;;�������M	�_�i�Չ<!x4�]�).P���U�֝�;?ݸ�s�N��'�~��M-'�Vc�-zl���`V����M��X�����u/a��`��ŋ;'�l��<}4���3@?�e?�g��_4��,!ϬJ3��ܽW]W�m���J�}D'���t������RWS�'8�6�J�j�~:ț�Y�uL�	�}��~=��	���c��o_O>�9x���7����{��Se��ʡ|���&�T����ޅ�m:�_�Ҩ��)�V\T��3�ㅄ�3�rkD�X[bd>̼J�=@��w 9�r�̲F ̌����zNqKc��!Kg����$U�3a˯�t�ϳB�����f�᷏ �2`��f���&��� ��{��c��z�'!�C��7�斢�o���a��yʶ�HsT�bu@���T��q��H�ZW�A};��ei@F/O�F1�<iJ�0����3�ҽUay��g�jkP	����yy�<O�|�ޣ1f���QZ�׭p�/��E+o����L~w�ɗWs������Q�N���c	+�9�4��ڈ�Ȍn��,��͟w�z-��i��f���7EJs89k�VQ���n*	�z����8&�6aȶS
?�4ߥ���}��Y�x��eU��cH�T����b�c�!Y���)GP����֎����1sK�-5������;�-ӦL;
/*��;v"1�����k��D��˦$�v W��w�c�f8H�3^���Nt�h}���^�A���Ш��hߊSV��0ъfB�b4j(�u�+��6iH8�h���1o���j�<��ubR�s�`�����UL�tu`�G(���:�Y׆��G|>����	�/�\O���/�0M㪼\��M�L{1ӈSΥQ��x�t���'�M��9Npt0|fʆl���^�#����{8�I�#p�P�������lK}����!H4]�;Z� �،}Qth�"z1-�������D�J�.�Ht<+��<2\��iw��X<�
�j�P��9�XL��h��8B椸�Ug4ܦq���a�6>� n6L'p�n_W_��9�W���:h�����V7�`p��&�WQ��6�x?q��]��[��e�PXH�˩z��:�����������+ߑ4^�����p��6g����V�{�B��9hG��譶�C�$�3���ӧvay��V\�3Z/}���#�O��x"ܢ�m�h�g�۷��Q6��o�s>m�n,�X�w�o�^����f���.��9�Kh%<T�i/:��SՕ�ּ���������MX5a;s���д3��pR���\�q78>D��,'�U'�++e �g%i}J,X�^���GX��X�*pG"#.I�q��OM��3��D�c�;���ud���n��ϡ��Vf���2�gh�g�)�f��k��yl�
�=OAW=D��g����P������ԁ��uD�f�2D����f)�<*�A�!�^W�V�H�I�e^wLa��N��h�a���M���
U����S��G�6�|�GH�bA�Ŋ'�:�ݪ����D�����Fܥ�'�[QJ3E }�@s��rӻ���F%�t&�\�*<�)#+�i#Wӆ��-�6Mw���;?��Vۻ$�$\�8�eL����;�)</����|ԏ��ux�Qf��Sɋ�RN�V9�6�F�#��}�JF+�;��8F�zf̞��;�L�_�۟F�p��?w��4��P6S���u|�15SCF�����t����?�T��3�^>�v�s��kM�b���C��:����?od�Kjy�G������q�~*��Y���*��I*�O�p��[/�'Ԉ�������z$G9�s��%|KP�������:�/._�m
c���}���EX����/:�੾m`Ξ���[թe�����y.:��`w�&�!��N�w&�6�o����J*�R�c��\�:)ndo�C�ǈ�i���}�'�5_q��(�=Ѓ���� �Nb4��5��9�ƁW��~���e�0iF��L�V��Ѝ�����b��)�n���Bq�+�� ����DS;'��/�N'����j��ժ�˗���iQ��6yw.���;�L�O�o�ܹ~�f��fZ��!;����M,ە̕7��(�0}�����4h�8�%̜
.�\���ʗ9�<�9�
�h�Y���U�^g�VD�h9���.[#J�=i%��Y�w?Qwh��2�5v�O18��hy?�*�0�|��;_e����'�k|�Ց���Gi��-x*7����zֆʁPE�y�4�/���]�=������l�@a��7��/�����~��Ë�pe���ai�넚������L�?J�2��K˜U�a^	���˟���{w�/$�)�hR�/A�F�Ϩ�0\?l�拦K����3�8HV������ o�1���VD/Z������3gf��{3H<��O�"�	�f=�=������V\��5��0�>
>��0<:{д����k;�nފ�Z,�:��ڊ#��mud&�Њ,Fz�`5�c�	�'o���>�UB���T�L��sh	}��7�VzN��!���&h�><�D�B�!7����1�3-7�v%|��c�;>?�y��3��SaJ{��>+P?x����~���q���ӿ��3��k񐕾��������6��?�g����c�	��MJ��j8�sӏ����iTX@�W�
���J��A+���o8������`�ςl�1ڭ ؾ��o�y%�y�q�Q�A��@��w�&���ÿ���´��Mz�	��~௿�"v6Z�'/�5��`��B����x0H#Ne|U)F-F�Sȭ��	E����K��sک���<m?����K�4���K���a+j�d��u�y~N�|R�}f��*��	w��(�:�Y��?����ֽj�i��m�t$͝�`�t?�`y=aO�d���FOU�y��3@\���9шL�|� ��_v�����=x�|�PO�X��ڍ����?������<H�@0�|��~�?_hlh������R�J ��`Si��P�x�\l}�ؘ6.:��Ai]H��Er��坯�.���U�1�s�%2�`��k4XR�m	M�ѻ��|��L y�(�;�Aa4�6���a�}�}�ɫ��/�dגSIڋpMh��Y>O��� ���-ݾ��ت<��-�K���U0Ug�~³zU=!!́QJo�U6�*�� ��v(�a�S�_���֮N�N�W��ٓ�̷�뗇����ܝ�I6)1u���5:dOėxBX�^�ę��I�-� PXq���~:�����)Z�%�������;7�nܸ1��8��_��E�$|X� ��Y��ݛ@+�	�!-��R��	����������_�|��Ŧkh�� �Dt���wUG$/x�jg_[�B��Me��N۹���>Osh{mr��jg@	���0������v�߷�ۯ�$�4��7�2-�L��Eh�s��6����<�ax�WՑIn��g2Y�Ê6�����G�d2����=׾�a4�5���������]q@~�/`��^<���J�+T	����B�Ⱥz��fl���u��rI��� .4�I��&��G�5����q��lfzdwWW����U�>�`u� o�<'�������`\[dP�fx�g߰x@9����R�{>}�X1y&#�a�Y嗑>��D�e���yo�n �.O��ޕ��J@�2�{�4�����c<>�hJj�_�N��0�����;�a�g]�h���x��'X1Z�-2��Ϛ�eL3�e��'s�Ou������PNǶ�˶+�Dm�Ff�H.DS�|�gjvy��0����cX����׽�cr����Qmh4}1�i�OeX�W�1���0L���n�{�e�b�-O�����*@�kZ��B���5H���⏼]ۯ��]lt��]�s�?_�����Q��)�I��'�%\���'Ѷ�~Tf�4d�v��=��J/�*3���v �JT��A��nӖj���	%l�.��̓�<����gjz_q/J?�/4I(����uj��5-M�6M}s�r�8�)OFP5�!��f�y��(�?��h�Q{g�	|��(�7��9�$�ZBI��f!�gO�:�Wȹx�zJ>�w��%f���^Hී|}���F�N�?����/4ݰ;��J;����SОc�y���_�$<��Z���^7V��y�L�n����?����}ߦ��q%��<Sk�Da��BxO<J�Hy�^2Ώd�q�����ۼTo�39n�4�f���/aHQ$��p����˩��?|�
W9C!#^���9�#	��1���zc��C�)Zx��C7��o�|{���n)��~���_��|s���f+Gˍ�>�����@6> 0�4�`$WGa�`�n�Y��z��_ڌ��G ;9a���pa����'�E�w����擻է��T^ � �Љ��BmB��T���E��ݏ?�)��5c�i-RB��y��}k��zv��r������'M�����q�S�~{^:m�R�@���D7��W7�o^��&�"�1��/2G[/ߚngh���>��}�x��I�G�m��_���$��&��
`�a}'�����_��6��TL�� E,��iw������S-ӆ�x�׀O�1/��?Sg�Rl<Nz�B[|xۊ���kW�zD�ǎ�J���1z*���O���b�1�Oh+b�Q�|N3vRf<�b���ں�)Ɂ_?�k-���|r���]�ڏ^�wB��@���д�Y ;٣�C�OpM��5`V2��@�@.l���net����5ؠ��`dL�Q"OJ}@\.�TJoj�f��$��%��79�@��g	��1薞X¡��#'jd�
b'�ɷU(�F�ɗ�����H�Mm��Z�H��Ƹ���lB�Wj*x�������kx�����1�f|��m���F����߮�[z�6ӈ6�D�{,�!Z�m�<<�fޟ�߭��d�|���C���w#C�˕��ԋ�Ϡ���o[l�w1��K�L�Cm+�!`�ӷ�˖!��_�o=<X(���G�p_�����K��+!Gy�� ?�D��{td"�d/��_�B��l��;`t���T�_����H�������<{��_�hͺt���'Ճ1���-m<,}m��}ny���_��wt���K�r���F*���i�9W5�Q���GŻk2�̣%�uM����_�D/��	�pe��)㯚�#%�Z�쾗�k~Idx��;x׫�`�^O���݋@Fy#�0�y�$�C�[����z���`c�#Є7�9��2rt?7����b�Μ�4�X3��B3���mjpb44G�A���q��>#.�}�b��啣��7o��q�,%�{�l̃T@�Q��sy;x�x����LѴO�Q�Ĺ�g9x��Ff�5Z�����\ޱ�� �֌��M/���\}��Yjb�8_��ѭs��ձ�(���'I�c��%,
YH�c��!Fa�-�pq�8�*���LWax�C|�N��c�(�uie��|�;'���J�����O7_������pr���9�uB��l�\tA���Cߞ{�_�;̃���]�.%S��X�8U���T�yF���AS%�TZQJ�vm"�Me�?��fj���gI8%�8b�m�/���Π��^��vy}&Xv���Hw�aT�|y�	#��yyI�y`�OF�7� \��ݩ� ��=}t9Z��׶㰂�g���{���{����RD�{m3
_?{/n>��ZFE7�f:�6����;|�j룇7�S���}��+�9GJş腢:�-n�N�f�0��SI�u-_��L��^^^�ky�.�.��'8I�9S�&�p�g���)�J<�����?ǖ�-V�=�� 5ϩEO<Qh�w�Lër������ѣ��/YL�t�Ӕ #����Y����1j¯Xm�]�)���bLyO"�vxXL�ز�<z5�h��!��6]/���;}�=�������9��u�R����9�xPf9� �6������R��۾c��WB&�6h<��@��Ȥ��%c��A��7��������,�a�M�k�+�Y�?x�e+ؗa/qI�ՃW�}�Eg������t���ͫ�wV�EF&�$/���hچ��`f��d��t�~����́��fB��m��Gl��&?y�6�ć�uS�m���b:^���{4$D�_��t�D�pi+�ms1�'ܐ���k�e���=�}x\rG�U��ܮ�{n�}��y��A�)�_4�K})[����oa����d�-��n�h{ۚI�mbf��D�X<��I)Hv�#O\�00�, =�c��V�[��w�
�[-Kq[�*a�*o%�8�v�y��z�߯�������?]��]��w�#�EP��K��3��7O���g;�A���S� �2)�p�qO��0-�L8�y���Υ((s�fx��;�U��)�}�ݜ�>(���I�s��Ȼľ`	�<izP �8�qB�u�0a˛����7�yx�t��ɀ��w��5��@N�#!�uض��\�j��w�<���x� E:#���Օ�:�&X��|EtD�z(��(㦐��qS(�ք�({�$A}���-V�n4���,�*t�#��C;ڿk�r/�x�|#�٭��"C��\���N�*�M6�V��`Yz��ns�(A��ي���:}���gM��h��6�%�[�p}�r{�ȓ�&E&�D��o�J��F�s<P��@[F� ��q�!��`C���l�W}u�TK��~����<��,v��'��ᵸ@�Y|2��}K�-�9�4��Ϳ��7�5zV�oR��b��5���pa���O���YJɡ���Ы����\�LQX�Rg@�~�|�?WZTb*�i����"�G��}a RpM��c�~Vb��T�q1t6�w�5\������'����<�N1���y{�R�>O�$�g�Jo�����iJhV�&sC��5pp`�)Kp��}jZ����ڴ�����tH>����/�������ԷK�E�/��lq�6�OJ���j�]�p@���f����I�\�?^�� �I7m�c~�yX�E���>(n���;��yM2�3��'��o�s�U�c7�^~����|��m&����� ��{�:�&�"�h׮�d�SfC�xa�V�����B�uy�g>[��h��c���'����8W��6���b�d'�k�z�`"B�s�"m�7��2O��R61jP8f��X��Y�2nN��Ұ>�V��'��*� 6�n�6�#���4��z�gy�}�@ �|`�i�i����C�l�� #�V|Xr�LTV~�����xy���Ѣ_3b���n��9!`j:n��d�/��l�o���Eg�0v/O!~���3�M�/��W� ��#0�y��^�#\'�R�ӟ҃��L'�V5�~U��n��5?Ý*ݥ����H(ӵ�S�������k�(V��o@�ڛ��s~��/}͓d��ݴ���'j&ä�f��\�5<DCDS���{8ԴW�UXw�{w�X�� ^ߞ��nRl��T�r�M�;����:�bWf�*�k[c��<m[ul���	�׼I6m�����]���J��B�)B�Ԍ��<<=�p��FeD�x�<F�Ý�D�Uf7���o��:��x�URźp�i�O�K˖�ӀQRȘ@x�����8ϓ�P<����?� X8`�"�/�%���^��b�܄\��	�J�!8� ��n�)��:����>+�#ax:�t��@���4��,�єʤ��w�Ш��g�؈n� ����^��k{y�C2����h?#2�)�*�|u�J3�>6L醥�J�6�r�`��?�(c�J�+vN��}�9�6�DSV�
He������uv����d��'�x֞;ʰq�xBj�tD�O�{��I)>��9������L[B�6}g��{f��H3�w೪͡�V�ݹ}�i�כ{�Ӵ�	���L�&ĕv����_�C�c�WG}����8�D3���d���3|nbJx+�2�A�S�<�Ե�!F�`�m���v��
�n�9
���]>k�-�ʘ�ج������
�]�	]�#l��~x8����6U}:o ��L�G�<aSz<U�m����������:ʓr|hz*�/�����z���͟���+���i�!}3�����Fɻ |^f��P�M����>�t�݀?�fm�Y��=~�3�{|�$��̓	��6D6��cfߖN����Tޖ?l���%����V@3��>�ys���>X�¼k�Qi+^����a�8]Z}C�n��Ctb|zj*�$��Lk7	730�Ao���f�u�!���=I޸x��ج��9�f�� ��YA�S��n�䓓���/C�`#��<S��=v��z������j@;9$Gp����fO�F��M������d�l��@��Q�:�쌸!t�F'�<�_�kv���V�8�w��	��ň
ox��P�����n ���7�N�Oިd��l�O�sM#��3F+5����e]1���0;n���h�v�2�1���9���{��y�n��������� @�Ko�5E�-��M֝�ҭk.S�ht���4���ݿ�4x��+�2��iKw��ךg�{8�@��.$W�۬.��J[�AV7���=l�j��6����6�.��1�7S�?��O�}v�>"�	�����x����U��{�����_ɕХ��N�*�z�ᓈ���a�>�_�#�0��R@ҏ�/ǰ!A�R�DHX�ARc�e%O���~�h���ڌ!�RƅV����R����a� 1��J9�s������ń�e��v`����dP^��e���͹��/O6�ڦ�ε:�~.�"�� 3��Ƙ�훂S�f�^J��O�
�dȝ����֨��̀:[�"�X�;[�TzFӢ9���E#�g�adF��R����c��a���;1?�=�k�`�@#Ɣ��b���/�S�yʸ~y���_~�i���}#şf���d�¦���/B�ᴼ`���
��x#EY�(>�n�`tQ�f��:y2�~�6�!#������[�_Ʊi"�3��Ϝx�
c8�n�)���׮o�g�\�z~s�ӏS�/�'Oj���<��IFȷ焅a���ʪ�>�Zߖ���'ɃF�渲��,1mb!V�Q�OX����)D;�;�A|����3^;��2� �y���Qf6�|����:l�5��D�;b����������В�qa�q^���[{_�jY�&�p��0�=�u�zg�f�l����`_=�8�?}���f���w̶�-lx�W�8�S��u�}���ӏ������?�.��FrV�(��ۣ���\c����A��8�E��J�����a�&a*�74�%����
��m����7�Z'4���;�1�r�����Q�v7_�~+z7��!��3D[��!y<��<@�uE�2�5ݤ����c�1��X�����M=)���x�����>�p�;d_����U�)���&a}�G���M����s�^!�:#�혊\+� �2����/dș�f`0��d�b�q6��{�R�k}U7,Z�������~�:y��V4�3e�ׇ������|��|48�?H#]g��۷o�0��v��p.g��.�\izR����e��W���Ͷ������+��hς�"���/N�cM��^ܛ�0m�N�p��x˙��h�kt���(c��1\�z��g���$�=�����S!���1�כ���y.�.?��~�m[El��7���җ.���VoA���p��rx���u\�����9����T�?�5�۩o3�Tfϼ��̵Һ]���i��y��#�d�⧐mޑK��e�V2�fD1��s̲�iΔ:mG��u��P���*8Lyܳ^u�3��*�w
��(ت���s�J:���
������a�Y���	9��i3ݘa4�O,�|��b

`��)��&�b$�:�)�a�pu*�#ή>āb����h�7�l]Ye@Z���� �(�����M�8*��i'�S5�Ck<i)�Y����Q8�;�l7���Z#h���>V�P�?��%ħ���9
�38��Qp�D��2z3!S��z����Dm+�V\�-7�u^���2��Ap�~���|��������iyyK��q#c����w��>`z�������a`K�����]���N���MW�C{5Y᪓{3]Y_���N��S�c���1G�٤�uF�ǵ�â�/6u� ��Ȱ$��v��٦��l�Us�`�鳺jVnU?��Y��f*,츅��>eȣ�3� tU��Z�8�me��<�ԸiB8���ϊ:��QD�3S�`b�B�Jm��������?}���4w�����fV�x6�r��3�"� ��|��8-�d��L��~�X�� ���O�t$����}�̃�����m9���3��6E�/9�S��R�����x/g=�u�X�y��}��v��9>�yUȝ8-^M��Ҕ�L�#�U��㬭}Ტ8,��	�#q��j�Q�T֯�2�g,�o�T<Pt˒G�Q5c��+W�Qk�����?�(\f�Af��VM��{p?9z.�T�5%#�U�~�Z��- D\�ZT�𧚴�T���d{�/�-<Ss텕�kpS�08]��[|W�{|(Dƻ#��̣�-/���p�s��t�C:�*P�e�-�a%��Q4�s�脷�Wx�=ئ?�����p�AĻ�)>���䓏;���LG��D��E�1��+y�Zq}��\�����̰0ba"�vi^ؙ���]`�-y��]���3{���ihwfVJck���'e��JE[$m�v�Aк]�w���QT�������)m����>�Qjw/��2V�y<Ԩx�(����|j������z���O�f��U���DK�^5���	����a������6�lk��ߊ/�gS�	J���I���KC�y�Ub7Q��p:e}��OZ�{�ց���ɶ�u�|L�_���~bJF�ߨr�.��5*�5O��"깑������nt��M��0|U����F8���鼘܂�	�r���6R�� ka�ڟ1�eo��S)�`�o%���d0�i�V�`���Gk�{��y�b�`�鳯�,�N1���eF�	��+�x��,$��)����ťm�c�7�a�&͢TX�J!F@�����ʀˈ#��08��h�O0p�yVc��'�gy$֨�q��0��Xg[ax&�z��+�l\��u����ۿ�|Sགྷ�Ÿ9��q+G�������8��ה�1:2���4���ߵ�o�׽X1����y �j����|�a��:Σ���~�8�X2u7¶2�bCJ����M�Ψό�/>�eb���<�km�q��6^��;J%\�r���+9��ݷ_n����1�,g�m/(�X��
ǝ�|�K�����}
n��
6bd�6�8����b��_�@<O�N�IlZ�7�NYB��ቡC��y�����g�����Ym�#�J^=�G+b�E�[��r ��;fy,|ܷ8e�P?��J�m�3�$�2�M/<[���0��+O��틶�g�!����
�O�j]u���J���>���zo�d�=�K����z�{�k�\yd��6hA����)�޹��L=�+5߃e��Ë�)��}�1}�;�s<����Җ����o��� H@���*>�@�9����x�woۚ$<h q�<*��|��oݸ\Lc��N����0X�����9*�4�����h��  @ IDAT�wp�2���\�)�# ]����+�X�����C�5T�|<P��\�z'���Y�	&��G�N��j!`Tp2�fɎ�	G�l�/p?�\�4�:�զzC��͓����������ͥV�����~���o�n�;M�PGK��P/��͍A�o��"�>�|W<سd�Qq�����uͰ���~�h��q���sB���juo��>��MGY�3���
��,��J�����P׎�w�%ݽ����� {��k%T���q鶹޿�b*���D8>s/��~ɖ]�e���>�3#��ww�\'Wh�7��J�#��X�jA�U-=��*Ku��-����;i��R�k5���]���.���LY�)�*���^ݱ
W���&�v%����PM�հVy+�Jٽ6��D>�l%�w뽗��PT��Ċr(�a��v��j��ۨ�Z^HXp�8����/����Q�O[6/v���`�1N��;�(��)
E|�^���9#�	�A �0@ĂR�<�w�):ֹ�y����d��5"���tJh�oB&�m�a����#��O�&3�����
܄����w���ic�AG���Q\�@����5A�#'6F���×z��5R��wv?�yi�����b*ro:�����ƍ+�o��������YE����Dm�k#U��y�����_l���HZ���/5e\�;�����6�[9h׵�W-J��y������lA�_���������������d3[x�0^�7V��1-J�����;s�c��#�駟��ܗ�Ϯ��l8�Ԟ�Lą�%�h|����1,�C6�FJ�c|���[�P�Qb����%��L��?��`.��8�������.��g4ϖ������5�rV�:@�U��14���7��P�˛���?u5�t�yԞS��J�N�e�2`�����)C���Ws�n�n�	��AuƜ����6O��>2-g���#�wnr A.0��3��Y�{?S;�	���?�C���w�<��,u���p �E�����6�rFD�("�tӔ~k��{��h8Е;3!��q���M��3���Y��Ex=�\��A�6��i�d���$ ��\<����!��D�;������?�et\on�}�V�M�X�⪡��g�����l!Ӱ轜z���'�{��k���e����'li{hU��[������j���2�N1`ЄO�5�^�* �y�x��pc�齏7���7�����3y�l�Z�<M����'�\{nݼ���ۯCE}�����~i�m�hW�nL��{��هmڴ����ʛ�MjR8�4o�	KCo��tXߙI�;Y���e0��uy�7�w�Hm�k�4�d`���Xx_y�]Wϫk�<����Zɷ���tJ[2c���Hm�X��9� �B��'9A1�5B�q�(����Q�0z#�-+dU���� `���j�W�t���x�P�fҲ�1�Li@���;���D<[L/"�+k���yW���3�#C�S׀Lh(s�<����C�Q����#�����wM�����Yp�$�ؐ�އ�7��_�����|��,V��>�1��7�����
��K���i.Ӈ{�m�
|}��s�2��c\W�(�BD�I3�>8%��t�P��w�}��X��	�Qp�`�WR�:lj�]��Âp.���8ő��bC�H���bpu{~�6�	��U���tJ2%�&Ak
m��邴��z��6�%8F��fSz	��)�_�n����\^G���u���H*u�4�E��a�zP��/72�v�BޡK*mk��!^ǹ�V���v�̓pr�ux��i��J���"��Q<���W_5���Z8�G��{\����24�������g��l�}�����F�+8�i����Jx�u����>��+�V�ٛ	ܪB"�f@��&�1(�+m-��g�2��3��w��2:���>�1��V~�;�&[��ŗon�ꘆt�:ŧO�U�L{U�x�hN�a�/�j���Fޒ��~�]�����:�
/��(�0Ė��V��F�����ԣ8�y�Z�C9p�'�C���I�����1�2f;���N]��x�L�1��
���ƣ�6�����	#l?�s6�웊��[����lt�cS[��r�pL��{���%���j'��� ӵS����}��o�U��ڮO������A�1^�%[�h�f��d*kg��}A�V�� j\swG<LŔ�V�]�w2�g<���g�5���nS�+�UI~�j���]߾z������kM�����ͷ_��w��͵�~��׎�`�r;"	�vl�$��2�O��#~2,�U�a6��D��ePb��JrȔ8=b��X(��=U���Hl��$��n��2��-��2�����Q�ޖ����~4L���lF�{dW�����5x4�z���������2���,�{�i������ĥU�->
�����7���Ō��<��o����͛tQ��!b�@G�Ay N��\\����P�������8'$�O��o'9O�<Y!�������p�U=?Ӛ)[^�ÿ�u���<Ꙃ�oԢ��O��%o��=3�X�]�5@Q�_򳲬ܮ��UՔ�A�zyEW�-�C@LV߫�!+���Ҝ�پ�_��8�!�q;e�w�n�q*j{! ����o�秄~,���=sޓ~��^�{�X� ,c�P�W�{���AA��ގ�@�l�/a�n)�����f�.�3N�Bߔ��^�Zv>�u��?�}��?�|�ɭ��c���2_�h�p.�w��X�a�����`���/t�⢲�"�� �w׷�<�rz���QA�)3#�D�[�<�H�Ry�r֏�ň�zG�T��x4�x��ƪ�2r�3�����d�Z�F�LգogS|/K�R1J6�n+�l�*H���ʹr��"pהe�ᇏ�4�-(8#d 0䢰�*�����hJ�����pJ��k�v�
��4��<{ګ�����IF e�m�
�]�ڃ�H��4I�_������ǈb$�i���ە�~J�*���}�1t�cȦ)� h�(�1@޴��/3%�b�b����\��0mA���!�zAށ{x[���wS��
��~g�:�]��h<8x�~���ٛ˹�V�	��Q�2b0hP��l9,��cd|�ñ�)m4��2E���ġ��FD�%��ffL���G������Yjm�Ϫ�bF�������"$o� �Մ�$�`�Z[�>M�;���<�;��b�r���k ��#�;eo�����};�@?��>���"{T�P�j��ch��⁤�M��ys6��c�y�\�;�a��B�2�.ğw2Vx4�wv���2�+����Ȟ��0�����V-�p���T}���Pn�~����P�NV�U�Qz�ut
�P��y�F[=m���Z�w!ژ��㷣�������7����?�3�����|�uq�7���U��R�k�+�8W����<ԝ���ǳG�(ӆ�du0�/f����	1S��ٙ Co���@)e�P�oMw�Z�Y���a�f��4%Rn ����c�u/��b�&�yT�ض�����w�������_�������N�����Xp ��\<�'*y��q�V"���|��Y�h�a����"��Q�~F������f�E���� �U��eQAy��|h��g����Ȇ��Wt��lM�+cʩO8�7k�R�k�9�y����=������U���p��zhk�[i�<|VfY���x�Y����x
i�`��=�Ap����)���Iӈ2NfH���}L��C��(�Rla�v����'`��^T�2�3��ۻ>Sn���&Yo��`H�f˲ʑ��tҮ��=���M!��u�{ɶ�D�)<�k�U���*@W�p#pAܽʆ���xc��X�ը�)���\��ۿ�zs/ϗ3�޾zMaz�T�1�'o����73j�|��w?X;�W�@H���ft!�7Bw4Ќ6�Fѩ�H��j'�H1ȵ���PWރeġ�[�92i;���:0��>��7u��Π1����|=�����07�E�������hۊY& �!m�Ja}��������{��4�U�y�]��M�7mLi%�KlӋW�n~����������0%_kAn�� /֩�W�-`��7B�C�֭mꙷ���u	he ��?f3�`����)�?�����݌�k�������N��;6�*�<���P�ESź�ze1E���/ރ��uG�����y��]-I�3�?�8���|o[%����p|*#�F�]�M|�ݟ��&��X7ĭ�8��l� k0�Ś>	�- ����n��G־a���)5�7c�9�U;Ű��EC��,�'�њK�u�N��V=����l	;��dʸ�3��r�G�6�1���'O���Z�b�DK�w�o�Ih�V0�֪Rm��+���x��I���f���V�b�3A��2��<#�El��c��jO�0�#�}
e���(ka#���JU�~��x/�'���6�~5[�<����%F|+����_���͗_|ٖ�R�y{k��~�fxI^%��>�j��t?�ё=p0ӊ�|�Mx��pj�n\K�SdeQ�Ξ�K��FC�A��F�����s
o^�1l����.��M���_6=������K0�'�~����ӧ�O�9M!9u-ϐ){�|���^kSj�ઘ~��ۊ8�{}f�-��	��$4z�ZE�Ó�����@�:f�r�tM�i��ƀ�Ry�����7��^�=�%�Y[���d�����gj��;>���曯�<���&��ԬZ�:���~�ϟ�����#:r?��&�n60�&��W�|P��ڦ"+�Ľ������y�� 
�����[��~�k���݉��-m��'��5����5�W�����De��]�����e��/�Oրs�|����iɖz���g�����0�꜑qhx Qg��7�����lpjէ�@?8 �*�D���j*Z�����d���R������2���z�S�zX]S�*l=[�laX�U\X��V�JYC1ǖd���L�2���²m㶘�����)�G��j���b��:��8�0�*��D���ʒ��|z�N�v�o��T�s1��Ò7���2�]7�b:Ҫ�_�W�{��ۺ.�؁��`$azj�"\mDp&���Վ�
	.OB(���<yK�`9L�0���q��t�p���6Ÿ����o�X}�	����O^n��3�~���:��c��j�H#Ճ���HxW&��3p�Q����ʦDv�����⥃�u�Z̝���Fj��(��� d���2��wc׾y���Ӈ�����P<F�W2�o4}ȳt�vQ��2��T?���X"�bђ�/X�.�N�9����Z�C"��?�p����:8��Qe���=���jcu�#A���2�V�LKJ�J��0[�w�d��AA�?���l�� c��F-�_����3�O����.��vS!�I�7����q���9酲)S�<���wS�ԃf��5�W���{�N:�f�r���=R�Lx�*R��n��z
���U��>fإ4?.C�e�q���w��D��_�g�մ[c�l�W�7_���f�0zy�{�]+0�b1+]{�/�1�s5�c�_j����/��n�����>��(�{�L�>[G��	���^�E�̨y�&��A)I�e�Ҭ)T}a ����B#f_�0F�v36�0�w�I�gd��;�6.M�D׻>c������<__3(�ЄO����AN�mۄ������F�,>:���b��-��������T���`��˟a��������2r#Z������6j�\�ĵ���a��s�����%_O�q�T�{0���=T�c�����VE+w�����/g@ipe:X�����p��6����F�m>aС=�~��_��b����x.�O��O�32���.��KC���>[��,���3��=s�V��	j\~�l!�vU6���Xhp�Z8\i�w�Өwh�7�\F�ރ�/����I���O���J_�;g�^�9�\=&>��~��څo�$m�fl!<��M�G0�%��Xl��Y���m��Qgi� �~����2v����<�v��Q_*^� ����<5~�8o�.��1o9R��_%��qی+żU���ӏ	
�{�%�;� ��S嶮)Ӏm�)�2g1}���S$9Bv��u��b�~g$�ه	�<(�����/����2�UEÖ��F��7�kJ�����[����7��ß6Oۥ~�ciN]��MP�"<j�U�ʔen�=ӦV���W��4j�1����L�:�� a� n;7�>0Zt���l,�vB5��+:@iwL�@f�:����?����լ���:H����^7gv�f�Ssc}��r��&e���ި������'�q�f�b+���~ؿ�Y�y�}���Q�h�Bt^�1�D��]��"��?LL�XuEIR<sďX��A�2���;eP]����k�xc�V4>�ɔH=�?�V��OE;�Z�^x�^����R_n)R������EƋ��J�wF��fu�>�J���" �1[mԿ㍁�-o����f`����p��B.�r�7�0���qG�[Z;?�-�U��^���m����qe���*��mh�i<ʳ5�sX��GGFO��҇7�[��O�֦s�.���|q�_��~d���gq��j���g�߾}g�>i�ͻ�0�j��k��o���8}�z��b������?�����Hn3��b��8��N�yt�69��Y���a��;�qZ�1��7ښ�z^��;m������-{�Q~C��M}���O1[�mU�K<!/��b�ӣ���@e�d����J܂�������bag����ǧ��Z�y�f�6m�ѦȂ��d� �W��l3ݛ!l�,����֤,y"����7_[��Rl�yX`�l��F�V�̫߯T��B&2v�%�Ԋ��e�ch:�F����4�\����]�ȭW�?D;IЁ�v?��6ɠ�o}�v��3��#�>��ng�~4�C�+ӡ�>4��(,^ߑ��1��^�M0��s$Ѡ�Tog����Ykc���ywӿ��g�9uM���4�#�Wm�<���Dr&Z���][��<33�}`�N;�F�;�w&��cm`���Z}C��f��P�?b�e�����^8���ɱ�0��)[��=1`��7�$�[{Է`��q��w��5 ��;�Jhy��juN��� ʬ�X�K�s�cr�s�ͤY��~���"<%�j��A�\*y��m���G`Wxy�)
�G��g���b�y�b��ۣ�p���K`��
������h���J�=b��S��1��.u����	�ۭ���2*n������B���x�Y��W�J���l���f��U��m�Q�q;��օ1�"4�S(K G��럒�߿w�Eq�+⍹	MH��s_���+��9Ic��b��2�7�%�wG��b�$�v�{�0��m�z����*79Ak�ϯ[6�E��Θ3ʿ�a�6| ~�q�e� cц�Gee|9ļ�;��A�Iަ9������D
�iӍ�`�T�r��a���[��ՆQ�1|h��HQ�3��i%���\K�`K<��&C~x�%d��l�XA{1�'e.��R�傅�bQq�`s��y���d�1XP+oݪ�P|�gd¢{};���ti��U&<�D-C���k�(ǵ*�Qk�A]c��^��z}1Z�2(������NT��Ag�mh���,�ģ��B0�����R9p�m` ߬��=7�������9�Ǵ��N>`@O�1�iQv�_lct5��������X�7���ڹhe�)��_�����~\l�s�)��9�<�3�?�{���O7�m꘷�⃷)��l�|\��Zɻ���%�E
�f�F����[PP����/�Q�"3�#��q'5������ϳ�"ȯ$:�h�J�^�j?��$۬�.��b�v�Z������C��U�V�j��A��T�����/-/���J/7H�{���>��|�AĠx����f�np�yG�B���E�e�j����ә��g��Vd��G��M>i��׈�f��xn�S!�Kكx����w?�+]w�6������Aw�I����H���S]ޓ�g�fVu��bY�G����{�̩\;c�	G#w��h4�X��6���Qd�����2��]c���������⹶��홫+M	)�򐯮�U9�_�#�a�&��Pe�4���8*�:�+�����_N9��4@` �p7�;�qig�A�`�����4�+�_�1�"��O8��{)�r�H8���~�M�na�MY�,��`�Q2�����F�,��^����,N�G�����oa���Z@���������e�+�Bt�|�!�F`�Qh��R��1Ų;o�i(�YҊC�B�XHB�3���Z������p{-b
~�:����3:���
g��F�r�i���/�}�}k��X�Եh:`/F#�W	:�?7�����]i���3Fas��/|���s��r�F�E^���$Fc��*I�m&&��oNw8khC2ީ��]bP#���Hކ��pKɜ?f��:��_��L�d�� �At�=!Bƚ���ښ������?��4�� ~3�΍��_�èUL������	�#E�`8�@�O@X�5�)���~��"qW��m����=��������� ���%�a
my����ٯ�	#��A�̈́3�͵�E�?_�#=�|��E2kЀ���;���a�Eo`Z����n0՟�N��(h�MO+�Vw���C`���r�+p�
��iW��S�ј���Mig(y�����b����R��>s�O�2<g �W�����iK�F��������f��(}���fqk_~i���]HF�.��&�P�0^g@<}�x��O?o���?�G����bp�}V�Q�bD���uJ<}���y�o��>������ߏѳ����^l�ʛ`�x��o��ߖM���j�(��=2�)W���'kWr[��	+�Ō�j�������E�Y�tnI�����tcH�{	�Mݔ��.��)y�n޸:<TW�0�/T��&�x���7CN#�޴@�E�%��"������ڔ��b��皭O�wz��^��773�����<�l����I�=����&/�s].m��O�M:��@��D����W3���Z|����1����_��y�1�AM�������i�=��S�$��?.���$#����	֯��S�ItKH����b�a}M@?�(k���r@�,�����q:s@���&��4]��h`bd�44!��Ķ����2l������kc�=����bPO�0��@�tt���	qyE�b���QZ
Rm���xFv�������8�|�v��C��N������"'�M֋�N�L�h*2�W[�f�O�u��Z&E�����x=�vS9�g�l#�{W���1����l'$8�}�Te������DFyƛW�!�Je�L����׌�/q6:i�qt����[��i�T��ݯ�`+�}{�ӨՈEX��"�!�R���Z�aP`ϧ�J�Q<w<�Ǡ��稜� J�=�!��Oi �a5B�7����m/���������JC$6_�`�e�I�r�"�C���ѯ\�*%���j��6����4A�+�(�%���)��s�|�K��;�ol����X��?8~ޑ9	�\a�9k�� �⤳7f��yԣ��u�a�J�Ι����3��p��q�CF�sCT̘ ��v�#bt>�B�+�npg:���-���cϭ�+&�x��-ϖ�R�+1sb`xg��VOZ�>�*�׃Q�w)qt��ӌ��}([te�5a��^LX�n�)���~F�0,�	N�Դ�[��R�hp��m<C���M�7���U���[�F8w���<�@�l���`z��l��w����(�����[w6�4�Ȟ�Pb �z��X�]=ک|m�����[�[�I�5�����nf$}��m{��W3Y��́��V���\���q#�m��6L�{c���w����p}��'��λ wSIy�W�ow|{��(~�'�����a��ַ>	��~ݟ��L_}������j�{�8�'O;�+Z�y�m ��/a+]���xq2~��q���٫��Τ��{γ����j<��KM�\,<�
O�(#���.�m2k�%�I��kx��2A�d�
���5pX��š�[�=�����S��^�˸~����x�9�'Zz,�6�"�w�
'�MǾ�䈧Of�}� ���=�F/��x���F����"�F,C��q^��`
�7����3ui��h�y��{8�)v�݀}�t����z�\���S_T�(�`_�\UR�1ps�3y_�ã��`�X���!V������Sϼ�^r��SFT��,Y�k�խK�3����4`K��5)>�ڞ�Z��L=��n�@_�<��*�o���㡯��߇�G���F=���A_��n>��vΓ1vz3�����dP�2a��~�\��it���YHI���E����� �Tn��~j0�g&,��^+� O�]�z'���rOgX��?4=�EO�ܻ>�?����fh���y����;Y�$HӶ��Mg���n�0ft���:��c����	��aiT����K^=I��C}j�ி;Ɯ^�R�Ww��=�c�o=WR�cdH_s��'d���g��PTfOeD�DBj���q{-�>��Q"#,t�!�c��wXI�w��\�����C���JTj�u��J��&�3ju��ٸ�\B��9��1�U'ehؽ���g��~���сq)�:�������wrb�\~�\L��ö[���oǅĦ�[�wԴ�Ayr��©F���GB#���픊~��5k�ڥ�W���`���q��N��5�a$�s�$�<�c��ٌ4�������)�ZV���hƈ��;��F�:`%�*�J�� �m �Ӆ�^�$728n$�g�� #ǹ������p6��'��n�&N�:�n/�J=*�LY�j�Q*��UhA�{�.#�U������<��]�,��o��a�8��F�/�C��|���w��Cyc�����4���LJ�t��_�>3�ǲ�"R<�?�Zu��+4n�Ji͎�^$c�p� ��r���>W���*�����6c$3���d�Z���Q�{�����K��Ű�c�����O�N�~��zqC/_ݮ[y<AuO ~}F�(��g�2��⍑=�A>�e
�!M���aft|�0���!xә��Z,"���'el�&��Aw��x~���cz�:�:��B���M����A�6×��8�5<O̊.�q������~�=�.��v���ί|����K�C��j(k|�sƤ��v�����0!ؗ*��G��!�s�&�a�',��n�p��f=���9V��z��E3�U�\�Vn��ⳏ;B�����
0=j�� gT�	ߏ=���K���ӧ5/�8̸�`���ن1�z��n��ڣ-���������S���,yp����-} 񰯯�:��W��]��ɒ��>��Ҍ�Q\��Y�5��}��i��H�-�&�0l��cD�7��iΓ9�C� 9�ԩgm35_>�M��:�x<q��?2-��t�v�wv����A}}�eh��e萝QH� &�� bx߻�c즳�'��t�+P��NXr�cT�Yڐ��׏�E��N�0-���������6�S_;/9{�U��u���iv3P�q��P[����9��o��W��O���~�N���@�ϲ�lG�|4�Vr잘��7�ŵmZ��.9�L�)єLJ����2���a�1|x]ۃ����:�l�^	�5J��U8��$( �zX/�\���qO����������ژ!��!�F��~���Mͮr��oD�+��m����<�l� 6
����=�A�X�X�#�QR�_�D�H���>��۸��mA��͎|)l�v�PLc*�T%a%&�-�0SB�pS#�a�� �s� �3�#���?��\W�uؕ�&��G{N%�Q�R��1�0iJ���.�ј�<�	GF�k��k��[�-��5�� .w�@)����A��C(��kD��~F��#8*@�B#�K�>o)z]8�`b�8�l6���V,b���}4K�����=@���u�iD��gmZ���\p�n�?{1�����eFy�%��B����P[������X�(��o*���M# p  ��W|Tѧ��-�T�J��=���/"�ĴcTq���4U;ޤL����)��r���9cK;�;�c�i�L��M����T̸��O�ݝ��zyyLA��z��.���]n�����o<:���.=�>��^꧋s���f�^l[�� L�<q�Q&���(.]�\]�9���:
�3ؙ����RTr����cM�c��s c����&����{g����+[JT^��]�h�����ߴڡ�V�kc��il��=ܢ+�Jٌ"��޳x}�/�vz�&�pb�|.F�póe��M�}����t}w��=�1�sEk��+x���Ll1��>�����%Nep�c����,��Q4�s� s$��
.��o3������d���΢x��
d����=H�|�=�0\����zs�g��k�ȸ	3I����m�V��J�P�l�\t#X��1m��}�g�\=D����	u�e�!�$O}�S��b�c�y��g��p��%����O�C�pm#e�39��2F'56ŷ��?�+�m����l��2� C)Át���Es@3�/8�FT	 @连� U:<ֳ�q�������ս#�F��=�M���m�Q�����wo+��x4{�R5>��y���W�pӋ�bv�͑+u���b�����T���]}�����gl�s�Ѻ�`+�@!�Gw���s����RD�ds�Rf���3T<�м_y�l��b<̨8S��j�^Dz�D�N��">�Q4hY#G���_�d)��b�*�|���c�;�!�vC��Mbt?FXߘpV7D����:�}E�ǀ�]1��3�2*��T�dl1�����腓��O��l����h�'x"���,x�/<���"ң�#�\�'�k�UH��u��g��lZ�Uj�p��c^�e0(&�w���R�T�CL�Z'bMR�#�����P.�s���,�F&I��E����+Y$��K%��+�P��e��VJE��=�Ẑ�u��x	��q�jv�'|��j�x��	ϋŵ1���m9�'vn���_�����ϴk��v5-{��O�/�����mmA�	E������[��ٳ'y�ڊ"�>��y���22N�0�"YSY�~̓�Cz�èu�7f�l���ڙ���K���u����Fsk�0<D��0Y�)Z�$>�"��?)��"&\�d �׷|���G���r�խ V�MH�k����X$�c��2zϢ��K�&$_tΝs&�\��W�0^+��0Cz��tZeuۙ���#"V���ų1h�����3h�!/O ��է��Q~��+'Ė��e��B�Sdz��d�ve�`�	������pxԿ��
��ӻ2��2P��2��K��@�]\�W�WJ�L�W�ų%؟�O<�.��w�+f���:**�2����:�9x�	�⊟;��;he�����_v�w1�[yԊ��;�}d����LY�W��5�Z���J,����<�%|� x1��ZX0'1���o�5;Z������^s��ap��ݻwG])�GA�Ds���X聁f�~���
�G�g�k;��I�56�gbB1|S�2��D�c4�|��ړY=�h�|c�����{��@.�Ģ1��"��F�A�x���pM�:o��=���`�
z#\���k<�A�\��Q�N����S�g�>C<>ݏa�2~���</>i���wM�h�'��tfP[=}a��(�.:�>y	�S��o\��I
f�������l�Nm���'��`��'���w��M��c���4
;�';��t�w����c�B�W[0�K�ϥ�H�9���H���>~�y��B:�8_q�-�8_<�s��o_��������5�y�܅�M�F�k�����x;�x�%�Ϻ�C����/��}�{hL��[�򒋻g����t�Vh�����"h�m�	3��uX`���(#/�i2��-���	^� p?������ә�����P��;�Է{�"���� �k�E<;U�	�È$�ȢFm2B:bx*��!����*�z��g�!���є�B�Jz�;0�:�;A�c�י'�l�<��x7#�����vg	�m���oM�=o��#mX���?���G��d�ix��t���eb��>�ѱ�H8��~8�6�#x�1ɧ1����n�$,5�ֽ6I���9N8$�������7�v	���0c(�iX�	�ک���O���� BOj��A����x��w�Ey!�/5�p� `#P�.Rt~_o�uZ=%���͒sK��g%.d������=��џ��lL�FP��ay���9mCq]���髌��}7�t���v�8�\����N�����c���U�n��;��a�i������J(���/S����u���m��.��/lap�R��F旯<w���`��=|2F�`�=蜻��`� oj|�.4rb���eLw��3SR^��|�/��%��t�:a�`�fq5�S��GAV7�u��g�F����YY)Q�%!Vy���w���U�g��?*�D�㍔6d�҂�D�΄�L��sp���
�"��<JH� �K;%�,R�����=��V
��g�N�Qt��և�X�h��_F+�?}�����kZ5��y��9�}��3����c�8&��89={#^�S��"#������������)���	ς͖%`tX5�!�Dgz4����M�����~Sx��OӔa���|�T�f���V[���_�@L�S¶C*k?�C"�P����?����x����o�DSɺ�7<=�*��Og��`�	��ωz�V<���<:�����.tݠ���-M��V�:K��ㅓ����9��$'EY�Cvf��5Pmx���{��w]R��_�>�(_O���U_���i#�o2=�V�SI�6>�OWZ�jk� K����j����!�?�^!0`	�x�Dc쪫<�r��*�S=,T� �M��Dd�&�Λ<�����5Y���r�:�O�o�'X$_�G6�3<�5'�G���ni`1Ӡ/�w���МD���;6.��ٌ�W��c4���}�z��d���"^���v�wA>���c�������~x|��}�j#����	Mc���J�s�2�jh�s����ms&���w�x� #�H***%b��wZ�c����^�S1���-5w�_��-�C�/"�l�|�L�u�v�����i
ď�{|��o�0Gk����>ވ� C섄b�T�qS`X���:b%�TS�D�Je�)���mt�Ë��>����ھ}�Z��F�=g�ɯ.��b���~����c5�� �X��q�kgx�����:c��`O��T������w��~s��OU��A�(�~*�����t�ѩ�^4��;���>=�9l������~��8��O�Av}�q�&h��Z?#����|6�cdo��U��}����^� {^$��?˕<��ǔAy�4z"Nׯ�"xވ�aA����<�"$h(a��p��m���.j���?U=�����(���??l��������S�bHfˁ�@SA˘�q+��<#b)^��;S�M�`:���	eP>��'N��i��)>t�3���n4�*�B�[�s�
OQ/� �/σʥP{�yqY;)8�qW�}��V�ğ�fo&t�B�XجxJ�,�iZH;R�=���@�k�gd8HXȌ��Of�qou�Nr@�,OUJ;�`0�ᾛ�#�K8� #���BH�ߥ�BQ��i�L����?E֪*i�ȶm�6�%  @ IDAT��â�B���I|�)����:�3�W�z�A_�)�t���SߚB+·��Yy�l<�O�x�7����m��A�;b�`�x!�U��O?=��h<M��ã_<�8/g�Woj���{�m�,�)[��m������qs?���(h�`Ĵ��Ĩ��A+�E{ћo�S��$�����_f����8t���o����޽�ɬN�EĪ�G���h��I�1
m)A��Fb�&�񚼨�X��0:I��3n���tr�\�^�)������@�96DΒ��|3m��q����������o�g��|d���$�+o<O6I�6C�2�NZY�R��#�d���`���&ތ�����U���@�>�� ��Q_�3F�c�xrdse�E9*���hǆ���;wnvR�W�v{�{�����N_�0�C��`M�^�����ǨP9�d���<���ŋ����o�>M�=x��sxw������HV������L}.R��9��ỗ�qO�9o�4�Iw%2��<��.S�>d&��@�������fQ.o��jh���fgޭvN`�crC]��`\1�`�1F��_kʱ��S��_�;exW���#�\2Q\��6=v��:�]��^�;�,^Cj�����(��!F����5��
@���Cp�,e�����r����V�#���Y���c����wUM9ʢ<���~L.�9cۄ��e�-���27"{�,9�.g�N��yĬd#�"2g
��~�}�#^�]�-B��챋�yb�+�`��1 A`�k�LP8ؙ\��`����Aڸ�։F0�F�g��
Sխ�1@9ᤏ����X���>8v�~�"	#\iT<%�S�����1�0��$�Ā�Za�aT��Q6�u�W��M�H	mp�f��߆�s�H@�������)m��M,�@g�b90��������V�v3C^��.����S���	5f����v�ה��6^���cl�xA�e ��pe$΋e
�����
��N6S�4�7�dJ記����X��ݶ�jV����Ԭ����Q&�;�׽�2�2�ԧ�5@��Ν����_�?�zyY�M�[�m�oz4�7�'��ד��t��l�)�~#��\8PƓB����8xƨ
f��������/�{�_4��i�)��������g`� u^���3xX�{���o�__����m����"�]�e����x��/�]A�A9�R�q�kSx~}�7�a
��������^�i:<z4����8n�y8�����lp����
�o�O��y����yM���΄�7����Q�˳Muo )���ށ}�1����:6�a�\���>��x�3m�IuA �c����-�*����b�R�#[�#wUO_)�!i0�pӅpnq���gy��C�M��О� sJ/��L�g�U�ܦ��"��9�HV�?<�P�	;R��gz���v�rh�3�! �}�9��J��3h�x����~��^��6�^�d&��NV�d8\�"�ꓒҮ���N����I�������#�)7x?��/�#�t�����ʮ��)��VSG4�?Gy�b����4��~/c��#E�gm���虾M)2@l�d��`@����p
o��pv?O���xkj��{�:~�������.m��@�{4$H�+o�rp�| �Jw�?R߶rr>�Bz>Lg��Xͺ �<�����m�<Q��'Oҍ�A�C� �z��v6z�k� K���\p����d����=��[rqktW�¶(?�I~Р._4�q�����c4�Z����ސ�zVV�"�f�T`vz�S����m{)e�&!@��ح��@��W���M �z]��j�� W~U�Ӑ0���%�d�)��	b��^ֱ3��t���Զ�Uz)���*��L����.n�QMI8���'��7)�>"�[��A��8w;��N��݈�/��t�,7�O`���[�Y�5�v%d����}@�	)U�q��52���i+�)Sy�2���d
��8��b�,zx)͌?����`<aZ�F��X�a��b2A<A���x���`��ʰ�~`
W;#���3JM�G�Vb�'%2<������Z�_IA���H�j�ia}�c)
�>�d1W~=��o)i1�0fe��#��~�o�V�ѷ[��|�'|j���V�ӟ�'g�_�أ+Ckv���[�*��N0�x����s{���.>6�\�OwA�a���ٖ �R�Ѻ�̖PG�p��!�*�Z���� �5�0}����߂�P���Y]\��Ҏ� �$��3���)'�#X�a�Hax��~���t?B*�F��q��]�'=#��W�Nù��L���~Wⴝ��n����W���|�|]hb�j�<��!:U��2#/*���H���;m�'Huj;�ªVqH���Xr����������U�D��tes�Sntw��'����y�s�Gd�����@�w��î<���?ˠ	�b�G/vh7+ѣ�aeA�0���>��kOy��GN:9�-�5X�0O|Z4qx�����U��ř�m�i ������[p�	;�â�X��b�g��w�3\�'dPBx��x�3Tj�s�G�X�i����U�7Z+,�NG}�m��A(�>?I������.����4[}�� �Ed�F1&ч~��bߞ�j��g�J��&ܛ�e|0<Є��1�����pI�����{dUx�́���0df�$
�z�Ȉ�|Sy�&��@�]����@k�t�_}�����b�1��$�1���Vn������ýR������~|G�R��5�*��jZ����|{�����i�����%�} E%�K#�}<Y��F^�0������B�˺d���t���RN�~|;ߝ�5Kk�RxOl}}#��G�|�&����[x�T8�~w�����F�I�P5k�f��d��t&�G�SF��à�X�]�m�J�fV�oȆ}�l���8�hzw��|JkFZ����������(�f(~�j:�έQ��|��H�E4�«���C�-ZS�B�'=\����̳�~з�0�g�_��[`��^.ä�!�x�鴦X��o��.~�$E�ْf��;���ԙ,e���_��j���cs�富/��u�yv�IvZ#��Nap�	.FF��sm�N�C4:�$32�	J����	���"ɝ�k����'���S��3ȁ��T�b��h	p
0���bӯS)"բ*z_�g������IÅ׭pb�1��y��2�Eg�`{��8�&�w\��|�:����W��M�
�&؜�y�7w�W
�?����[�P%�rG�L{���ڮ�x�������T�^c��/R[��M�={Z�1#��^y���Ǚ�y�!5��ʟ%�nJ�������.�Kf���׬�]%��Z0p���X������Oy-[}����@]���0��#��?�4��,�v�g�F�]��	��@�_�^Y�Ͽ�N��Q�w����w�&��y�口K/�@����׮�yԟ�ˇn��8t Ô�`��L)ۮ�&�KZ��7ܡ���I1u���.^X���4/�޿�������B�mp���yO�67:Jx?-��껐�{:�U��$��~�>oޞ�]�b1��m6���O�� �=2�h�����㖂ON��>e6�^�����H~��9|�f�M['�mq�QF�Ŷ� ���%������-Ph����_L
��}=��61�^��uo*��VZ�)C����޽�����O)�8��6���F�6�!\�M[�WC��go�^G��gb� ��d.UYY������߂=����U�{��������gnq Y]�ĉ_������ͷVl�3Ƿ�"{딋el�tB�-�Z�ͻ�c�s�3ᜄNJ�~ �r��6���e(ѲϺbB��$h��d�%�ж���t�ݸ�G�3fe��c�&kJ�c�r�M.�J!�İ���v�����~u���«�|Z���?W�]��f.H�y�q����*.gtH��!�g��(�iP�O���ͦ-��m��c��2Z�|���?Ŧ��(�(a�9d��:�x�5�m�L�N�ɛ(�~[g�o�{/;�^�u������o8����*��g+`��&e�ɴ��C)�ii4�*q*�v�	��o�e��{kTmc��lQ�C] ,h����GOS��:GG�!������$<W3Q�R!�0�O[���r,�J<zPӦ��P��a>������	F?�1Q2�S�D1I���!���w�+�ql�&�C���x���R��u�`"��:c��0(m��Z��?eN���B����O��o��g�Y�ϊw<g�O�=Z-jж��w
��̷���a�3�u�0���N��	����&+�
o{Q~���;�C�e���Tx���O7����|B�'> ��-�v����G*4�������^�Pj�爵�l9��c��uT&a�/)�Xp�'��¬�U|=҉.�� M���o�Ɋ�յ�ŷ��®��}��d��EB|�2�ɛoi�^Ӡ���U(e��_f�$w������>o������:J�C.
t���/�;���9���<G(82BG/u$�H�'���<��2q�ef��l��8����94(6�_!�a�>j�r7z���U���'�Z@��5=9��N�6����w���a^v��x�ᰐ�/�����m�^��԰�^��Kܤ��
3)����7�=i�γAʓ8��M��*O��!�����A�/.�9 �������ΐJvw�"�­�RΨHhe���s�A�������C�G(�gX��X�w�̋�}��.-2w%���iZ�]D��iա�<'��C�����|�x��.����f��O��M�xޫ�w6a����~��X��8:Q{�Ne06����𸕲��'�|WZx��*UUFl�T�^Sgޢ8޼y�����?��Zt% ���J���Ac�������?�������/WN�x�Z�C\���x%K�~ji�a"�@P뽞q@���7���"/ʪ᷼��}�'�N<���^���{��oQiw��d+����0g>k.")�આ\eiG�t�L~xvx�6��i����y�	\���ۏj�FZ ��������+m�0�ϔ�����@	�Fc��q_3~L�vĬ��p��BFu;f���1S6�_.von����|E{��}V;�Y���S�I#ʳtԩ��c�2��I�S�+�ՙ䓴��s�ܢbI7�C�Y�n�Q�m���|b�M�F���Hy�!�w(��� ���#8��Y�v\n�{��o'dut��� � ���4m�Ԃ��~��������bV�aȤ�;\�F�:z5p'���Ap���ɳ|�l�b.Z�#|��Mf� i�dñ���PX��(,-*`�����<cr67���/�,h㇠@@�3�m�	�DA�@�uŞ��:����!�m�����d���_0�x;�e�Z!J����{5�׻M�>���Yq����N]gR���޵�i<���U��>2��!)��r�=��2�?�,u�`��`|O��#N�(.�6t��I�RO]�FƪJ� i0�p�h5��ʸ��`c�٥�9~!q�����q�Ϋ��PP����-��~�8��MxR
s_��/�a�[��
,,�K�pQṁI��16ƚޟ��e7����P����&|-��LV���d���ǋ�=^<{��I�5�Ǟ�
|{���g/���(_�Ǎ}]mkz�^�C��4��*���D�PKuf�_���CӼG�8��Rz�|�g��}����k��0B���FT������R@P�͓f�k�+{�*Z�ꢜCK�z	�|[F*7���E8�?�!��eo#U<>H��J1o�%������P��=- ]歒�'����ю�/p,�-یw�6<a��L��M�o-���º�!{�03)��\'O�)�Ic��x���M]]��**"6Z�v��f�cz�3l��\R{˦��[�8��yb���e�C�$bB^��q<�]��5�]���OQ�>A~9�w�a����z)a����-��2 ��q���{��`���)��x�6B��ޞ���y.EbCu�����]��7���X��޾���j��o���/;��i9��ʠֵQ��OY���Ҿxǧ_���KGy��rT��\��Uxr�4��fBᮬ7�q���k?��$$d��)G^�5s��~V�SG_y�ߟ���ה#�R��r�*��B"�x]����{T/�U�҃�	��+�!)%i�y��C�c�����;���#�F,|�������&<��~���ho�̆�k��b$YF`�Kht�z���p!>�D�*��%�i�P$ 3�>�3��Sh����5�CB�Ќ�Z��ᆛDQ&H+a��#o�CZ>w��޽�jsFB�1`)��1�B�`hѝ�M*��c�^aۉUz/���`o�{�V�/L@�fNf�_f��e������
/��(�12�Uw$d�x�c�T»/�y��lID��Eʆ��4$Z	4����|�D�_X���o\|ϲ�x�d�s
�\e,@������`���&�}�i�S��� X6�U`
#�&�UP櫮~���:n\�&o��f������-�6�R�I|`��\q�>�}�W�ȓ�՘��G^:|?M�J�����.��Tn��[��?�m~�XA��vO����	<Q�yFH�G6�*_~�y����o�9�q�[	����w�Ç����p6%փ���ܽw�Ɣ�F>�O8:������/"�H6v�{f�u@tp������ַ�/6�����q��S¸��b���L�;G���9b
�6���̳�����o9�	��4�*�v�\�� �/���4��K�������8��0���Ӽ(�D�A�B+��DV�����Z�˚�� I_�׷x(���2�Sˢ
J�4˼@��&p6j��1?>�6<x�C�&�?uD+�J�e��|���Iᤒ
|�k�N�r(�� ;�(�Y�b�4m̗�ĵ�l3�|�h=WyU�߆�ᒛXU�����7�ŝ[�.q)�w(����!�P��;�ȹ^(觘��;�q��m�y�n>�m�~m���)z�����)�
O9/���'�����Ҡ1Iy���y'�M��������r��tU�QY����������p�)��PsA�
�Jq�m3�����x��4I�]:�{p�H�	�{XvP#�I�33��ĸ�_���(��]t����ӝ��̆�.q�;n���T�*�k�,��]_W��e��k|:Vȹ�x�Mx}�y9���ǁ0���s�+i*/���L�>O�#��Àȱ��	��0����y����5)��V���X?�_$S�n#O�b��/�3��3�X�6]�����<E~#?j�k�!����H�U� v��,[r�J����
�!\��+��A(K�uH���^宲�8#��[TK����s��[�o,��q�V�"����صw���4Pwd�U69��q��#�������<�D���l�̳�@�\��-�&��μ:*J~�)�y��@Gːp����G� C �
<�[͟�������8o���4nZ�v�N$�y�g���|�$Z@�,q߰5�&- w$^��)auK�D�!���+�xW�E��z�N����qT\u3<��%�Lp�z�i�=`KC`�W�y�*���g�����E��8!N��#���>Z�a��	��շ�Vf�Xv��4�z��*v��חz����w��В�ʞ�2Bj�<�b�8���חV���`R&p$w�$�*y�UlT&N{�[}�5���9��s$ﻴ;� ��
�y��������l�ʐ�
+i�Xmyv�VW"�?����[�8p7������M~�e���#��(�n��
8��\�B,ޥw��t�>.L;Ҥ�:E=�+eK�K%�F�mL�F|B $��]x,?漕�.��Pײ��"���(0��R�Q
A�����LJ�Y�����4)&|��&���#*.�)K*��bXa%�����I�8�����Q�
�(ٖ��a6{�Z���k8�Ҳ���O�Ļ)3�1�4g�e����*�[ޜ��@l0�
T�8����D%k�6��7ن%�����&�Y����yB�g;�g�au�<���z����
�t�ʗ���¹�8I�Q�(`�pF�-�7B���|�ܚZ�hY:��$'kر}a'�e��@Og9$D�]�s#��ȃ�s�+-.�i���,/>�2�.�Z�J�U%����
�@Xi;�/_�}*���H��rŪ�3��B��,���弔'#إ�K��[�J�]z,�=oE��)!^�I���@M���M���Ͼy�R��x0Eg���C��r���4�I����w��3&��V��"��w�×�/�c��l |��c���6�mdR'��>�ty�}V;�!Ƥ ����Hk�m�ت�̶�9���F���-fdR��k��_$C�i���N�v����TV9댱��eU��<����Fg]Ep��چK�]��K�b�q�;�|��a��Bp�5-|��N"��%�
yQ LJV�����iŊ�>�� v�,�A��'?�#��6^ߌ"C��vN%M�,�!�)����Z���?�7��o��w���O�s���l~H�̞�gN��9��N�x�|9�U���� y,pm5[sZ��-������k�d`D�-�p�69�-T�'y��tX\�
k�G;�)����(P	6K����K;|�	�D1'x��;wz<�2� ��k�B���
�]�,�4��e�������A��ٻ��k6�!��2� q%�gR:9ڭ9~�Z�^b&v��V�è��*kgC!���E�R�b^x*���EC}���״�`�~̞N�,�u4�%*��@���0~ʾ>���O�?���s6Z�c���3L)���Ќ�MVh�$��2"�a>�t�0�ݿ�y`��L�u��!"�Nߡ����H�h=s��7�������7���@p���L��Ǭ�;�I�^��A !�e-�(��F�"���]��C��%oI!�H�⩢q��f�@�+��+vA���&�<dnTP�Z��䰚����wc���_dڂ�':�����}�\���A��
��sr	���(�L
t�
����0S"���-��?	o�O9_S"�!g�`�Wу%3���L_��V54f9��_(����E�"$I���9��=�2B%�V��dG��$r1v.�ۛ�?�^���c�l6_�%��;7�,Pi���n�c[�J7e���Z�i�!`���vº3�"e�Ow�͸���F�y5#�W9�[ʽM�#R��O/�͗�Y��x\e� �O�s%�
�o^	�J����?j�Ԗ���0W#�r�VV:���+��׈3�����g�q��%^hA]�x�XY�S������v;�vfܞ�c�.�*c����{�������'��Ғ���1�
�{>?�pwNBA9�)[�P��P"��P�XT2;�N��oO�����<ڋ���l��"���s>��=�,m�C6�+��7)Kp�p+��e�N���W%NO�w$dc��z�����FGގ����m���̬�I{�N�ݦ�Z0���J�f�f����w�8��;���2e�ᒍ��5�"5��[=�*�ʙn�?��s̲���K�<�W��uN�Cltz��R�r�!���`��C�����s�#̥�S&[��w0��g��=�-��"���Sm*�A-~�$�yN#P�2���;�5^/�pm5焳�-�~$|�:��iz	���������"���o��n�g5bSO<�4�ʯ�GtҘv��<+�D�>KQe:��#��1�����P��p�?T�\���Iϵ�E*�a(Hf�m��>��s_���j'��bU
�c���<����c� ��dC�e�X²��8'k�[6�<��(hΕ�`��U�\ ��׿Y|��/7�IX�v��s�n��Q|D���IB(��� 8Si����g�e� wDWʮ���7ro�nC�17��U }fn�A��@Js�S2�O9�,q�\���?�h=Qq�!��s���+�*F�}�{YiJ�������(�)�xL�(#�������r��
8�I~�=�(g98��&�*`�������!6�9�n���X�m疔R)��\�N�P�Dߎ�e�!֙6�ކ~��]s�ا��a>��7�-;ծ����� �(@,f�i�r���S%��Պ/Bt��f�R�T����������KY-^6��FWlD��Ҕ�3(a���3�:H��3�C�RҭG���c������>�Q�z�%H�yJ}��ez�K]��~�C��x�Yƺ�J�K�s���K��O\$Tt�F.�Ot ��;P2d�V�ʿ�}�;��w0e�'��
+@W=Qw� ���3���One���~�9+m��'Ȅu��n���K�[��SZ��pO��X��1�����+{�iNop�>�x�V��n���"��
ڀȈHL��a)T�ڴҽ���o޾S?�QH�c���\��X1Nu_U��B\u��6+��C��ڃ/~�	��9ɀ�"�:��b���_9����h�6N�����������ɢ�(s��*�`N�'��o,Բ�5ː˂�U��HL�V)ʤML��!��!R$�?�VL�J��;LR��A�/�	T������3OTG�t����Z���sOY�a�I��a"'��e�`î'�bO}i�"�*y� �B,f�g\UH�0l��W�+ƫ�g6�:<O_�2������]0�p?<(wX��F�bj�n�6�60��a�|w~�A��<�^*W�ˊ�/nZq��"l�H;�������� *�S�`�m*��O���!��ơ�t�����a�t5֦c/��;�$iӴG��*�o�c���e���4\Oݴ��Ĝ+�Ex��y<ZI6�l3�Cga�㙮s܆���u��A��Ϟ"�%�fH妆�{�[g��p����/qs����#o^�Wv���ܹ�I�Χs��Xm��0��E4i�ͻ"��a�`��W���nO���u6��� �"�R�i�4 ���K� �[��#)�Q<����E>��S��=����F5O���W���l�r�>X��7mo�=�^�OZU�޽Ê��q�G�����d��RlI�������E3��^�e�3�(��M��5��W�Ħ��_�dՠ2ʽ��-H*=��!�y#7�Av��u�<�dG3�����>ԑ��צ�|m�]e��z]����?d5��NX�6*�n.��՟�(h�P�T�܂�z�b�|K!�*�8*���_�o	c9�� U".u�7��2 �]v:��5ʻ>>��?��U�����}��O�f�W���;|?gA.9�>��������ac�o^˸E����g>�:|S�T�O�:$y�Uj��������\�g�������9ּ.;�*d�p������N�s�ӪJ�V �P��}�%�����l�U�?�]�to�(y�U����)h'�#�@cTb|ĝ��2Ԩr�N�[pt��Z�o#G�A�w+�U�q�v��|��p.���m�wq �k��QH�|G�|��)U��-dLd�
F
�����0�;�ӧ!\��0^�T���T~��D��k(��U���A����R�*<�	*� L�u�/�+~��LA����#q\�F��<�������=<�98�%�i������ ��L�Ù�T�✰>/_�"�,
ڕ�������<~*�>����n�п���Ϧ{����s���>����"��[�;�Ǒߙ�q�|��B*ƥ@R�R�3�*iYH�{��)JX��@g�Z���榌_>���^(@LzV����`���pV���BpٱL��<fsU��%�k�r!ȏ?����?/���=aN�U+������ K���	�
��36�VTii}3�ڎC,�IyE���Ug�t�-0�R��`��g��$��tţ0����g����0���8�֍��b� 	��P����Fx�#��$�=˲�_&Z�����8��q2��x� �%��og��_p�'�PWC1.�aD��OJ~��OOp����_�WsIϙ��^�����ա����/J��2>3��~�#y��/�fcV�n㣀���u�j[X�6�\c�S/\}�����S~*�A��=袼l9g�F���)_3ԘMJ��i��Y��F�p�at±t��U�?psũ�+o�ϛ&o�b���*�%�H5�g��GG���߯<u¨�)�yha⣗�1�ĝ���
]�������2l���?����&y-��t���p1|��S�^p:��/���8ᦜͼ[��:�B�j��i�)�'��}��M_��Վ_��s�:C�iC�c�� �֢�f��"��v��=v� v#mQ�"y0w)avh�j����=��MX=cX=��Uh	��Z�&@G�tJ��#N�F��@�~X'\�ș�qn0���qU�Zw������M�皻[QTk֙��M _��K�]���c!�kK�
��܄�ɠ�^1?���o-4M3k���F�L�����y��V��<�=6�Ԍ'rJ:�ƕ�<��������8O��G�؁X{�s�g�${��1�z�g�����}q����ٳ�`X�,D�����7H��W2���"��ɟ?Vocz�U�an_Gȗ�%¥��������G:�0�,6��W�]��q���K�#�pm�K�)������/E~�C&����.��CdP7/�_Q�HR�;�_cB�fm����$}�D�ߠ��Dq��p�ں��*t�9x^�r+�N�Hi}��5,6�ԗWXG>|�����s8�s���]f�ȳL�a{���Uȉ� @�PS�8<�j/^��q��U1�HbD�#=�Y*QP%���p��gg����t�" MT�S���aH�3{tn�ꕧ!��$X��2OUf�3�7Qo�L���$�J�ܬ�Oo{��:�g��N�|���2VR�W?VI�g�gW�@�����.K�he�e楃9)�۽jd�0x'gxj	�^��(}��q&ki
?��fȻVb9�톦��,s{��r��S� $�{d��' �b"�W_|���
�=�@���7nj�"d7-�陉XM�A���9������L��h���L^X&��bP+Q){���Ooݾ���n�Xm�L11�a�o�{a�$��Ն�ZԄH�ã<m4+a-��.H�@�Y���;��r�2�y�_B�L-0�]�W<١����>��_�Xz��1
nd���2a(��q�P��p���E�\�n��S��s�>�q�g�7N�e��ɆKX�h*u�S��?Zڳ_�s&�X������{���e~䗬z�,;��e>�s�冪�7?���M�^����p�Ll2�/�x�?�O��4u�圳S`i�z�B������mW�ɢ�FY,9^�gi
X
�W0���&ݹ�Z�8}K��zL
����6$fT]�mbV�4<�� �~5g��U��.���| ��$�d3/�$��j��^1D�D�"�"mW�8Y�=�l�l�2�ɍ�T��53�#&̉ŵ��dd��-���K��ŮV5Q�5A!�a�0C���^bO�>&������HXď7b���n0���]E	*���%Q�zK����7*f�)J�?t�Q:��[��_M�R0fH_/�w�>s[R_G�M��.�rm��aG|��8��P?��4��2V�����(ԙ� u"7��vO#��D:{�X9�7Tn�Rd6�Y�2t��9=�c6�<d��|e�I�c���&�vNNU�H�U�>���eGCK�[���&_yN�[:���bt������� F��p�V����s�7�QD�)�NL,��iU��_�F^6?�Er�c�wQl\ �Ɔn���<�3���5�/{�N$WI(��J&�����b|�mK�[�t��³�����R��Ms���yJθ�o���0 M���ߊ㯁�_���
8�������4D�_ߤ�4T)���<e7o0WZ�_k����a�ٴ�:��&��u�cˁ�)'�B_�����Q!Q�⎂��o>������s�C�m;dC�41'��3e�y�.�wk��sW���p�<��o��`rVy2?b �f�%m�)�~h/�<�_8\��Q�5�T<>�x�2z ��~�]�=;�G��������p�&�byx���L�R�y�]�&�C�\��2�SZ�`8|8X,)�B�­�u�JI7��W�믊��2D�w��{�j��O��bT�xu��[<��}��K�~���J�0S&���7dT)�f��R\5�ȑ��Qt\%y��]��pq�Òvj�}�{�R�܌x+��c|Q��:5ni0eڴ�7�h�$��u(W*]�mie?��r��T�;�x+1�4��d*���_���z�,U�ۙ�\apݿu�:��+�y�lVQ�������<�F(����Ҥ�ɚ��߸po*ܴ
9<��q�}E��
fEz���>��D��I1�K�텊P����N��9�ᮣteO(��(�v��L�L�F�o��S��z�D�7oviD^�4Rı�W![Il�b�'���?���4d����=O'��D��2��/m�H���H�w���"Rp��h
�*ax��w�-��oJŐu]�tD�,A���]z-a��t���U������2�Y�����A�&��Kn_�ef�LK(��6���rU��<�9��#:O˚q��?��x��-7�� ZS�w<�H%�-�7���B�'�F��F�p���h�z�uW������&M��B�S��Z�Q�tٴ���mq��§)��,e�9����-0��=����/��{ Os����؛�X�W9ңC\Y�P�C�'�7#/�|���d~��B�$��4dڭʧ�[��u�x���+��S�BҼ4\kk]U�G�ñ�_�%�u����p�G�:�UeJ	������[>�H����W�p��[�}�ٹ����a����p(�ɹ���LC��.�IY9�X�{�R�����U䟛�~����-���z�P���9�ȕ���X53	>֪�C��a㉃vT��f�vӫ��Jn��r6b,�>���a�;'�͝ǋ�W���ll�)'v�=[�[������왜Z���I�g�)�7s��VJ�D=�,�4\��i�2�%@��gr���4�},�U��6��~����y^^��gA�ݗ�?��w��a�4��}��S���Ê]=+�a�w�H��2��;$-��v���� =
��ݛtX��W��n�z��Z�ϯmɷ̑�ڻ�u~�M�a*`#
���B��U�l��*�� n��b��Cr�=�Թ�d:T�X,k�E��Z�d��������t�6�̮��X_�.���'ቐ�� �皚�9�̐L���٘��L"C��\�,+B��1�U�/��w�T@�&�Tv3@���nA� �B����q�g~ݠ ̔?AB����I[I�db2�W1�3�᱊�\G��As��zm>�Ma(\����Y?eb�C��n��n��l�SBf"d�������v�<��LC�У���AD(���z�W��.��E^�[ȕ� �P�U��Z!;VA���1w���������Nhr�� �q͡vP�t��u
G<����� �y���Y��tw���)��!��bo`%p���R�@a{ű)>���P�w��EU�\������e)���|:��<3'L~���'C��0�>g�^��2O���<�5��P�ޱ8�]��Qݹ��.᦮9��	��TȠ�ֽT|�W	�C��a��%=N&�2�^�f��Bj^��;�?{����ˍ�[Y~��U��5V�O�y�Rp�u2��O����꥜���-ΕG볽�ethŌD򮰵nw�G�d$�T
އ��*ԄWBV�Bw�$��:ր-�{B,4(	�Lke�"kP�����]සu��{�,>{����G�S��!K��0a��;6�E��R�F�9�2�|�X8\��b���5��P3���v&�g����['��sV-��1�ˆD9�c��?�z�0��Jw,��'9��Fzfۡ�>,X�
����4e���  @ IDAT6��x��\<t�U]�t(�����Т�l0	��j��I���g�L���a��k�cY��L)��o�-���c������e��g����T�d#��Ki�;�^�3s�yM��%��c �����k�Ҩ�^����y���x����0+l�#ec�r�7
���w�̢�u�6=N�����\QgxGgRe����YFS�q�\�P�偺�'޿*ߕ}�B\;w�ju��3�*�yb=A~��)��&���������A⪧ ÎX���*HK<��𪒙h�
�	`vu�������ҁy	re��uzł��A@�hz�yhXOϽ�RA���eHS�En�Oƍ3��,�i��S!Ķ�/
�����|M�I Zii���#��+�}�|0@�'M��;���aήr��4F���KM��LX��N�*{.?�lAK���t�� ��7t%Kg�$��U��_��wA�[U�~�V�������j��vyt꺵��	6�����_��F��x�m�jm�������˿Ӭg����oP�D��ա�<�*3X��l*[4dQT�k��ɓt�B�q�6"<K����6υt��T�}�>���q�|�q�F���4U�ܕ={�Q�6�*礼� ho]�O���Ж9���w�×�7��N�zE�h��rrƍbf��}�ȇʝ��N�}��Q��6n��18���-{<�ǥ�	uHQ&�u�Or{�ױk�z��yp��sv5�]�������m�	EbQ:J���Q6Y%�zg&�G	�*e�Y��H	d�A��|�թWm1�7B��΀�HS,�+�i�v�9^�8��4;h�S���pb��ӟrn�-��qޓs ���/�������*\��g$2��	�0��!h:�(`[#�}�GI}�駋?����M��(��� ~{GY�!fNq<�[_<d���y�z7 f^�rq�,��#Z��4d%9�у[�R{��پ���\��*b�en��ŷc:
�[���\�繥���P��q��;�TŒ2(	�̱�苷�%��>�&��o��sqD�EW��L��r�%�J�Z�e$s���.����n�WyTn�_���=����<���*</�e��;���~��G?��]^-��:��O��,���3yr�nm
�fD�<u��:�$��ZPŞ}m˕�2�irܹ:MQi�<�_E��z,,�2��|l��^j<���iSN�p��5�O]���G�j"�z��e_%Q�eY����1j�}�3Q)�&W��T�#��` ���@�� �`2+n��$�=c�N�bO��R��ͨ����d� ��k��������L#�{2>��c�L��I���P����@0$�����)�Ril��`i�T������jR7��b����T���`��R!�m��i ]ӿ ɛP�A�����~�[��o�\���o�gm*�����XZ�%�M���u�D�$��t��ׄG}~�!`v�J<]/�L�y�6�%P:���"��� �Z&fTU������tX>�R�Y�p n�H���`�t9!�����WWT4E�sq��
�ok��Z����KxP]�9�\��^*u�\!S��O�N&�R�)�XN��S�"����T�����"F�km!�e+2�Ok���O��i�%{DA���K�=��35��՜���2�7��GI���ᆯ"\�{գ�dxl�E�):�w2�R-���d]������U߫��U� '񕕽xO�	Z���"p��4����6J�;��9+h9�����t 9t������O�����?�e���3q���%N����㝃K�(�/�)�*΃u�Sk�u�����,��`o��l�o�uO٘ȗ���q��_�����g����%+]M+��\[@??����s��w�dU��1/wP�\Ei���N�Zf��_�8 �}#m�,�^5/�'��4��l@]��P�Ky֟Ԗ�va��R�ߗ:�x����?�E@�6 V�
�1
�n�^Q���(���t�9�v��i�/�x'��3;SA!|	-�o䮎�5c&N�-�*���P���@�$�i���>��*=6 ����^�*ܨo�t�/�]M�)Z[�%c�ڹ��I��HX�x�>�����:<k�E��Y�9g�b-u�^b���1˓m��dC3��JB:6�?d���d�5��
? t�W�U��̭b��H�����Z���І0K���<̐B��d�btA�S��inx�LH�3��U��5�y$oe� �[�G��m�q����{���GL��R��Mh3�a�T1��[;�T@W�Q�Vj�>��Ik��x;Ds���ISK�|.��y�1b1�p����$Ӎ���!#��c��=��E9�k��K�j�]WU�(�
A-Z���Hp�i%�F}Ĵ,�1T���9�-i�QV�k���$G�黗8z52�,��V���2t��t��姫Jl����J�=�ȏ+�lD�87F˦���>*���KN��%�������7t��Z::o+�:�8�SL���a�/����#;�SZ��@��^�uJ�\�\�~҉�N��w�Wyb?�P��-����|��S�me���a��zF� n�4뭼b^��0Z~4�
�P���O�+��.�4������0�+�Q�D�Ǉ��]��_���<��μG!u�H01�y�w�yF��`��2��)��F:�ΐ���R�p�AQQ�.����u�Ղ.E7-�����0��-H���{,`O�z�h���ᒡ(%h�745?)#��)�˹�nu��h�9g/Xuyz|>�Փ��S�,�x������/��������i�H�[n��9&��M�,�����^g��<|���7_q��7i8�O���#��Dξt�\,�����;�4_ ��t:�V���(�2�P?�2 � \wHޥ��|S׼̆�����_�/�}�]��n�~�8�#��(?������)P�kn�n��I�&^�"_���
eXW��K�l���~)� '�xG��2�0_�]�A��E/��ϕu��L�\��s�p��`��C^Z7�E��)�����\���ov2���}����g,�v�۫1�;���0z�=C{����X]�';�kL���t��+|
"y<ʆQ����uMk]�b�v�`r��P<^>�V�f�-1M&�&��r�b��J�ӌa�{�k��/9[���0 ��2�̀�K����ҥ2����r�� M|�$N��g`\��c<x��8U^V>�* +�W`<��\�Ɛ��ʜ ��l��k+�| �T*���\
�NY\RH���-(�9P���]�F�5]Tb����piLm F���;o� �J�]12�D���yA�i��\-ʾ,%X[Ζ��>c*��j�v4j�69����O�ɔ�쩛��G���D�c�_��a�ӏ���20��� 9��U �O���\+�UA,��s��(;�k��K�b\L���ݟ��s�қ[�+�V��I�$���|9��'�B�нp.�;�'�P�[?X�7���F���$�y�{�xL�8h���ȏ��]bsAv�ʐ�s~f$"}�"k3B˿�i��-4�BA��ȃ43�	Jĉm�O��Q��/)=#�����4����)f=�a]�0�ࠜ9cj$&��һ�7��8��l6�p%̕U>��d�i�-L&o(�t��H~�斧v(�]����5���Ȟg�اWl�`���AK�s��WNDP.�
�;�1`h�t��+��9c�?r�PU���~@����ª۟P���;�)�����	M��c�/ߝ2iQv�F�VW�$6#�6�*��
aû8*�T�jx�W��AF����|j�;��_�p��4�]�{�sR�o��6���`�_ϊU�fD�#��<�A��������]u�2�<\��1�]:�<���QB�_���#�ڶ��}V&T�r�썌E�R.��14ilw�¨�%0<	��9
-g���	o"�w�Y���1���*��=�
�Q����u�,q:�6���@\��&{��skX�9�� �Z��?A��n�Zb4�x([������&���9��g'�'�\�Gh)G��_�C˂:�](�l�by�#t���}.�1���8�����x.1�����ߞ~�N"f�yTlh��-��p�L�S')1-(MtfV^k׺�2���3d�9T��#�ze��v�a�j�6L��[�#��}��	�!M��O����C�dAxd���
*�:?#'IJ��M"��WR�.�Q����&/^�M�5U�]�`��������G�b��c��l[���s�-x���d��N���b�킁�id}�B�R�b`őa]��ńnW�n2,r͕+���P5����[�R��^é��_Zt��2�0�0\aY���u	]�\�[<��E!�A�?CW�خ(<����o���Q�+���+c�?
<�o�'��$a�:=y	��L|�C1M��R镯2�eͣ}�3{&9,�^�g'lZx���pX��U���1����_��A������ǿ.~��{��%������;{{y>��=]��?�3e��<�u\m��:��� �B3�'�CIo�H�Q$�q���Pn�R�a��T�(��M�Jη���uUy|~,�� �'�?��)؀��x�e�}�<4�:ZG��^�e�QIp3�s�\ccR�N���KhĿ�?lʏ�$�WD%I>">?6�Q��w֦��+})_�����][Pݰ�9X�o�Z���r�.?(`QB^�/�BsK������j��,��� ���@/k�{���_��!�vW����U�!छ�.
�� ���/a��}5�X�X٩��Mh�S{z����&����x-������\���
�͌��nܢ"�+�"R�?���u�-��="�&>��K��T�:���CZ��n�^p>^�8�7����K!N�UIt��Q�Y�S��[���<Q���,��\`�TڨN�$��J��G��H���<�\M-�nq�������'�#����l�Q`�q!\
�-G���\�V%LZ�%�X�ۂ�Q�J[]VoЃ�*H�m��#�pr�h^qE�m���z���u�ѭ�g�ѣ�����c�aZ�-��)��a�}"!�
�ƪ��������B�01��4��/��1�Z���e�"��̈́yU ��@*�+���^���U��2�iZ@��/��+�u�j�ߟ8�^"�\������`fxJ4�wf�èT:Vq)D�"j����kf�D5�E��ʒ5-�;@�J��ΟX��Q�t?F���	��a �=�����Pf�pC�M�p३1fa�-�%��Aw���P>�!-��J�v-��- t%=�*,�m1�p,% ����F�[�K��[�/����s�*�_��암M?�0����w�`���P���`�S6n�*U�g�fo '����K��I�.�h� ��d޴���dD*��_}zY�,�/�
*��l𝸺�C�7$��?�U(}��ɏ
|���S���W��Bd#�<����Fx���ʊ{-m,������Uh����
nm�;P���̧9�(�A�&}�ǩ� J�kl�	����-V����r8���nOIC��ζ�j`�`R�-6ۼ����g4��l�qȐ!�d.�����I�C������ �Z�Q&\������A�z�*6bU*���cWJ*�L*����-�ȗ�:��t������F�wc�?*Xg����G���&h�a(���T?+m��h��!"8�a�鰾��$z�0�ZQ��7��*���^*�|'��9{�g5�V���y�ٶ%�w�8���lrN��
�6߭R�2��)�t� �|�L_�j���qaXo�uvHѠ����8'�Й�ҳ�E�S:u.ࠞ��V�ꉝ��V��!V������r%d�a�P �|�\x��6]���替�X)���}��z]���q�VF�[���+d9�]�&�M�����+O�vp�޹��:�uS��C쐙��_��|%]1�?ū.eM�^�^�W����1�o�����<@i���m/Q��EChK>U�;�_��V�#1����w����C�����.C竑����|%-=�Oa'��S#L�J����A�CZ��X�F���{`X��g%e����D��w�#D\�L ��q�,v*A����HC�=L�L9Vs�u<�x�[Y��BI�5.)�mJv�S�v���ZM�d(�A�-��4?�𹎤�E�u�{1���;13�%�7��:U���H.�AQ[$�"�:=�4A#&_��z3;a�Y����ѻzr�D�j�$�ƣ��ߒ���iNȖ��R��5�h�F0�-g̽|�!�/�$�9:X�\����p*X����i^V��[����!Q	�o�Vެ��'�JXS� �a�#z�kϞeW�٣"�pp����< �U��C�q��_}����]w��/!������G��CO����F�F�3E�6`6hN��	���ְ�yE()�m���ս�6����f�{lv����◟~X�z�A��tY�-��{�ك�7������~e?/������&򌳞C�f�Ф%�^b��RŎ�{���wX�Mo��>VF,h�m��n����;ٳQ'�����H���b���<l�g�Sw:_�eyXF�S��I�Y�H��(4���i��5^r�Y,y��*��� ��$������21x���������2\����lv�;y�o���j)g�+���d�ql�����ϓ`��id]1�+��^�΍��g�&��nw���Zv�^�D�t,��<�HG�ź&uL_%{��j�sfM3�,���(ʯ:n��rp���e�w��5�v�܃���D)qt4�%B>��a�}�8g�,�Ж��&]��R�*t���K\i�e��M+����2�'���R>���=�n��p��(/��D�\n?�싎W/��z閲m(��Hc[�$�qGx:,�ޅ��v�"� 8$�&���~L�Iޫ��esћt̤K�WRa�����L���>�Dy9t�<���|�p�C��p���9����z.��4�ٲ݁����yfy$��I��%hũ�R�������#X��P�$w#�*L�uQ�47W�w+(O�Ȧ��H�ņK?��YR+�>�TA���'^�����?"yխ�F<�o}��˖e`>���^�^�#T�۶9����:-���G�y_q;rG� 3�·^��Y�#C�9G�����)�������#H��ne�Td���Y�'�n�Px�]2�>Y �\dP�6,"�b+př�P�y'� ��zR�'��Y�_�s�(�u���]�l R)�UE�A�,!p�ƙo^�x.^=e��9C`���+ĥ�=%'9�kr�$B�t�w�<)��5��4�G�����u-An��2����k���`�����ryW����"�1����7���ob}��~/S�.�/><܆;��s����%P�ܢTQ.*�
���qk ��b���C!H��Sz+8|Wzk1��!w9����D�)����Z"��q�x��}��^��������X��P}�8|f��s�)
�������^9�o���Ӎ�@�z~�z��6�*!N�6_�	���}�A��*��������2|�Hy[\
�p�;�����(���s�&��#��Oty%/~�D��~, Ì��S��7N�Iю��m8�K���:���v.�(c2��-��C%Gb͢ᯎG-��ׁH��y8��P�ni�|b^��"ȽB焓�P��-�6�f�bk����v��+���xU:ƭ�T��U�U��U~R�J%=�^U Y��Z�Js����[n���q�,#s�K3B�`�Ѱsx�.�C��idxn�Ky>���I�'�����{��c?�{�| Y�H[����w�`�$��W�������iǫ�}��r�,1=QVt�N��e�έw�l#�uJ�갠ʅs���MhCc�~���h�%(�^,�<�� �);B_]}����3'��V;'�훷l z�Dr���L�ϼB]]A>P)3���:�+��׷��T3�'J;�&���҅���	<'+�`���SOOk�xz˓��3�1mA�o$(�\�]8����{�!OS�DZ�M���O!��z8t ��su�V]�S	L��#*��h*_��"t��͟+W����W�f���A���x��W� -�A�4J�9C��Dw�!�2 �����(ad^Š��+��"��bYi����],�U(AK�z��u\�ܽ�`��l#S���)��JQ�r�Z�F4��,%bB`i2���³�a�K��l�Ji^��Z��=y�8⸤�G���\ ��=q�2w ��cK�7h[%��L.m-�VtI�h%�V������Xb�$A{���,��e�l8�7�>�����R�8��Ǯ�f���!�/�h3��	�BJ�H?ũh�KR/z�\�/�]egpq�_R5@�`���G3��~ϣ��p��a{��j�|I�'DS+%L��`��[�|�7�"����'���»�w�}n���l�y�3����������m��`�B[e�-yE���^�����
�v��}[Ň�8P��1Wloo���]�]�ܽs7���nk���u��@��&�#V�)�z~�iT�J[�T�alT�Q{�Qo��y��QXwP,{e��,�t�W_����S�K9U�
��;N���W���v�X�E���o�i��C�����ź<��T��Ȥ�Q/�tC�Hov]�t��U�N)���{~�Ë�7�P�);�7L^�z���]��a$q��Hi���`�[���<O��}�,#�/��_q.˵�Rʙ�7XUƂ�q#�������i��R�����F�����(���W��s��-'`����(��y�
�����َKM��J�5�m<"���Ѱu���KP�d�%3��/�����K��*>�K��R�G��By�7�8�	R�w�Q�sAs,S:�z)ە�5c�V�E�W�PV�/�e�fc=2?�I��ռ��|�_�CtX7��b�nr�UY�<��M��X�yxzxOK�޺����8�����OG*���':�|�"d�����MAҐ�[;L`/ͬ��P�AY[�VRo�0���̓���0��Wb� /0���HE\���FXϫ��߿@u@�
�t��G_���|\������QJ�So�w:��������?K�}T&���4����E�gWkr6A		bV$�L�Uf�g�¤xF�r�Lk�;T�7Y����,�7rhIMW�m�������
p�*�L¯cQ��2��
37j��wZr�D��(c�{yiLl��.��E1�4�&�����Mb@K1�C҇p�ojz~D�c"���c����ԑP��Ps$
���Wo�/'�ۘ�\*(RAR6�W} r����@ ��,&�����µE÷��ޠ�NO�F���o�.!{Ea�8c�'#�9~%̍u� *�L�(t�2��RCq�S��g��i���0���h7Yi��P�@�� i5p�˭f����^�T�@,�q��u���0'�>s蕹V�;,a��4߅�*@?�B ���䜳�d�i����GS7����2i;Dd#VB�s�(2,�(���@�u���Č�qY�I��+������(t�K�ep�(
_�TI�~Iy�tR�ư���uﮆM�ɾΑ���/��(�*/�����ϳ���+WXn��r
y���UO�V��=`w�)�u[�ȚUN�XǺ�S�ɽz���v$�U$; �G���2�iz�V|��"��%����ڪ�@e^I|�,�(���9�(S
�<J�trx1t�⥂�I��:<U+��3?ţ�,cᩀY��b+!�]��4�"�ż�{7�?�K���+н�����uZ�\e]�&��ʘ�_eJ����V0���Y�$�HS�RSK�1|�[���?�h��ћ൏ҵ��֧y���bQ������e��?�e�P���z�U�mbW����( �[��[�e��Jn�];Zo�d�Rf^�-pt^�{E�kSڢ$��S<ʭ,��;�q�ߌ	�ۄ�Ǜ|P�ⲵ�"���tW�SZ�T��Y��o;�;�,b��ְl� �HW�j�)��;CXz�Ѡ�ڳQB��H�+�uD�O�RT\�/�']��:�N�:|$�JX"��#0r�M��{8�=CSv�����?��ߺ��E(餈���Cg/Ӻ� e���7�ô�f�_�<7�N���k$W��*!>p]��ܭ�U����0Cd&��w��Q���R0VL��ـ���#��/�@�=+��H��o�zv�e��p@��`�WXCHhb�r.�-Z:!�Ϸq%n�4���O��D�'�rSx�1�q3��/����"ߥ�B
:?酽bu���3z��W/v ?�7F#�⥐���
���x)4�j��M_���?�����u�Qb��
T�7OU���q���-v�FP� �o0��a�*1J�[�>�"���W̗�{�wp{����X�hj%����E!W8M�����D՟��Wk��������4D1�g ܭ<Z����[�^+���1�~}�$�����t��;CC$l�أ�~��G��wDA�ՈBt�K˓y[&Z1�O�k�҈R, /9DDcf#9j�,k�z��S8�̷�ʜ?���%�
� I��K�({8�r�!1y ܡ�~�g��í;H�������*~x��e�Ӿ�ܔ2$��^��Y`�`}�?�]��fQ3�K�������ڰ�q�*d ����L� 4 ��(p�I�K_˩px|l B/��BO:�ཥ�2º��"�<;�p�{��*Tt��v������~ܻ���,�����}��V�%���(���t7��Eٲ?q�"�s���ݻ���[|�����#'�`=Ŕ�̡�5&�on`�b��+�׷�ٶ���.?J�B�~�`eU9�4������Yc�WdA��u�\��ꭵ��RxXE����mO�*��F�Ӣ���l�P~R�U*�r�p�?y��O�"�u����G~�/�l�v�$���~�|��Rv�#t!����nr��>��,����V���^���_(S܀����<$Ģ�H�pDH�2�q���J��E9��f��M;����)Ǉ9Ty��{��@�h1ߧ㷿ئ�܈�/�����4*�X��0w����R�-O�"x��2�w�T�E���Z�Ko����ޠ����2\��BU���D�(��x4"�^1;��~1eF9���S�UŴ�HNBH�H'�LW����}�M�~��t�G����>�4ؿ��)�B��!D�Z���(a�crD�Xˤ%�� L��+�=�^���#�'
@�puL+f�:j�3"#e ����1���k��������q�xN임�Y*�*6X�^3�K�ׯ��	�����V���R�R覷��B�VZ�lޛn|\����61������8��I�7����}�"�C�r�aI���Y:f��׻g����0X�z-�Ml �Z� vʮ&Ū!X<�/�y�,n��(Ȕ��$=�
k���~����(�n�Z�r�2��XbM�Rq~����N�2�k��J{4���s@�����C>H�4�EV\fn�{'�;	�td��ru���1ʷsB�UR�#���)�/< 	𖞱���0n2����΅x�$U���Q�ax��&U��/���S!3�\�򡫼�KP�R�\#��[?瞦eyT�<1�m"�D�(F*�\	��	���y�	lD�`J�\����G�x��O��M�x6�Qb	UJ[geH v:NT��*�($������.�6���J���p�|���/��a(E�E!��zï��5i�U ��tn�c~,6����0e�xm��߄�]h���%K��C�d0֠tNIO�F��]�ֺ$?�麈�M���ƫxر�ئ:�'���X���VC�X�,�����
�I34�fj�u��L *�����ʗV�3�\S�~*�vD�[�W��c���I,ᓰ�Rx���ܑ��3<W�Hy#X S?��{BT���Y�H����Ͷ�\��JT�H�p�B��(�nUS<���<x��6��� 108w|؀�(`j���
�7�͈�!d�@�Q%����|���>A�c�N�kC��rע��i�z$U�/�J�g�V��-���，�Ui��L��=�	l�O��S�7��!��|!:���Lu~�#
X����{j�
��v�t����h�����۹��:�;{2�A}���k2B(iآ=^}�
�8�6Jw&��S�hx|�6=�"�a��=4S�B\q5♮�����^��p!Wj��T���R�=y����G�r���IO_��MΫ���D�-��CF����0l"�6���x�A\f�yL�����1�x�Q�D	@HyL��G)�:��5.q����7*�� R)�ͽ���``= �B�"�zȧ��8MW�Oq�䖠U�%�jKKx���ϴ���p�|I����Dju�dix���@�.�;7��lX��r&��7�{�V�D@����q*q'[�c2/g.*�����(�X:���v8��٘1w	���2dc�d�1������D�A��B�ɟV�chy3�+G�
U紹�{+i6��p���to�W�����cn����)��ż�0����"hea{�w��fL!~o�^�0L���5��S�Pg_�i�����eڦ�γ��t�b*\��#�Z�T8|�c�/�䗆�zg��rV1����ʒʌ�ڇ�����/�+�Z^,/�����ݕu�5<C��u�����4�����2:[��
��M�-��+�b��?�j���:�[�1O��Z̥��m���o�	�����{��S6 ��F~�N@뻊�~�$� �R#5 @�z��0]�XY�-ԇ^�К�s�Tj=]@�m;z��a�q�C=�mEvJ��%^;j�6���zn����^nr�y��`�a~e�
�J�|`�� ��ʏ@���^�u���r����F�Gʪ�1^�:�����5t��Tn@;��^a�v8�U�'�L��N�����T�@�֍�B�HK�vpw�p!��V�����Z���mL���x6��&=�{"�,���@.�|C�0�-L���(R��F&�.�����U�y�w�� 
�ֵ(�ni�6����j"���
3�-��d�
2���?���i�!�Ay�v��<' +���r���)�)�D/�'��S�ˀ7�D�R(PF�$R�s��F���Ty4i��U
��) d��Ir���I���;P���0�.fy?u�a�0��=R'Կyu�8z�h����ų�ӳ�7��^Ea��*`;Y`yQ�ۨ�Л�Q)�,'�P�2
sϼ��k�V�Y ������([�]N
P���\~ʼ���h �xv����]�Bfؙ��{��,-h\x��A����H�R�0V�J�J˲�@R(����h��Yxg9��lр�p#��4z�Ғݫ�qp�}�@Z�R�J�{%���_�t����V���V��b5�
���ʍC�*U�URny����4��U��%�ҽ��;X3T���A�L�?<�~��p��+�28xu����fCb���e�+~l�c}��L��,{V�sr~�bx*Ч�mBM��Ͼ��{9�yn��RJ͘;�=u������W�G���Z)jh	��S
${�QG䳺R���sj�M�x�DE�2q2z)
�B�5�I[��{�����oW�Z/8��#`)O��B{� CdB�V.�,7޵��r2x����Q�TĜ�@�8(�\��L�=N��+D_bA{�Ͱ��6I�h��ˣ�<�{�=G!S��"_HHy@e|�1��ӑ�O�J~"Ky-
J�8'WDȃZijEa)�b�&�*˩l�3M��Z.��3��/>�B3S�C���[b��:5�V�jX��
��W�_(^Z�H�vH��F��Z�2>�~m�V'��i�I����F:�r�}�:
f�,]+�?��I˖������)%Gk�
�uF#�/��������>��QI��[iF	K�d����̛�gĬ~5J0'_c�F6�㥄��N�Ys�����r��~���s2F��p�D?'��^W��v37_G�0���S�.ϩ�{+��OX���n<�o�
S�k�U��z��/�������S������<v�0)���@̸��[�m<�jdt���Mʆ�{��~�K���w�S#/�����n�VȜ 0��r�w��|�{nS���߸]���1q�ͫ�lQ�+{K����=fe����k'y�)�:B�]�ex/U7im��7�4��Lz��'N�wl��<;��N�,U;iJ��_O�VW<��&�[I/����=a'�G��f{VZa��ۿ�XAaKZ��@�i��5p0/� �Dީ�q��4�_ e�F0�0巚�E	�Զ1��*/��c�Ѱ�:',a��B�x&L�_|���NQ�n�`��� ��pEʼ��i;:z��6�[���X�`����;�5��orf��?���d����q�u)f���W:{�Z<��rr�/-�)0�E���X��3ZHܲ ��w���7���^����*N@v8̡n'�7���,���r��%D�����~ژ�i����74�𳊍�߭4�]f^L�\��_V��eZ+]�`o��a����0Pv'�6$�2��މu�**�ӱ~��C�e%���R�.������\���s�\H��J�����
�<d~��8n�b�L���,��EV���Õ��b���ca�Ppr���sx��F����]K���tM�:�ę�)��h;��SJ����ʛ�8N^�]g�'w�Î}��W�d�
k���7��B�J|m�cu�,�O_s��K.�ِ�v�A+w��p8�oRJyf�,����d� &�����k��%�����6-&W�*���W+� Iz-�F$��5�H/\�OqݡS� �[�q�s��=?�t��ǁO�Y�a�V� +L�W�eˏ�2L%#x@?��ϱh�a~����!�u�(G��3I��r�"df�W�(L��*�N�����2��IJΜ.�K���!�ӥ���W��mf���8�L�t\���J��{�ip+������s��7�^گD�)��ʃ�Z9��B�eDT`:/¥�6x~{u�Z��c�$���#�� � X���xjP�9�xh���RyQ	𛻘�O% ��l�~>��U���x��+J>e�!F-_�X��K}��/X9^Gp.���n�x0�y*6p;&쪐���m)L�Jg�K���#�1F�nV�ѯ�+	�$-���0b���i��"�Dm��ـ���r��`��˦Ũ�e���u�VOCT*p��'<�L�/s�VTo_��2}g`��P4ƊA!�z�2���dg�V�p�p��[>��Q`\�<]�P͡��"x
�|�X�d>�J����al-~����/�<�qs�����<pVZ_�����^lv���ߞ������`�U,��s�l�]�����̄|�;4i�k#~q��;�=�$U��O8�
��R��D!�J���`gi� MD7C����C�Y�(V�����rR��j��*�������V��=:}N.��+�0��A��0�Pj)�=���x��J�� �R���5�R��j���V�H���ل�a��Ⱟy;a��<eX� (t����וz6zu>��U�5�;�k%u����i�Lw�wU�:/9��mM<�*�;0����q\�����[��d�|O��y⎸ �XN�G�y�]%L�߼dr?���c��nr��%�S p��2��Yo`v��'ߗ���rV%NE�f3W
~V	�ᷜ3l��(�0܄fz�M���WC�����X-�6A�q+:T���D��T��D�C8�໼m�؁�E"!��Cx�����F�񤻂,��[��Ǥ�w̔�x���������;�Hr$�&ɤV�R]�fG��[�������nDO�L��,��*j�{��I��������p8T
�}H	�E�=��<\����;��%�ն^���8����s���m�Be�ނ�a��7���W�*O��f�y��U�&͖6�f'�	�H]P_M�ti�s-�k  @ IDAT�VK��+5&W�c�Γ������&ao���N@C��J�)���)�&�;ڀ�<I��ݍ7�6�@��Ԥ���ڤ)�u���W`镈R>xû�U�à�
=��Z�,L��:B��^�|��{�Ya�b����[���Ϟf�*'�ګ�`v�5ad]�p����sh���^$`R5�46�$�����&P���A��ʧǻʨW� �B����bpr�p�NF��oP\lp�YΐG��;����!� 40s	?�pٛ�t�E�$�T%
���-ҫ�o�*�����0��;�(̜�p��A:��s3/��·p�$�x4^��wp���E�2D�|kXִT�c�_�eN
���<FޅAY91�_��w$���BY=fחlƺ�\��bs�mM��׻�����+�Sz���Ѹ�����˹-��4��K��yh]y�����U����D��Cm���<#HC�P�����}>�F�P�ӡ,����)�-P�RT6>��O�^�e^�K�V�P�$� -��#��$ �^��H�Ǐ8L߆����̙ʟ�i�xz�
�J�t�K��~��_�~���E��(KK��:f�8>~?z�f{�˖*�L�G0y:�ֲ�X�\�;^(:CԖ�J|Z
��A����!��q+����"�s�N�����D~��F���L��pIG���-HPǧ��%4��w,�~"��s~KRq.��WI�+� ��翞(��J�ܔ���:d���w�����0q���w�l˗�۷P^Q�L�\X�{f�� �#NZ�m������5�v��BT��%/�&�1��"�t��^���Fx����~1j`��ya�f'ĩ�����٣L��M
50�N���3��^�a��n� �0�_*�$*=�vR�߲�~�S.VR���
�(���� /��� �9ù��'�v�&ca q�K�yUڷ��q�O��1	�k�>��w��z�vBP����M���k��{��G�π<��zu��UO��P���tv;�
P�R�_���,���נ���+<��bL�C�6�aJ�,�Z��(ǂcoc�?��w���4���o5Z�B�O�`0��ן������S���/�M��b�@{��� Q���\�ko�#��Z�T�r��3ٲ��
Ga%�-�$W�̋�P��0�� ����EP�����|�<�4��[ܸ��,hSa�C�*T�<��z>3�Ω;@0�}�2Ddc��C0<1 p{6�.�W�{���]}*<��� ��������%7-x�97�9򦖊%0����� �EE��1��D����
�y8o���Jc�ΰ8��a�3���C�����(��a��%���uy���m�u�����ڃ��X�h<���l�Y�Ó�uiS	3뮂s��l)aM�rqHj��\�X� �7�̪=��J��T�����U{�O���n��`��]Xw�[0�)��k��D�\	���)Vy�	�@�'�*��W��~{O�X8��}Wf��M4�����к[7��]@k��Z�ww9��r�p6[6X�;�}m=�*ڀg�/So���=��و�;��-le/��bgO�4b�tK��@���I WK?A��3�߽� ���YQYC�CI��o��(�_OO+��F�a�[d����<y�����h�bQ�ٸ����Y޻B�|���j��/34�V�S��HR+���d�M��q/��|s��v���jճ��/�R��Q� �9D��̏o�OO.�ۥ_9�[�Qs)Y+��R��'�(� ��܄����7��f}-'-1�]d(���V���ʨE�-�,x�b�.���.����	{��th��c�\y6V!�$o:U��E+��X�?�v�8ٹH��c�,�Xq	?�L��QІL�OC3o��ӥ��t�[�L�I;O�N�	窫D_��ղ�QD�"m�y��.@ed2�kJ(9�<�f�a:]at�]H�,)6�0�2�T����P���Q�u�p*��(P)(a�k�٣'W�Ex���X������2dl��n��߅��R�U��n!DZ�~��k��E40�{����!_2o��`��;�b��b���#V�z��&�`vd_���C���}����kx��QZ�
 ��;t�K:����b�Q4|<;VQ@tO��}�+.��W�'427ѽ��攡��6�E|�Z�⣅��:,(����%�F٤q�!Z$��Ji�aV��\Ű�{�췮��ȓ����0nP���H<9yP��9��!Ģs����l��{����6b�B#��^�8!h�wd�Nh����a�K�fGs��,��v��"�����U�D��Ao�����4�|K�T�EAҢ�C��h99��!ʻgt>z�(yQ��§R�&���m�0;���q��U��n±��GS	sXҡ��no�O���~n�E���v���y�?��ϔ���%��D����!���tX�[���㗜�%B9�ox��������c�ݸTژnV*:���qˈݝ��Ϛ��B���{}�
��V���2�Z~���C}*�G?���|;a�>}��Ud�{��li1�Q�E��A��w�'�G�Z������/>��͹�p����3�*ܗ��|��F?̼L��E�S.f�����*�<���O]=�3
P�7t�G�V[4pLr�i�4�K�6�}����)��#�o^)�2:��{9Ɓ�}�N�J�q���v�c��T�9�N~�D/e����b��~Y�r�?;��TZyi��{{�I�:��}V}#d�SդMLܴM�cG�+铿 �*{�+s57�h�(W��n4�6�ۯG�-��'��{���~�O�?abn8J_�<q$N�)��"5��!n��'�!K�P�߽�b.�SO�p���x{�sE��h�L��L�����/�U�Sn{��e�p�CҐ!8D�]��Y�F������f������Q��(�*��o�*�b"�qh�/&��>8�L1F���!a�kz�e�lC{P��*��ƣr8�t<�2��4V�O���a3�<ͳ;��
����/q(g��-!�����(��!�0a�v�Ɗ7�$聑���d_�����/Fq`A�U��s���X.j��}C��*��k�o�Ǻ����ɳ'(_��^_2���g��w�����t��t��g%��7�˔gAnA|�8f��x�S��i��=	I����+��Sm��b��r�K�~D�wF��y�
��ʨb!ݵl��{U*�[y��!��8�p�����>wI��֗�Y/+#�|(`	��ևX"�P&X��|�����:$�moО�P"r[ �-����D�r3�kzM�4tE$�b�Rjdޣ��@/�o���9N��n�(��/O��H5��S�ڈkaq��'O9S��ߵ#?	G!�ܨ��QH��Γ��J�W���D������M<m���mK��?�a*8��e��n�^�F�+���ͅ��V�' _���&qpk���-z��r:�Q���T�ޢ�5���bn/Y�z\��(���ƺr��$_�2��g�cZyh�Pj��WI���r�:>�b���շ��2���/��Ob�RN>��v����X�]�<U�ɨ��_~�����nkc'���*c���z4��m���
�8���.��c'��!88f�C��8��H�$�#�R|[>�q�B��U�%u��-�+���r[ƉD-��<4-.���C�ݮ$���1�I������+��'<���
?mN�7�M/	�W��YwR�ɷ�^=���u��=Hhb�ĭ�����S��Y��I=���j��u�ƭ�ƣ# ?�PV]��V�;r�\[RS���#H�M�xc��Iò0���O��о��y����C�U�^�c����ʢ�W>�6�\S��x�)�؃�������c�M����@\��ǟ�l:U�%;K7(`4L�����a��9�K��]eP�+�V]�l�.b�$�
��x_h���)�?��]\+`��N>+��#b ̟sWLI3oV�x�ڥ��X�T�'�D�+C�<5;���`N��ysfB�!V0��Z^�z�N̯i9I�b\+\Q�o{* �@��_�/'hf�
��qLCIK-^4T&jɉ�q�]��G�D��i���*`�g,�����w{��7z����ٯ>�D]�{�!�,����������4e�I��2A��H����¥�[���OÆ�)��\��0* �Ex�.CS���kl���g?&��_|������;�c	�qR`g����;o�J6̌o���2V�{:�fp���g��\�T�TV���4�+
q흹{���^��Tr�MeQf���e��{*6�(,�1	���2y�����
�?���y'��sN�֫�$�����՗_|���l_��ʒ���1$� t�59!������	�n���u���	��W��(��RK�"So�Q
��6�Z����{�����	�S��?�Y�s�So/i$�ĿdD�;�Y<U!�ʖc
(�*��N�'��sH����Q��|P<��W��S�hk����;���w�}���D>8�K,��,�b�L���ЅKXc�BA�o��h��y�ܔ)�*�N���|���i��&��Ã�4�h]��;��ݕ��|[�9"Ӏ���ʾ|I���Ip!�sN�F٦��d1q�	�lZ)bY�O�s��m�}���M�w�|���]Tg����❖��ȗU�qDn�a�Ph'��UEѻ�@�E�Rʋr��y��P�%P���u��!�>�G}~om��GVZ�TzsLy�HF���&�O����ϐ[�%m�������wB��]�)ؖQD.�bs˟����c�7��w��x��+U]��:�J��Y�+�����-8%y��W\����R7�u.˸]�2�3��W�u��@ѳF?<������l�b;��`�N>uu�,�
��摗���I�4��n��h���U�R�A��m�c��M+';H er.��Ѭ5 �g<��sN1 g]Aì�N���V2]W�1��<ixW��r�c�Ԙ)����fh�*��T�p}7�$�I�Yx
+A�D�WĨ�6!�H�xs��Y	�T�Dgx}t�Qqv\p�$N��č�%� T���{���!f�!�WX�-�x�����Gޭ�=�;)������#~2<�8�	���7�>����\���	�XZ�j����G��K�� !��g�M&.w~ZТ��7d���la�*p�@��� �$�5	�Π��h��wH��ݷ����C�� �?��dVᤂw�&�T��n9M�jB�ʩQO�-my	��U�� J�,Ow�Uɹ_�X�<�u�E��J�J��#_)��6@Yv�R	���ws����/hT�FWX/$��/8��dc\���������š�������K��"�H�̒}7Ѵ��5�52⑹;Tp��T �ʳ
����a�kZ��ȴ[�T�|'D�T����QQ0�Q�'����S�O,�!��O�;|���pQ%�{�1@�U��&o
;��ҙ�S1Ml�`���a"z�-��5�qغ��exW��iJSi�oY�E�xO�cͅ����R6v>3�C$ R�;dN��+\����K6\�XT�/�?Np��an���B�]x���5Z����m>�|���@�h�+�]����-V��e?�����4[��4��S���d��C���c�~�5�{��)�q���P���V~�H�]Eٔ%O��y����{������/T{T���@;#��6�2+���L�έ��˸&U�y�? q��/|$/7�w�&����V��X�&��`ʤE��U��4y��R-G�1�]����I��3,ݭ��'�3W7/e��e��N�S��]�[��b4��,��O&�|��N��h��K�WV��1� �gȌ��Rߨ��Mnd�O!U2GH8�݌Xb*^(��q_���r.�>iS�$Z��I,񒎱m��S�)��M\-]7�-�3�ϔ�t���*�u	_\�����}P�R�:�5T �����G��P�ڛ*�]q,�܆7L�+�����0��Ȓ�4jFBsW�[��`�p�jÚN2NfN܌��BT%C�Cѝ\hc|����sr�'�zz��K�� ^:����5AZ���[�cV��;��Î��:e�b���T���<=v�ˮ�688�w!p���LO�̙����G��7q2�>��(c �Q��_�"I�F�Y�a�(\�黣طfw��W$m<x��O�In�I����:4��c��f^��[6t^��QT а�p:����\�^����
�0��<�!�'9�ט9[��K�}�g��Z�@\�����G�(l�q㬽����]V��O��!_Ή���U��xx���C�������#�.�7�1B,�P`��Z�����{��c!�͜��3'ڻ����FS�{2���<�M���j�����`�D�u��b( 1��*��@9�w��t�ot���Q�~ww����$��ߔE�x���s_4V�aq�d7���jd8��ݪh���+�C��G&s�Pf�Q5gثO:��Ƴd,�ye�~��G��?7�`�蜆K��9<Zg���%)i���;H��	�m����O�J�K�s�lΦ-�Z��'tİ�N�X���t���3�eg�X��B��k���Ͱ��:ZD)Q�y�������W�/��� ��O"�c�	�c�H�G��!*�B�� ���O9j��s��D�DZk��L�`>�&O�*h�����%���$�(�։�-��<�ܶ8wS�!C�Yt��ޜMz��E8Kv֐CZ-{.?d���4���oxϕ�_��X�\!����s���'bI��<];�.,*����M�j��P�����0\T(W�ʼ������*���� ���<�=X��Bn��O��p;��)p1{ݴ�øЙq�ˤ���p���:ǷIf�M�1(f�f��p3ޱ�EĮ%�V V
5d[����WL\랸�3S�p@���@2)�@��:�E�����"&���d� �".v
C��H��>j~fU���Z�6�Υx����d��"VJ�4���T�V�{�,�~u�Z��I�k�{�����O���!s��u��C6�t������.Hl��"��z��^n�����ŭx�d_F�ݜz���4�^D0�la�&'�;ܻ��d��a²���=�¨�C7�-솏J#	�qhec,�')�G�\��xXARpF�ߎ�
�/2l���1*m�Ţ��pw#��]��3w��3�q��z�}����=&T_d�Fk�5�2���t�A>ج-1$m���Y}�����J_۩4O%@̤���������E��8�@� � �yV��
�`Y#�⥢f���,�$� ��-.�����vv?�.��XwA�����(�O�T]�8vpݥ������q�&�\",��J9�+�Eⅆ��8@�?�[�Vv�o��i�.�B(�;Z|T����9%*Ȉ�P)0��S�6n��Z]QN$�J~����AX^���iq7}f\3�tt��˽�*�� 0�8V�]���M��y%-�d]�g[~���g~͵rNi��'i��b}�rh*[�0�*=����#��e�zj��2�h/ߔs�4���&r��24��i�m���+���%|+}����7^=��&UJ�ބ�yWy~�C���+trϳ�?{�1y�n���B�je�r�Όf �=�D��������������(���pI/������e�R|��SN#a�� �\He�LYj]�t3�0*nnp-�X��m#R��-*��x;}B�S+~���T#�"���ٰ٩.ų�/�ݙD�<E*�b(O�w�	�m=�}�Td�p�8tK�m�"8�o���.�ER㪄|o�~�$���ɜ��2������n��^��N����Ѝ�t��f�/���Z���b2"X�юA��,	^t��:4&���d@_����G�"䚲��݂�������^�|M���?���"��S۷�j����g��������z����m'����{FL�g�/�~-�|�� %J���P�晼7��t�iz^�Y_�ې�v����xj�+���((��(F�;N��g�x�r�:c���=���抽���sh'��~*�ɳ|�|OJ�!~`�`U�U����l�+��y"]���nЁ� �����0�ß��E�a��n��q���y�`�s��i��UҤ1�̑��3s�I��M#�s�kk�������Gs����ba���<?���b�B��)i�K��'�/�^6z{:9�ygZz�@��@�D� ������P��
b��иh��y���l��#.d��
?�V����C�?����E/�޵��+?�g#����B_%J%UeL����?��%��,WA�AsyH��*a<i��u��#����9w�$af8�@V)�L���%�M5]�RX�����qq�c6�W��g�T��QЛE�4���U��5�4�\�{�PK��`~�se���4�zR��F�x��de9�!�CSӆ�ؿ�r� jŽa^�4��L@�M�.մ �H72��0�L�t�O� 9'͕��e�<��Ţ�U
OP&��L��������+b�\��ԓ��5�ʯ�<}iKטΠ�
Z��ECo��y�^�2�hY���ӄ�/"�>x���4@��hΌ�\y������ud���1�8m1uJ�<#Ȭ*�I�NC���Swp��mtbiS�Q�:��,#�<�,��7�E?�ҋu!^���/J_z��.�dȭ��I�F���H�j=pچ������V�1G��JY��&ə���6Xn�b�&�dL�������G�rH��}G��1��8�f��:T���F�	�J�thNZ�A�eI3�%ڼK�y_�xZ2ٔ�]�I���b�$@���<�T-5��#�
��൶eW^R�r��s.��_�a)?Ky��0K"L�JǼ�*��
@�
�ִj�s0��D2����á�-,A�@s���]�S�ZU�=�O��LZ�������K(�,<��\�g�K/�k���e�~;�y����昸i�'����?�̝a�#ă-��ɸ����y/W�)�����k*����.�Y���� K/� Ҹ*d��;�-���P���{�����Ɛ����99_�����p�bw�R~�o ����#W�Q�\���L?1��"l(��U�&+[[�n�� ��5�f�p�aL�g�
-��䨙X��W�T��� �1�6��W�B����	/��5�' �b{��aă�� �3��"��^���y�=y�cR�����Oڟ-���on��!o� ��ʷ�6d�<�o� �?�a)����n�NZ�UN~�y��P�K��r�kG��i�K���5
7�1���A�q�z�ՖQ>@�PJ��ﮬ�I���*�0��H�:`��*a*�I����*��&�J�ݥu�NA��`���P��������'������	�O��80f�'��yX�ώ��|��1�/�ۘ�(RQ�|r��d�>�l��4:.�UK�����(@�:�օ+��p� ntJ�si��ᑴ?�Y�3~S��=�*� /V�@w<;	y���ȥL����:�����=�1�+�F�z�1Z�|+�W����2�KC�內tpb�e�]i)ϵzyڂSJ�T)�r�	���g�	�x��j�������U��!��u!��U����d<[@愩��͜RGQ����cat{�=��r;�OׄD�Z%� ����P����&���rYs�/� *L��i��;���M
�:�5�3���R��������X�,��o�ïfT5^� $�R�ˆ'<�����55����C���MK�����^F�2O��Ȼ{��?������'�1����P�F�ppO�G搝dH{��\�[�g��fz*�Q�:dY�!���A˃�~�L܉�Y�g��B"� /��0�(�5��3~�$-ٟ��^�<�}��W��~%嗞�ow�J��r�=�����ٳ0��쐏�pr���6v+#a��Z�S�_֣�/�M_
�Rj2��k�YZ�k�V@9�Ɖ��^f&G�9��b~Eo=�r�Jb�o|xX�W8�?34dZ�����S��������^Uh��҈�S�眰�b��K�(΍��)�h��_���O�|G��dʡ�ț�Z����'�G��(��!/�7[a8W�Mt$�rou��$@�~�ޯ�w�&�TEX�6���Z�2>����L���
��L���'>�P��&�p���Xn,�B&�/�2����Cna]*� Ro)����m��9EA�ky �.)WKA�H�����l��z�A$�d}�ғ���d (�U�S�8�����"{��;�p��!e��M�C����GW-����o��re�<0{�4��#v��*�.��w���a����7�$~�r������Z�\i���a�R��c��.�*�u���8�TYk�N�+]t�ca�<�۠D0�F�`�W���`<o_�7v|���%b(��C!ʷt�/^f�AWGopV�[D9Ԍ�rN;ky�}���:\(@ g�sh)ϖ)}&���/ݬ?�I��O[�3T�1����x���������	����?��_GK�iY�@�Jyj�E�΢$�!��j���7VN��v]��=4'�}����<3�Š$�r+�����[�𰹢�#-��w�i��!�ᮨK7�c� ,>w��*f
�*_��f1P)[�}|N�g퍖g+��*��.�� M3��+�Q��Kًd�k��/`i���b
C��2%��fF�z<'!M�,~'Tp�ך��F����C�- �s5�J�8�p��u�R^��а*}9P�e��_�}��s����1��DƨX%B^	M�)d|�.x&2�44�����Z9���u��?W&�\���s�֨���8�|�*/�+��D��a�7���S�V��K4��à�]X�^E�4�=�×N1ݹ	ce�g���!�n"��|�=��׶�[(P�UEp�ȭ[��`��.����xL �Y��TW朳ב�r5���^W_@8��+��+�e+���~4#���4X��S�s�nG��Ҫ'Xyl�p>=�(��X&;�Tx�B���0NGk��� �����x#|���[,S�U�:���:e��>�"M+�5L��:��Շ�,��E��HC��-e
��w�yB������׭[�`��<�烴��o���^w���¨|-�$C'e`����;۫��b52��R��Jyѵ��C���
��Z֌UF����yʏ�ՠ�ʪ��S6-�Q*�B<�rt�
�C˦UP#��N{�V����u��-�����P�5����H�i05T	}�*�%����d\KO 
�8�jG[�Ͻ�\�i�x[��*y�*����W����i�H� ) ���u�J�$��?m��i���{��_t��ex)���=�eGuV֘�QC>��h�	�֭��0q�e&����$#���~w�-�Z~ܝqz ��?; ��NXN�tp�9r��˷�5��!��ڃe�5�ж��Wy2;)g��P�Yը��6�o�tr*�r��'��&�E/�� ���$q�	�ϼ�Y�%��e􁇜z����!~P~�JlG�N��8^��L�r뭱KR����J�JD@���jN�Q��<� b�TH�>���$�]������cD��]���S����஄S{���f�0\琝qc�l�ާ��Dm��Y�{����8���_L�T�`h��Ĺ�{0���ߌ��毣�ovYb���9	��F�zC#{�F��a+�xz�bO�H���;O�g#FW͹��cV=>z
�.6o�MӠJ�VʇpI[��2KaӞzT8���״_w�ϭ�������S��<�@u���;D5�5���t%���>����[/w�vʇ�>a�x��"W�1:�_��<o_S�G���;�'4�����s�{Qd���~J�k˜�ʃ򛛲Z/RW �7|�p�Yn�{rr�������<�[7��T�����=��@bJ�8(b0��������W���,0Q�9D�p�,��E´I8�"��^�B)�/�ym0�peu�e�X�T �1�Բf����-��peȞ<�h[��vCk�<Z���o�Q�M���e	N]�|ѝ�߽��8�f��އOw��D �q�s���ȫJ�C�Z}7-�Ix$����h���ƅ��f�|�u�Q�f�e�"+=�<� x��E�o:���H���(���CfYaIPӲ!S�1��>Hj�,[��[Qāc'�9�<�R��3.�*o�\5�MZ��v�mhL�4(W�)�\H`��f�0��I>�������;�&tҒfC�B��<*����[�^�涽WyI����+g�z^<�V/ e1��� Y��tB�*�����KKS���u����*6\�r����\#�EG�`����/a�Z^rE���x�痮r�+� 
���We�l���
��-��tu�*�����#� ����iW=Ί���e�.ۚ�z�Kҿ�����w�}��1+�Rn}Ρ�1؄-�A�V__/�Lߴ��R�*b&�X���P���%��~��7�L\i���E�oX5t���V���H �%7=�`f���lo�N���9��h2̙Һ�T �3?�
�reM��t�N��
a@8�Z�
��r�d�)�4V~h�i ·B_��޼g�g���) �l��W#\����5�3����=��=|( z��sK�����_��k��X���"ܵ\c)�/���%`�O���y'-r�I�� �5�\+���[\<�|�F�`
w�'SP`�>��'~P��D�
oӨ�;�-_�2@���Wҙvh�{+d�D
t�V~��ɛ-�����C�|2%�}�(�����e�p�>��DY��<�u�ZpHH� 5��$P�o��8 �B_��ݙ�h���yD�g������Ջ������-�~ @�Z�`�+_b���4����!�G�����f�Q�J���&��!�X��G;�=�{dӋ��~�E�F�$6��)T'1%���R���bA+87��zFn�+�� Y(�݉�o��M�.�x�L=+�H�Y�P6�'*�7ZK��7h�����%񈳥�s�~�[?�9�i�J�D*��}Z|��(�x&����^�A�{sO�F&m飌�ܣ+y�4	�ÒZس�'���V*M�Q�]����O�q�kE$����".:���2�,v�t�:
�7yˎ���ʏ�9뢸Ha߮������Hbõ�/����7i�F�ʶ6�Xf�L�[^T�t�Q�JWAt8�tEDk���i��M��)']VK;�*����!�탑��*^�� \�Ϳu�.˧�ށp¿4�#��#�[f��:�� q��v������������2�"[*&���6tK��#�����y�����Z��;�[g?�)G˼h[BF!B����e�I��tQe�m�"EX����8�=��ܿ�t��W(�l��H=EN~���
p�̓�Y=�=H����7�p��'\ɱ�@>�l�7��#I��}����|�o��7q�]�Ɲx>e)[{ㄽ|3���4�+�j�R��p�q<�y�$����S��H���n����f~�}��4���(U�U�8*Q��ef�o��WF	!�
��B�ޕ1ϭ�Z���U�@�%��E���(\V:�Q���$Z�C�nR�{�|���o2���}p2�V��y�U`X*0�����lU�M�c�����LE�)(a~�u�*�k�u��f�zK+��z��n�@�(�	�$�@���D��/��_��-
� �K9�Kݽ�}JvX�i�K6|�R�TB0�Ok����)�M��%*a�Vޫ�É�M#3�,��M���]ivJU�+O7V�G�� �3:l��R��U8*^�����/^�^ms,��F�&��:W!+�H5[�a�ې�D�=崢]�8���dç]I��|O/�g�.�C��w�=�z�"̻֯�T>��@�'}�{�
�4����!C�ۻ�Ի;�l�X�ĝޤ�f�n��bp��r?��$N�bL��1,~ֳS���S���)CU�J��x�i�|�}��x�I�-R������L��f*��I�6�LK�
��.'4�o����������vYᵆR:�����`���>�V~�E�ݻ�A��Rhd��"�1vr=��uz�+l]����ÃR>\)��lˇ�������)��K��t�13�t�}v`�E��?��-����9>=��3B��	�+y`�"S����5�m:����e/;)+�i�u^�J������ MƮV[r�~�����a~�gʔt�@:����c7��i��]����z-��e|��2�Ľ|����~���{���hm�t4<ncڳ5F�ֱ�#�.����{�t��|:��8F�}��V�,� N�d$�PA4�P{��OǇ?�/m|���i/;�4c��%J�1� ��~�z�/���ѯ��<��W٦��Q޴��Qހ��N�����-0C��]�f��0�x�N��r!<�Jgl���ER�U�p'�!����g�����C?�e�3��������dqW���EӰ��e���n�JŰ�LJ�a��*���8�����;.>���|���%&�~Sy*2L��͐�.f5�+��Wq���x�p��Q�HLah�P����n҇X"��`ٯ��+Dy��sh&�1�"�jP�"u�d�g+\c��/��|�5)ZѫR�a������y�� �}-1&�0w�$U�ϟ+�d��.s��i�IZ�`�?�� �
�"��_0:�z�c�q|�pSi�ԋ�H7�'�;���ʐ[CA�e��(�h�T��u��i���o�ij30�!=-`I[ɪ7N�E匣�������G�4�GX�\�c�9-�T��t�:��!(Z�E�.�E��E�(�}�h�,}v
@�%�(A�p(�j��g��k��]��s��e�0=ARP�JZ�O��G(�[�QA`ݴa#d3A;J�N=�8��m]��Q�ꢑ�i�I t4}�����(�O�
#n����$Jkӱ~�&�*_s"��L��6r58� &h^K�>�o�8�]|��E���� N<%�y
�}��������ha�8�62g9sF��&Y��N��~�iΔ\el�&T�0�tT�r@���Qv��$ ���#�>c��&�Ĺ��V�ݝ��ﻗ��u���l��>r�	�v&��������1������(U���O��b�6����O�Wa�U��mvv��\��P�zE��CG~�Z0����/�������	���q�i�]��� ��.����FM��A� �X�p\@F��x��E ���Rגps����L���~��n��?�=�Nڄ��X����-߶�^��x�[*R��x\bN�ְ��)��k����t"�/"�dU�^
̴*'�:qM$W��rh2!s�(��8�-�`�k�� �V�#�8���i�Je�ۗ��6�[8�U���E�pN���'u�̅������s2�X���7Q&O�����;O��L�C9�pL�澒W%/Eu�8y7n� O]��Y��y�Ŗ�m�4�~���#��0�E�;�*J�CvНeB���
u�LO^)����04 �P�%I3�
�3Fd���m���B�D
5�,	o�:�[����A�L(N��.�Y�أ��=<�x6�gM��_������wX��!�34��s��3��ظ*tm���ڠ�0����M;?<��R^1Y��8)��!��L8��	����-�W�2Qv�69�Axa�zJ���%�$�|%�/����c1�c���N0�S����^�;��:�����k1���bp�n���a�z��Ui,�2�~-��;A�g#��m �47�>�2Vc�<q��
����2t���@ ���5�ʞg���P���?�tF���^��T���f^���� z��
���zXs�D���sb��t��� ̓�pI�򺊟�Ϫ�.i��s���!̣��X9��[vT�2�Z|f��1U�F�ɠf7��~u�x6+X&��|���M`��^�������Aw2�g����c�#	lx�(pt�N�S�5�"y����t͓�˕Ӭ�c.��̏Sv+�G)��C�	  @ IDAT<�������g,�+9K���6[�`u-K�ꡂ�:������eY��)��w��Ho��;K�����׿������㇡�~���/_����y���S�����P��$����Zg������a~~e����S�U��VZ�r�X>}�p���<�2�S�(����bE9��<Gvy����c��Ő8��i8�B��Iq��!��N1��s�|\�7��Z8�bꈕG�H#hӋ1|R%����#��>�K;��	���՝7�~u&�[�H�.N�
��	;	:��o~Lc���wW���R�&���+��l?拓�~�s�]�{Ϻu��&�	��.9��T��=��
1�C�o�֢Z��bf[L��>���rչ@'-�c��2v�z�J�|��h����k��&g�>x����ӧO�I���<2$r����D��*��O��2�������xW���:��lKQ�$D����U��P�U�+� �������K.�s>���r������a���(�A�瘫�Ɨ�����gG݈ w�;�^�h�]LOE����P*\���",:f��f1�=��W��%���\܆Qrs~�vA;�z΁�6>��Y����^2��}&E{��V�*�J�L�j1�
l�P�2�t���9������~�w�Ӛ�#0A^"��o�T�X��.&�+`T�[�0G�#���P�O�\t��V�{K� R�Zt
|��&�C�X�����<C�a�u���帹��9�ö�.�y�3�'?&_>&�\��4�ho)�.�����.���gh_���3��9�������L5�|�"��Ĵ_Ӑg7s�
��S�/����%��\a�Cr��%"-��3��T]L=��J��=���eM�!H���!{�kz\Ē�^�iCZ!�"XȜy�p����y�a��!���)@s��������jA�G��)oX��Z�Lg)��c�o�E^��|C�L�����\X���V�4�
�P�|����M:؛UIU�WKUmX!+U�>��3�5�K�È���c�(��{ד�US�g���Iў�1C��54����>�=~�š�OG�<�x�2W!�j����QW_:�̣h\��C�*��T�:�"�vcsHY?�
_qvύ���hk��j�{��'�,�NЀ����1��G�����#�|��F���
Rk],�22�h���B��֗�2�J˧u����I�B���
���(�em�C݀.�U����t8�ő�=T}���~�s:��͆��R� ������l����aS���`G©�u�Bfh���n�̴�[����>Ci]�I�3�����"b</�R,�ks�#g�矋���0��������Q:"�Y���<��E�3����	���c����l-��HW�LS<�¿aa!�y3O|��P~Z�)�.j�A���]�o��P�m�ܲ��P�*c�lرA��)zQ��PR��\�Wwi.;!c�r��N߼;\�݌�i�n�d�I���n� DL�c�M\�:��)'�t�a;��d�ૂT�z4]`QT|�������Z�4��Qp��wW~5zE��-���cX�0b�ӎ hV0� ]�w��ez	�Q>�A�8w�'��8���*/���.G�[ˌ���XT²�u�$�D`H-�&J�K�dP��\&1�=��o~��U�A��
��!����(���9�P�6�*�68*�N�?b�d����\��ByN����>�"�,�W����U!�B����r�ڡ"�u�w+M6�L��
��,CL(�(#)�.��U|��b��4U��J/�FNk���$�9�]���!u�	�k�z��5zӃMHUM����y�k�X�i��?�ՎcGX⭻yrBwP�>i>y�9LZis��u!ʗ�%x�-�l�TL��){�9g�f>�1@��@Zu��	Ap�LI���.]�A�w�Q0+��:��uV8|3��W��t'�U`W�L�������+�l��"H?Y�6��!;�T���y��RVq_R^��5WM�~�:��\�*aUlVQ����0��)'=��8��;�g���ڦe�'� LG�_�:�(ǽŨ8:�F�'(Æ�--�t�鈪�9wm��~zư$Ï�?�����9=f;�S�� �}�9:`J�×����x�]�1����*�'^�NɄy��F̹9ީG�\�	+M�e���tN�e��E�,8��K��*8�q�Ԧ�����w	�>��[h���g2�`^�6�y�%��)��{*�j��rV�^�;
c�G9wX\�b\��2)�Y�-��w������D_|�#��1�'�����Nt���[����!�""�J����%�F����O����𼷰�Y)<�3)fQo�&���l�bE�vb���Q�)��$�b%�Ғ#}�%iTu׊W#��]���=yDE̅���N7���<�u�k �8Y}e�m�m*�Ѳ�@A
�R�Q��J��_��S"2
�X�@*DIHIP�NL2'5F/W#��DmU�)�����I���3�)B�	�ni��s�s��[�VP��&��kCaf�8f��"fMh����Ƃ��$#b�`1_�7~�q�8�H��zƥ����KD��Yr%n�&��G���{O&i�ܭ8=�����������j�EZ%p$.���U��-��d�Fd7�u勓�ܰ�}�ΨO\����i�%��w]z�
�z�!S�kY�/gy����x1�NX'���w[
����b��bv�<�xše��I?���n��UP
���Q.�4i�ŭ��W��w�l�^�[8�y��������9'�%��6.�^�Q^�*ssۄ�J���̈́yE�VmJp�N��z�?�V���d#H0��l��wd�q�zQ��� ,�#����3m�r����0Oϗ�0���EFp[�آ�9f~+=Y'���'����/�l]�8G�#/�A�$hZ�Wq��3}�c��/�Z��%�I�**X�Q���'�;\��Gly��K��YU��h k�S�N��}�E���r�7�Qْ��S��9:5O�xX��f�{df�k��|�����cM��Փ�ig�0r�_���F�O��nZ��%�KgY1���t
��	;�ge7��E�1Ws�]!O�𥝓K���@3�Gd|.�-8���N�f���\:�rNY�{:Q��&�g�x`���i��ƏVN�2��KK�<'�*�?\bJ�lX�#F��8�����9\�]���M�'xqjmr�-�e*|%���L��z5\�M��"eĔ�8܆S(�X�o3��Fe���ֈ�LӸ�
�4p���o2��z3�[4��G���㌕��U�I۲�U�⛄h��U��������/M>�˦������w8W؝*lv�K��GV���~�)���c�Wo��y����{3bx򌥓h�N ��I���$*��^T*�ĶBH����LU�"D���k	`�̔�2F�N̒�������s�q�p7���,�jP��� &/�wނ�4��3!~�M2M�U �����"c�2�%��V���gኈĝ<��A&�P(���c!渭^��n�^L���-]�)*�1��(�����C�7���}0R2�Ҟ>l�!Q.�MhT���a���O.r�['p���Q�Ί{e
(��A�d�P��˔�VU�$*E���:��*]z7�F�Z�j�2fe ��Zuo�z@c���[�����������6?�����ZD�>Û,f��v9���p똂H��#)f�vl�.����/m�>u���OG_|�	<:7z���4�@>�<y4z�Dl�����!��X�qϱ�����������ҥ5:����Y][!I�C6v���=��I��4OZLdmu%�ZJ9QH�\p� W�!r�Z�K����c	 q��
���}�݂�-G�;�+��Z(q(�x����E��'��'t˺�_��
GH	�,�¤e�2�~Z��]^�K��
֟+�]f^ز�C�SxI�Hl{�5qbvx~�6�R9N�>�F S��;�X\��D@��g+���4c8���[\P�'𖊯��i������L=Fa�����&�)w�����[��G�Oe?(�龅Z����9_o^�ʞfN�  [C�8fu��I�"O=�_�hص �|iͮ����*�6Ş����u�Q!�-�l���	-X����ॷ�_-{�c�q�r��X��'���-Z��G=�k�Ja���kczz	���r�uU�[N����zgR5��o�ߍfI#xZ����tΰl�?���"��3'X2)����h��p�Y '��htK�M�_��>P��/�R��#l�����k��"w�2'B,��d̼�uŜs״t*O��<��^����U��"Pf�o����/�+D�tSo��(�'WDL6>�T#��D��H�Um�w�=�{_�E�'y�D���N0Sy��R�������h���G8���DY�4�Z,B�0�b����oÕ��X]�&�O\>JP���-&MAH0~�bg{�V
�8A˼�0-xfT��M#�۹Fj�N�u��#c�t�N�g�3�i��lq*0o�
?�vf�9c�V8��?h��R�����W3��`]K|C2�ҀO��{�k���3�ӻB;W�Ѿ�����p<~�3��E5XZ�N>��)+e�6D\�Q��ZrK�Syi��f�n��{ϭϡL�Y���
!��Ve�	�0�����W���m��;�'�]�fc�p��2GIq����=��L^����ȡT��{��}ˤR����mh�]�<�)a;�a�Z����+����ѯ�l��y>
�Y��8���W��3lysΩ
�b}�:Z�w��0[G�y����C�aK88��ˈ*����8��I����0uΞ�8Rn��{���\���CfdH��^���B�`�u��X�ģs��R��AE��^�� !��I��N��R�G��=�?r����#�����]����(8/qqޕ��T��S˖�"
�|���S	�Z���9��}�a�����
U�$qRΙS5{��Q�+G�c8ǻ�=6�̈���UA��rK�v��&�./9+
���~S �`�)��O�X"��t�z��e�P�MCK��{;ƒ�<��G�̑T��#m:���Q1ss�O?I�Y�'�1�c�(y�Cؤi���U���݋�n9��uGG�-� �
o D8hW��A�X���Y�zm��0�t�NZ��g0 n�۳#X�+Ͽ���,���@Z�$%?���;N�?��Iٺ��JEY����iJl��O����bM�itkI��|,?+cfi�ń�΃�-��.�pջܑ�@X4a�/��ʁi���UgJ�6BL�*��aZ9L�.�|x'p�o7iIG��g�z�ş�P �#;�s��Ӵ�#W�38��B��"��H��Jd*G�����y�U���bf�Ƈ�
N�	���{V*���"�|rWa��W��8IB\C��B)3�DJp������ѿ�Ht�֍RH�(�vo̼� dF����U�ăg�;��h�C�Ŭ�"�$��o$�^���&����t��@
`��P�U�!��#�!�P��+o�]R1A���7�ׯΨ����|S){�$SUv�������_�PvZ�WP�4��⌛���ZA����$�'`C���Q&���*A��8-<V-WǬ1��&￧�X�=7�ɜ�0b���kVm^��1���'���3V�=���ѧ�}�5�X�s��Wf�;�t�d�$�����������F����6��o�隓!�x����P�z��R����Ŝ��T� ~6Yt��c���mg��`Jr�-6t�5��5A�m<��pX�Fv�g�l�e%{LQ��sz��s�B�1V���|��P�|f���4�|G� �+����/ӻ���Ď��=V<{�I���9���;K=�U8Z��@�4-/� 8oK��p�T�d��"hI :2 ��#h<"<�òt�]�'hC�Ρ�9KIS�+ݲ�=C�*MIj!�V�:L����_1�=-l(�����U�G��0BN�p���š��RI��R�w����y�|ߺXr@��t'�K�����_�\�	Ƀy�r'�dI����u"�ə�Wu�q�ۭY��]`���";5�K�\	�a��R��7%,o���Gv�W�P���/�����=��C`���4���k@��0��O������4��
��3��
M�I��v>���ڎt�����8�l<*��r�I��T���Quj�2w�(��	���|���%��"Y�h�/4�Po#��ٕ�/D��w��m;�m�>���]��M���5n��I�l߾�/
o<g�����2#[X)������;�}��"q�5�TÏJ��/�CtTAaR&�����R�";��~!׸Y)�P|��-�~�)Z��n�s���հ"��⭗�����h���U���;� d�J��T�6�9_/�-Z�0��-��p�E�/�N�`��k̗�Gu�ZB6T�]Dy~s�hx�0]|+D���2ż5�~u*�ݭ��F�ig��7][��^�-x�7zt��� ����s�n�͵He~���!�1�/��`�n�����n��|	���/q���,?���h����I������y�-{�����A�Z2<��YW��N�]%���Z��8����g[~�!�1���_}��m�_�b�ڛI�d�ek\�(�Q�Q]u��!C�Ϟ2��$B��Is����p���`�s{-D������C��|g�I�=Jߪ��0��)/��$O��S�ɡ2O��8F4�FS��J�d�r�ޫ�K^5ꭸ�@W}��tKX�q w	n�u�$;T�Maw3�q�A�(�6m0�
�[�d��fcN�_� �,��,1<�B6X�Lw�"N�Y˷
��[���z��K�2��V^p�?7��X��-,4�$�ȇ��In���k�=�J~ĊE���W�:Qe���F7�-����G��Cn;}�Un]9)^�8$�t(�}����`�y/-3�B���7.�0۰�	*z*c�_7��T���q�v���c
r�̑j�z�����uZk���l���EVNn��J_����A����"L�Cw�)��/�U����k���쎼w珁ji�N�T���$����ݹ�����;�^�!
��L���׊å8/%���C�a7z��^��#/;]=/>�*���W�(S
�uY��M��!l�'%gy7q_���&��~ϋ1�{��x�I�z4�ɏ�n��e8�M��7�3s�PҲ�
�=�)��,s�ފu���/�����3��NQ@���I��r��;���%������z�x��2���E�dG���څ<O+@�_B�mn�k�F��FA1�������a�#B�q�+8�V.2�2�9f�qn�%���*��L�ЄY,`�[�U:�U~��&<|m���6�^6䮂HO=.��|����ܥI��q���}۷3����u7���ۡ���r1��z9�r�G�'��VPT���K�TB�(4`s���>�����/�oJZ˨?�5��6av�lfP�M׆v�)�br���U�S��w���7V3���+L�ײ�0l�����8����x�Q'C>��Rxi�1}���ĺ�𫍺Ã�Pm\�H��
�G6	�ߘZx��"s� α)�C���a� ��PVǔD�
������<Je��蜠K�;�����A��Xj�p������(��vn,����3N��ED�Y%@7U�`��t��j��N��x�(:�&�������@�UiގJX6vl�[��U��_�f��{&�GX�R�L��J��-��76S�(s���"O�s�crw��{ǔ�1Ri�#
�
�d���3���<TȴD�ܤq�"�Ȫjy����y�e�ZΞ>y:z�VXOc���T��E۽��r���QkH�9:��n�c��R�JYY����^d�]T�6�s,�.n�����cxm�|�G1�ꫂw��z-9��n0vV�k��sq���+s��rʅ�v�J�u8����ȑK�a8Q��(��r.��^���`�����4K���ds�m�/\����3�����v��W�;q���S�ihtߕ2�ν-��I�R��<��"C����{p�]�zZϝ#���ey;�?�Yv��2��bqQ�[X�9{����Goa-I�F�%nB�L�*K�{^�/�
W���_*_��l攑G�e��4�?	�hɴ ��B%��3
7�ޢv<����ė��7���!��DV��
f9�u���_����˹��b!r~�)����� l�D��On���F�5�J.��lȖ)_�Ջ'�+��3��:�j�f��C[�*{@�FH�[i%�+/~�h��a��V3�v�w��B� �j�N��.�z��MО	=�7C�O/���#������}Ѥ��XC����~���B�~��[\}����S�Flh/�vƤ������4��.���w��ET�h�G���ִ��B#d��ңEC{���#��.�_3�����WvZ���q�&WUڨfxJؤ眘U`��։�b�`��o���Ӌ2}"��X����E��J��uIEjJ 1���Ma(�)��݉����2U�֕ޱiÅ���'��\ƪ� ��e��]�[ښ��U�qr�CoZ;l��E��Js�&�U��R���������Ai3v�*ʸ᭵�+9�?*3o92j�{��v��r�L��z)r΢x�S�$	�4�0��<���l�������B��7��\�@�x��w���ٞ�y�|��LR9���M�������J��"J�
�:s厗L~�$x{��D椩 ڸ�n�"���ʣ�BEʺw��=-���JV{����!V{���8����ڲ�E�W���������a�W��JeW\ݪ#��1<%��2�"�>�\���#n�3/B�������O{X�qǃ0���O���!�ƭ��G���[x׽��§����*�=!��qO�r�x�U>큄P�m@�W�Mz+�����Bw�9�Hݸ
W��Λ8Z7oڐ�r,�#q�%�QnK'��*+�KuU�i���pMֿ��x����?��Q�_���8�^��Ɉ	U9M�J��Q߁��@@e����M]�J�\��E�`�Sc6�:�fn����O�W���/Qb\-(�/9ت{J�����{Ĝ����i�p�)�Z�z�;a$Se�0E4�A�r�g�Tx���	�@�b���k�ڙ4��)<b�9<W݌�*��)�n�x����2&�A�a
�����N~� ����d��7n5���{�	�{+0�
�tϜ��c�?��!����꠻9V���C���i5�5�Tx����ع50���z�]b��Z�����d���	E�F�%�d�0��v�EũJ��}>��������6�n��q0�T4+���+�P�2g>���!� \��Fy�P3_%����!e��bxR˖�}�{�/�0Fc8�����=���նK�����]^ƛK�+���k�l����E,~6�*K~;�f��� F���FE�׏��Q��9�1mw�I�X���uRZi�����:�n�"Lc�E+Op8K�`���b�q3$ʇ)�c�o��֯mҫn��.��n�r����r�������f9�p�H	\+�����y{_}�U�qX�����Όx@��\<�G�]�,��&��Z���g���!V�2,���ZOQ�aY;��c,R�"-X���ꐡJ�C���uL���ZF͏��rq�ۡU���d�<.�>4]h�W�L)����)�>�O%���C,bnY�Lw1���(�P�<`^��"im�?]<�̆x�0g�vã����m0T�s�xd�e�|��G�\ }�1�)�<eA^��´~pM�Sw����[~�&������\?3��)�~��G��j���8O�=�׍,��,N()��0	X�0�Ϡ��Ʒ��o<�OK�s����x�g��f�#�ұ���0�2:2U���:�s�%�P:	*c��i\�PB�}��(JU���(�(�Z8�=��4>??n�HBʜ��z�¥���u5�)�s%���w�[�̀��X�T���fs��Œtɸ�%C��'��
�G4��!᜼*0� E�2F�U���Jh6��$[��q��a|�u��%ါ�ˀś�B�T^2_�X
5ܢ|�s��q�C@8A�PM��Y5*�1ްY�Lǌ��+2��������K�����:��>>.'�|?q�b/�e�ƿu�����ʵ`�����H׺�b��{���S��?<�^��y��wOa*(N<�]��R��R���c��;g��y�~c��ٴZU�����^���ߜ;cn/��?r�=����X��L)X��t[*��g1����|l��<�H�|F7�]��k��c�����z�d���� �*PX�b�w���0筩 F+��ʃyQ�9������q��Y��Uw{(]�ws��[�0�d�
�JzQ�+4�[( 漀���� \Co'�GY#X���D�!�g��-��^k�sM��_��}�6&-�Q6yz���������kaW	u�O�,�)7h�"~�vږ��� ?�RCJ�o�
��7����y����!AP��6F_|�eVQ����_��mV���������&�o�2�,���
X:�
z���)>%�e��.�5>|?�<Q��ێwyM�t�ʛ<��G�����wD\�#�*\�_�,ӱ�Qquޚ��8�G�`%nǈe�Z���C��i��[i��XC�6Ɲ�аk�d�e�,rIyI^Oߒ{qK�R��O|yN_ݭ=��ם�w�ƻ0�eq+H�(���Sߺ�t�=�[P?�)����Qh*���%��B�mh��X��7qr�(*`�<eG�z2\��em�O���T��o�_��YzC:�$����B�<ʰ)0e����Q�R��˻��T�I����D�#fӗ��mrKG����U9@Z���s�<�(��)yx#��}�����H������!�����f��?��y���њ���;Z��ū�p���
�~$￱�Y#� <��3�
�ʌ�[6���V		^VPw��Ԑ#���e"��/�!���M��A���k�ořh�� )$�5�?r��>�
��%7�kx�����?}��\MG�w+h�!�|n�ƹ���Cp���O�:D�JE��d/iŕrh�oU�u��������⶧}�*�����2���>�>�~q�er����@) dZ�W�\,.��W�T��T
 ���s�JH�6�<�e��0�%�۩�ĸ	��܇�4nZĚ�E��ə����m=8e����\�!-��X ��� K��1�FP�	�w���pс�����R�V�D&���z��˾h(;*����aGt��R	�r��ƣoQ��V��*�z�:;]�M��x���-
�>��@Y닖�(�H[砪�ZԖyd��m?�H��y�Ù��_�x9�
���+Kq�n�0���$��a�G�Xy� -<���&�V2�$5�(ʔ�V�t�:_Z��G�(��#�����
�
�_~�0��>xo̠0��0�8�T�ʒJ�2�-�X�D"�3��$D���S ;*/�>O�o�tu8TE�y�%�Re�vC*U�[~���?`���h� �;��a%頕0�i;d�6%9��=�C�`�?8����b���8����rX��k�bQd:��!yZ7ml�4XU�{}��D��<������ýWB�S�Mwrߍ�c��%�?��u9E��*����{�����=�I�n�������y�� ���y� ���H�����&,놊�7�`Qx�p�h.����I?��≿B�����P?�-
������L��t�t�I�l+C��F	ғ�8yU84u8�P�������Pf�_�ބ�����&�ZJRI����zf��y���>�����V���M")�~�@�M^Q*Uwό��̛�@  �@`[�B���C�T}�޸O�ENk dC%�4��jM����P[k�cX�TH֨k��7�([����`�Y�U��4�+(ꃘP�$N63��w��tX�-���"�D␫���L C T^D)��N$X��Vh`��#l��RL��-=�L�K� n�If.�ڣ��~��w1x�|��t-�No�i|��$�q����MJ����k��?礟���NKR|��6ïO8�ރfݽLsx��e�qhǣ�d�7Cz�	bѯ��7�Nx��U�K`�?6���訴�yiup�A�'����H-�m8h�_�p�V˲���m�{_�]�07	v���pV�Q&?�g�(����O�c�p�iq���n�z�~�D�ȹycA����6�7#~�!⏰�<��c�۹Hz�B�匴:J�Qnғ�>�WlӪ�ee�!y�e������?܂��([O�R��ÇXi��@Qʜ��աXP��G�^�0`\�B���G��P91>CR�,��d�L���e�Vh�q�8��+�~i�q��]����О��"�_������ИuQE�"�&�k̡�~�����G�vJ x�w�N��,�d�:�W��[�Kˮ�lr���cd�nv�=)Ak�:�;�/~'�{\�gCZ6/��@áa紒��il���D�s���g*��x�%o?ePe�C���?�40�E�lܿ����}1�^����E�r��ʺ
��.y#.�W�����{@��<�/e5�Z/���WƓ$\���4�겔��~Z���w8�	��.������ʿ݅\�(��n��Q!NÞLF�W�i��n�6�U�V��-�I������N�f�zaS�'��4�ַ��y©���L� c���H<��d�&o��=xB��Y����7V���<.Y�jZ @�js������-lp�Seh�-�� �?.^�ֳ�4?��д�� ".)�=_D�|Q	sZ��Nb��棢���i)B�Ըk+}-lS����J�L��y&�;��JzfT4���H��:
�-�4���4.�Œһ�O���|4��4�O�8��jC�R���pf��x�Z ͥ<� I�',T��K�|7T�9Ay����3h4X#I��hK�tx���R������2�%�"%��G���8���`���(N���aa��i>
�wi _��|�*�'p����(�@U���L��l��� � �A��E����Z'�8{q6�/j�B����Vmi���FNE�<����b�2�{�QX�X9r�;��C+��\̿���h�t�����_�e�7V�V7��e"�CC*~�����]"��y�Z�Fc���(jwƪ�UW�h���e��J�su\�����|8�����(_(#�+F���]z��{����������Z�����#k�UH�`��@�Ų፲�����0��!
��:��ۙd��M�C�. �aL8���e�1Q$�W�rHԸU��d�qF�^Z�����,e�8-	C�U:�g�$e�<�l�lo��>%�SB\� �O(P	��OQ����[(QQVwsF�{hş�졸܅ZJ���o�5�4��{w�w����/�0jQ$��I���%�V-X}��6_������8?͉�7aw�����/�ۆ�tA�)Q��̈́��
�~�tOZ)d�9Ԩ��9lX�\uk��`���y�p	��5�w�W΃Tv{���Ǭ¼��IVc]�ynLL��G�<4���o���S�n�-x������D��A��^ᛙ|���(��=�u��c��uft+�|�K�||����@��q$�Oma��n<R��Ye!�,���=�򵼚&� n�_,�K�7݅���*;U�*=�v,��2��ÐD	Ǻ�+5�N�t\�b�gT����qgVn�f��vg%�\6Hd����90,�9&�5掹9��Fk7j���^B*Aw�C,��ӈ/I��x.�!�)<t�������e����WD,i�Y>%�XZ�DW背XG$Gz}�Ϗ�*���'�1��,���yDI� \�h��t����䪸 �ѵ�w��
n+x볉9Ư)��^��1Ij��>�fI`�=�rU���������˥~qOE	*�!���H��0��l@]���ee�%���!�]�Y�m�z|��������������qC��@Ėg���
w������x��PE�>�;�H��]���]g;���,�p��6{���1�	6����l�n������Y�#NSoi���%\�A��02G%�9���~*)9
k�gɩ,(�T�乊��Jў��@�;�P-iZM<�С�7����i�6��Ul��H7��ѐ~H�ߔ���PN��=���Yҫ�ʉ��O��EY��N���Q����)��i�H�K{Y�k�CY��Ή��Se�H������6���nݺ�4h�{���S9d)O\�bYQ>�~-�Nܵbޙ��[>����X�\!j>	�,��`�T�a�zDZ�P�%�eS�t �+��B�-�H��Gn(|��6��-��ӑq(Z:Q(Q��n 4�0j�d�Ľ�Ol�J!uk�"��k��.H���<
��q��Ni�|�p����K�~?'GW�W��6���쯉�vx+���;��6�R$xJ�|�	����/}��,>i�T���`���S���ԣV#����Px��I��I��׋8*��}:��=u:�'aD����&Xx���d��)*���t���?n�ފ�'.�&Q��뭺�D{������jt?�0;��Z{�8�`�V��4#���E�)&���J�PL1���̏0���	d��(��Vڦ�T�DW�|欱��B5(O��N�Y���sq!$x�����?�&m�����І��T`�^�E�I�Y� ��o�G���^�&_����]4�p�a(�%�!�����3@sG��g�^���S�^�˼Q�P	P�p���cn��^{rm�J>ʼs���0���B9�F넸����?��0��ǹ4/�9��������5Y�1�dk��Xe^�a(���+�����qe�o�D�������[��^e2�CAY�}���٘�Zo�mT
�N*��l�L����k�{ŘсCG</^�j�`��>�t�	���**6��g�SQ�a(�ź��̂��!/�rh�\�h����9�빕���!	O>����R�͛�k��|	� �B�C�>��W��D��)�
I)��c�U´�E�D~9Q>�λ���/#9��r�����ý������a�W��¿������2h����ȅkl����A����-��%ʞ�\Vؓ����ĭC�
�N�Se���-�l�*Hy��eYq��Û>���٧�r�(a7�&�,]3���V��P;.�m2�h ز|`O}��ҵu�}�vXA��������#/��C��O�_����n3�G�֛�����^	8��p��~�i��7����w]	��T�	?�}5���^� �5��%6ߪ%�a��-�'LQ�O���7:�qt�<��JO���]�X�b����2�� z��zY.qUX��]��	��4���! �*�
~tz�-��
Gu�s�c��-�<�������9A�������鯛�a���(��h���ʙO	�5g����2οAe�ت"���@������z���p7WcУ���J��d���-�{�����:��d
z��+e�G�e8�
.1���W��,��`^I	� ��eP��H)rW<�?	p�������~�)=��"6>���k����3�3��
��$IK�Ǭ��⶟�R�� 6������6��a��4�P��s��<��7of��74</-��^��*⇖ z-5Mjٰ���9���Jm�b�C�1�ĩRᐟ�6}�
WR�Ӹk5r�����?*d7�ب����v���b "tb�:�h�Kο��yb�Җ,6�.m��C<�L��%ånș���8'Z���̕2}�ByUDeb6����J�O�d0�
N�94��k-8�O��2�UC�:~�)Y�/�|�'�G� p�k�.L�8�12y���Y�ě�L0��X��F�  @ IDAT�p�~:'L��ʀx��a��>e�C����l��ql΃sQ�s�]�qa��(�*�Z�\�aNO�8:�9e��r|iϮ�(<��e�T���I��3��������믿�*u-J�yh�P�����?�����t�j-�������Y>��/{�1�/'ؗB��1Z_P�?!Ml�A6tx�֝{�WvHp�Z�e�Xo�_���g~�k�=��+��Kl'B��I�)���^`�o>�[+�)�M��2�:��o]s��� �p��3@�B�W8��^K�|���`��)�鉯����SѢ;��B��\�����4�^᭏*�N��n|��AU�w�ѝ�޺ǕG���-Q pR$��Q�	R.#r���;��M�
�������@:�4��N 1����2WÏ�B'�{9]��\U�0Ь|S�s��o�`~�G�˩�|g��<鑃%g*��d�0l ��V9�ŕ�~ES<MV祙�W�Ya�X�.�2�\�P�z�S��NO�L;g�E ���KJ�]t����Ygn"6�Q0߁��%��i�B�#��p6v�n	��8����u�w��g���8�_g�?�R����e��lX>���N�`����u��Bm��Zb�F�ñ���6�
?w���ok��ȹ4L��6�&�U�f�T� ��а:��I�{Z P�ldP��@KT=s�"և(_4H6�$��ĖW.�0G��C*$�(��}���)P �<�G[��Q�Tشܹ������-~��"�����S���~O�K�!Á�X=�4���,����ů�{���gX��CT���c�Sx�Z�vݎ�D~���2��f�W���>gx�%s�ܴUE�kQ78D���9{�<wR�
��^K�a������w���Z��H-x�\���7�8�&�.p�SEˡ6-3*�Γ2�zB���V��R�Ѫ��'77H�a
v(V>��m�}/0��ϰN2'�2�6�s��Z�,'ZA]P�Z������&��Z�� �O��	��~����������/P�v���ǜ���%��8ܭ�s���������_����r�	7:gO넖2Onp����l��T���Z���]���ˬ{�����������?��Ń'ϣ|�cΰ
���.w$��L���|Ew�_[c51�We�֩/�2�%�wv@��M����(.�\}�����}�����3B�ZTe����"4����\?+#&Q ���/p�.e��i/E�8"������;ﶼ�q����<ʂ����z[��^#�U9�o\}�+q��{��,���FU$���?��H�x������
ݍF�b��B��+ɦڎ��K�Q����F��g���I����~����{�j~��4�TztY^�w������	7 ��m��$p!I� ��46.��^�P�����Q�w^�b�o��yq�E��La�XH��ӿb0�x�p���?���!;��o������/�׻���-���#Ԓ�UI?�)_��t>���HT0�Q��Q��Ň|I<z�G�f����D��ү.��2��㐏�'�Լ({m�q�l��|��k,�?`Ɂ�Q/�2	Z��J�b�),Y����zw��h�T�T�T�ܨ�vHwWq6(�|���똰/c��쓛l����L��}�F���o��%Ò�Cl14���O+8�$2���K�k�`�I���t�eycC�&���<���.2č��3��3W�V�ܼB#|��)]�)_�@��� 7_1Dec��\����NW�,~��obIy����Ⱖ8��x���<�Z��a8��?��b-����<7#�ƺ�^\n��*W�^c�O�H�6�1Qn(���'7� ����wc�R	T�VqR�<&N-x������4�U�TԜ|�b"���p��WV��_?���bW����fn�&G��×���@�HD0kY����6J.�dx�->�6�����YA�Rm��r������*�*��X-i/�!�^uk�o��k(sW��᧿�aU�kc�s����@��;�x���.z��O�Ҷ���ᖢ'���I����C��_�7��x��(%<����i�Î�����8�iy��y�˧�ے��K8+�����l~Tv+x:�z�|�	���оB􍷡F����<#�>$`��DV�D���L<�ҡ�Cs"�Z��,���Dk^�Y�ŋ��:ܒ����)��M�5\:��6m�'Y�xq�򦿰�4���'���YXe�P�/��{ß
����#i�'���b��x �?!+;)��k�
����f`O�1V%�M��6��Sq�\�Ξ^'ZȪ�Iذ���(k"���*Lpb��a#)|]���*8��%��
tk��T�B��J���)\ϸIIe���{��	Y1��q����-f�P�|�a�'ĉ����J<N��F,�n�	�̭����0�|܇��G���?�Gz��w���aG�t��Ӕ����'�u3KN]#_T>:��*	!%�*=�H{˟HP�h\y�@�a#~5� Z��w�n�>���˘T:�6>-`���QӒ�'�����i�n/�PD�*Yc�hy�v����]�0J{�[���ܛ������r������ɷ߁�'�&���A��x���x�d����(^5g�yKXa�֒g�v?�pk���{�^aZ��|�c|l���E}wz��),�C:f���kve>f��!�p�m*`Mr�l���mP��ˡ��M��Z���9W�P��4��\�M{Ncm������&��6�Zh�`*���w,��ʯ�T�`S�Q�se�e�<}��Y�t~X��s�9,�0do��<e8�yx*xʉ�u�V����;w��{�p\�]�8�{�^^W�S�V��D�G��Dy6��~G�ց�ۉ�
�CޗQvM�!�S-�wYT��l߉�(��g��y��V87|u���;L|���Xl8ja"P�gEK���<e8��Т앇�3
��<8w���m������Owa��\Tj��6�l�0q5.�S���EڴcA="�'�j<�.}I��+���r��W�LW_:p��|�,Օ���k�3���u��8��xW�&�)�Ͼ4�<���O`� V��aN���w���b�_�H�q�l���4\Q"{;	O[`��9��(;���#A�qXx�n�y*B�/*�{�կ^���ɋ�I�;ʚ�Y'}xv\�7?�O߸D_���I�(d����(��Vmu혮�.۩��	��,���|����i��X$Q�(�FS��0IL�HƷ~}�u$�8���l ���M����er��� ܔ�@�g��/�U�x�~%&�q�0�vT�ߦ���q��5�0&n�}�E{��\��8y5]K��G�M@g���&�8����+D���<5��9�O%*[*4*)���
1�<�S��rR<#�)��5��+T��3ɗ���N�ԭ4�@8q>+(�4p΋��mx�mWz0���0bO _մ�,�����l������?1����Ώq�����u�p(H"�T
i������͛��jt��� 6u�T�m qY�c��V���ݾ}����Y�D��t���Ǭ��gb|	����w��
5��L�[a��8A;���=b�WY�ش�5+4�_`z�F]��|s+�lG('[lɱ��0�JCx�XV^�xAfX^�aAS�p/�����R�~]n������m?.��}��e�}�^:��<��w��D^8����E���Z�T\����u<�Ws�ӓ�������'��b*�*U[*��Q���֭#^{��YA�KX��Y��c6�e��m:T�,����aA�Czq
-�C;Z��g�=��5N� l/
�s�<>j��K�P�PLQ~�,xƣ�� ��mqKO

�e9��P�:�B��W8>���&*`�YU{�2�{��-����>)`ơ��E��JE,ï�7�B��9��C��Mg
�uI�w��·PK��j'�4��+|�I����:=�O/>�r�s� aS��q:�󙯧�z�S�o�^�)�������v�3�Zv.�jr��[��T��$�5��`�S�q'���v��*�CT��򐐌�Q�H�/��������e�;ބw�I��/���²�������;`ó������R�(J��4�<I��-32:���%
Xi�
	��.�IA�r,>g�1c?Fh���C�.C��x�I~�p^Ŵ���S�o�v �4�q؃6>�%l����,��Ӱ�����A�
�&���w����JQTnNOј}���R{����!���sB��l�t�0s��w���k��n+O��`GZ	/�1q�l�/�����*L-��2b)����X+kF�Ɣm�7�h�lx�:a�܊��F��Y�T��Wq����:��[��X���g/�c���xV�y��/�(mC5{K^�NB~���5r�3_g�	�6����)��=�T%�b]������tT	SIs+�K�!�ݾs+
ح�h�Y���k%A&ʣh�T�!�lJ��ELS?qe${�Qvm,fr8R��;�굖/¸U�u���`�p���X���H�(��b���"��]e�x}+�EA����[������.��iv��+��r���$�*)��#pK��c�D1�lyARu3}i�A��Q^J��O��yS~�b�QiFH�tk=��(��(+[[�bA�F9�~@�(\m���},k�6�s�#,�O�<�
�H�ѡP���~w��>�"�uU��i9��8����Q�$��oP�?[\��uX�iN�H�1+X-�empw{�`������o�t=b��SP�c��}�9c��劒kW�q�Ӕ��J�Ve��T�-cVͪ��pY���;����M~$3�6O����52p9��;[��-�������)�3�{:5-M�_7��x������rbYQ��]W�Wa;	k�F�d�G�8���}Fˬ YHTr�F@��RV���'���C��x�Q��&KD�0(]nʭ��ս�&4?y&Y`4� �ʜ�c!��(�p;Fn
d����v����Q;�L�BB�g�)�����RF�d+�LF�3���Rʉ�!����nT��%���A&*78|VP:x^\�k���
���� S�Hd3f�n^�|�þ�AVV�CU�h!�M@~�N@�p�x��#�q*8�
3���r�s��I?8k8Gv���������B(��+��ۏ��;�{]R�NAu�����d��+��q���Y6֤�J/^�[J�X�02$A��ir"
g1���`qy0E���$9���^t�4F�Y�)�qU �E9p�J!7O�:
��6:�{u��	�	���{��b�f5nw�e�N�RX���Dn8h=���WlA����Aq������:��,C�T>RW,s���C�zp�MX�^��o��M��ʃf���~�+*����D���
b�� z���-3^TU�Tb]�G�=r(�^����+��[$pv%n$1�(
��Pţ`pxW�n�&�k(6��J_wpTXT��*[�h���1^!��÷�/��-DQ��9 %��ґcCxo�b��O���\�)?�Pän���Ǖ����ft8F뛊�Cݖkϴ|��.�Y(yI��]zl�v� ��%*��w`�tsl�t?������7�gU%�
��=���NH��1RG��[J8�z�����p����[��m]��`��`!���I���[�	�P�Kv�y�'NB�G�����,��W�����m�R>B�[�ͮF]��q.��@�X;��S��h%�r�+~�Dל�6���D��,���΃��ϲ�Yg�-�"�BW`)��?�	����'ˣ�Xu��r�Z�4���������[�N�/�W/���_�L���q˳�l\�6�?�-��Ҹ��lWf�2*�4\Y���яL5A��Y�X��?QyE���iv�Y�Y�@�������	*%b�J8����.�~�6�V�����	�� ��� ��66�t�;*��G��[�0�u�Ӵ�ݷ^�ǭ�fB���_p�
3�UN8��~�qR�j�IZ���P�"�������#�3����^6����M�}CC��`�u9H���z�Ͱ)��% �W ���*|а�ҴK���T�lh�<u�h���*S�q�l)������L���dx�@�<YU枃��}&lcE8��>�26��WN�/+3
���M���@bB�X�W�?2����ne�峧�R���{�2Bem�yX*e!�wQ��z�%∹
w��N�;ԩ����T��^ZQ0<�5��**��U��<���(`�\����ل����1����'ʓ���	ƌ�0BX�F�:f�'�G8�Q�3ᡑ<�ğ=��^��\�N{�7o�g�L���:�!�P��C%'�1�Gě�J�
i���f�Bɣ�+��Nx�՚�9V�O?�w�P�S�����SV9jIt1��䧧���+C�yxAyj �_N�ת����p���.�0CCV�!�s:��37���,q�{�y^�G,0��n�~�o��냫w�Gv���*VY���#"��)�r���_r��4{�V�s�a���3@�����&� �/^��e~r�1�˥�p�u��z���|�̰3/��������G?�A���{�X-��Q'b���i��G���l�"� /떥����K sҎ����ɶ͑�*y���+�t��rI��N�z�7�ÿ��~q��Y)(�Y�y�LC_y�g���z(��2G\�������Q�I�iF�C򑿸�!��0F�+7>#\���M�Z܊i�AR��hBu�WU�%L%">�r�E��pZB�c=����_���A���
nҮtg|6���)�*�0O�Gn��E��o�A��(L��68x���I�%R_p۸�U`(�Sa����Ib9���]���n:ϺW�;��<�i����ӵ�y
<u�{b�.�;C�b��n�6 s�ژ����ݺ��cbx:D�¢�JcL�y|��N�fp���� i��2?�F�\�+���ccE�[�ǲ(�Ղ�9��u ���pM�i�6Z�,�i�L���R��S��?`PKH�S�m�U��~��������Ty�GW�3���8���Oq��M~�EI�XZ�^
+.��.�(��|���e]�-���{���6��3ɷ��?y�R N��#VJ�Ϳ(�
�
�0� �<��D��l��(��%'FZ
v�d��kq�!��^E�FA�2�0��[*a/	�ҥ�"�B��|��E��r����:��=�:XT�%3�H���X�
��h�6U�����9b1�yoQ�Qz3��ƒt8���&��r�y���uQo�'�	|K�A��=X�Q�k�\KCҥ��cZ�i�~�4�Ls��?� �<�?(�Gw�u�:�W���=�;A�)V�=��;�k�IK������M��]��z:y3^�#L&x�0� ��Z�A��q:yZf-;���d5��&�x�2%[n-y-��M=�L�J����M� �PE^^|/���\ƣw�%���O�pCC5��:Zc�d+K7�ӹs*
i�FTQ���O�
U+V�dű��4w	2�)�ॖ��C��B��>>M��:�=2�g��MG�jz*#!^���(���@���ƻ28X�weX��(��t�o�X&�`h2��S"�@~q��������p'Y���pJC�����2a}w�����n����$|+�@���K���?����mO�7_rmC�淍���O-{�øX�FƆ'��*,�R�d2t��.���Ғ�V�UC�*b������ʥtHr5��-�G+E4��L�~�e�
��!�����[7�/�b��p�C����8��&��L�!(L����4����zU
A�~���1|ʐ�����{�.�g����R,����n#�B�aS����c�q��l����T����9Fu�9^�
��:͹Ml��Ε�ᑤ�]��j�I�qFi*E��n��i��`p�L�5��lw[
a2DKx��9��YR�m-��so���+ݖ�'ls����mn��5z��k,S��c`�s����$T���ا���b�����{}]�<q'�a��ǽ���>k�N�P����Th��e>�u�����,C��#��o���*���?�,%_j�6ρ-�Y�R�a�\�2��N��1��nf�Rj�<��N��ς�}:XG�s-����)�Q��78w�(��2�U��3)/����r?󣰞����2AR��z��*O�Ӽ�[�;��:r��[r���e^:�c�[*5��1����EU$uXݻ��qD��a<+.��I��z��$-	cp�sb�xB��1�O<ˍtQ
�:���p�f�vh�WǬ@�d/��h�:�*��iyh�S/0���#=S=',�D&Ct $�̐2���[��� S�7�>���o?˯`Sq���q�R�@+B����g<�&Nv{��+�����/��8��o^��|~������ſA���6̸��K\����\�ZuoZf��쵒H�~1�~| Φ�AO7v}�g�V�T8� (:	���������4|&���S�!x+J�奸^� ��(X�U�rWy�5ҥ�e~V��QB��%_���Hk����78bq���	>�x�/6�j��,ĺ��IP��jEc�f�*a�!�<��
^V+PXwUv��/��?*eVR���C�<J	�y��e¨0�0�s���s��l�����kV���E�vڴ�Ty�gþ>V�*~j]r�ù���.������>�#y��y�7�?�� ˦���R1Z;��Ω�|;�	�R���T����X�WYV�bi�N�_�׭.���|�a�[c�P䱊�c�EQp�QdQ@���A���E�RT�Ǳj��`�˗/d�{li���Z.�Q���y�C��!Z�7*n��e_}�y6a��F�ң���h/�b�r!�,��*�Օg��<@J�4��G�Z0������ye~!Q�Op����,E�W�SGC�NQ�$����ȋ`'weܸ�k�yu��;����B	�0�m���哕�+��Ո޺*��I��ԜJ4�"��?����Yi�e�F՝�?�e�v�P<�ps�@�:8����J�f����̳>�#�2f���&��Cʎ�n��2�<u5�t"{� Ih�Eh��o�3�u��V�������沼���`^FL�hy���%$�R��L�C��_��x�=A��uB=r{�-���y�sSY
��f��L�hf*�d%Pb��w������ 5�IX�L�����Q�D�/>�4����L��D��7�[07��K�7|�B�7P4���\˳
��4U�v��!˗a�4'Y<��l�W6=��[�h�+cj���⣣ �����	�g_:� �����lؿ
`���1Q�t���|�@_�	8w����֠y�k�4��ɓd
�g�J��w
�V����~���Qi}P �4�����@�o�[gl�kxK��K�	G��q~X���� -Z�Jy��7��@yl�	��X�����8G	��7}N���U�0.���-�6;�p�;s��x�y�G(8�W�wI�
T-Wq��/҃=Y<f�}V��f�r����K�N�ʀ��g������T�� �˗��X�(-�!Q|Tf��*!�ou���;bC������@���5�2B���W�&���fE��
�J��R߹�-i@i1Z�\��9X/��n�����L*J�	���<��u�![o0����\M��T��L��a�t�`��o��Ƶ(N�F4?����)C������a��p����w�P��~�������7(a����\���|��%��ǋ���(���0e���\{(��ܟMK�u#G1��X�RJ��"��t:�ϲ��h��!:)��d��:.��#��zeD��:g#bp�|�
���:I��Gd|�mb���3iI��@�����w� [Bvrj�v�0K�����h&��N����A�P�������Y��+(���s��h�:��p�Ӂ��|\�*��sf��/� �
�����jܒ7f���21\�s��0�v.��Y��%���Խ�C{B��-���������eX�-�S����*Dd�u��[��ܮ�zÊa��;��{�����Y�6OE�ڥ0 i�t+���0Kr$��k�vK�e$���FabȻd*�������W<橽O|x�8:s7a��"�M�7^z�^	Pկ!|��u՗�SO�ew������K��4�0�:�
~NM:4}o!֥��4M�[��B=HX2��g��-jq�@�������0�X�C^
RM|�k�;w��y�梬�3�G	z�C�`�Ȯ��ͱ���z�2y��[E�ZT�ܰ���Tl���0�thG+��7@A���7�I^[Nަ4iS�r�9?��c�#�6ܮC8z�P6\ƥ��0p�稘�����hwzT
b�A�rb��|R�z���I�孲�s��lnzT�u�U��a�����/�s��R�@��<��*=�Q�/����eGN��+������)<Л�`�����9WJE�����
�;�1�K6<Uػ�t��U��tD����\+��r�'�A�T�o���Me�<QΩ�2���Y��+�%��3U&7�7��'l��f��#?L��f4�p���-�
D��0���y��*���g(_�jw�g��r �����O�F��b��0Q��q�	��>=}�h��J�#貌_`��<[�h�۠�E�=����V8-u�$�:	W�ƂFy�!^�QF��km�3DU� 4��6`��5WLn�'�讏|��G�o���򥲛����9i"-������U�#�<g^K�
!�D���ρ�����̙�9��x�
q�M�}ɛzO�l��sI��������XgގvO�&<���g8elջ�te�:�Re��6��4b;� ����/� >������Y�x�l��w����\�Q�Z>��b�K��!����'E�r�;0���h��SPƎ7�2�2�@7d���{B��8�2p�?�`ۡ�Sx#MM��H`H���HT�7�~Oܿ��f�
�ińX��2m)PC�1��3�ebK9)������G�T�>���^^�c��c����L(�0|g��� @��_��'^�g��-��9>�X`@�Q4 MC����W��>��t���rx�MIC��=��UZ~��*�K�u~bi��.�3x�i�:{����.��"�3Oc��8_�Fʽ�^3dv~�)��}l@�bA��<�P) �������D�ȡ[�����g��&b����2N�&�(\
�:)txɊ�cZ�w�����0�W+�b��"N�]�vy���ŧ�Q�d��G_���7�DYy�6�c���������7����/?���.�Z�T<~�c�\R�� U�4��׊v��5�/�/���gEr�4�����U�6�*�Z�đzMj�Q��i����O����9;�I�W�|i�vZ��OZ-�TD��\��Y}�������Q��#Z����g=����Ϲp*��>�yV�!ʖ֧�2�f�G*`�^_�|�f�N(f���S�A�%���ǯ(G�_��+���JG�*R�T����� �3�i����Qs�T�y��ʭ�T��1�+[HP�?���:��<�A����G�����_v=ʗJ}��'�j���R�A��z�P|7��?�WX��#�n���[S�D���`	"��#q{��{5K�͇�Ao, ������v$�Xp���(��(ܦ�:d&v\��U�݈�+��7��
$x���D�����_sXͿ?��r��Y��Q�˪��TЫ��T�[�pZи[��gv�j�NU�=OXT�0�R�OY�|�M�K?�S��L.P�������[��/_��%�s��ᚮ�S� F�����/z���6���(��u,{a���{ϐK��F���`kLЗ��O��d�E-�$
4˅Kʏܳ�qznzjG����`�~c�քۋ��%�􊵁3CB���%|M���tEP�xMt����+ � ��2�2S!y�w��H�,�T�i�B���>�мMP���OT�����R���w���Zi�;�����*@A@�Aɏo�ud����*8��[�+��>�)� �w���ұ�ah��T�W�p�3�D�θ�$uY��zV$R�0�P�(7�ŵ}���3Y=漣sL�&�D&-g2=���yAW)`*/�u5��v������^uq�������UA����L|&n���Q��Ė,㫌fV<2�F����*.�8�"���r�Y�W�\D��j9��n�lx ��{�.�m���|ʈ@�W�������_~�a�CJ�.;�on�aﱇQ8Td҈*@�럖.���ə�7np^��0w���;O���	�>>a�ED� $�j�V��9����՗�!�.��*��˳�/2����l�p��#���5TRTZ�}á�>�'����G�e{�J$/I�tdU�J�J&n���9���^_��z��#�5��(�C**ΐ��j3�Bf��]���V�l�''ol����gˈâQT�w�g�KŚ�Qeݡ]礩T�WR�h����ST$�r�%NE�U�7P���7_/>���(�6r�,Gl�1)Vs�ך�u,J��	��9;�sﺝO���a��i�#��e�i /#��h� ʎ���'�N��(_4&�c�AY�E����
��|�*[>�۸|o��8v��������8�� g��ȟ��x3m�:����~W��zLxV=��n� �Sxo^+ZT��E2igg8l�-�i�)ON�W/�qEFy�0��	W
����r�t7�tK���쪧�W�I����S߇G�,�� �΍G�~��2�ď ��H��2�Aݍ�f�Qyy�ԍ�;�.0r�B9���vډ)�61�k���C��G�Wap��!+V^�9�=��#�`r���*��d�z�������i� i @��W��������� ����,�7�4�͞c��'
7��0�H����
Ҁ�1ݙWD,~<q�Q��M��R(��o��^N�|�ು��Υ��T��y_��I�OC���N�M!:�/|���iR7���⮂M���d)�L�s~���.Y�]��\�J�j^I#�K�[&{W��WE�F�F�9S9����Ν�2T�!�?BDe���ci�<g7� ����v�믿Z|r�<
yO�6ܦ����KH��.i��L	�&�8���� d�1[��2)���q̼�������(_W/�H��_d���A����ʜ:�9t��2F����P�d���D}L��⅋�/�9_6��8�zA��*�h�������(%]��!�78��~��{�8�R�kq�:�<��أ���5�SSQs�x7(u��g�}����c~h9J>�,����x��(�Qc�b�������k��$e�J���	��o~�+�V���.�	��P$ge�.~��j�$,w6
��h+ҠJh���dk��(�Z�g湏�,R)t�I������6b����1[O���>�\mj|�_�V��ɪ�_3w��/���Zl���2|��<a�W��Ôn�jG����A�Md(rK��EA-�7�N Sa7Ԙ<�:�ut�ג���>�9�j^�
���o�D�@�o��Z�=�1)��%2�S����Â+��1�����:����*��W��~��J4�8��SW��r�����s%"p.�Z!�S�P�(W]|bh����zGy&@�_��q���"㎇9yf�㎬���R�	'.G�c�����ݔ2^ZV���#m�2�)%	S�X�7���E�Τ��j��A^n����P�����g�M�*g�Ȃ%p��"	Y'��<�Bc�;A��fi�!���c��z��-�U.�Ċ�3B���T�0]�)H���oc�D�LV@�ޕ&�J16���mc]++�͞-Be�D�~��<�8���E}�, ac�@����n�NKb����w2 �I���dbeM��N!���&���\���
B�'^߽ƣ>��x���l��P���v#�+�j��Sq/[.BZ�7���=�O��e��K�e������`El����ϼu�����*��g��i�g��
�gZ����λ�V�QB��N����ء�9_�]��WiԾb��o���:�-]ک�Km<��!JY�n�
L�+�3Ј��}�D,�(�(\ۛ�!·\�*��F�'��\��!sXgCL]Ъ�7R��>���
�2�����E�<~4��oOl)�	�L�5}�zƠ���|�8Ck���n���"U..`�e̹u��x��x���M��a�(�ĳ����Қ祕FA�u�J�>�42��ɐd����C��Ĥ|�F�q�rp;c"�,�Rx�u���C��u��.0�L%A��!F���d�Su:r�Q��I�-~�	Zy�qLl;�1P��n�Q��4G�ܷ�y��'.��)���������9�>FI�! ���/2��4H�J�sU��΢[�Ж=�|��}w�U�W ������m��
O�*� �w(���O�g��E#�$Dxb�����9��V�Iy.���H�g�ȇ���"h|���os25<�iGtl^*����W�ο��Oᝃ6��N���;�O{�n����C�>�8R
��}x0b��zefy�>�m8�z�Q�-`.�Lӝ���-�}��e
7�b����R4����"�e�@��I���[����r�s�ʤ���Q(���b�i�>iɢ�;�XE�	#b��z�+e%����ۆ��G���(G鉸c�	P�r5�n��aʚ�P0�]��a�k����R`�����r/y�e�g�j��� #�I�\�f
���2�DÔa
+8���wb��#;�KQDd�W��F��{W�o�1�V���k��$T7H����[���|�QJ�䐍�i���C'�J�1C��
�(���8p�|��%�^��������P� ����q
І/l5�}��W�T���`a�,OW	ǿ1�O�`��c�K?W#!t�`^�w�JyU!���'��Ub�����x��V̲j	B����b�����^V8�P��-����e/�13�(�yc����46N��KEYs��\��<�]�=��O���}��.�6�Z'<^&�m2�ᤍW�9/�!��۞����PM
�fr-)6�ul��u?vö�(�Z�WH�>w�9a� k���6
��&��ZG]�X�X������C�M�@�@KG[l�#��*�*p�ӂ����m�Ӻ��V)�ާ���a-��/o^bE{�~Y��֩,�DE$�q[�@[�1���L��1Ƒ�g�b�Gx�'�j�´��X�%8p~q�Ȩ8:��}��m�[��|e����70�<}�b�~��K���o]%���w�ֿ������]�/a-W�3�����CQ��ǔ�^8�K�a^��Z��\Ս��e�e�F��3�M�V�Ë����0T�q+�ħ[]� �&y��^<uˌ5��Z a����\��ny�v��=M�򽂋E��p������Y��2�5���L�5|?��sN�H�)�ʿ}����W���!R�c�!��
b!��Z����?n�Ͷ;�#v��
�4��;p��T�ðҔ������SJN�c���ie���z�Π:�2������M�5́�YI1)ӁLx�h����h���IhE��!�e�1c��0+ ��%8���.�+;�{����t���3Ƙ��I�6=`&�mp�uՎ��l &��XִX{��p��b�G�81"��I�*�+y�E��"*s,�_���\���U3&Q7��I��5�˺B�JC�$\��@��	�	gì 0�)�V[cr<��I�Ao#N�
��M	cdNz�ſX�2�3�� n�O�����2K�
R]��+�q�ޥN^��ti7�2x���⟆o�c�� ��n��U4J��D�w~:H�O}4�O��%�3���a����|�Ƿl�K:�[�n���  ���M/�􍥞�;��s��.¨A�*ÓBnWڌj�w�x�GGɡ�6c��AWoeO'�6Q&���9;6����^rȲ;Z�3�1$ �,�0�bHR6y&坻wP��0h��dm͢�R��jf�  @ IDAT�Щ�p<g���[��X��>}�����k�ߤ�R2��w뤻�?�o��w߆���3�%L�>f�
�SR7�SG��I&�3<i�U���y�nL:�ܹ�G��{���Hԥ2Q�<���[zH�^%mE���q�1��Py㷗����G\f��/�&���O��[?݂G��h��T�
�W�I�x��M���s�
U��{��A��8dX��1:RW;>��C��8����b���t`ﱠ�!'-�i��~��<	?)�ۭ�~���ӫYͩ,m�}����=-`��U�TX��{������~��3RrJ�V��w�Cҁ|� Ϯ|#��+-c�{GGh/R����-��,�rS�����a�X}���Kˡ��d��9�2<xG,�K�7�n�=�!�Eyd�(̐\2���+���6N����8�h�����\�RG�}t�������h�'�~�]2uǠ�/��B`-L[lu�7yQ
A%o:S*O:��rū�ĻJ�|��P�4�lb��{ے��W�����n�O�?-����0B��I���j/��S��@:|'/��|U�)��DIrQ(�|S��2Pu0��r7��4񝺃�&Ȳ���9T�PKG�Σ����QÓu�*x�t)�Y�.4M԰�%�
��:�L���P��	x�k���b���$)i(	�Ĳr�����&���L#�(3���	k�'��(����I�-+		o�e�JMR"lh4k�KN�{�%�l����s�)z��8�@�skÙL�m�r�l��6}��"�����	�*,p4 Q����.y�U�b�Y��\��L-w��5��3�ɓ��{�T��wX���AA-����s �s	����s��(�P���
]��KPhqQ!��yǢ(�Fm�3Su��O���4��#��WaTx������Eٷ���]�CU�%�R�TZ���1,��hx�^1R÷i�z�� �Bּ&�N���~�x�Ʋ����#��+x�O{���aϗ(O��8o'u��A�E�R| ;6�a��\�
�2���h)1�nt$�O��J��]�ٟ���3����e'�?c%d6L�p2���e7�5�l�_��_?���{o!|��hh����=�b��E��r�'��,H�J��'ԫ���z��]L�t�����t�	��BY��՝!5ʐ~*�������KWþ!�x���1O����c���]R܌EO�q/G@��/_�!7+?�ߡ_(�"~���/8O�6���pa��ټU��i �DFT��]��%���ߓ��Q��E�J��ü�(iҐH	���?��F���S�Wx���l
����%�;\�����?.n~�y5�v4����&�*O�������;I���'D+�c1�|W'ú`>О���z�P�ygʈ�[c��'K�C�Ұ�Ӽ�S�%���p�C�sAs
�a)Y6�"��X2�T �r.�Rp5^}����rk0`u���y\��,���Y���:@a�`��$�5y�n9�1ܖ�bE�˲#�a���<�[�>t�	<�/i�]%_�ۺͼ�Ȥ��bA�x�h+����#�UVE����e��)E�#*_Zj��j�F'���V�䌲bG��֑뗖c�e`���W�ј�C��4���I�Wh�NT]��vu&�;)��e��Ƿ��6�X�r
E��rn����=���+�Ҙ簎��9�Pn����mcG�1��J�$T53�,S>�g��c��@�O� ,��|2AB�*a�G�eƚ"*/���Z�L�&K��Li�'
]���M#��	�o����� B	O�*e��f��R����f��7�/wa`z��J�*���A`��^L�xo7��Әꍯ	���w��p/��]u-�e�~��,4Ĭg �o C���<WҜw`̐��_3�:<�Y��O% nK� ��
��(��M%���Y��(��)�"m�XN���vyZ�D{��S�ʢj�Ax��QA�UieI�Q�*-:�Ð�L�ܶA�»���6�r���t�5�O4ȷ��j�m� ,T�PK���Oӝ]�Q"�G�,-(���Lx��s6)��U�s���' ��_7�6��@aCf�܏Pr�@�d8짟��NB�y�U�Y�_:KQ��Q���sU|��1	~S$�G�J>�`Ԫ<�x*'���v��iAq�=ғ31�� ����v�Q\�:%�K�������n�t$|�a�g���{��V:�>n�x4�m^�x$��2Y�U|�B�V�W�YA����<�;GVA�|�������)R�o9�B\)h�Ug��g?�A�<6�Oy"�vY�P��J����ɻO�b#gx�����'_��>h[;��Cʱ\�ti����
uq[F����K�N]�쎢���!PL7�uu:,I�1'm,=��[E�d�����m���:�.*����W�m�1!)zW�L��g���|�4+�BF~��:�
zS��;~�p%�Y���gd�Z������ ��̐���U�L�rD���\Lf�ݰ�������O'���@��=Gd�:.�\&�k
C����U� �Co�G����Ȟ��P*��z#�2�{)�P"N���>�!f'ARGS��O~{�)-I�Գޝ�1�0�x�r<���,B��@��SI���Lv�n�u�gj� �θ�G�}+�ǲ����&=�LFe�;p�c	5Lᣩ;K�=6�
��ƿ��7�u��K w9 �&J���_e�~����2A�ZӦ�
��X�l2,�\6���se���F&8�d�ϱ�L��>N��3�T�tT�R8���iC)��2��s	��V���$@p>s_
����:����`M�[�g\	��at�k	3s4�LN~r������6�z�9�/�ج4
<8�`70��Wo�cCg�U���J��1\�s:�3� ��b�R��JEo�8������m�^Q��'m��U���Z?�os��6c��<����&���c��a��=�L�����-C/�Z`xV���Q
��k��Qw�n�چ�+��<:�ʂ�bf8�p=`�'���F$6�
\�lؽ*L5�6�*P����Qx�e�,/B������k��!sĩ�u.�8�e:Xa�&�'�zk��Y��+�!��L�'�R8LJJ���[��|�	qJg�Zm�,��v�p�-�R
�i*eݸMG�E&v��D�BHx��W�z��>�E�gV`_�<�:~������G�}��*��K��*���D�mZ|�=�ي��n���H�<���~�1i�~��EN/X۸@�e�%�!C�nw�^gY��rF����E��v-�(��Y�K���%�6r���úC�͊���R�a��$E&*)�i������*��*+Ĉq�F�u��.���w�7@��H������f�팞x��v��<���/8T����6r)Q��[�k�X� D��we	��>@Y%l|t׋o-Gn�lv�����I���O}���Q��'��Gk�&�������X�/����n���Y� u�:��PO�i]�d^+OeTV�4��IN�4m�wp����V-���!u�@A��}i_h﷘z�s�
�L�8\<g��:���U�m����F	���C�9���a1��h�Tt2q7m�Ϩ1jR����H�(h�u5��3��7�b����3�fx	�l �G��o	�&�7n���u�FHJ<j��:!�����W�f(ԥk���3�1���;T��j���}��[����Q��*fq!J#� ��
����.
6p�Ln��l����.�7��[@�b����o������#����L@R��
n���)�3�O~��Sy����,z���Wb�!��ma"2��ʂ=�!B�ur'q�{;�WE��k�UL��p���(]<���J�2T�0��fT�lЎ]�G�:���5Y�$X��a�3����(�G��@��*Ji���R�����
�+�;�p<ġ 2=^%T��*�U���O�[p���͂��@P�'����',$\��=��O�?�v�
��P����Y|�7��g�'3��|�������������W��O�a]�:zӴ�&O�D5��gP�i�C^j�l>�<��U���4��õ�U�Ze��`�U�V*
Fx����^�ԯ��átX���� 9�h�v}��_��rSˤ��x#O��|��mC���w6���/$�2�ܳ��&����.���#��pS���r��!8���V�H#�U���Ip���ߍ�T��я��_��Y�L���@�$���&�B�H�;7}���kNJ��_�"߭�>�_��]���[��q�[ڦ۲�l���w䦝L3�K���(�y\�\\a��<m/Z�9�\n<v�79c�E>��u�цmV%)wk�e���H�Oq����j���7�Iws����@\�=�]�r�Έ���'��\\O���n�r��G��*`8�խt�Pڴ�g�����L�*b(���δ��*�)K��=�cV�ػ�r��	�Z&��	�0�DS��D���!�\2E!$\�-�x� ��081!�aQ�hq�+�hΌ����fV�E	�C���+���{j'(e%t����ZH4;���z���´��BN�4�\��	�=J�JoE��3�0��D�˫~�+�c� ��"�3�w�π���k�&�S:~�Gv������r�T�Ls���T�����nEr�����0�!�q�<�B����<��.��FF
ˤ�!�`�Q#(��[��;<g�w��^{�*�}��!<��Cs՞Cx������n����B����ť��j�8Rj���ue�!����W�#��O]���&<8U|��Jw}w��a]�+�ĵ�"�q6��u٫�6M�φײ�ݗq5Ά��0�R�]4Ls
���E�^�Kz_����Z4)vJ��Kv���[uV���*ZO�i^�&|�a|���Ti�t�=�ә���j��Y��k�l���;W�
�&G\1:���6�lZ�א��F���7l�ˑ���ۢ�2���̡!����KnQ��f}��˚uH�D�8�wSe�r�_�_I���ΆK)@\���[�1�7^n|��.���k��8�cп�5��-�?aY͛.���Y>�k�w�9e6��G[.r��`�%�ct����,N_�	<y�*a�*���j�6?�'�f.��+�o��/>����sŘo��W�7�ÑZ[mx�	�ʉ����~K/�uF�f�j�x׭���]�d�J��#E}�b�#W�)��wa]�*�Z�,s�f@�BC����(��[�t�[w�y�+
����х�{�2�®,ܢ����,;��&1���J#���LBY��TB+�76d�H�[���b��C#{!{9T�� �����u(v)<	��L%���8�W�
@Z����eR��/( ��cp��#Ih�k�i`�x��lD����AS�����,/y�,I*sB~�l���PM��4��4�П󧘖�
�*��f1΃���3����R94��p�!�)8a����%K�t+^xba%-�	|�ߝ��҃�Ca�P�\���9�)��@�Q���T�����wf��a�V��/r�y�xh��������5�V��}�Mv#�+��wW��W�����C��udY���=EZ�k˙��-s� ��mr��)��2 �|E��2X<�͒Wg�����xV�k��񶂡��+b��a?E��;����:\ו9L�~տ���9ny�"eݫ���=���_|���K|6H�_��C>�{�w��ո}z��w�c��p�~�]��x^��J�TG��\)��w���޴�*�K�J�V);��?ʈ
�OWM%M~�P�+�W�/�a��.��Sc��<^��͓(j��/IZ��j S?�=x=BP�h��JM�"�m�i���|�����l��ů��_�X����F�5�X��_�/������� Nen�D���)	�����Ӂ+n3�M����R�H�n%���%+G��nx(5�?�z�Ŧ��W|����?|�ŗ��q��hw�b���W�UFh��
n�	n;�>�:m��j�
�;t�z�_�I2�C9+�W��������GÓ�(�uZ��p�$֘���._���J�V�Q��X�0����p�˱��㛋/��OL��ɱZ��X�R���0n����T7��,A��Kų�ݤA3s_��!�*FZ�j��ēB ø�w���������c��۬κu���	��<2�8:"Q�6�� #���n�0H?tP�^��u4q�ݢi�қbz,!u�Ca ��.OybCZ[�X�B� }�c�G��)��!x�_*��.>��X	�O�����pg���\�/晗a�g{�'c�8ˡ�A\�ժ*������*��}F�xt�R�7+�4����`|�GI|��O�l����uޕ}4㘿����=�`���3TÄk�u��lP�2��+�Qi�a�e�rQ��sc}1��&�NM����<�Lg��x;�O/��dX�gh�]��sp���w����xc��]Kֻp��*m�Э�o:u�xۭ�U\�o��0�򼮂�5��E��i<͋N�S��ǆ����2��p����{��i��a�/wd5"�a�S�w
����M�����(_����V��[y�ߵb�9��0�F��(��i7P�\���eD
���g/��h|�J���dm-��)H��#����J�#n�}ȇ�]�!��"��ora]%l&O*
��M�ėH����j���W���x�[�#2b�!-��t�J�#%�S��I>�a�.�"�3%G��n�uY 8}֛ς�{Гxt���_�'h1z��.�f��ѥ�o����W_}����u�MD9��e�Օ���x�M��WNQ��W:��)���f�������΢�d�`��,`��7�+�̡}�%=.�o�Q:�(_�@�ra�2m)��7n˼z�@бWq��)k��ʇ&��c��~�Z�c_�aqC-*_�b��<#�d�X��[+N������21��t����Y)�ƁVX��-�ff��!���4�q�T���WXVϹl���=�P�=�]<~�yrh�J���h������4㻈��2�8��Ź3���7鏖�Sˇs��3W��%��X닏�i�|� 	����i��$KV��<+�ri�:���{~͓V� ���̐�қF�|�G��2�V!}�0�^�G��S�����:��,iY�iŭ2�0b�(���L�d.�+Z���ӳ��x���S�/�l^���tNT�����(!�?����{W��VĬ+Z�7�ܭ�����7�#u!	�_���F�X��	!6�iX�|�n��g���ϧx}FQ����w���L������W�p���<(��N��2q�^��g�.ejT���H�p�tU��qTxqV��츌�����ns8a��g���_�gV�����f�CgJ���X�u�t��9��w/��bƨ�ah�ߠ�)*K֎&��CuU��в�����)k������p�E�юA���rGZBny�V��{yiTH�4�I�$���$߯�u��O�	����S�\�pw����G��w���>�5�-����Pǯ���i�A�u�wx�/<�"�t�x/&�Fʼ�6JX�Y0����$�o#N\ƾ,��"�x�Q;{9g�~�����,_���z<�1S�ا�x�'�'M�[L쬪/jAꎓ�����b��� ��M��w�-�Ϳt�֤���l���u���E�zʒ�,G�R��|�t�~��u�+��{�Q�tlJ���I����ɀ6d�
��HVkOܒnK[N��#DBؘ��po
�B �s_��rk5p.��E At�I*͝Xc�!�E��	�ٔ �ڼ��os������?��%�l���⇟n/����#*r�C�u>���=���7� ��9E�]}5YP9�{%;r$=��L�ɝ����[#�L�{m��a�F�h����o���'N�{�4cBf�@ �� <D�e[�#Sjɟ(}}�2��8��V�Fn������VVu��pBc.<k��4fZЭ�c��{���jO`�n�� �O��a��ߧÒ-�U��6),b_�����nJz���t

���s���cr�}�-���қ��_�S9�x������D.��5h��G�H���4�l���z)�[�H��Q���^p�M�5��%Avc��B|��(��6=�[tR��c�}�jۛm\�͡�3�����`{�0�)g����}�߸8'��>q��8�6�ٸ��x��{^.�M���{��9�Gq��(���~��+�1^��WUe��a��l��g��"l
���72z��a��g��#~�'9�L�.�M\Gr�5bl��f�hTt�j��s\�M�,���gƸ�a���?r�٦m_��Ƶ:>ᘷ�,�ŷ~눱�
�ʦ�X��*z�;3�^�����U�U_v
���X����k������{�-��/�鏍G���Xa�I�7?��a���.S�ë��x��N3�q��q�#��{�=���m��!��p���"��TE�����}`Ia���������|8�������;�u�ZZV�c?�({�.t���R��\���.�����]�ԾG�k���*[P�~�~���i�4ý9U�fg�mXlKs�Ic�M��;�؅C��y���;oH�(�{��5�3�{����۽�\��0���¸Bgf��mw��=���ב��/��f�N�t>±���M������hE�ǡF�*��'8�8����6r�/Fp��[L�
ħ3��m}��S��@+�My��5�{w��L/������ș�;7�Ə��;Ɂ�#��GM^�B��_��v��E�-�׊�Ѯ�B\ߦs�3iw�u����7v=���s�4�=���P�'��>�?~�`���O���J��=KB/f���X�y��pNG�ue4?W`t��Ic��3>���q���w�-U���`�|���u`����::�x���8.����R(�O}��McȰw6|�bC�|��Vg��Q�q��� ��F�e�v�bQ0a҉�(�*� 6��;��=����b��T=��z���N�-'k��)F=���#�EZ�?i������������0x��#�S�I?��V�O��2KI{�4ˤg����׸�ane��ߧM��fΧ��`sbЋe����v���x�}��51o�<����Η�pg���ٚ��h(X�C8�8�Ӧ�@V�o����o����ƣ&q�g��?O8��0	�h�R�Hc�����`�1ÁL9V��>֛7��eI���-Z���b��h�0�<n�I�7��Ѽ�9Y���N�)������:���6q~]�����dH��җ�7jZ���4�X-\GW�$Q�6%}
?��ϴy���ط_}���-�h�&�1g��/I8)��������r`����~|��t˫ïv����v��m���~�KI�7���)��t���'�-͒�e������T�����]�G��y[�����k�u��ͧ;���7y.k#p:�}���/���9�_\���ril�`e�v��ϭ��EV���3�(�V�1�;)խ�3%m���Ç���J
-�;�̀@^��(�7�P���?�#�7�??���`���������<��0�Rz=�n:��#�>���C� �pkAB��2H�,����6D�Q9qb1$���TX�cb����2ן��)��>i��;���V�A�8�U+L��t�hl��ѻ3��Ĺͦ��F�ɬ�&����z�6�cd�S��c�
�.�?�A��;����<����±�n�g�,��(��Aĳ�9y���.��;w\�{7�Y\�#�K#6�+����Ғ?����c��k��f�CO�;�� �Y�C�8��4y���M�[��|�5}h��٧���"^q��j\���N
�3��z�����/���Q,{^�G\{�{�Sޒ�sƍS�5M��\����8�`���[7�y=�1����ǲ�L�#�1��a1y�!p��:�P�(m�kZz� �#e�L�~��/f+��v�+3�:o������K+�q�$wv�g
�n�E��y�r�|)B�̪��Q��g�R�*;��o�4p �GC�IG��¢����M�鹶��?�Jh�����	�[���DI���g������h�tC��"~��m"b��������W`���S6�Ã�K$6���~~�o���}ȣ����>|�z��������`�3<�lO�:T���N��c��D?g�-_��w��?vm���ڇ�v�.)����u�� ���5�9��5�7���s�w�݄]uUa�'�㘵�WwISbL�.���57~���g<�+&��O�elF�t�RÛu�;�s�36F�+��"��5x��u�xS����y6�̀�.k*����2�3фBY5�K�W�^��\���̎ ^8�
-�z�
7oE�`��[�|�Bz�>qp�Ba��#�@��ׯ����6�hc>��:
r�{���狚�u�3{�[�<G6��[y�{����2���mzw��R�DuT�\�+�a�Ux՗9�o�ȼ�f@��Z!s29_ķ!��{l�aN( r� �t�3ԥ1���I$���ۈ.`w{����?g�F������PN�e�����tzhg턪���Դ�}D��kx�qai�״7�l�/�P�s8��i{���ڗ�8a�ױ�;����:����L�4×��#���,:��ZL;UF~tjn�[z�<e�|.�	�mꮃ�9)H����Ǡ^>�A�΃i^�!�Ph�Nwa� {�Ӈ֜~_f��H�����F���G^��q�W5����ڄmݾc?6��d(<��l���Py�g�u�������fOiU��C�2Kd�3 ��,<�������9��36���0���*�mXy߁��W�����&ޛuaN>�|[;�_x�AMfǎ����cO0�s=g�F9�CZ�h�ݛ������i��ɟU>�.�6pr�4sS�u��O�H��(s9?cSs��ϋ��%����S��s��M/� ֟7�������u�X遼�3�>[.�P_��~������tW|1]��6��&:K\��K�����_��T���o�Ue����m�o�n�����)�<c�U�;g��[�oǹi��S�gۯ�;6x����؜2+����5���u��SY�-�r:*��k���|1���}���ҁu�p��><����R�kgϾ��x���\o�����]~�AEFe�A*�3s����a��&�
\$��jU�BV:ū�J^'K�Ё�����6�o�������v�T�V�Q��<�Πx�&{�p���s_�:����8?��;����=��|������������i��7~G�Y���T�q�TN
��-�\�&�IX��Ұ���&�֨��c��8�?%-J�.���lb~ %����BR*C��@��R�љz�u{�������O��/^��љ'�����VeZ�nNą�;並j7u�q��[�y�*��w�nG�Z:`΂�r�}L�"�[P8����t"�q��n��.�>���K��]Iz�2w?6ő�|S'T#�H��ZI�AS�=/�pΝ>i�.D#�0I�̍�ّY�A��Ya��̓��Q	�Yf?�ɓn��EO������?gӽ�<|/�2�e���Q<u�Na��M��M���L�.��w�}��]�.�a�ZK��r��'$��#7����<��N� �:`����R=�F�-,�X'��Rof;c�6ވ��	��[�@C������2��ԛog�F��Yg�җ�F-Ҷ��:_)��4����!��wtM[��zɹt���mUD\�E��r�-c@�k�h��9��Ie�0�k�<��4�9��N��~Zb�9E�%�r�B���W��+��U��U�9������$��~v�5�]z��~Vu���_�Q�hۋ�"�O��fu���Ȋv���>�������������~��Oa霹?��W�9׊{����~9�Y�7o�RN���Kj�Y���`�L��ø��v���or����}N���X�7�4~�}0,\hsd��͏�gM��s|g��ܜO���m�ۼ�u}-�	8��C1�欝��=�}�s9�L��D4��5�����4�N�I�E�*6��� ��*��:�a1��uz��������.�4z�]K�u�0Oӆ����O"_RxÌ�G>��Q\BR�P��}�؉x�v�&^�5_e�ձr3��O��R��4�b�#������2��ߨ�Z��ʍ�r�H0�9�e3�����\��O9/�v= s��s��sx����v�V�'��VM��u�ҳzNI�6\��?�6��Kg0m@6>�jB�[H���s�����km����{ =6,�Q:|`�����,:0���Z�a�V�S��p�6�f�l/�x�y�޽� 8������s� �mҒ���4�5+i�[��=�͜6l���Am2�?r{o��'�y�b?�-La�t38�����+=�_�ᘶ�(���2^7}�m��u�n@�g{&[�j=k�����N��S�8\ا|����ۿ�h���^?�%@;�~�I��^�}
���L���9h)��˟���E{��n�M�]����㬻��:5y��\�S�Y�y��Ù
_X�yd�`�&��
��%���WX
o�	�XD�����]��U/vB��ů��n���O�9�۶��\p�"m��!���OT8�˓�x.��O�@��_=��T�)�W���pb�S���7��x���鐸%S�m���C�f��e�m?R��[���J;�B˘��Q�m��&C��{g����7<o������ ���.�<���e�Zݼu�7�Y�~�'W�D�����3m�|���L|�G�di	7�>J�$K@h��U��+%�)CFH��y�����'] @��˘�sx����{�9�U}��<e�7����}���È.�.�)�W/�����U<�=�m�թh�$�D9������>��4|�rϑ�5�vX�r#KP��4�LG��ǝ�=�A�" ����ƣ�i�m��8�x�J{�g��܌a�{ϣD{p�;�`�1�醿�X��o��y�B����u�T�5!�R:�W�B�@���CS;���كzt�q��g);�]��&,Մ'�j�\M��iF�ςug�L��a���@9}#�P�!�<��� :
;�2��GƷF|䌙0,9��~b�r1�y#T.gL;��c���u�`�>�����'�ЯP��gf��o���M?K��_�~}|�*���l�n�j#�����_�6f{��S���r��h�>��t	Rxg��l�,�轈��l�Uv���L�q�'�>i�W:��O��	;�<O����r�ܰooSF؁��e<������,'�Mͻ��	�"���Ÿ �Q �8KCc�ɏvc��N�h���G�"�����9|,�	3t&����u��j5�
�M}/;.��5g��چ���/�n��i�_���Kֶ���k��Ug����/�#��_���v8��ۙoB�9��[n�P�����Rț�	W�.�\�su������������C��cB�6\s�>p����3�Qh",�ѐ)r������s�'�^���d���~�[����C��?���}uP� 'T\��S��>دה�g��1�Ȣ]Z_�a'[ګv��>O�\g����8t�|$�S�8���љ�'g����w�3Y�w��?���`f��P����`�^X�B��4��/��:e񟿹qx�X�����G�Y2���_�V{�Չ�чm��O|��ɡW,��q㗼\p�ͷ�}S�����wb�aNu���LO�
N��luVt����n�L�Ҁ|��p槈T���SΔ�9ˤ�������h�Ml�7�a*�ǎV���lp��5(��Zn��Y�!��w�f�WM���x�(p��|ƕkOWx��g�(�WWU�Ӆy�C�*0����{wٮ��z�wྜ-��CR	��E�t+�-y��UPgѭ<�p^���� �t,��ˠjK~.�6�%7��������4�=k�>�-�Q�y�W�ez5e�78�D{I�O2A@�y�Gyq~u����g�i�P٥1�8�\C]*}��}�ƫΗ��wf�](씰S��"�T@j�uņοN�e�6�Ƞ򑎋D�b�C��w��k+�>}��eg[��8L$���m�I����1��EEL�L8�Ϥ�9�Å�сy�<K�z�PP_{;*��&q�r�ևV�jC��1�'L����a��G�������gR
7��|�
�|�K�9�r���q����[�Y\:'sC���\j^u%Qm�C�z�����pFlWʑ����4˷�Û�U��b���ݾ]'�A����kՄ]�A_�>t�|�ț�̞8&�~���:_�u�X��M���:m�"���͋|X�ɈJ6s�iW�la�2�.|��7J�:�#��r���E�ʥ��+4z�\}�Kq7o��@�(�z�<'����'�B���&p��М�Q��=�6�؆��ɺ/���'3�:^LR���N�:��Z���w����-�;��ԇ��9n|�K��k��9c�����?�O�#�5l�[~ģMJ�-�n�x��%,�l����b{�����ݨ�yM+.?>��F��|����&���~�0��84�ƪë��t�|�����?��	�;�nY+p��3�ʪ�������x=�N��4`��4�\�������M��R�>��Jc�r�l�f��C̢R���$`����3\+_�;��'Oy���ElWy��~��\���j4*=�Lߥ���� �K|2�{�b�$ڦ�߹�.%w���)��yQx��À7����.;�_�o��f1D;)�E�tfK2�(EN�f~�"��8���k���f��/�ʺ3�%���ςF*�4;�(I��̤#���ׄ�
aJ؈Wy��ν���̂���~pe���4�"�ڋr��2ϰ�$� L�~�سE�Z�<��Ɯ�r�7���O`�v��(9�P�������4t�֓|��b>���tL���u.]Ϲ��2�Y���L�p��I���.VVN�y�TwnX�	ѡ����%��[�#�uG���|k�������f�V�{yMk��)3j��i��䍓��2��|4����O|�,��-)�����rª��@~�~����rC�7���z�K嶼�8��\��Y�����,G���N�f�/���^ԣ������_ʷC�0���M��fvV�:fu��Y|�h�G�����X����eĲ�����a��kr��r8�޴*�os�,�Q1X�����j�:_���A�*��
7���vB��[kي�~A�qPAw���S�u�l7���.3)��Vkʠ�?ꁿi�d�4J�dP>%�v�}������#R9v�{��><o�Q>�"Ox��Е������1U>�|�����s5g�8�S~w����?Y&ɻ����1�L� �u��ٟ�<�zϘk�ۯ�]�M�)'���{�N;�x֦�����o��妝�  �D~�'�F�fO�j_���u7�f[�3�~��\g�%�8_�c�GhX�[�ŉ�	� t2�I���I��x������3n��O��-��/Q��@��K�?�p��f[c��]&t�n0It	���;�iK�'�������m-1�[�)cs������U�TO�gʾB�80<@J��\ t�������[�0y�/G���-�^~?����޺� ���@��|Ya�����A!��>���PW�+��{��v鸠��G�O۩���!3/����B��O
U��!JS�U"�B%QA~����E�N��(���8�W|�&}΂� �<���`�ߥNT�ڇ�a���/�|��f�MH�Lt�ަ�˛:ױ1(F�(�tf������3>Sq�E�:`s��@�SXz}A���'�CO=xH.Bs��Ӡ.c�����,�˲��Bh-<��Æ޿��G, `����eP��7��������t�>L3~�^�|�����u�6�����@{N=��u���{�g��γ�<)�A�<�Ԥ��(C��a��.���X�=����2�1��o�������Ƈ���&�t��J�  @ IDAT�q��I.�߁;��_|�HR�Tf_ rV5y���3�������R�Tn�SC�tqy�	//�L��c6gu�'�X��f�B��,��?�u�]�˿i=q�K~2[�2 玾��v�;3Ut�W���z7�3�F�^�t�>��23����;��Q%��ǈv�O å2������^͑�H!���g�uq6�l�.��MeG%���j���{%�I�2e�8a�CN���`��8�L7��O��b;Is^�[����ї�^��Kmlϐ�x�JmK?@�u~�\���8�)�ZZa�v�E.���<v�"�	K�Wܲ��}��Ն4�Vt��a������댧`�\��Q�F�d���0;
�;�Vm�2bo�����v��-�v{�ef�KpS.~����e��s��]emZ&x��� �M�S'�m�C�p#�|�pI�6#v0��_��r/�A�QP���qZ�i�8�g�`ț�2��R<g	p���㧬AC�k<B���GO����,��s��2���`��
��&�v�p~5:��.������e*6S�2E!=bw>��y>��]�:�A����~�����a��j�Eo9g\ԛw}>2�]�2iX��2�p��h���G��c �ȏ����^�w��h0�(άwXuh�X����4���1�J��:�gԿ�Tt���_�Y�x�;�Kց�=Xw�.�Q�����&}%�dZ:���C�8�����`gDSd���蠥�� ��L�a�����-Xa���e�A솼P���Pf;(#|;���RI'���9S� ���ɟ��\���9�"���c֙������&���^I/�heH�<z+��3�ߟs�K��_:GJN�������sf�A���x��4x�e�ec}8 �>lˮ�rO���$X�:2��q˛n������4OmӅ����z�j~��������!\leo9f.��ϖϝ>�,: ҞS[��|\���d�e"[�7#��~EĮ����u�A��E��p��n5���R��f�է��W;�t�ȳ��֞��z,�0�6�����R�Z�6��ЯdLs�2����^�R`���ǎ�8�����iɋe.b�4�V*��z6�KA�gg���B�QSw���'<m��
�:<yى	�+�[�{��mꀱ�6�^�4OK��`1�5�W����-�֍PqZL\�� �l��~f!��4��1��BP�ڄv���)��)�WK]��G�����eO6#ǟ+��R��QY�yv���e�O����˔�Y��r��� ���NzA��΂2��9�^f*X"�R���~��
��^�[N�e�4�� 5�Kx���`�i�6bz���»��3�[wY��oTF�Շ�:"��;��@�oa��d�C��y�WށXC�2_��xޭiQN�v���G�>2� D=��v|P���
^g~����'Fh��o
��Q:#wY�(,6&�$�D)P�*���m�n�{�����>�$��z�Z?bK����A}i
]?b�z7i��y/�zD.��=��=[t�=b�Θo�ܹ��p�:�n"v �����補SHV��g�҃I�XƎo:�>��ŧQ�u�|�ӑ,�vp�isө�(�;(95���o�Kao<\g�5�=���4M���~1M����2xSb�GO���S�KsAF�����ʌ�6(�8[3h�e�� ��	����&���]�[�?4��-'��Ws��E���zh��69rW��߾��><�nً�堿�����2^�i;:X:O�;�UG|p�&�=����8�5�͋�q�vh����	����NI�dM��[��k�זI�F���#N�}P���]��K+7ݰ�A�����,�D�E�.�ύ8|Z�>e�/������>�CJy��#�rH��G=��[D�E�e_�n��,��N��+�k֖�������5�Ŷ���͸��MW-��ۓ2��={ݰE&!��sG�cz��[r{��w�9|$�E�:�%�R&�;��(���5o�����־m~�q�%H��O��v����.�{� ��P��O��_���5����96����t��������'��O�$L�̾��^N4sr���/�JM�;�Q���*}�|��:0m.��K�����x���'����h1�CIj�8��L^0��M�e��v��	8��r�f}+�g�8:�h�]�7��vj\3�t�k�[���2�w�O\?������3T��wbH�<��%h+�+�)����]���X����9��y7�^'�3o��	��(���{,���Qlk��c	Үve�A�P4�T$|x�w���������7�t��g�u� ��W�T�z%����2i����y�{�l�~)l��K �tꅺ��>��֣�Xl7��%o:Z����月[���1�9�#�����X>��[9��;��}�rF����,�a���+y|0����oA����˼}~t���7����k�b��,g���N'���Z�1�j�画n��ȍ�ܫC�r�}Ӊ׋�`���Do�<J����"�n��y&��z�]�s݉���E+���e&��-�q����G,\G~����2�_�Ţ�Z�mXn�ޱ���i�(Ny�������씟Y��8��G'b
_��r�n�% =K�u53��0��Cs�gNz�e�2�����9��w�3���S�i�\� nCO�n��׳�[�-�]MQ+�n<в�E��V+w�����Sf�_�S��7ȿ�/��L��M�BS��:/׌NtJ��ei�<4ex��}��orP7�Ora���%��Ǔ'O�+�]������(�\�8�K)�� m]�E�?�t�-a���<M���L����.�J �b+��5vt� q]%���[��z���s����3�ЮϘ�q���;����8y�O����1M=T�/!�	Ǽ5�e<`n�ϣVyl�85�c�eH�3bC���^����92��b�R�	|���Y?g����	�<qr�NNI�xiq�~2Ê}�+�B�GB�pmE�+��l�1ABE�6Xa����0FIJn4X:'w�����Q &wP���iGSɥ�w��
v��u:�q��1���L�e�O�O��˗��JW�s��'o4�Lǡ*��)X੡^�Qj^����?��#�y�iqLSA%��.���� +R	\�s�G̻1?���?e�vۅ���G�6��~�8h�,>��$I�I�����*��vxǰ�S���)��"zը����\(N������:�[�l�����!3`/�;����nb��u:y;�=�6�U��T��r<GY^ʛ�� [�>�H��*:b6;-�l=׹\��GZ���B��1F�:bm?���g���&? �`�+hO$/\+�?����P��/ }��J��g4䙮Rw��o�ڕ�v^U��O��>��&��Ƨ�<����#����]t%��>f+��:�\㠹<bxY�S��/��9��ѵ���,<:�.:_��F��C��%N���ӗt^t�]�
���*o���^?�>:��}���T^=���6c�Ö:��>��p��.�ԏ�A�sڲ{?�n;��tK{�yt�e�oUf˼a\�n�:�`���׺���g�LH�����-^�y����w���IH�5�.e���@7h>��\�x0Y�:��N�va�����4�!ev0Ҟ������7��ܡgy�y$ɍ�{�v|;n�pD��܇:�V"�µ�7n�o!뭜}2����� �!����>s �b�x�-�4��/���g��u�6��2����ͥ�A��iBYU6\��/�']8e(|����C?Ot#�xq#�֡ͺ�^�4��
�q�߼ ��.�آEF�x>�J����J�ɫ�Ks�	��i<l�e�|d�7��}G���؎#�Es�]�,�;�s_��9pp��#�C*/��	�W+���Q�L���Tbų)_��DV��Y��5oq�·������\X���QJ�p��E�l>�DF�ӓ�kvk�ip�u{ɚ�sh��)���H2�ͣ7��0�����gW�FOC���<2�-$��������D��]����<jC1|��g/2����P����_}u��[�̀�J������dK�f�`;���cʮRw��cZ:b�����8��YPn>�ϔ���aU�3�\0zT~��[#�v��A%uT���@�2#7q��I�<�7���oADbm Go���c,��}����ć��}�V\mo���K��Hse��:�-~�[��G��n�u&_L���f_N�O����0��e|p���Z>��1�a�x���{��U9��X̚-��<�1g��x?n}����k��w
�!�O�6���ڠ��x�|&3q̣����SL��@��I�5l>�4�i�ä,�a_���{l4y�=��І�����:Uὁ�^I�B�C�������7����b�![��R��C�y--�r���xҿp�}�K	XN�s��/�0��e�g|iC[�}�o���qL�`u��!O��
�,��C��5
?�ô$�x��K��/&����K���ɂ݃$��O�t ��|����>��/�<��vWWXä3t��:�<\a��e�b�á<�^r��Hg��d���9�ߜM֞�/6a�K퀓�XP'_�O�[|��.D������/�}��g��Т����k���1cx����-�!�����ӷ���:rKt%�]����q֯��6�ri�G|[�H9� �\��F|����օtJ��W��sڐF���������׌pUCJ&ia�|�qjnA7G�ұ��PLQ��۹���m/��]�V��λ�*0�j\}q�������i���ʶ�s�ۗ�����:�L�[l�LC��U�Npy�q#-�BH�u!m#N�������&a�=�R`J��l��ӣҖ����_�W:4�)~1�3�w�?�����᣼�~����}��Wt,��@f��DL��D���t({[�e�_��mPN'�-al y���ǕW��T�W���tή��[�,������K���wx|��-�>Ju���:�g��6�|U��K������AF���d�f�JZ�緃��b�4�&e�I�t�V?s]z�~�q�̠^�ű/3x�,��c|�>8��Y�It���=T~�k_�X�l+t�pC��g���ym���F{=�w��~'�ِ�P�Aa-o�p�=��^6��g V��_���� ��ψ|sa�]0Y��9�h}���.����c[���U�y�6�5Y�fsdn�m�o����*7�<�1o�+[n��m���,��r�+m��{t!�A���Z�+�=��n:�:�_��s��[8/�1����|y�
�ԡg�3sD,M���*)�6#L��
���d�yp�zW�$}��<p=G��sm�VV;T'�E�����K]�����:~_ױ�9k�^�e�����y���&���q�rë;�����P�K��@��aa�XmF�s��l���gܲB���';({�np�BGY�������~1,>&�3�u��E�|����6��-�T�j��q=��S����7�CdH-)9����Z|G�候�J����j��=�m\o��ZIu��i�k���x�w�\��:/�=��b8��g��X}�
�٠OC�r/ٷ�$C���m�kpRE+N�Z�&߬r{<�gw/q�� zɻL0��7$I�c�/ʔg�1i�5*6��|�@t>j^>��ꫯO�tx̣�wܙ��s�3���T��G}�E��ӑ�^���~����O@N.(�B�ӍsD'���b�:�ՙ��}��G��w�$���ß��=[~<�S��c�/�}����缁ʝR�z���6��Q^�Lj&�s![�]�p�s�ԍv�f�4��$x'�zF�ډ�`��8D�� w��l<�]�ݼ����=�Y�����A��V�ؕ�`p���#�x��o�9$�J-��d�C0�s�H_�)�Y@o-q�3���s)��_t��r�Y�����L���y�4����i99	;�1�~��e��6�BL�����EZ����Ô/���x.�:K:*�W�љi��S~�ӡ����S�q�);��V�^��5_#>�5���_|c��B��U���Z|:�Փ����O ���_}��������-So:��lXf��l�q�2���?����?�)���ί�o��V&�ʺ۽7y+~��733���ml���&m*o�)�v��f��!�1#u�b8��m�{����g,k`h:��/�=��E+�Ooq"{n�1�=(�LF�o�::���Z�NY,��ʞ!g8���~p�zqLZ��y�I7�}�u����ӂ�S>�~͍�OZ|��yT_��ߢ��������@�7�6�_�U��X�<m��.�脽.���ͭ�^ڐ���6�.]Xwډ�\���-�Am6�s���Xn�>�V���3*�p�%T�mG��xd��:�\�1:�׫���3-�v�o���n!嶫�4����2����y^�<�N�b./���J�I�4�)�%�3���=c���b�ҚC��W��n��ޤ�9�S�x)��(Ϲ;s�����
r�+���<+��Zl)�Ԋ�q:���*���v�����	��_n�3�,Lm'�����4X�� ���]�4W@�*����1_����'�@����0���j���#-�� ���cԨ��Ց��3=�k�k�ܬ�ż_|�M֔���GitW�W�؏l��;L�S�[�E-�l�F0��H�jt�#w�`��S�%�8l�\���{w7وO]�p9k��7_~������M�|���z��L������_���c�?m�5H�k-�|�@�)�&�.by��ߟ'^����[ƺ��ci�o����2ρް�C�2��'�*��7��E����ܾ�i�1�91���iy�]�Ŗ'��f�5]�:����s�?������q�tfԹ�e��2ny�=[�C::^nn��œ�b7Ό�/܄�&	��i_:��,���>��o�}�+h���@Y�O
=�1֟p�=zx���x�37Q/yĕ��I�#�,��.����6��V��D^�Ag�2C�����~�wCd�0\	�rN�8{�.h��5f����.gLr���Q$}}�l��#lxu��/͠�@W��|H�d�;f�ذ�s�oNp0x
6�C�xZJ���p.�kI�v|n��&�~}��5ov���r����sm���to��|��&�`W�0�-%���i���W.��ʎA\¬��eێ���m�������:'���H�HM�yb�z���F=9��,[���D>'w��A���+u�x1�����@I|w��*czt=�gG~�O�l�7[�z�hAK��97�sb�ą!��^Q�+�x=���=SҾ�:��ҡ�� Tx;�zɹ�S�͙a������b]̕��J��R�Ѩ������@�)_�:�ߩ����C�G���d�g¢��%@�9R��t�Jr�O� �w�ٗ���N͙��?��z7"�ų�-���;4�o0�HŔS��4�����"��Q->�V�)O��kH�����.� �А�ۥ�ٝ�u�������':nf�XS�#�o���������*jt�e��\��W�* =*����/��d����-����6^re$7����[�f��������;��y��8��W����/����7�=��3欦��?���`���Y��W���Z�r@Mۛ��7�4�QDL��,s1lm)�]J\���)��Ói�M�A��(����?|�e�b���~��N�iCR<˺���ʾXnOc�c����e"�u��7����?��t#�=�N�p+�q����n�3���}����ǡs�ćOU!�x�[y����o�ʇ��^>O_���O����?���O��c�pt���S���������	rs�-��c�4̍�#���<߮t�X����2)+M:��f����'������xlj���<�T������_�/w�]���6�btIC+r��C�%l�"�O�'��/�"5o��ΓfƦ�[��'9:�OY��ca��|�<���_��ߺ�����������M��2��	,���~��$��#s��)�)jq���3>vZ]Z�>8:(.g�x]{F�G
CGv�{rdn<rQ���I��ˇpp�ζ�����ڐ>�&�b?�Q{�$�2sQ���Yw�b��M�*T�+�X+�B���$�"��� 4\?-�E�
͂��?^�N#8�����M쯸�OR�4���>l0d��¡(v�"�(3��E�L�r���Њ���#2H�h�E��V�Թ.��8�'\ͧ�.z��a>$~�&oKy�˴}:�����Mc��J���|�_Q���]��#�S���,�!��ȚK��\�<��GVg��њ����!d��q��`��H�����jf�X����_�葩p:a��f��Z����%_�ɡ�mrə�����E쌃e��:�.��6�7�6,s��u�������e�y�o��_��,OR��z�d�V�A����l����H܁�v@]�,���hbs�]���c��b���u��l�8����Ҧ�b�Û2���ҙ~���"����k�`�>o�oϻ���Oᘴ9�6�~R����e=��O�0��㤃3�.�9N��<����s$ΔWfΰ+�A:��ěE����)�$f��ch���SZ�?>���H�=��{�%q�x\��������������Ol���ͥ#��\�v�.�v��3�h����Bd�$O |�[{�Y6�j�ª�M�^������W,�OvR����M�H:<}��Y����U7N�Ο�4h�+7Fbl��� #�|Cɗ��g|�E�V���<��M���EBA
[h[,?��䍽8^�+n~�[�:_���{��_oX��i�&�死�s�e��7�2L�`PWo�_D�ώw-�4��9G�j]��<i������Y2&�4�~�f�wc� v�Zp����J���Bc�B�L=B��N�u%�i��<1^*���"���U��G���d�Y��;/<�С��]�v3e�#N86�����C��F��D<K*���\��ď���ij��رۂfJ ���LT��G�v2MP�UQy���c��r�Wi��b���`�6��9,���X�t��8�z�j�H��k�FCg�L�ӱ�I�ȯ_�7���Ŗ���B:hy+���R��إH���::_��X�5�������=���	��K����NZ�q�rvλog�|��bft�\���G����7:y�����_3�u�]��|W�K'���;4�����O0����F�sP�k�ox��`}���ʇ��8`z����;���|�˂8kG�8+�>l��AC������;>�
�'�y�}�q���?�TꇇH�ӚT�����3��Q����w����E`�M��	�`'b�y70�sq�Q���|���I��{m�2ܜ��'.������u1}�M�E:s�9|.}L9g$c�+������ҟ�ֳ����ۊ�[v�s�����Y�:^�zL|蚦���#f9�p����>.9��I��n-�$��r)`j3k1ŕ*ڰk��G]�N���nsCᛋ�z����n�'f�]Ю�׸�̓��%��o��v�O��MdxK?�,�a�5�3��Q��ζ�����״��#M�\h]+��V��P���>�go�����Sf��xxq��\�e;��g&���G����ߖ�A��RY;n�'�]lCÑ��Ro���*!��Up�q�SF�9�O`׵�E⾵שׂ�����S�7l�����?��S�4�&�]w��˽/�9�~��[���KU$�_��B��&X�_І)��)�D��O�P_�9�Ү�%���1^�Z�W��X_D�^��a���|�ߧ_�N��h�ιM��,m}�Q��>�4��Mx,�[Z"�����r6�]������`�q�x���⋛L����S�aގa1/��nC�[)�����oO"

&R�̱�b'���D�X��P+���'�d�L�#ox��,��OC�\�7�tr ��n#�:��t-��s�`+��<��;>���8��v��)|a�vSE�K(�('א_���J+�%.�{]LG�� ͓�ʟ�M�t�����fC� ���2|��ɣ�,�����	�F������o�a������"��v�A��{�F�#����D\��7g�<�+��e?�K_��ih?��MU͋:��������\�u��z�C�3kc���6�c~��!/Y�|=�n����\�:3�ؿ���/�Bc�߻H; �k��AV�ZW�ӱC
���1w� M����ym�����Aۗ��-WX�E.�&߳i{��'q�L�����3������H��ӝ��=G~q�v��E���~�:�A���1�A����d/�i��8q�� ����f4?z3 �4�g���{y���.�G�u>�^]�x��/��w�!_����d�_��-��F گ9��cE��ə��\!�ip��F������{ϫ4m�)����A �SU@���M��@���8,Ϟ�f��샶~���n3`��$iӬ�N�L�Xg��\�H�h��.w�ٱ�^o�FL�I�?uZ�u�q�]�7>�cڮ�rv�ud�d��z�Ƹo_������x��/�|�#�������������FPF����$����ʰ���~ɿ��:~�r��𥞣0����K���>�xlRR�������#�k���1nl�u���(ȯ�$]ļPoE�?�����Of�N�X�CWa{p)}����_<�F3��L�;�c-I���m.~M<oǸ~��k�3'6\+tU3Jj#� 1��<$iP!� t�\���Y,ȣӠV�E��WT	ӣ�"��B�5���	rIɎ2�fi�O���:7ʑ~���/������/�#���wםo;�v&��@D
G��� :N~�����?g��0g/�+l���r�����y�a��B:-��Q�#�鬿��s��/���c�����_}���W�������޳�c���~�]�y�x0br���rK"���8���+�����-�QD��u�!^=��\:��,7�y�*�vx�Qn��}���h�����{����^��|:C���J��Ƭ&q����k#�X��tS�&pa��qԔdF�^��X�mq�6�� �i\s�Ӵ퀿�� �p���6e��SF[1�SW���zmhd�~��N�OmN��o/O9e�Q��p��e�N��Ҙr��F����T�wM�uh�F@'ݙ��?tG&�=,ӛ���o�N�7��C���%�o֡�N�^���O�~��ۨ[Cy�~��Eɮ�-Lu�,}֟Ao�-o����'��^}���ŵt�FA��=Ə,���U�`�C� ��Q���q��}ڎ�`����|����U=��mޤ��yx�@�}���^&p7�?{��b��V/!�o���)'~�%�Tޖ��.>4g�t5ra,�0Yθ���^��ϱ�)6a|�n�菜!��o/x�����:_|������d{�ܷ��3�����*�Q^��#:�+�R+��=�0�n�p���+�g����K~���/vhJ�#�^�����ȅxS���d�5�8������ O�kz��	;���Es=?�P<�C�xd�k޺FM�vzN2?q�H���p�L&���-υ�c^;N�h¨�	v���*)������r[n/)4ϪҮ �y�o��џ���x���c �5��-1�(W���ԉP�ͨ�N^4^·w$Ί<�����^���_bA��1�O�P�V�/��h��k�ċK�֕�eg1δ GV�H�t vP�ƭQ����kw[~΋O�<ς�G�|9|�da�l���x��u�G�!b�Й�W�ZW�c�^R$�p!�i9:'M'�)���q��w��<3R@�l��<uL��茋�~�~�0;s��y�B=e11�H���@����$Dmc��	*�@�ӈVJ���-�d�7�ݟ�!6z���/������ڂ��r��f��㙸��K�-�� �`����x�G�m�^+S�x�7|Jlp��4��ڲ���E:�ۗ-�7\��i��,P�G��i|�˫A>'�V������,���ɲ��E�ʬ��8.�W'�Q�����C��Y|d�lP��G����Z羱��u[���#W_Z���������DdË��Y�2�)�"����z�~fti_�4����{,+;%�X0�'�lj�O>:��ty�N��2��J�3���=�]S'���(�~�v��>u�~�7������BHi�"��s�}�i�M�L��/y����6G}�����u�����z/osSɣ]0�A�x�yc��.x��_��=�2�[�Y�ʋ_��^��9~e^����������VD:�"�F�-�ܪ���Y�T��>H��r$�t�����$���<�'Z�-r����LX�o��@&�{��X`��|�yKم�TS�a.-Jj���Gl���hޕ^Hկ}�I=�X-i��Y��ôHMe��r7�r�D4Hi�"����^PC@8oEW��XUS@�������l�e�N�!7��;�B6����9��"�<*�q�\��C`�L�i�ȟ:�m�߬<�	�滏<��ŧ�~8<�n�;��4�,���@>z�MR�X��R5
��c$Vl�J3�_�3�2�F�V��MI���O�tB�ʵu����<�Sv�v��ÇOx�3y���_�`��W��;��#X����S��\�_.čUw+�e��ަY6#��e��4x{�+أw��|��(l�ӭ'��YT����G������5�"A�����wv��wP�q��FJ\:�T� ������:�Y���*�	������Lj񅲸ũ�� @�bZo^	�3u�`��u��S>���ȃG;� `Ay�H'5smy���)\��l3�r!�����5+Y�L�i�x�Bm�ΚGJ>s��ύ<B�����:�ѳ��V6����ef���ҫ�8�9�':�MA�2�"��G}ȇ3F�z�[�y��8O�Y��
c\�����.�$��]�G���Ǹ�ʦ�kg�Y�t��:޳Tm��o�7va|l�]�1���i��3��q��3�ul#'��#��"t��$�~��-\����+�aO"mu�^��8��Ug�lG��H PBm�h�hJF��9`���X�ئh����K,F����;�b�q����?��S���@��cY�f��+`(m�#�8�x���N''�ܴA�/A�m�1��J7�N;l˶|���x�i�郩fP�`5��bڤ6���L�~��ƣ�x|��Ẁ�7��|� ����!�1D_�4۪r�� (|R��'���~!u��&�1��C�;�1�a�����h�N�Pi��%��Ħם�+1)��9T1i�fc��q6�'"�s�&zH�=�fC��>I������NI{������z9�Y��ęԡ���&̓*!�0��9�F.��\�D�Y�\���!�r�@^+���1f���Mـ�S�UL�;��K<+,��:2�"'7*�F�Թ�dY��5`4RɅo�˯�F� ��i��P.30�T|�����a0�V6��k��9���|�������g��ө��z;��GLr�iYy�#m�����ʣ�ѐ?3_ʛ�}ȶ՝4���s�=�����g�)k�q��y���ן���m���b��/��5���܉!mZ�zS/2f��n87�a�$��#��U`���t^ޱ�,�hʠf:T�a�3�w��[����S��~��X�ʟ��N��w�l�Z���!)�� ��Η�%e�����,b���@'�䜶!����e��ú�clͨ��H���:�L`���B)���ha7�9&=�,C��������@��q
qҀ����<��9��u��UQ(�
�әg��# .Ӵ�����d �8@�K� .'g�<k7�\98�=�u3f�NV��VY웪��v���#CU/-�νk�޳����t��az왴��Յ������5O�:��h�Q��{yR_��3��QƤ��G���׫�t�l��m��30ࠥP���d�0X�, ��˒�h�����s^��i���MN�B�x���^p��c6Ⱦs�m8X���8��oI�MwlBG�~x$j�*�\���'ɹ��f{@��N ؂�*�u��姢��̼�l��%�=�֫Ns�|���̐�W�}��>;ܾǓ��������؃v�Z���tV��pL\,mi�iŋ<U���>\�.�x�s���7g}�6���V�KWؐ����ˡ;�!!~�1TDݰ������/����VG�~��R����N��e7�	�{�v�Z�.���Y�'��@ؘ����b��~����J^��	�=�iڊ��Hõ������1��ZvX6���	�~�Ȅa`Τ���:T#�l�z�6�:_��\A�B�5�r�)�TZ�	�@.q���/����˨C��,g�,�W�6X#@�!��/�Wg�:�xr����b�+wO�����[6Ht�w�C��� >:��?ϰԽ�J�Ngk>��[W��CS./��V#�@�X���ܙs�3p6�}���Gޒr��o�s���w����oY��'N��r�}`'f~���H�+������1N���7^w���T&���%\k��6(��j����S~u� �D�ջ~�h��w��.��,u��wr�f !u-��'�M�U��V��`�i;��-
qx��ܴհP[t��E3	B���k��ە����0��{��6�X�N͕?��X�");?��$��73guxjS�sy��uz�^��s�۫�uvv�C��㚿L�èb-��i䷎ZO旦����7�მUo�6%�9,�V	qΛ�#�-�E�&�C{��[vf��4XwH[|�BkiEk�޸Ξx6��QB^t�>ӆJ\�������0����u%α'pE��Y<t�}�l��_gQ=��$Pߵ	�َ6�ЖG�UN���<�����&5��I�j�IQ�XUқ��9��!��m��c �7�^:|�@�4��ow�=�_�x���v���<|)j�f��~Pg(vо��I���>�MO�H!HtC^����
O� $�#3D�p�|��Y/7�΍#z"�q��or�ӿ���/�d�/�4x,�zg�ԅJ�TP����k�zt���de<��+{�d�������n��9��ܤtf�-a���z�NBMn�5{�\-^%i��԰/�iXɂd0w�a�#��}�z��Wǎ�����&c�e��t�3}�%�	Bv6c���["���kr������P]r�R�R��0Ha0E���U�0���l���:Ep�
���=�3#��krbz@��f�*iV�`�9��p����Bh)��-���Rf�쨗!k��Qk���M�W��r���d�T�7w����|�ٔ�x~�=�[{g9�G�tXP�Y�[ q�K�b��#&,u��l�j���8_և�Y79�)w�;����S̯��z�^_�E��­{�>���&Xl��7�Ϋ��t�|�quҫ!�0vaƾV��Ja�)8К��ԜH0+�$�6r)�:�E=Xs�v�IDn�w��!=��og�m	�ࠑ2��rV� ��7W^722W�@&�x�:0Q^�8ez�^�3D�@�@�`ʥ=���m����?j��������$52�T��-�$f�ǩz7��/0<�T�ē����;N���K�N��ԑR&Q�$N������x=��Q�1�<�L������E�mc!��c���|�mhy�Y�qN,;���p:�CO��t����^��e���hY_(ɌO����a?#����7�z֦�ڞ%kЭ=�[[ɆIyQ_G}�O�hm��L�4p� �Bj�Xc����\��Rz���i0]G3>� �[�k�/�e��{����q_e�X��"~3o��1q6���N�xՉ}JdF���֫
������.�f�c�u�Y�Io��M7�}��`?\��>r��Ue>	��Rߪ���~Y�.[n��뜙�|^I^��Wy�l��tX�dP'u=	mֱ��U�� i�T�u��O�[M  @ IDAT~����7���!?����|YO�Mu�'��3���Zބ��h��s��&�ϓ�ů����gB�Ʉw��i�O$��������+<١��͙�O-a1�R�����	gz��`���~'�p)v����uy�\T]�/CB,NZ&�5��������G*���ش���>���#��i�ӹ�8��i�V�A�J$64��l|�U��6��z�tt� ����y�a M#PW픳&�4�G}�շ�p�S:��̂}Ϛ���rgv�u&�8�4E������1'�:�^��,ro理�r-1���G�<����x�Ѹ^�yx���x��#o �F�����;/�����͎�7n�c]�9��{�ȸ�V��AH�}1�iC�T��P���e���PWζzt �ެG��Y��H�l�`G��8
֑H��K�}�Խ[q�|�iί��|$`'���w�����:a�6��8�˥��VyS'ᷢnyx�o�#�G��)e�N����XP����h����O���%����$?�Tvy�#�N6�\�-"����;~�;d��5�HN'¼�o��э����>�St�YJ�v����ި5�(�!r�����7�h|��8����P��F��|��a�ʈ��v�=�|�B�}3���7mh:��@d{)��o�M���Gtg��*;���`����:�>����r��\��\=v��~Ŷ:4���:��$��������X�t�Z��#��xGފ1+���,T��>���C���[����-�B�a��]�����r��H��aP��(x��ߺ0����b�(w���3���t�f�:K��.����Rr�ph�������].g�|��&�W��R�7_�r�
7а����7?խ�n�|�@��U�v�ur��(�K��0��VGŗ~�����v8O��1v,�>�}K����O�wo�U���1-oycuhȄ�e8�@�c�;�]Jc��j�����	��6�RӀ�ϙF����_3��6�wu��z�D ^�B�8g9[�Ԟ�o����e2\p�*�x0I�G��-^�^�dvA�I��w�֝�6q^4�2&�<�B�����,�ͽ��v�����o��G�L܈l%M�f[]����3)^g��|/y-kЊ�/^�9Gny�٨|[��i�eFL���[$,gk�W�>>g&���>������Ā�#��*\�?��1�1*�K��K���Hg@'� g���ź�X;񂽃���1^y>���l���7߱�!o;���
;0���eF�QB�U�2\�+��Ea�M���r�^���s�HdPv�8\�e�I�q�����
���H{��6*b�"t);w�q�a��ԁ>75T}�S�],>��+�2�!>`��EO{��4�)�(�r�2ɘ� ��`�������I�"0�<��$�r�-�C��6q��Υ���S�Z����j�ߧ�BV8~�i��}�:p;Tx��ɫ�9�olbvA����*����U-�=Y<��#]����2..���C����e�2>�,o��~�W�*7�C_xym��e�$���@������n��ٲ��a�\H��\�&�(;}����U�?y椏�ϥ�f5N��v�Y�F�P��Qpj�����0����,C��f�uƵs�k���nw��WJX8�������w+׆]w�Hm�괳�G��$~�oH�h��anh���8���᳾��o�>�	:}LR��%��3Ɖ8\�F�u_7x�3/8e�=�x�ޑ_��.w*�6Ԓ�xn:e.�DUJf
�@����7�}S�J�ӑ�>coD����������.q+k��"�]_zJ���P��֬:m�b$��7���+���f�"��7�Y��x	l�P�Fy�O:.]b�3�ެ^�wa,���C��yjy�c�x�H��z1l��D'=��٘�)KN�
���,���:x(X[p�8j��ù �	�qO0���^G�
!�sl1D�����u��<a�i^ٷ��aK+���/q�D�Av����uUG�X�ԭ�@>F_\��8�����H��pV����e��ec��sq�V�̞�F�/O����eQ#o^1E�B�t�1َ_�H��9"�BySn%x�f��띃�up(�ޙ���{\�୛�8\Yh���l-A�b_�s��?;��?~��,}ㆅ�l7q�]���%:*{]�D�]+���%����z��Du���&or�����w��Σ3`�֣2��3����4�:�������q����5be�^� ;u��������7��5 g��g��I3Ծ���]'�%��_�7��[yD�_�B��{��p:�w�6��uXr%�Ⲅ�-$.S4*a�ܕ��&z,���M�B�5O�Cu��8!`ne�V��p��iG��e[��[���K{O���P:*��PN��Jc�͘gW����~�X<�c�����p�eP��a���8,���Aǳ4\��:V�̗a��Hkp�V�4_ܮo�~�>��7�$�i�k�s� <��z+���mG�/:����ᚦs�͈1��S�����a��8�I��hg�L����k0�xe| �����NfD ]�h��/s�˽�]�1>���5���ǒ?���G,�����yK'��"W"�x8�[�������̞�B��G��·D���YV�ȗo4�.��8�s>+tg�N��v~��q.��I��S^o��_zT��7�W;��s.�3vsL
~��.1+�+f�޲%�z�|�z�������?�6���oQ�k�k����M���w=2������д���e&Pe�8�Fcw�-�����G��طng����S�g�A��^y9��vs`i_n��$���|��q[ہ�f�!��#Y�Bjҟ�z�Q����Yq�K;�����*�jB�8a$R9�U����i��E9H^�m�5�)�Y���p�"�K�4B����G�u������ |�[�,�ف ��#&�wс�rd�s)+�b����o�W�%�x����HM�axg|�#���W�m`N�fm�k�@h��A���(����U�:}+ҫ>$��ݛq��	��:w&]P���z������w�:__~���׿���x��8dqٻ1x�V"O6���֌�d�ѕW����g��"���v26P�'������7ƨ�޹�X�#e�DTX����G��ֶ�u��9z7�'�ĭ]��Y�6D;fg*����p���Gq�Lխ"����cʆ�cyo$ʔ��0a�9���\D�����1^������:��0�a���#C@W_����Al�����4Wg|��x�?��ߑWq��5��KY��t�t&�e�8\���%��q�&ϊ���޴ˮ�H�=�A�I�V�����`���Z��D�$�U@(��yߌs@���Ϊ}��)2"222rع�,ﺁ34�\��G��7L��*=�q��Su�i�[�/�őB�3��<��b&�8v�?�ۂ� �e�'3n����F�� ����-����c֤���CcpO]���I<H�HI�@M-�B�}�3���2�]���^�M��c���=���v��������Xgn�|���������:oV�����U�Hi�[t���n��xcӤ�9�!�/֙oc�;��NwYr�"�#��u�L����w�#�}�ȯ�I`�\����M���G�+_�����Q~u@��H���y{͋YW����8K��X�u��n�b� ��S���J�t�?/���)��	("Ɇ�;m;s�W�7^5�D��l3�"�VΕ����mɥJNH�I�=�/��B���)�h *����Ȫ���p�Px��)��E��>��
��l�!�s����g��ҡ-x"O�Yc����8a��������Aص뜌��!�<+���t�EO�L	�/�eeh��7¯�`-��ܔ��<S��u#|� �r�	y�r�EՆ��g�/�㬠(��6R�o�}[s ���]xtx׍�_l�x+��[/^�W�_o��໒�Q�pU�*�|�ƫ��g뷍[Lݟ��vV��B�,Ɯ��y�RLg�Է�J|����s�2������H��2M?yR�0Ԣ�僒���}#����l�z�z�����c�Q�mdv��?���%_̣�KGH��h&�r�m���.d#&�sƇ�?��Q(K�yy�t6N)S�jy��p�4�Z�r�uN�9#�?o��C#�*����	B\�5��\�aIf��)��.��UF���������F���c��ep�/\��<$��z��:e�K7iRO
�gU
�:V	w����6p&���)����neEg��û~�^��X�w�˳�]�G��8���t�Ng�I'�wqʌ�z�ۃDu�JC�|;~�'�A����3a���3dV��=^��|�W�,�g�i�9���O������󲞽�C�7����g���i�ã�H���
�Q"��j��F%2~tN�vY����+R^��V�K�'о���[uQ�ʵ���O���/�ԋ�sζ`�0���s��=x���_���g��o�sΠ��T`1#8.��x�A��_����UjݙNl�+�@"�� 3,~c�=jw1���u�*C���}S5���Tr��J����9�-�t�;R?����{}�+̉�}���a��>ξ��\�Gyyy���w?�ǟ2X����]��7!��SF�5{w��?eD}{x�@�~�|�]Zx��|�o&�EF��T�X.�M;瘑�|�������.M�Q��)�Jւ���߿���d��"�7�_���'���8�>�%"Fj�'n�[�h�NM|�,@'�L����,�A�Ɨ3_���f6�]3��	�\"��Lѹ����ܼ�A�L�t�"_\�X�U~RN�9�]����.�4���%o��	N�DS�>�-����4⫅>gj�l�t�c�%g���|��*gk2��4Jݠxי0�=�G_��t�%�c�$Yܼ?zy{�^�F��\��;�\��C���0i��+.U�tT(e&X$����`����f�'�~���W~H�K�
�3���H���^��"�T\�B�_ʷq���Â����m:��8���(֛C�$8d�I��Ȁʤ����Rj@��K��D��3h.�~B��ůXr� �c���!��1u��?>�7�<6��XU�R/������"w�Xl�*6��{�~`A���NQ
w&�u���t��Mc�ܷ0ġiVJS����oe�#<��й�!�}��Y�q5\df�8��^�8F��?6d�Oz����D�,����?��Y܇�ⵛ�Z�D�45?��_�4d�k��,���Y-~������Sy�i2G]a�7���j�i|�����|��7�i0΂kx���'�y����o~��	�y�k����%ߝ��T�b�į+OJc�n�U��t)3V�/���`Z�u���9À_�U��~µ�ȃ�Lq��o񞰍��A�}����2��{��|�c�=������>�;�+�8���v���ن�7�ڲxB9�S9�x���/�~,�-(.�z�q�*�� #�����޶%�^�J�_e�-[�V%���1��L�S#�MH���耳�m����B?�vM��(:={��*��	2ǡ��*Zf�җRХ�~�D��!���}0�	��E~�H|S��
����%��	pp��=��IJ��O�±���aip�� ����o����$&-�ɺ�L�X��R?�����-�+�E,.��h|�l�5vh( ��xͨ�:�H��7�
�Є!!Zw��(��img\���H��d^IU�d���N+L������%^�7S�S�(@�#������l"�����8�bxn`���T�4#	ՎBS���4�T*�F�	12����s@)�G�~�m>�!�a=�@Мb�Aa�7)�3Yy6�is��W�}�Ye�������pr���o�9��]����͝�*�ӳOHﴷ#+�(=ܕ`�A���I9M���J��֓�����o�ZΤз �C@�w�}�����K�V���Q9̡��r񞷺F���1�� ����KN�~�	o����F��.�5_~��ͣO����~���tV?r���ͫk>��m�شq��E�A{���<�1IM��k��(���=@�G��2p���Rb����e�
��O�=�(@&�1����xW��l���yȒ?Ϳji�tMՎ���<�6�����A�ez͖2e?�K���V���sCg�r�Cj��S�i9�/ӈ���줧��_�pl�83\>:���v6n`�#/a����~�^�_3�����������1�zDO��o��6�L�m�?�寛?�៹��Y��s��P��}�=G%���ci�bH�cB�N�C�9�}�q�s�nM|��r9I��˯\A#|e�S�>�86�KKwٮrt� �7�o0�n��X���{�|�գ"4Z/��o9bֻ��{���u�I�P[z=�R��D�
9�3��n��T�l�	<ed�*��s�=e��|k:Y1�Ê�M�ޏ��b,�	��8�Y�)J_nL8Xx�f��������^���=��v�%�v����K�<_�g=̞ghqv�-.����Q#����f=x���,a��3���A�9�#墘=��/�lS�ҤAX��?I�o��=���3ϐ�#pJ}��mH��2ox���ȯX��0�~(��PP��5l�8{iir(�K�\�J;ˑc|�2	H�T��I��
B�=��i�u� ӎ�q�!��lk��pf�3���;Ò�$?���h��''�"�P�d�W�C��r�]AUX�E�ĶӰTI��7��ܝ"�2~s�$���|r�f��f�)�]4	�t�ࢸ��K{��u��tfD�ŏ�y�$��M�(��Y���|��R�Yξ�93_��)`R��;4@Oh*QbH�8K����y�& �Tʋ�}����~��&5��8������f�L�nO��j(����lP�{g��ыw՛�҉��Q��s���=����bf	��G�>�|��7�˷��� ����穼v��~�q�[Y��q�G�e/��A���0��m��\Mey�}Џ=��Cx�h�Nʌ"R���?�g�c���mg���e�(;�O�)^�ڪLp��M_�l�VM/.S�,�ʮ��K7��^�h��M�x��S��5��N������5���ih������Or�2��w���LAi��d(<���]��9f��,_�������~Ɂ����-3��+X`��R�uj{��*q+�9�3�����x��mn+�	o��ޑ:p���['>76�5S�����/1���
ZO���{����I�e:d�9}�y�}^���Y���5�탤�x�2�N�k/�c��agЫ��E8��c��y�?	�U�?��89�!�HB�Г4C��i\��-�	N�	������H��L(m�:ֺ�z� ��Ebl��?�P���H�9�?;vVJ�[�����?s�D�H'��jT�c���`�}�]\�֪}{� ��O��-#��M����]
�\J��D�_nK��(Om�O��<ߨ�4��5�����h?��t����O�x�y���Ap��+4LP�٩XB\��-�`wg��{�:���q>.�)�27T ڊ���)<׹%[\�y���>��F�O�ɐ��/ح�p�4|�.-Q�� ��1��ڴ
�N8g��������
W�Lc���z
��Td��3ari�Z�����Y*��~�Jb���Ĥ7W;�����b�+��(^���f�����c�!����ʽF4����^<������ZNG`�C�h����xi|Q�Z���=1`"^܇�%a��<�e<�~d��ԕ�z�
��׺�P�pO9*��Wy�~W��5��7�<nå ���C��5�����ͯ~�EF[�;��tX.���*�u�xɾ}�:D&Z�%�����M�w���+�c0L��t�UIi�Q��"����g�UeȦ!�W���-70�_�q��`��}
�8��i[��e��kX�Ƅ9��E��o�Jޅ���g�_��?i'|�f�Qz���?i��+�H�=�]��)���o^�h@z9 �/�I7i�C�r��8�X^��	����^�AH��X8��qʻ����i���s�!_=�����}4��\�i��W�6f2:T�ճ���>��;{`�S�IAgf��2�:������T��ȸ]Ч��]d�As�Aa��a�C��̀�)�}�7'�i�g7���7�{�5�Z�7�-�֍y-�0��ȟ���0K��V�ֲ�HؤI��&��@	N��)G���<� )�i4a$�/�	��q%����1��o���̺ʢ�X�^~��:wō�O9?�����q���o7��{f]?{ >�e�q�����6�#K��3���e�e��ϒ��9����/������WԎ��G?���n�� �p�ؚ̬*���k|���A��� a_c�h��b����6z�GǼ�!G}r��^淡TB(���t�
Ӟ�=_4��deZ ��{O!_Z����"����ְD�4Y��%P�~a�����M�]�tv�hۑ9p�rID�$W�0�.�ʁ���b7+�Y?��1�Y%\����g�ӈ��-�(Ǜ­ņG�T>�'0	�k��QA�׬rEaX�3J���NA��yL~��,�0C�gRS{F�eiֶ;h|�1�i���	�-Ii��p0���6����[�f�n\�'PW�}�4��/��N	��	�M��
�����S���]~=��[�W*9d���b�[d]��#7���Rrh� i?��~0_B����,ռʆ�W���S6�rn�S���"��)��b"�1��S���ߦ�s�ŷ8��<�/%��0nܶ�кʝH�Ӡ-,�d&M�g��t(p!ńq�>I+��8�|��Jy�(1i'�ܻ������ײR�(|��̂�r��"\�-��^�ׯ��	{��7�<���U6x��t�吁�Y���78��
�����1��o�{ĀK�.��v�:�=��1�t���q��z��%����,��̂y,K\l/���x�w__�g�����<�K}c�2)F}d9ʍ8e�+��<�5ħ-�A\��鵛qm��nG[|	�(Y����I��h�?yl3+W����VW�g!,���	n���s�=�Dޡ�"@2��>�Lq:@)�GBr���W:o�O|���/���J��u��O
��!Ӷ�ݡ탬��!�Gg�4�Տ�h] , �# ^�|����.rs���7��<��2!�:	�)�c�����J}�]�K� �e�o�*V�v�~�F;�x�pm�Q�,�[��c=�DRD�Ӟ�g����Q����<����X�����1&�)��z>z���D�8F�L���B���1@��b�J��:�>y��\a
\���	�d	[�T^�b|kƊ?�{fJX��H��ٓ�]��8���fM;a,Ż�sVNFc�[�-'KN�:����XvB�*(&�uM�ДD��<��hd�����������4$�I�_\xV8"0�/���*��J�O8��x 	�0Қ�k�`RL���>A����F���-�����2
#)i^o�8��e�������~��R6ܸ��B�P�D�Q�s��6�\ax�
���*�N�ǂ��C�������'�4n��Q�N���{g�Q�A�s���Ğ={J��2��N��|�G�� @8CK�#읛�yB�����S:��x�ϳt{�3��y/_L�ո}����y�C�|5|�cJ˔���϶G;���x'շ��h� r.q�YCżg�v�5���i�i�3aG:�c��1��%��ye~�2e�ߙ �^�1�\�y�)�T]��'��-'�H��7NMx���i�L�^S��3�z˺j�{C�^^e˂o?>|��R�ٷ.I:��
������A�o8�"o2�U�_�x4��O�M�s�a�syfע{ҖG��,��ܹݳQ�����"�n�����P����m�@��#3&+�5����������̸UV��&h��"2��:g�<�
��J/<�<i��^��~�t����z@Y�i�x���m�ʸ���@�uE�#r���@�(W�s�y�g��9�D����#%{�N�]'n�>?'��,	^�����>]��Z��eC��i�_x.���gB�!�ܑ$�3�@�n���4V��6���U2!v��#��lf�ɫ�-��0����&ixc]z,�G�d/1�3�a����gi2S�[�~6����+,K��-R� 
�*�( �L���I#-.l=
Q̃EI��P��;����
SA [dG<k�zEaс%;t���=l.a2B�ܝu���wt��:�<HJʘsEb0X8�.�<�C��T��g%�J?Q�EFpGw�G�|V��!N�Yy	H>��5i�0:��&��}N>����+-b%
&&<��"C�r�$��y�'����gs5��)#��2h�`g`c�O׬y��ۈ����ƭo[ҭ�>�|�Y�q�S��u-��b���ȫt*X7����G��;�o��gD��6���ExNf��<��������:�0��pF�?|���/��u�dCc_)]�<�@ȸ�>r"� %�MX9�mx�йM#=�k~ӶS7_�WE����[XF�<ɇ�ߡ"<J�v���A�(9d~h3KK%�4\�=�>a5$��a��{��a\�.�	�4:����|���ʴ�j��/9;%�xGa�3��S~��[�&|��˻�:q�6�����kݰ���D%����������52�p�gk���`b6>�pC0��7N}[:zlO�: �_�-}���dk8���L7k�(3?�].8
�V�߉+߷���5|�"/y&8�(��I��oxi�fN�p�=W���- �/:�	�4�)q���f�2	�C�J;e�*@Vi��q�LR_����TPa�]���e����O��9��[��j�3;��_`�]�/I=c9r�f�K�]��7O�s���&P�w��ס�'��+O��T��<�m#���?)B��6m����>Y_ 0���'64}����g�-2}�A�3����c�������7/7`�F��%'�s���_r�8�Pj$�`-3���8�K�����pߕ��,n�#�����p%X6R�|��
Bm�f�(ꈽ6,?�i�ڤ�|3ʥIq�buZ���09e	:'�ju3k�ѹ:��fq q*˼:+��&i(�������_�T�9I�$(�pf�W�$�j!A�8�#0��%�
Xệ�d* h^_�3��pR�q��#�o�@[�~���<`1��yAh���:mjb�i뭴�2�`�����>x��gS�?��n�N�E\�~��e@�[W1�hW�����rNXLQR����j$`��f�|��5K��~zҏ�2�����B�k �[o��Zh˞i�eh�)��##�U^H�s�la(�*����?n#���Y���"�堗� W�2�\y����P'�+o�_�JϾҲ\����L;~��X��w:,��*C_p0�0���0���4�y�Y��w��}g�|���|T������
߻�ǐ�<q���Ѵ7�>��tC�aCM��8�NtFJp���=�'�1�f��0j�W��C�e�q��z�fw������8��LzB{�=��0f�ԩG'��]vr��E��A��g�b|�{~��[ȬH���T�.�ST+�	V㔛�NhI;�I�SF�
fbc���Hp({��AH�k����K�E��`W�ܶ>�l&σ�ǩ&��b�3M�ӯ���B��7E��W�ʌ��}xV<		?�0�r&4|��b@����#/^�6I�ӜÏ}aC���a}4��L� ʶ{ި��W����6��r�S�_�����ͷ���W|O��oz$�e���	�[��5�ӕ�2��&����b�����91v�Bg[aI0t�@��=Z�N�ы��w��^�6r�$���c�L�������6�F���=��7����幛E�9\�U0�,=M�>Sd��dܥ[F;�g33o8��l��%�A&؋1���� �vl�vN�'��E�S�(�=���f�-
Ԏ��5kԑ�<R]�u^�?�AD���Z��|:$ʻ�S���O9��gX�á�5��ŷF��@D6���ӂs�GT>��l��EQw�G.u��2:b�����T��;#WW �)Y�-.P����vQ�31?O��6��v5�pS�C�nBJ/��"��m��0�)��9@�>D�;�|�o-�Rt��t
������e�\3Q^se�z�������p�S!+����P^2f��+ζ_V��#O�A��(��<��P�	qa��HZh0
'������O�W�ͼ -�F��IL�r��Y2�p�����l;��a���]�i�����C����UqӺ��+������14acH��X�4��,/	�D���I��8�M^�'��c�X��u�u�6����)�pݔ'��?�E߬L��|*v���|-C|i�'m�Ƒ�	O�MoYſu2a`8p
���-(O��?���e(E_�]K�r�M����+e
��q�0y�q&K�8h�Gg-N������3N��qc�M�+���w_�b�&��>�[���Цc�m�� ���b���&A�@~I��l��ge�� ��DJ�JТ/��ʼ0ŷ
[|��3	�7<Z�CM�:�u��_����Ls��ҷ�Տȫ��o���U�̄��W\���+�j����߫���K��x�cR<T\�qD�|G�9����ESՖg����r��^�7��i���|�+A\$1
d-m��<�� Z,����-~lܒ=`��3���0����\w��;�M;����P�g���:��; @�K0��F����V�~�ե�k6�k4��h0�A��uZ�v֧؃`�Q	��{�^�f�[ޔ���ҽ8ـ���M�Lo�0-��@�:B�L���/�)��G��d�S:�#_7�a����>�{^��y��
?��o6��ӎV�y���kig�aQ��Hl���Z���6��th��C�&N��PJd�oq�h|=[�����5 p�h������(0��('�e����D�@B�pMR~�k��W�3�,����Ԧ�[�w�>N9	����������̿�r>��͵��4&��F�|��㾁C�Gi�Z0��̿ƀzŲ�F�O5�i��q_@��q� ��p���#@Ҡ�o�,I�`��U����~����X%%�qS��S[�[g��E����6����W>>��n�-�y�𲳗*��0�"Ò���nZR�[�u�
<���������0�t�f��Nt3C�8�ƹ�i�f�#�uch	��-^�>Z�p�f�ʻ~g�t�ohZ�X[x^�u��+|��2eN:���,��Ѩ�&s�i�'�Z�8� u���S�r_�8���3��	��,M;�e�Qo����V_f=e82}�w6Mک3x�ۓ�{�L_�z̀����v�GX��,N˰͟�|n�?�c��_�"��x�Ih���KU�M¤�y�S��gx'ov����0��w)?~2����;X;(���G�����_V� �y��V��8"���ꍁ�3.:�W^�J>���/�Bs�����GA��ѶB�L��֏[���K{y���+���$�T���?�ɢ�O^l��O�����C���C�~��/0#v�L�ݧFY���n�'ʓ��훫��EV�V��:5��A�<�����<�|	!P�o���}����{��W��;`����[d���xY��>������~��S6O���O+�,�zN��MÏ6׼^�>��P-VRL&�.�
�LӤ�X])q���ۻ��sȹIL@� ���Ɛ�����v�z�jv������«�̃�&�m,Û7�[`s���S�_`�^�1�k:O7�R�p8ܖ��[��j���Cu�����|;�6me����3E���s�/����u?�lc��J'��`B��7�ezQ����7��q>7��O6�~9I3���\��p}�Y���;�ﲑ~r�r'd������`Q/�|���X9A���H��*�5H4J:{���/8悍�6e���c����y�z|��K��b�,�V�T�#�H �*��w�{*�7��(����H�I�����ȄY��ʀ�¨3,JP���"O��I��P���`��CM�2-��|�g���Sa�S�k�I1&��� H<C�$4�eq�a-�6���-��v�eLg��`ڙ��q^�+�0�ʒx���(����3����s���}zL#�u��rvFQ��,d���a�Lo��q�����K|]B��Y!H>u��8�)��cXD10�����;�0�N��#��7_��[��H@��'��9U�s���#a�1(v c�r0z���y�8QZ��r����o��ۘ��^�Є�9HN�{���*�<o �A����r@���i[����t�czq+����W��vp���F: 5`�-���{!�l��oԺ���j�C��*������ �^���4���#�����5���7	9=;����O?}�����C� ҈G���1�1�L�`�ҁ�2�~�'^��cm�Ѵq�P*l+��3��������{�����j�:`��9�
����E��4l��"U�=�S����..^�<�r��&]�Q���v-C�F����/�%S�z�<u��c�ğ�H��S1�$��&�x��:&��C@Y�:I'��Q�J3<�rB�s�[�б~���|F�%ƗUp���G_����9�ţ\͌��ƓƗ^+Qh0���%�̆�Aw�V���*���J���5$�_&���R${K����A�٤��%i	lY?k�%=){O��&�L�
����*��m��^��5{�.������"ѿ��b���6.�� ������rV�5��/����sF`~k�p���?eFԣ#<8RP�]6�" ~��%F�%#χGԩr��p�Y����v���%�x;�P|r�Ͱh5_R��>����U��/�%���̙����!#E�I��%?  '�ԁ�qD���E�mWc,�|��[�0����k���mI]�W�e�C�+��5\c�=Yn��.g���2�:�2^g~��8�ޱ��c^aIC�M�1_���,?T��#i-NQ��(����7�#.>[�����:����9^�%d��5F�i�����i�6��O�'~�X�~��q=�\	�9��s�l��u6��1�+_�)զ?`�SxF�'}e�G����Ge*�"�����3�~A{�����/"�a�z�K�r9���t�6���z.-���v.!�F'��7>��XKN�˲���&�DI����)u�+�/�Z�~��ه��{n�==V��K�5�����ǅ[h����l�\{��q���Q�׭Q��˗�	su��s��{=R�s�l^w�,�Q�V����4Z�wMԋ�.G���?Ğ8F�U��3l���'������2���分�>ũ��a�@p���[�ez�Zlʎ-c!\��S�$�k���Ĉ"�m�H#��L�a�!�1��1e�S��x�+_�g�����T2y��oY��:�Kd1H����r��YU�����9���+��6����Op�@K�,G>�z�+��_���g|@����x��6:Ox?Ā|�+\e�B>�s��5�ҩ�Y;�:C��+(V�|���-cZ�<k���-����҅����Q�N�k�q�z`Ɩy�fj4�n��r<n�/�LT�2I������(l��$�٦��ᗠH���.�����l!�ɥ�TRa��em�a<�V���7ԽˌO�����2������1h=h� w@s`��b�Q�tj>��Q��� ��PG���������{�������O�8�i����Tv�⣛4�B�p��G�
�J�S�٨�B0�6l��@J�l6���9kPV�	ǭ4 ���G�LG��%P���m+q�	@�ᚴ.[�Ԕ+�d'˝p��1-�� \y'^�5��1�̫�t֍u��'�1���mz/�BE:���k�οnܾ�?�T�?�D�/��W�Ieo}-�st  @ IDAT����L���1�p�5����ǰrU���Qy�=q�6��Z&\�}D�hK�uU?��׎Op��������/�7��`���>�f�����N
�a� )�N>'�	��Ji�oJ�ֻ� U͵���]h���$f�:�A�0g��+a�1�� ��3�/�'�#_��M�y���8[�<������L�02�B5oK��c�I�ʡ�8t�F��~\^��:�l�����LW��h�3f�;~�gg�����Y������+f�<w�3<G�V>J���b+��_D�v)�_�O{Wv�.��o�P�C�t$g�s�dUf�4��i�ȺMD�@���5Dt/��	�<�-��@�lh&:as�-@<����������F����5���4�z�L�PZ�u�Z*#JЪ<��$��(1N���P��i�aT�� �X�иz�>����b�yP�{��4��'���wz��b=�K:@�{�N��^B�&�O#,]F��ª�2S�:�I}h�����JR��SE%_T`^��l˵�$�G��%˥Ё�B|��yB�w#'�����S�N��^^Y�"솏��k��jǄ\��
V���������Th�wO�|Tx�wa�;��YJ;T�����S�ǅ����1��bH�J�2��@;�c�K!�C�,֙�?�� ���:���x�c�1;���fU�>wÓ�� E7N:�G���Gˋ��xӑ�0�yH�s�ӀR�ЖT�il���M�օ3~0<o��n���y���� ܰά0hX[ĻuX����*聒��l��P�姸��V��|֙~��F^��z��K�n�-ď����3|^:;6F��7�K�3��mY�}�˰(�_�1�sʕ�S���_�q��f���̕r~$x��1��տ��	ø�Q����iۋK��)5ͤ���s��R��q��PL��J�;\$���Sv�.�,?�c����6�s�����r����Wꕳ�M�4��ƚ�k�>�+;�����Y�0�2�1Tms�G��m���������q�8�܄նyV�� %��2z���\��#�q��ƥh��7�����MyT�z(�}�%Wu,�t�1W�0G^�%��*r᠐Ze���O���l�(��줌/y�C�!<Np��]���l3�y
_H�6$aʏ2�,��;��Qѣ�W��RG�<@ǃ �*ޗ��SJ�/���EF�a����`�1��H93xB�
M�	��-�~q����F��v��K0'mb���-3N�dp	�P�4�6f��a*/�Ӏt��dv�!�:���b��#t2�N��%Sf2�l�&Nq�T�
�
�
{�����؈M!�;02R�SW	P����K�6˷�x�H�i��;w�x���Cʸ��AOI���
�H���
�0���;a	%��&��S.�����א�M��¬=�齖�f�(]�`qo�m꽘��RL+���&�+t�[�I��#šp��#u�௿�Ӹ�2&�O���f���DR#���7�|7D�&�����$�t�Q��(j���B�̚Ldnq�23T���^���z��|k��ѓ��޶}8�Rg�?[7�ǩ��8�-�$U�5�|3ӳ�$��
?a��d��ж�~�Y|�"�>gŤër�mg��<�9���#r�a��@yO��S�����*����n�.v,���'z�Io6�z��Y���q5�l��=�ŉ�k[��y�K�,�P'��6��c��0Mc����n���^���R�I?q�c�g�1&�<ioҪ~�޵)3�2g���7�Ҭ�Uv�����i�����4Ts�_m;7�՗�~�����t{FX^���Y��$~v����Ù�:� ���7�VD����^�� i�yZI�8��i��Rv"�«��V�$0q�|\�@c�$�,���_���Eְ�9	�w?�Y�XFL��W�Ջ����
_��?���36�0Q������ �E_�E�Z��-��-�v���4)�s�$�|!�Yt��	�����!��`�"ƈ���֙#2�B$�wY�C�Z.`a��j���^�O�	L�G�=�+ļ���
V�F�apQ6��=Ub���G�1�2���OhY慢 \�^m�w����~���={��L p�O��#g�:��b���ѵ�[��#��ظ��yè�I!�
�B�Zn�	U;e�IWL�Ya��,A�4:�(�y&�3`6>�X����-hqz�8�ё�t����2k��7��\��#ъܝ��쉆�:ʡ��|PyZ���蕆�*����	�xP8Q�Ж��#S �{5��.=G�N�4���%L�n��#y1F�r5j�8nE|/���
�`2�>����<Ɨ�o�pr���I�3���_�4��ȡ��|f�:�k4I�vLy��:�B��t4���ұ!!⹜?䜚;$�6".�xf���G��hP���b~$3��� �F�P)*�Sf��a����k��Y�gG6�	��5V�Tm+�H崝}�[\P��߀Q����^ӻ�*>��㌛#>g��z"5xL��T�\j\\!�17�ov�$�O��?Gӻ3h>+�12�@��?�d}w�8�RW�R�АN:#p��i�����6�,��<����WN�����f+2����m:˷��4Z�N!Ӿ��|�vҖH�}�
kA�/㽦\�x@@.�u��8�߇��\#�e@Bҕ�@�gW��:@���\�8�;�����<�-3�i�	/aY����Q���S.�x�_+mۺ�~d]Q�������sɎO�!e���ˍ�ѱ�� oG�aeP�I0���7^�C�9dAC�j�8c5�f��bt����o�~�`B�b�%��r�-�-�S/)<)���/���Hn��.A�X�n��6����<Q���
�|���w`G�|+8�-�k�� qѧ��h�R���m[H�\����Ǜ���n'Bп��R׷��@6��Ծ�y��`5��_�����z]�I	��r<%��dW�,��M}�wq��`���٬|�ǒ���K�4I���EF�(\��j�ۇ�G=XL��B���7_��7�|m�U|� M��c�U��f�nnT���$g�(��qtre�FZ��{>j��l����B(�iP<ddKD�%-D�lQ��|�W ̀�s,�	��.�T�
(����Y�2Z�S�ԩ`��Yg�~�I��,K^�A���9Q~-Y��a.
E�+e���&u�Y���	
��|�Ε.��q)UVdd� �7K�Yz��Y� s�eɞ��J*(�d����`�̶ �#x�!�a(L����������_��h��K�b��.B��5�^�|�۞�ّ��\y�������� a��l8��-?uoan�Lc�g�X7��5��rΐ��и��Q�@��X8�\��Ɋ܄���ǲ�W�L��{o��,ـ�;K{�X}s��}f�X�ޤ3�>�rФ�8��K2�ªIZ����Oy��^p/��[q��#g�p�3��-L0�i;�=�q�Ǝ��b��G��<�o�1 y���C?9��gÍ��QxG��9d���7�x�af7Js�w���|��g�R�S�a��f��g<�Ã���48}2��j�n��#��~��z�3�1�V�5�w8	cg4���Ӟ-M7�����k�̣�D�y�y/�m��0���e񠰄S�����`ˏ��q��}��8���/�����2�-_J���O�<������Ů�ny#Ȗu�2�w��:�/��L��z�/��.���8� n˖_�\�L�.U8�.8Xs%Ԏ�Γ;Q��+�$]��` ����k��'~��n�$n֕���J���4!���ؕk!Ҥ�֧�'��\�˛x�P��v�&P8��O�\3@���~]��l�I����.iI)����-M\ԣԙ�hQ���[m��s��37�n(�
yu�I6þ��=ߠ������KuP6��Rs�����@v`���$�e��W�y�Dq�;�>jl�/�Dw�Ft�a�q�Y�O��qO��z�ǖ�je������[0�MwM,��[#�e���['��Q���0��1�ҴȮrH�1�;l\�p4�t�a�:���ʡj����k-�0��]�>�Ip��'�3��{��#QB62޼��%8�.��CA:�;i��:,�a�/��8�>L�X�2s��u�y�ۑ������x�)�<��^?k`Gs��hGL�HM� p�-h����
ؠ�a�6(��ȭBT�<���0�8+]C��%I�����4�:�i�^{W)�����D��y����L#�h�5}����'x�Z­E���������R-/�<���B����T8�.sx��ߚK����i-pR����-;(��Te��f��Է'l���O��k;�D��P�,G����t	�"�#gI�����J�����=>���g�p��'��R�?�3s�@���G^�����ΔZXn�:޹�����M�ֳ�� ���i|˿�!x�7�3^�#Whݫ�"��^��S�Z�m�%�⊜��4L� 3\,����0�PC���r�1�愶��_"ۙ���l�
������5�O�i;ޖ!��a�ď�S/�S��Wq����@0r�Ѳo����e��3�,�x�������ǁc�ɫqd��������g���~y]~�@%I�cY`L'�2^�ʿg}�E|���'��K���4\�1������w����������_Sv��=�0�'�୶?��/�����o�]�o?猣|��Rl1�v��3�98\EęU�v� ��44�Pzd���vKq~�zs@�A�Ȍ�[�Y��O�o�4ʇ�g$�0���8#��z�ᅤ*��T�b��������H��*`'i�ZI���w/|����[w��y�ʻ��K�^#=8��w���o8���-�����Ke���U��@f
�K��_��z�x�(�N\yz�C�2�񞉍w9s�����Vl�,�_5|����<d���r�I��fReX�~4��?�hFj�e.��5�r��K~��(yE; C~&?i��a���f �uav��i^�+n��l�0�' �;��k�FU����y`������Q:};S�L�]kՒ�V��+�@]b�h�9�sse�R������l輗);A� a�(�*�a�"�r�/�ۨ�a�!��_*�p�?��<��0!d�C��R�Fؿ��ϱ���ͧ��A�U][��/��0:�w�{P!���)��[��ۉ�N��N�.t�2���|ү0�F�)�����.��M�*2��
�
�Y�ܩt�n�2�����"dy�|rw���1���J��*I�W𖡛t�o8�����+G�t��1x�|q�(�_U����P çDXL.hd:5�Z�*_�t
�}�y6�~��(<��'\�?d���~����:��`����;�l,��T���S��|�����5�6��	G�ؑy`�#tF�����ӟ����?��v�9N;�z7�p�&E�G�]�+��u��?*Qg����f�l�w�q�"u��8+��m�&>>��� �vb��1�]�Ҷ�\���9Q�{��-Nm�c�E�#�ޓn���[�	�k�ӝX�#�M��g�����ĭ��Nb���5�ܥM:5�&��'�|����|:�u�����&<��ƙ�3���3 ��'x��S��r-gp�4�T\4�./}�Zݴ��/ܑ/e��Lp�)�8h���6���}|��sfP,[�>����1��z��߂|��Y	�/�١���t�2���/�^0����s�����3�q0��w��>��+d�r2 w�P�9[�1�,��:u���W�U7�� ��kG�����啳����~d��	P�^�n.�[7e'�	u&�x�����y\H� �G��� ��Ҫl$�֑��f;?�1�+�������)��FX��3ڨ��=.ľ�R���K����c�̚�l_�p���[1��\s�"��3�2�ň֖W䑖w�|NИ|�A�R���6HN9pR�2���7�����l�� ����Wu��T�h^a���O* طR�a�ѓ�)-�b}����$����7���岼K���5�0#|����{�&p*Rb\[5�C;�4:):G�׷�Φ�7l��kN�� ��\d�:��-C"<4Ĝ6N9�ᣒV�M����1\&�`
[k:밾�H���<`25���;�u hNgzd��Nx�k_pF����k������?�f�__p�}2̄3R��	�=KJB��9 ��O�VFZ�F�ޙ�J�/��hT<�0:�|��e�$DAW� |hYQb�S����
�#(�sP��޽t
�(`�h#HZb�Q���l���(�;"�6�����![��H�Gy��@4}������/B�c���92D�$W. �`c�s��n���Iy�w�	�8�1!W���`R:#����w�}�y��)�}��+��rz����C��+u�Q�ԫ�B;�-�Q��ڱh�m6_<z��O��������O0Ȏ6���l������i��2Ҵ�>����1?�3;��[�2�<l�ʳ~ɰNxH�ү��O�:!^���_���N;��NHO���/3_�7bԛ��<7�Ɨ'��ي��(.i�"�#�ڷ޳��l|K;�.p��"���5�K�����ӑ��.�$Tf�&Ot�`ؤθ�rD����4����2�\�����|n�i�I�h�r�?���!��^�~��ҍ������<�7�s�g�ɧ�8��<�*cV��V����ن�o�]�2�e�C�[����{����z �kF�6��,��8�����d���s>s�`����i��5�Ϋ}�оU�a�=.��<�9sO&�}i����3(���>�RxD���JD��!��*�Md�L=�*����G���Su��W�ؾ��>*\"�~�B���1��Odi�|��\d��Bi�-�C91�[�zp���	PU��J�8R
�#�P�>j�Z�Cv�۱�*\i�������|��>Yٿ��Q�ٻ��F�a��Ҁ>:$T^��8m.}*���B�s����qT�L�m1�|����mI//0���dF;��|!Z��A�BO�D�|�7x�/	���qB.���L����=Oe�ϫM5�}��+'��F�)�1��xv�$y���F�å%a�'ܣ_q�Kc���eti[i����*@�.:2�K!�z�frXv��/�ݷ8�C�}����Hh��ک�s���`H�3B
�HW0INʟ©��X
q��ȿUD8�8��u��mF��&7�ޙ�F����i��';�K?���/ן}�����r�[����7X��r$��Pj;(;�Lg��E�A��[$%,w�3�^H+��oc��3�*�v��$L�_1�F��g��0�&w��ǥߨ��X�g= X^��qϬ�8��8��hgj���f;z�(b�)0��T���3��2�Rw�Q����%�tǔ������*���\J����N:�0F0ʎu� �}�;�%]X�6,a���������\6y���[�6�9��ԓ�ƀԅo�o�*��5��ю��7�UV�������-f��<S�h�3_~�%{g>���UTm��=F��ܵ�&#)7�D��>YL��x��g_.G�����G�S\��-^�p�b����k\���0���X)~pٱ-�y�>P�p�g��Rr�g ��J�Y(h�7��$�؏7�&^�� ��3��`�a\�h�F�ǈ0�񦟻a��U��e}�+�LP���a����s?�M^\q|3������4�l�c��G8���9�4]�<uuɇ�MGО~�7��y�/|�0?�q��?�s��g�tIv��~ÞJ����r�FE��z!�8��x����%HZn�	���}q � Ɓ��Y�W���7Zt�o/2x�S4��Y>c�F��H��D},-������[F8(�ʼ8+�y�$y���N����� ��8>�O;�'EE7�����/Y�<�zW?���k��oX��O�ÉYw	�z�i�CS�/�����r"�chrw�g;zG��$��{��7�^9�EF+N��6q��1���6�����a�L���q�=2���E���G���9���94�-�DD��+��Q� �چ�=ˑ��k��E��Փ��j�ҹ��xX�#�\ew��뽼mH��Dˍ�YAF5��7�Wf`s��^P�Od4g�� �΄mD�N���w1��;/
Z�0h/Ca�uF�«�u�~>½y� STP>����1�سu�A��->E*H�<�Ԣ��sx��%/'TΐA20{�8��#����}�zgH�����H��)c+'iҁ�lc����c�byzv����������?��cv��-�)ʱt��)ShȀ�茑�P;����#�ħa�}�}�4�x�x�6�o��48ff�}.6����nd|w�lR�i�*27��<O'�{)����Ox���*	�s��ө�5a�$)���uw���պ��7p:������3G�Ov�����y�t�y�.���л��v�(�7��d�b�t��-��z��y�R����x���9:��8d��#IN=��{���)�9�;�lʃo_e �߻w���t =������0����ٳ̾��@������h]{�ڍ�X%�,�RpI��^Gb+r@�wx�ՙ�:�dh[>��v�]x�+˰����NÙXgyb�kx�� p�4��*>�gh W;��-,GW�}HrA�Zk���Ӹ���N.�v�	/�����Y�#������8����]��+�Ԋ3���C�8����r�~y!�l[��oZ�錷����s�=0װ��
����o�L:��
O��N>�
;^��û�C��&�4�H��ozq���La��wJ�����%�YJW��<������,5=g�c�s�2+m�io0Ag9���_�/�z��`��=�ΐ�F)�a��B�׿�������'��>���}�o�_Ő�A�A�1��.�A�T�5Z�I���g.gy\��qmƶ��C�Wu��9��Ph��:f�t@h��"�P��W�����a�V�-w�hoZ7r*0��:����iSn\�:g@����v�,��óS�8����yxtM�����'2�w���m:�S���|�m�i#�w*~P����O��E|�����݇�w�ˑlG�u�r)���ş���Cgì��f�y|�	q�`��GVm�4+�|��a�k��S����Zd�l�4���}� ��%h�?a��#��ˏ�Ґ����wEn���LҺ�%{�G���vx� {� ��e���� ��C�9�N�9����ێ����DM�[x�����,¬򶑪d�$B���)���H�!kW�D�U�0�p
����d��ă���3�;=�����շ����u�)���F2�C![4�Wy	ߎ�ƪ��v@�x N�m�ĦR�<7��C7r�t�B�Ғ���2�lҚ��Q����A�a�zъV9Q���U���?�{G��u*����zF�"E�(߭���|�s`	Oځ����x2s%�K�M��o��0Gi^*y�9;�a�'��t`��-o��n�%-��L/�Qx~�+>�QD=|��a��/
�oi���eq�����8r=>�İ�ᰊ��c��@.m��!tz��)��y}� �ۢ�����4�������S��b������a=��63vʧ�[�X-x�W��)Ox(׀�R���_��s9*ƪ�3��3Di�#w��V`;��=��uF��Q�Lf��(������Y
�Bˊ�H��C���i�(W��IyQF�O���/��[��#�cb"��`��Qa|-�p�4�n��8˘�v��O��)�W�xn���I��ؿ�'<��I�Wa�@4��p��ׯa��qѓ� �y�������?�~ʔQ0�4�˪�Nl�I��y:v�gT��4:���o��ټ|y�y��S��ki���"�Q�k���Z�"��%��hп�46���C�3~��"F�	��3�QvL���ċ�/6�h_�0�������bI�'m�r�7u�}��'ԥTg���Ȓ�'g�Q:R;Ju�Ƹ��1����=;�P���[�,��9�Z����7�?e��:�3����g~��5���2��s6�ιG>$~;��e��K�����MG����� %ϕ3eU?|g��@�K8�^�M����[�6���y�N�EHN}?����]Q[tWȢrg!�[��<X�X^�y��p]��Y_����\;���� ��7���#��]M�8k��[�R%� ��8�!�| �Ě����럹�W@�-p?�D"���5�.�P-��u��-6���X�("�k� Cm�G;4����"*$�n�T �L:�\��{*?	�8GV�B�]���1��l��'M6>��@����C�!Brz�*yc�s�n5��yXzw`�N)�X��4�����F�HBN���c��l|��jX�o��ܿppl#ng唹o��x�7�o٠�e@H���*��^W��=<��1�2�+O56\;wD�l#bKðq�zx�=���kDA+�Dd���Q��:ة�i��\�W=�E^M�R���v(e;Rt�5��Q�̌YV�H��O�`��r`�p������=s*L��}%��,7��e��%�U��%�J�`
��+>?�+�G���,a�᭯�{�h�W��;�a���/�剗���9����<c��o��[�݌//i(E7��f)�g;`�(���P[VI�"�H1\g�i0Pԉ�F���Ef�!pug
�_5��ޞF�o�T����ٍ��wFg��e�&B�Lqb��6eǩt�QQ�.�w)�ـN�_i޵ogx�&l�U@�נ���gg(\=�vf�6-l�5�H-�*TO��u���^e�x�R��bh�)���7lw�Q\��s���!��.�tyJE��a\ۉx�x��F�gX9�����|�-j x�v�E�LS%ݎSx�=N�:y�Rϸy����z�_��MX��*��wp#^ܤG���3��lxp�o�9�9�]Y�'�?��!uo�0�V>*�ֽ"�~�nlߝEG���Pգ`�U��:XDV��_4t<�ӽY����:z�^��<t��$KV�r���<�Q~)��m��s_/��Y#C�\P�o1\��J�{���*ɑ��z��;��cy�U�	�=����+u�����3+��[eJg^�@��ʣ��|�N�q=�d��:�!T�0�|�~=�wIA�bջY$1o�����߾1�<�<t�W*1>R�J �ge�S.�4����-��Y�l�.��KW�H�D���)����5�a��.�"-R �p��i�䷍Yu�O0��	��^�N�*T�[H` W�������K9�w�i\ ��g@��4�oB�u&>�	<B	�K̘6*&���� �CS�-D^�E�Ë�ٛ*?���1&��*G��T��	�
I�b�)�*L�f����xiV���I'�<�H��Ί�8+�r�K�����/iMO�TS*�
ѲFP};���s6f��<��Fs�ޠ�^(�4fᙗ��6�T��aO��PS�<;r��8y`@���QB"O^QV92�(�*)R*Y���X5�F�T�!V&�|;+��2�@[G��"���bN��]!��)��I<D1аT�1�ds4-qȀ��s�s�	�+�S4�o(1�0015I�<a߀�[�pT:�i|ppui�cOJ3_t�X1�Xj����B����6y���/$a�Dv��<��o%B��FÉq��0`D���umr
�;K2^��Ӿdi���U��e7��؉��8�fK=�C��K�����0��K8�i�:��ҐK�`Q�& ff0Q�~�E#P���;��s_���5Q�N�q@[
K�ʮ�%�5N��6Ki��t0�tt�9�.:��N8�+���[����v��,��|>ﻌ����!%Q��	�� �����	O{NZW궕<�:{8��|��(C\w`�c��+c�4��+��<�*#���j�jͥM�4�e({�=Ï�;�� >Mt�m��>��"��Y'���e&���0�5t���<.Uwc5KL������@Z�ۑ�Q��s���'��W�	�hQ~�� 3��A䠙=X���K��o�/�"q���7ܥ9�B�.s�[$���̜d�3s |b?��Vg�a��;a�ڣ�4��Š�_Tx�ЁAp5���	�R�Jf��笘%+�i/�6e�.5ƼZ7ց8��3$�@`���}P���S�WW�LҎ��/0��5�r���@U�<���mg�����#�\�MK'u�x��ҭB�&˦�#�����}�M�ʀ���c����ҟ�o��~eb��L�:ɯaJZ	�y�� qw�L AP�\�Gn|��Pg~�}�7%�Sl��+ρg� ��т�ʛ�,'�%��_:)���tX����`'b�t���s �Md��Θ�W���0Tpn] P�dC�P�[�@�t	�@��T�~�����I a��ݳ����5<Nf+��s�'F`�9�e�6�?��B�����;�R�|�U��:#�����b�b,�hC�	%ܺAÀ �N�9���V:��5o!> ���G�W!�`Bg�P6Y�#��s�����"��SH��!�k�̼1�r�C�D��ƈ����de�A&OT�c�ո���3y�'�2���o:+��u����5<��G0��(,�G�-�廜t@'(�c�pp��NDe�[w};��@yr���%�tT@���rˑ
��4|d�Qݽ��!y�]Q�B%r�U�E�t�����P����4NF�4�Q�(�S�?����,E�z}����!
^�@P�H�-I�0P�<�B�rM�".�x���� @�	']�#�4��sv�h0qp&F��6j�c�v��3�˴���w�N�{�
a��,��R�޺���0���1a](o*��x�������;� ��rk�	�|�>���>a��/��'e�fk|�������ɫ��򕳈�-�<lÛ��N��Ik��0�#��/�ݺ��x۫��^ۑ�<�[�C�L�����o�1�B�_u�&
.�_3I⚍��5�p�������4�r�NI��p��j{�>� )��(�3��j����v�4ִ5i���ap��wpu����{�Q�>�ޫ̤��o=� �d����I�aٿ��=[�15b��[�5��9�]'������G_$<F�,��\a@0Z��ZW���X�����cg�䙙���~ ��%��Hg�#+�vF�ȆsTw���<�HR�8�-�[̾�v=�l���t�����K��P�·mN�8����@
j�}��;o�sA����%�h��� �����Gt��8y-��xt�Ç�%N/�� �U��D��:����ma�g�/��Ɖϔ���7 I�w+8���7�4�O��@<W���	�w`ʅ�ZW��e�EQBn&����s� �Y�K�>ԂW�!����XA+�:!.���;�
�k�h�D���sx[2�<\��o�;���	FvG@c�f���?>A�8��A��6��n��y�/>����P�O!v��50$lH��ˌ$}M6�
�x���<I7� !3W���UZ )Y���H�m��״�E�?�PZ�����G#��5��e��� !��WA�'ql��όR_��k���]�I/͞2o3����/�gxKzZ&��7:ʃ �C!����F<����Y8�*O����o�I��+)�l����m.E�9�G�\z�ꙣ�c��n:MFe*#��/p��|*y;5h����|�A��;%	8:��l=8���y{��ǀO��N�@�K�����E��v��w�u;�}��CI:���V�کa����>e�|�n��u�/����_ͧ"���^�&&RUw��NCX���G��x���㌜H���Ȅ�~;��2$��_�����5����������&�����0�|� Q�LǷ�g:ydϳI�[��j�����[�b�<\|����+nI�Ϥ�\���C��N�C�<�#�D���� w�n�)^���\�-�����(�LC��j�F}�S���|FX��Ի��l�A4X(�g��w�=\g)�0�33斏L�(�S�5����=�Xk�;e��Ç��gݪ�k��E{GO9u�>�O���>�?տ7^w�����%=f$�s���ͧ����_a��R�y�)xY/��V��ꫡ��,�����쬞��u���)�W�bH�C��,�`�1��1�"S�.=�a��֠oH�Z�Ϸ��r�x�҃F�����ejx���K�왳���4��DXD{'����Ϻ�^���1{6O��i֏fE��	����K\S��/UNx[RӪ?K�m�
���{�ĳ�$�1�=��$��T�� RM�����HR+9�S��1]"V�ᠥ�]"�Ʒ��s�|�nf�&2�����t�"��(�@��*y�œa]~�c�1<R�@q�+��4���}�3,!�Ҋ�R��o��W���!�XM������°+�������l%�+��#������?�ǿ�|��G��qF��lM'����:9g��pf��su�w(ˆ��jy�����XV� �D���q�f5^�uv(K��gC�	�ӎ��r3��M�Qp��j�]~VԠ���o7�s#'x���UvPv�4�=�j�����@;�+���XLVD��)3��"��Kן�]r$	~�A����Q��L�G\�������R93�]ݬ@������ěY%*2�=�涹����Gt�b^�~};7;��_��s0����O����^���h��fj]䘪'c�����;9_���p�;�ۚy�����}y�!7t��̋�Ąfz̸鄻��X�@��u?[Q3����O*��k�ʬ���8H�xрm1�3��=�md�]�0��܋r�1���_���ơ�7��G�#剦5��(�H�i�Y�vv
ȁ�uLg�O�!�.���J�V�Gǎn��pT����'�3@/�:����S��9:��+��8s�Pe��A�/����ٳ�m��O[��^p��|�{�����Y�N:]+w���=���pp�>k,+�<��֮t�Ҝ����G�C��x��8��r�z��g`jw��p��f�����\^���g�I_����f����7m���'JL�����d���e�j��G��D����8*7z��No	�i��VN5�7�GN±u���m����i�g�]iͧ}�f=-�B����S�����=k�A��E�p���F��o
��~��ɘ���}�S6���%��q��{9����q9��"����-�`g~9��y+/m'�J~��z#��G�t��qr�p��+'�snK=���x^R��9x�{��ڵ��k������������us�+���5{�(�ƨ��+�*�K$�WYf�a�������Uh_/��=N�V���%�2~�	�}�cz�Q���d�7hR���uO�9�t��g<�~�������O 	h���`ͺ��I�x^��4Y���UýBO���>9�	�,����L���-.���)&�c��x��2D�Po�Ǩ$�:]
1��)3�(XؒΗS��Q�Et�s,�Cx�̹�Xp�_�\�~�z�{��o�W��B㔬����X��z竿�cz�����~��&r��{5�:Q�W��s�=i�f�z�;�<�: �U�}��4��zIhq����°'�A{-�0S�۷7{�2k���|�(	�'5k���䭝��̐�Fگ���sHyu��ؤ��I�_�R
U9�Tg������:O��K��b艠�$/cX#5�������sDQӈ8ZBn��YE�N����h�?�dMT31��W���m��駟������{��oQ~�hgP��Hl��:�}�����C��)�+Q��=�y�5��+u��1�ŠƷ��ּq�Ffь&<��;�pJsvY��k�����4r��>��td)G9���d:0��R�y�� #  @ IDAT	'z�I��砄�����J���\���>9ӇՉuH9�$�S��&@��5�4�H�X8ԡ�q�k�<�Ì�uT��zv�ެ�Y8:'Q�u�N8:��o�4��.���`�PX�J��<Ҏ�Ó�`�}8`Y�V��|�/\|�:�.{�w��g���n���p��.y��e�F����W��̷O���\��}�ZK�^�ܓ�Om5��O���%�P�gM�H����]�xh���}������"2���U�9\�)�%�&��a�/gdk9�^1�;��x���w�74x�z�^kͳ� ���2CƱa��,�c�0��<��vr.~zh�[���^����6o�^��7�E��g����d�V�*=��^�^���Eo�7��G��^ۮ�vɉA_���@O�[��O/�ة�R/��t�ʙ�mJ״�%E��J�Q��^g�Ǡ��]?5X_z���ޅ�y8��\�����Q�7�\�fk������٦@� ����to����_���|~��G�S}ݖ�`N?5y�]O�:��I<jv7��ΦP��yv��hp�;�샻���s�;�;���gz���cѬh\�YOδ�50�PR0����N�����`-��I����{�ŋI`@C$Ϣ{�Q������+�O���n繎_�	�7�=M��tU�?aDs���O�s��ѿ>}��jL7Owq߸s/ƶGO;�����rhz� S��&��|�(m�1]�i�C6ȳMC��X��wx1#ʘ��]0��ٯeBo�v��N�sdr�tb�S��6�T~:����ߒ@I:��W���";��ȁJ�ð��3gޯ�zP�����5�rL�%:�rd��mR>�n��@��>ݣ��2���٨N����)�5�����\K�9�댈'"�:�ւ�����%�Q|�!C�C��� ���`3h���cD�W�5Nq��<h��zu�h���%�]�nݛ�0-]�D�8�u[=�:�P[y��������>���c�~N�������_W���ȯ�8�ވ�A���:"\o;`�G��2e�~x֩lf#^:'Fw�"Yr���X�QgxY��	��ˠb���!�T��CS��z�+��i�-�t��Ћw�}:p8�0�'�q|��m܏�.�=?���q�o�����f�g�����Y%�����3hﹼC���c��p����ﵫ���$/���hv@d�F��q����.����`u�q��[��kk�x!j�djj"�!2��+����� �I�N@��C�[�BM�8��8:�'-,�mK;��e��������,�xp�V9��W��b�Z&���8?+��^=�g]�}x��x���M�����Qk�o4��n~س��K��7sَx�_�h�[�hi;k����h��8[���m�Z�20R�����%�R��]��� ��C&x��h�S�{�i?�Y�r���ɟ#�sن㵶����q����Oy+���e��<ܞw�'��\9s7o����[�Ӷ;�������5�v�5�����"p�ݝ6Ay��K�ηs�iR�c���EBBݵ�q��G����"wh��n����0g?�W'��8m��vF�>8�c���9e�_ ��q���p&���T��9Ø�iF����{6�P,�@
/p�ո.�m�&ғ�U#q2�o�a��^��2x�1��Y��pJ�i����br���0Ω�����g��	�S��[P�\%�<K�6Z��_~zz���������d['SCx�V?=y��' S����ߔ���>�:X���&��Y�ݛ�;]����@E[c�:7����m!P_�;�el헲LN�>ǚ�q68=�+J�?���zB�{lv�{C2r:kS�1]��|���t�W��r�*�<]�^���|�L����6�Y�-�$o6�7ы~�áF�:�th�0�<�e7�G�鍨K�6��}���f�L�	�����񺷷��w�u+-@x�F��::1i!S)�|���3|Y}F�����B������[9�C�z���x�x���5�ț�a2Y�=�R���n+X�c���໏�p%_�8��E3����1M���}D���)��d�Y�i�~�����"������%��}#��2�U�=g6��!m�B|\�KE����ш���D$�ع�o�����T���;�����1�oih<�ɇ��N�v32X��k��gx��۴���iXOy�����m�=��u�+p���(+���W�h����r-�m�Wnm�gce����.u���%����;u��i�w��-��t�;��q�0��b�K�r�g9Em�~<���-A6�n<j)��^������^�k��Z2q��0v�V0t���൛/g�糖/<o��E���y�,(�>��^1GM�o6����_���ӟ�����P���7�������-:gWf�6v�mZ����D��ٌ���� �c����r����T�A�U���6pFxx���#z��eN��ͮ=�lQ)��V���Aqm��A����z��������|�{��8Qn��RM/
�we�_ρ��4rӱ�1����s�Q��}������2zؖ4�^����hM���<�������M�r~��L[���SV��iN=��k���H��mm)@�����NJ�uW�R���y�j�����^r�‛?��ӡ��8�u}�L%!'cDqh�	OXc��k���~'�S���=0W��0[D6�
\�93���$���sfj	҆���]G�r`�2�@���?�=�3I�[�+�:��A�sz��Q��!n|Y���o�}|��"}�z��I���I��w%�
,z���mS�3^�����F�w���V��ܹ}sxv�����x#���I1v���/��E�P��ְ޿�Ti�в�6��MJ���>��\�D0�ã'�_�/���z.V�Ck�6��-�~?_D�A�rp����ZSq����D�ZU#����ȡh�Fp?���h�� Xt��O�,��HҮط�[���h��duWo�Z�Y���;��+
�^�8��� �aG��U�:?#oN�Q��F��O�F�C?����8C�t͵�x�4ǻ}�g�|p������a4��w�뻐��A���na�/J���0�qVM�k�dDI�ֻ�5����q�
�X�{����c�ǘ'��6�F����2��_���C���֚�T8^>Os�߀͈|���DZ<�]�cx��я��"��E�����9@�L��N�
�n������E�x;�e�m�s�qp��L�8�)/<w�8�����haz�q��:Vl��2Ҏ�`k[�z`��<���'�ql/��`��{e\�(�Q~}W���Յ�Kt��pr�ə��w�K*���G���l��k����b�t:���L��p�E�M�Ygt.����;u�:���x�+��	��o��C�К�V�~���{��������e�� �C��P޽{�z��۾m�ܠ�ru���fkmW�1�{�U��~x��o&^�~��O������k1�����=뛭,�x>��Mī>0��xr'}��"a>"~�\�����j60�cKk����w��O�]��o|�;���͌Fm�#e�X2%c}Ë��x3~;�R���p.}t�Z8j+��&�+���8��Ëc*��ܻw��� 8��gv��y����Z�����kڧ��mC��ק�}jH�$A��ágE�t�����1Q�IGY���%~�{�p%/(tÿmW�=~'�n!:��G^u͑2T�[����-�N�{T�k%x�({�~%(U4��^n~EL���l�f�����Op}&m�����YD����uHu�:�1�1`���e��ǁ��A�`�2���IG����Ne�ï�C\�N��w8^rM=tx��z%���D��Y��N��M��L�֝��S�����M;޿�k���5d����!�)/v�@������7��Fo
i�y��H���,���;��ۗ�[D���sR�M6�2��3 9E�3fuz9[��0�`r���x��Wƪ��H^8X)*��Ƽ���ȷ��;�,`͎vd�u�3E��s�j���e`&U��1�l�Ҍ�x!a�����"�#��ѴA��Ԁ�<�'���l�������>}��Ftތ�F��;����W�Y������#��/�g����Ah�D�1�j�G�p�4�6Yv�(c���3��!�]w�(�]��ſ�����{F4�|��>��G�M���RA����KDBc����	S�ciZ�L���V��&׋E�=��ⷎ���k:��8��nb���������z�Kb\���F�Ө�'y��%0ޱ���S�h�k4��(��@vN</����f�3j_�$�	W��"�X�j�e����Y��9�S7XSO���q���>җ��|�!�8�=ל �ڀ)�c�ڑ������������s��[t�m��ș~S<+�AO��zq_Q�%�S6�8��|������-aԭ��}{���;6����ճ��5iK�]�o�d�؅'��e����b�Ѫ�À&��ahpڴ�g��s�����h�/9\��ZO%j�D�5��bs̼�(��h7����'-��1�w�BN�n*��U�rp^�I
��J�/��D*��8�K�ڭ�bW��E��g>�u��/��ڱ�rm�=�l��([�S�/v�F�-��ިL���{��E��N3#	&�v#Pb �!���0������-G���@�g�ӕf}nN��|��������OO����?�,��CS�߶�u�u��ϭ��T�1�
m�B7�<�����,����@P��v����u��#A���cq�����V� JC:ڎ���BG��x�����:��{���cJ��d�g����kmk��D�����I�~dj��+G��)1y��RJ�w��|�Ry#%yT���E/�:�W�����3/�ܥQ�)7(�<��Aُ���;)�tػ�M�)&m@"x���"���3��zL%r�P�\(�qΎHط?<�y�Y����Ӽ�R�k��V�jM���4�z�Y�l�Ҕf��<�%��������
Q?���FK��[�a��I/�b��Om���;O2�:���!�ۋ�QV�FX������c�˧�QW�e4t�I2����q��[��Y��y	/�U�i����j��8�FK�'�&ʴ�@ƈa>7:&*h���Q���~f�[��\�����x�c;<OH��kS,p��h�޵�7�[x}���p�&�pr9��X�����3���i #�x�ߨBt'G��02����_���G�>��^�u�SxuܿoD�h�����?�Y�{�b��(7�̈����A��s;��^��W=C�D}�����L��L9R:b��hxU^��q��X��s�4��B�QvG�{�|G�u�~��y�8�I�vt��|u-���+;��t��s0t�p�gh���D�Щ�8�{���=���}�>���G�~x�5<8A�o��k�`�vy ���l���q�z~\�w�k󿑵�|����-����HYp���,W�~Y�/K�<��-x��j���_�r"D"���V�A�_����ٜZ���x�Y�n�]6i���>6��3�M5�&:
����!��M�7��u��/�1/{��������q�H����x��n'�k\�D�9/N�6�f�v�5M~�I������YCz�H؋l��[�,��J��%��A��u�}���=$��dt���U�M[�ߝ{����<�>��{w8�7�B(���Ev�7��"��9��Y��U`�'1u�<;��Bgo_1��?�I�ɲo7���h_����w���<|�������i��D߉w�Π������v9\�~��;w�ލ���>]imܫ�"bW�"8^�g_Gg�k|�X���>�q�ȥ�M�k%Ѕ�yP�u��c ��O�`Vs��ca.�`��  ���x�]�#Û�S�"�?��:z68ԧ�`�q��9��GN��G�[0|�u0e�΋�䮚�aH�N�7�0��1g��+H�W)�|�)�W0Q��9�[(`:���^$Q�5xG��cpL�#��o����V�C8��y�}�Z���8��M4�x��^8�ZϫyP��RG�������wN��Fe�����O��D7n<�h�v���|t�xտ*����s"ne��ܽ6���������ӳQ^�x���ӻ}T�(� z�9Y��mB8�s7[�45i���+9R��(�\��۲:����|m�'b��zD9^p�� �xfd{��ae�f�ܻE��w����{-��M�vl�ի�r�^��I�F�9�����jp�e�w�Q��Fx��,U��9'9Q1!3H�C�pށ�j��巑�pֱ��9x�a�f����F����<&ݰ���3��Ǿ	���Qn�Nyݛ�x��ոFD����t�06���u83�(�&�j��v����M�E���C���H�~�%�DK+o��8�խ���r×x��jq���!�G�;��c�Tv��t��;��/{*�i]��I�<R���Fp�vh�r�0�ԩ�S����S��#�_x��upV�\9��t���P�qώ�o~'��=z�4�CX섴*���s�XT�/�����~��lK�}Ԡ���ߟ~��ÇF�Ϸ�������>6o�Ϳ�u�M}��ݣ�<�;w9S��)���3>E��Ýh�cd����&I��o�9tE��O�X;�;���Wٔ4�u\��x��������nQ�96j��'�n�j�#��u��4&��N�D3���Tr�"l7v-[P�ed0:�Sv��kE��gfI��6О����y48�xR���g�����V۽��h��8��!���t����ϗ�Q6D*ߧT�I�~8/4Xo��&g�Z��r@3�ɵ�[/
X2��ڞ�`W�n��An�w�[�co9�"�f�8`��#�7p�����O8����Y���C�?��=/��BH]N�%\��E��M��
� �eK�g}j�9��|�S@6��w�}��c�;g�2K.����EM�+����uX1�\9$�7c4�	F!����R�@4�7�*��p��ԅ��=!N�}������Ӌrn妆�W�<� e��{0��z�SN�Λ'��40��7FF�A�;9�8����DZ�\n(L��V��X�nm��:�+i�� X�/�>�i��A��:�{�Z��^.Ϟ>�{�����6<�����g�'?������a!��J���<}��5O��)��Q#ON��B�܈�y8��I!��ơ�'�(v��jF�2����3�I8Zg��5��! ��O�Xe����n�x����zS�.�}���7������Ek���������5T�t#C��G�����վ\�z+�n{~1�Z�x��� 8�K2Y��3l�A>�m�������}7���K���~m����?�K��ӿ�ͯN?��'�2�h���:��_=�F���o6�-��o�]cő�9�^{!#ʈ�d���x���N�Z�y�}�d��S�N��0J�r>~Qqt�ov�/��F��t�uD�ۧ���h/�96�@b:��pZ8�o��ę��g�fӏ��hO[�:g�?�?��-؁'��WݦNGǻF�4y������+��~���K�G9p<�<��w���O>ц�au,wʷ7�����|�v���Ӆ���K�8����u��e���Nx���;�|�Iѯ_�~��_�>��:ZQ��7��Sf�O9\)��Ͽ<���������?����ʃ�/��ر)��"[��ܨXHu�@vD��y��[j@�ŢC^�)���e���!���ׯ��gk�C����4\ip)J�ێ'o�/��;9�m�Q4�u��/�ch��Y�b�γY����Ho�81wr�n�i}do$�hZѨ���7ߞ~���/σ���F��"K��C��]C���iR�(��ė����wf�fPO�{�goL���J`9WE&��ޚd;������K���O6D��������m�a�缨P���E/�c;i��񊜏(��*a��� y)��gBv���}+/�@c�4v��>v�'	Φ�w��@���,�e��{*�YOϰ�ݫ�1�$�[�$:ҡ��y��\��w�^�m�/��.�~:<*S�9�����C��w���\(T�*�,^��&��gNA v���9�϶�l4 >��ￅ���;� y<���.��]N�#��}��!�?C� ���s`Ĝ�w�MK3Gm6��k�q��Dg@Дb����W�D��ye:���ڽN���a[�����G�<��&*�l�Wi?��}��楾����~v���<}��_������O�mV�RC|^���szҜ'�?���F�"i��͂�(����h���f<N�T���U膳<�L=_��z2�2<^g�(-���L�D�!�Ҩ0��k1'�"��~��Ӌ^����������sLS{1<�ݟ��M�l��{���������G����J�MM�/�-d��\��r�� Q�s#����v˾�|�tI�K�c�����9b��X��>�#`�2�[�j�B��cGy�/�u4�Q���g��1�i�'�B��+3����Y��|�x3��&W����������/E@Eqk<�p������D�X�e�#kDnT��D��^��D�B��T����*7�	�kx��#v8e�8������u�H:x����G=e�X�L�\WV��q<p_�Ҳ�I���S��s��x��1��;_��W^>�p�%iS)׹������-Q�S�Q�-ѝs$-���>Lo����1j�\��t1��,�*� r�{vV;e��ta���:�ɒKw�s~��ʊ#�ʺ�2��p�5r������C�>�����:���! Y�sUÜV�M�GY����E�܋���},VT��y!થ&��ԾiTӱ�0Ѭpy�MF{�o}�ǋ�|r��H�0�j��`��]��/�����0���8$��o��ȕ�?9���Aof��`/�+Q��g�]Qj��~q�����Ot�WOvp�$+�8�k#�� ���Dp<,����uO��<=�W98��z���� ���Q*Pt�8��,X|�����o%����9�0���Z�O��q�)�Ӣ��˜��lz�r���a^|�'d�u8���ޢ��j^��ţa����J�$�������_WS��N5�s^ÄE�r�� ��[��-ܮ�֨�aZm�r�N�F��3�M�PfJ�##��,۔�����C�pxz�|.(<�E����M�52��n���k��3b���7N~x����T_��j#�[��|�R�� �*�`ِw|��|F`�+�a �� �����#�b���8y;o�X32(a�����{Fad<a�]��p��x�!�2D[#��ԕF�>� ޸������?6��h�S��>e��l�0��Ŏl S�PÏp�̎�2F�ɗlb�����I,E�{�c�|Ft�'�����|�t��5%�Ua�?��铏>8}��G� ���EΈ;:�aC�W���m��\/=��0lsF�Q,\�c�.�]L'0�&��u6�¨�a�N:'i���Η��]�MW�xNǁ�_����Ct����!/X'�E-�/�a7b�|�޶t�.�^W.�t���8�-B�<�8�(����#��t�������U^��\��^�M:��U��������s0'l�r���CY������s�x)8�����j89��e��%k��)Rá���?�e��Z��~SQM�U�(�:��:�ױ'���u���i�@(%��P|��Ac��-�{.De�0Q=���q>�[e�k���hSaE�p���i�`�6.�uo��7�Y��z�k|b����9{k=�n��椇���
k�øt��e�B���X�8m�R��T[U���㬭[��AӺ7s\mS��_��}�7��CW}ǧ~,�nV���Qn��<;x�pя��t�Ν;����^�N��|]�ت�w����M��>�@�'jf�F�=�q�������.�P���� G�8=�Z��������*�l̍���۱������x���g�i'�w{�t��q�F#�Vg��爓�wٚ��湿rk�G.�k��5�.�G򖶛��ޣ~��D?��a@�D
{a�{
�~'�g��3�,C���7(����9�$!8H�	d8e���~J�O�ʫ+�Y���(XP��2έ: Un���P�b���Յ��X�P48L�7
9w����@�:��	}��o�')����\��Z�3���m:i;Q�l킊̷ߺa�;u�Z'�[��<��]X�"b@ա�^����K�a��o�L�(T�2�|V-�F��vD*q��lZKq�t�7�l|����䠗��v�s�D���3J���R�Rc�ڭ��O>������cE��ѷ�%k����8y�N���z��8���E��ix'���tְ+�:1���I�4i(�o��ځ)Zہ��So}�}N�_���6�=�-�~����o�i�陌�:*��>�ރ��X!����Ӓa��=�Y�N�A�L썒�Ҟ��.�Κ��B��1��(�܅��G�o���E߬[\��Mg��a���Vݔc���K����#�q�n�0�2k� NgZƣ�Αz>y~��ׁ�������\���YT�sԥ,�ݥ^�,����q��G���j	�=�9�;�<��.�A�j�=i���w[g�<_�{[�`�5����V���=9������k��Eئ����������7�Mtw�����񑽃��%��j/װ	td��;�=��e[�K���%��6i�7����E�\Z%$����3�6z���4���yt;����2q�
�D��?v3�����ïlS�
�|�5�i fo�q�g�A�q��wӧ"���KsN�3��l��mS&�%C�`�gn:�9�g���R�p���t�m�'�>�cR&�H�9患�� w/T<ID��}�*�l`�o�:0/n������\���|�Z�i��w���å.Q�LJ��	���+���O��E�Ǧ�B��Q@r�}+dw�U�����o�5�k��78�kH	������	��3�}�������6�sSg�=���a섚�e���1����Ax�u�[�h-�}f���Q=߼K�=̆5��~�����oB�ԩ�L�q�6�/�_���Σs�	c�PhY�+�l����A/3�o�(��X��?u��	�Q�|2��Muǣ���xqLC��<�����?��Q� t|W.߉��N��\.f�덐.�ӱ�;5�w�N���8h���&��ِ,<vp_M����08:���},M��+�\�8Fc�5"�;�J#���0�]��3z�o���*�ń9E�2����MK�𽍤S����c\2F�]��h�!��F�/�P�nGj;���Ȳ�ŭ��땉��<�j��P�L���'�Տ�c��sj=����t^�5�uz�����[c߶���������u&�T�ut.��>:��&|~���1:�G��9Q��:�(�0}R�pr�,�_��� ��]y��.ã�y.<��8od�=�	�cI�F����}���i��%ʥK��,����*3Z��3��n�*�������9�s���y`��_��h9���{�M��t�۩��A�_�G>��9�����>�-��'����0��"W���:ԋ��w׎�����<vn�:���Y�uhx�4u��s9my^*��p62*"jO���;-�@��A����M=�����iޘ7�޹TH~���0���A�w���Y5.���9Rl�V&��*[0�X|�;8S1����]�OJ_@YK��Ǉc�?i���
٠���fV��y#z�����쫦�*�Y z���K+m����{�w��C�c��m^ή���=MK�W������d��M�-��#��N�p׻�Fd�.�fF��|NGjm��-{��@� l���{��#����Jo��t���i[m��}��3,�n�����䲲�o'���$|�ζ:�<!��N ����K��n9[%ǧ��5|�>�%)\��%��S��ʱ�"0z��e��X�-^W��(ѷY7e`�|�{�1�V�`��| ���Ըw4��BT�-(���	�2�WFI}�(�i��TD�0���h�~a�Z�~��X���W�n:)��GX" A���i>KS=2��>||\��0؁i�O{Kd���qpo����a0��< /,F D��U��rZ��>K4����|����O�0P�4Xj�N�#�:�e���0�+#���&�o:(A�؅�����6�<�sX����E�C�v%�	�O���_���~�f��� Vf�,Pmx��i�2'�uDi�r�݅5X���1Maǘ�t��zk�^f$��"��V�yֆS�?���fn9���'c!M/�s��W�&���4;6�Gk`H��o�oㄕ0��dɤ�&ʊ�����/O_���E29]_~���{f�4m�Q��8W]���ѥ�f���C���o8d�ۣ�i�2��D��xk�ƀ,�GǏ�_G�vg.�m��~�j��6D�W'���c��a
�N��n����o�M}��s��g;򊦩c"t�m�>����'>�)�n�@z{��;p>��s�w<?�����mSo%��������C��h�c�����K>'X�����s��9�oߴҩf�61x���H}oNx�����:�ySq-7y9'[�!�ܗ\�U�m� �a;��kk�����|��-D$rʮ�H�W�z=�8�Pں�ѿQ-�N����S��y��pljy�/^�X��7�D��V�P��5;�~S���L�+��aс\w���Y�A��<��]�i%�L��Л���f."��û�^��$��!=j�&�9:)d��q%|�qp�o�=%U{sFd�W��ľ"Q��7i��M�6�Y���DX��d$�}��E�>�XEy=W���r�wNZ @�\.�/�C��q4u����搧'��=�K:G!�(��9����T}��ck�$v�Qفu�p��8����a�68�.���M���ڛ�� ]��&��� �Ǖlݥ^k5�����.r(�3ߗ�Q�����׹
J��TP��>h?�'u4���73����i !2a�Y�����3�G� ���
��S��M�9�O���1_TdF5�	Wz 䨓��W�R�hFW�!f0�t�TF���%�q�ʳ��2��Czz��=�p��#�s� �:�����sW�B!=7-���ƙS1S*��� fѨ�M%���NI�/k&_��FILA����q���c�:8?��a$��I>����z����o���5���X���S��V/ظ6�WF0��Gu\5b�h�i�x	��E|뵷��\r�K��f�i:�`��� @]����gu�Ρ�YC���Ag�/^�v�ETs�;�\z���j��*IsM�17�N^��"���F�3{��b>l�Y��7ꚎU��6?���������UN�f!�,	��q���ap�a���V.=w��J�&�zv6��Ql
����'e��O�dؒ߱@|�z���޷��*�w�v�ڽ�જ�|�����8����{��;����������14�8�����;��׉/p<��|:��p�t�L���h�A��	�{�N0Ҏ�5�o���m^-��Nux�^m_���Gx���/������H�ܥ��þ�փ�Cw�^[,�8���Zyv3;s�����MAM����[�]���3���J�g�@��ۖ��Mo�$UE�xm�u�cYь]<�O�����'�{3�بu`�c���^ijt����"g#�u�3P+}���Qvh#C"`h���ǵ7�:`و"c�bK�̇�+m=��uD����>v�;��>����r��7j��/��	W8\ɑ\l�G����ѭ��t�|��Δ��ѡ��3:h�d
�t�SFp��=� ؋Cm���}���K"Ϲ��]��nFw�������T���Hᠤ�@���X���e�׷z���,�x���l������~s�JNث	|����/����̦���[2�����.��L_?�������� ��>�V=�Szl-8������;�Vjr*�;4�#�Hp
ݭ�J�5��i�գ�焵)g�򚇮U%7]�Վcso�17*w=�;���:FPex]c�p	��}�&��L�Ӣ�0	�z������I_7�f�����Q�2'�-�w�lz�C�<��b��l�:hMœ��`�� �>��������������Z~|A����k�l�w�oG��N��z+sV$��bS05(k
Bw����a���S3�$�i��C���)���oy�:+��b����>�u���?�|�	Ѭ΅�fnHpч'5�í�<�Y���
F��֚��zL�����j0j�3�#�s��i�()�q��#����iH��|D=�/�L�Z:�d�	����kG��7k/Jp�gS��)�ީ*��,�$C�[�]��s�尕6�P��wQ����p�Dg�'�:��@��u*'r�e���� ��:`tm����H�7tw��6y�W�Xc�88���	o�:���H��h�����Ҝ���q�]ε�~�k��g�s���z<[X��^/\�<4:���|���gp-c��3}��	���=� ��Z�/y����ߖ[}B�t�u`o�e��^ݵN�%�l�i
��6k��-^�\;HP�'lA��}��6��>������
����M�D�)W�F$�p�7�\����N��ÑR.��^[�}���gP�C�ӯ���Ի�T��e:�NN^L�3ч�-ҏ�ã돯�T�A�Ցs���ϋ r�f�٦z�I]0�qG��r��A�s�f`��צ�w���F=�M�����f���Z��hX���=8�n��� m �W��� ��<�\����m����`h���_i��8��|x��W�� ;���^��`tB�Q�m����/OO�$| %�}�����E���{�o�'�:���W����1XI|�Voɖ���ᩍ˛}�2[��?�!�L��yk����O4���Z�7%W�5m�)daq:ϱMH����Z|�g#�h�5(�n~�6�0gIBBY�9�F��3%�0W��z	�k�z"`�J�A��SBF35�='����;J�� c���˨�?̨3f3g��FE���� mp|�(�V��v�`�s��AcTh�R��B`x�ty�����rVH���Jt��@���N�w���s���N���4 M�n ��>�����p6�#t���7<5:�Է|��留�k��q�d���r;�m�C^�fկg���:sS�� ���40�*C�,ae���U ��������$�h��k<�!eSׄ�{�'���)\�bH���-Y��J����d(��sE6�afmG���Δ�%<�̛���8.E�шՏΉ��
�t��x��0@ә ��o��	���#��S5���0�{S���V�5�ъd��i�.�LA]�g�22��%Bى� $�螷��Dw����֡�+���?�x[fe �.v���ۇ�c�s�m��:���iҏ?�sʷ�N����~��/��ci���q��4��uh�(�i��a��m���?���(Ǝ�'�/�&Q�I[�&��HǤg����i�Ξ�
��-xhk��ت�~,{;6f0ˊ�`g�+����c���B�|��Z�hvI�Օ\��6�3e>O�8m��k��녃��9�-Uj�
�p��s��pt�������q�!�>�z6/<��Fo�f'�y/y�RoE�9P� }��Q~�E,>=��=9U���(*8�h
[<|��n�*��36|���(e��F�rӾ^�*b��x��~��f���r��<#s�]o��/ǖ����e��6��=�;v��8�fou9/�#���
9s9�6�Ӓ)�S[XH�&k��Ӌ68��y���W?��w�����?=��o��>����rz�ӓ�9P_V֚�l��z�p��� �i3�X�=��G��<��6t�*8f	vy��W
h���A�-G���Wsت�ٓ���2Kn"_ź:�}���[o�Ns�-��	{к���`����k�  @ IDAT
��ϊ���9h����[v�5�����;+]7�G;bA�6���D��28v�G���l�s�߽79S1{p]��b�qxN�_�(
��\`R�*W��~)jW��>�a��¦�g�@�1��Zpj�5`����A/	�3#��C�S�]���ְ�f^?vZ�6�atTX��8����H��Ո�P"a�c웃rI�߾>S��7�������rK�-A�$����%\��)�8��dv0噏k��HM��h�3r+#�t�ѝ�͹#a��Q�}a|��&����n�wS��CVg�!z�<�^��̌6'�"�tr~7��4�/���?t�M���I��˿-7�{F_z*g��oLg������tl+��=����d�2$����p��,Lv�`�#�u8`�*#r����v�P���3r	�|&�S'�>�^狞nG��(�@�"��)30J?�9"�:���}�@Ӂ�g?�:�g~u�����حS��|9p�:�����sx:�z��#�=;����q_�mզܣQ�`�w��tx����ۙ������u����w^��4y�p<u����O6M{����UN�CyyG�/=�ۥ��L9���I��UؿP��-�g9_�q���K^D��){���,?]oQ�0cG����t/��a�]�Q��>��2c?D�v��h���T���1���r�*|��S:rF�g=|��wxr��Y�[���x0���:mO�;6}�O�Ms��e�v�oM�ȃl��
L���n�x�!���>��E�2=���x4��E�|J�e6e���j�`3������8A@J�is�8'VT�!�@'$h������9`�N�w�����r��^�I����oo�[0��m-��˥��_�����0��U�q�k��%��ܲ_9��ӿ�t&��֞���_��OD�l;��8���3��wM��F�)Ho\.Rt9g���>��Le�x�G�3s#$ZHx��^�6��ˤ��32���)}O���e�5�Fi	�TM}L�IY��ǋ�0�@d'&\�ٕ8�S����8N\�	�XN�����}j�٭��YJ���(. C�4��A�[U�z	+�ퟦ!O�F�F�`�	�Ӆ"0}�����G?}�i(e�귋1�{���k����/G���Ֆ`_�3#���Ys�2�u:��`�m綆)�(��=x�:cS���#W���z8:;OܟA��b�8x�_/>̜�k!�6,4z�?F,�����p��r�C5�2B[��/
��O�(mv_./��>8�a&z{���1\E�з2���F�<rp/�%��:6?��Tjz1GŽ��8��a���O�W�a���3Ǳ��Ę��}�Y�rLU�:��������i�:�F����q:�4`sJƉ�؇s2�.	��ҏ�������9E�8������>}�8��4�0�J���my�F����3��3B����'KY�:0L���
t��^>'����3�A7z��<l^�ހp(��sL��1����)}xsD��zL]�<�#��Du,�k)2�Ц'��?����s��3���p������Թ�cj��=J_�����dZI���6d��a��Td.'%�O��66�B��t��i�f�Sx�耭Q�������2S�W�}���(�wg��^�yK:�9��/s�;���5�70�\����,��l���O�����y�����̋T�U�o,zAM������j��f�W�p%��_��9�^������+ߕ�[�O,���S�k1�����7_��Gҿ���~�]F.`gM�����Z���>uN�i�%f�Ȗ�`��Km�6G�կq�L(L�]!�[nt��V���8�Iy�#�i���̓��B \����`��B�s�D(E���z/i�j���������ὖ�u=x�"H�X��?�V~"�K&��	��|Vg�	>��!+��O]����礮���۷ �*��{��Z��H����^�>E$�C{���ɞ]k�����"ENy����Q�g6���7׼���|����c\GLW�0��7į_�-V���}��e��e=�I�>�0�C-�K��Åd@�/�&@N�FZc�,�&l^Q�0���ה��!K�"#����n��:�4�[��ncTi[�C��t=#�c�͵�i�?�(�	��Ż)�z�� ��Q��`ME�*�t��1-�������8;�s��g��7�z�U��g�x�?�3����x�����f �����rlm�a6���c�C�<��DB�g����?���}�,�iHr5v�.?R���:fsW��G;̗b�l���|x�`�G8,eHB�Ps��xr�W#� ���g8�Iipvߟi�,�.ȋz�@;���JTv�w>����4U�;�r�!����\�H�~R�����S��e��N`��弭#��ʐ�h_����&��G��ј��/j �hrs�;~�)��l��O�aS⠢�ы�1؋�{u��=��Bs=�2��p<=;�'��D�{������ڟ:��;�J�u*ǐ����D�n��8u����Tv�r��wF����8嚪����v���	О����\�S<M.K��H��!k�+�3�.oUzL���>��b�O輮���M:+��c.=?t6[+gp��wQ��ٮ��\���{� ꋯ�9�����Pِ,@H�k�\HU8v|(���R�B�|�%��E�����ӟ���O+=-Bs_�q.����yց�#P���B�-��;�ZGB]��U�>�w!9��E_�>�s$�_f�ɅsK� �=Qn��I�ҟYj��y��o������;������l�!ĩ�8�`s::j�s�d����w�O|�x֘�9���5^0�/o��K"��?ҁx:�����W�$�G��`�7|���+��zM�v/7���j�~���V�;\VN[
q/p����?��OKq�V�շ���_�������X<϶�pģ(8�����
����p�vit�m���{a�KW^�;#����\��P0���c�B�O[x��n��I s�(���l�1/�2g�#eO����s0�·��.%)�y������������i���iILH5u�\r�af4�ԞX�������������'*�N�1a�"ҩ;ؕg](Nw#�i�n&Euc��ᜇq��54�6Q�����1��R���U�x0#���`<B����l�+�Z�������3d�/�3�������nο~P����y0�3�m�ɿ(�\#ه{�����eXc�.�1a�/�(�T�S����DS��%k0`��M#��#a�7��+:�ù ��ʰx��+d����_{����8��q�mp��W��TG�hh�0�mg��L�e���z� �������o�*RjQ��Ђ�!c�џ9���쁏a}R�Ͽn�!�,<05zǴ��zI�8!pq����Q\Z:NF��	?���+�ժ���|�w�26�.����ښpma5�16�o�T�t�=\�隈]:�?��3���E���Y�~�>����D�73]�{,�Ao��F�;d�\{��:S��[|K�I^/�۲tz����N�NӚ%�z�;]�������v.�<j�:�<~��i���xq��v�;��f��3�����أ�94�ɺ�g��+�Էxh�ڡ�tŏvQ�8׫>�v��z��zn���3�U�}"1k��gMU0kJ�c%�O��a���������<K��^o�Ă^B�ۼ��2`���X����Q�$YW�_������v�O�����_�yl��+v����ޠ�R�0Q�.�܁Ev��r��̝��NN��_#�k�G?2�����ع���8�Lgp�I���I��Y�P9��.�_63���7?��s���o�>��~�b밊�h�֩����g+{:�ķd6�[��c=�q}[�0�o`*G��(�2xuPs���?������� �/r�)k~ɋ�'��"a질��=n5������7��M����,�����?8�������Y_'yh��uXޥ�l�`��8n4Cxx��N���'�3�9-T۩��h3^ ��9t3��n�1���@��֎��/0�dI�h29B�!���%fԡ5Bx�B|R~��v���?ox?�[�5IJ.��U�"6�02"���/VW8�C��)S}��?3���x�m?��9� y������AW}w�EG_�.-�Z$,e}�B�:���M�xvz�$R�r6�y`Fʾ�Y�Q!�Df��������t�ЏY ����鋞�9o��ʃ��.�!M��G��>G������q�0��0�^�����HJw{�D��28�?��]�:�>9 ���j�k�Գ�hyi�O?|צ��?{?G&xS��U��b���c���ʤS�j���� �iw��I��jp1�^7�Q�D�yi��7|B�H��[e׌��yg��̆�5*+�s��<���N	s0=�c���;J�^5ʻʻɞo�$�9�>�>�K��D�e�4:��}ϏN�������q��N?*+g���co/�h�R%�6�H��Zmv�tc�ϰ����pf�Q���:N	�.�8GN�r�O�^x�8�=?p:i΃~��s��sx���m��s2��W��.�G�4�_u�����2!�u�ӯ]U+�܁7\��Q��]|��S�����p>F���q�Ǜ�ނc�n7�����ki0���v%�2�Ygi/9M� �ڻ�]R�p�hl����ϼEۧnr�*�
�?�o���w���Ӈ}T�˧O�~�ׂ�o��:� ���$��Z3�h�ӾPQ���?~~�ݿ����?}��h����5010h@N�<�`z�"n���������꙽%�3Q,�{����'m�����<�!�1x'�'��(�]yi�3Pw�]e�7��Mѯ����o��~���"C���Ӗθl��hr;ς�x��-�||���w?><=$w�NN�b+�n������Rݾ�DS�T��љI��6�n�Ѧ��Z3u%o��۷o���ӷ�ɞ���G�n��f���A���sp~�٧�{m�ml_�����F�(exm��6�#�ck�M��Δ��o�$6�zT��ѣ����z��#�{�����~�i������^����l�M�K���C�����ztz2�)Eٷe4
�	�B0�f}R4J{2W�̻w��VG�����m��M�PQ�u�t&�Ncfzpx�C��Ή���1�:94��l��K��D�LER��՗��8E�|(�r�g����z�6���j���T}�h;���sF�p����r�o%E�<j�h\���`��SGO�+E��뿞���_N�� l����k�).mtl�H���,�ș�R���1*�.��uy)�O�����.��|`����\�g �"cdXT#Ռ����_�n������{w�6�mT32�>F��U��Huft�P�[��h�u��L�g(���_N��~w����)C�\�mx�qt��`�ò<h�9��K��6���Ot)0�6*�V�q�ۮ���i�����H�K#_C�.6Ч�5�6*SX�qV��<�2tx�-�;EOt`�Ч����=8:�u���.������:m�pD�	R�X���B���%d�n��F
y=iSOߔ�f���F?ѭ@�������s2m";��x���ҫx�=x>�x��E��|8��,��p����Ɂ������W�+��Z=g,�)s����W|��p�N�r��c�&�d��9Nep��s�U���#T}��|��*��@x��e�d�ި�M��.�X����Z_��vK�)���8Üuz�m���UM8�guQ}��@	?�dmm�����2~�4���hjo��o�{p�����qz��������t�����F�m1f�E�����`K��z��ǜ��f~��-R�}KD�sb�9��_�m��Y�u�"�%�}��?�Z��,�Ù�)c?�P���v��D{0�L$t�
����+U(]��ZcD���ԟL�i���Q��g�����^_y���E��/cK�
.)�����ux�N?����˯O������:}�(�%=h��i��){&��)��{��;���8���a�ҫ�~Q�����E���J�{���;}���"z�>ʑ|��w$ܾU��<komVN����b'��O���X�B{r�K�w7m@9מ��QF����Q�~^�#�zi���9��{w��l_e�����,��O6bF�!4Ҡ0��J|�������������R��m��u2�,!���`:$�q�f�͔��"}ktx�4=�鲎�Y��s-ZL7��l��?�TxoG�Ôg��p(Jj��H&�l�9~�mF��1G�_��Z��ej`ι��w:�\{v��o:j#�=���ĝ�u�W�`���V�1�/7*Sc�K�M��zg��S�Y\����g�q�h�{"�i�(�?2����Zܟg�F$�_;��u�𘖅�����25 ��	�@Tg�:�a����:aX�I?��d��X'��d��� ��K/8�]�Wr��������fd�����?���]��cЭ���������g��L]��`�'S��_�x�/���|H�N�^��r礓��I�.��9b�O��JE!f���M3�܁���ov�>ݿ���Ӿ�w��ݦ�n̫����N�)�a`u����������4t1�q���y�󳙆,q��i[|�u`u�xTi�V��u�{��`L�]�50�e�����;�(������������Q�����=q媶�����D�z��gx%�(0j%s�x)�MN0�:�>u�+��=w�2N�Ҝ[��Á]xCG�%�ͣte��ߑ���|Nuu�]�(�3���![��1%:���������];��-�e��<�RߤX#[9�M^����޼��Ѽ����O�0���{�^Ѩ�NT�:hS|���Ш�i?ᨾ�O]���5��ȟ�4tx��'X�,�^�wK�A�ŋϿ�Y+����{����/�A�gGۨ��i�h���_����"_���[�������E8��`�%��K!�+��'�v?G$�c2dL�ي^䣃=�n�U���!eo�����Lv3���e��i��ԩ����>��F�D��=k����8U�����o��q��f�7�������н�����{�������A�y��v}���k�����m�[=�m�[]C�( !��9:Q�$�w{�s6w�^���xf������n����m*��g��$��~�Ͼ��Ř`��6:
1���1��6½t�z���t���!	�ړ�x+������v�m���[�N���K+ِx�tVw��|�k[Oڈ�������X�*�us�>�Lh1m�f� ��"޻�������Ӌ�u� Nؠ�5��o�@4D��C�������n��]�刕��Yh^靈Yx<hJ��_�p|�����C7�vF����Mv#�)�=K�� ��1t�����b��u�9�9_�T��#[�;*)#�����#��da�t��"�B��=}p���5��_[�P��o~֫���C��S0B3��o�5IN�&���m�/�G����?�,t޷���%��{e��+��J��oO{@yu��:Khn��ԯ26@n�h�~�Htγ�����zd̹ģ����Ɔ��_Y{YT���9c����(RX�t~�G��h��yT�����E�����?���wu?��\�dTnAcɌ+��e=�.���ꙺ๸r��$���@�Y4�غ�x�;y���G�_�������ٽ)�����_ݟ�q�ݷ9�?���/�6��5��:���p�J�8K!Y�7���Y���`�1^��[Z����`N��Ik�tL����Q����Y�<�o;,�(�#�o;`S�?t<8ܣ:�Ku`��㙚��l�E�4Ù�%��/�a:������qp,8/�k�L����)������'��u%;y��7��鼗���y�3��ӈ*��ˈ/xfpk*p� 7r)��ᯌu�~�Y�8�n"����*��:<��yK3x�<��'z���OO����R��n��_��T
��_���������?'2��~�.�c+ʳ/��쉲ѓڊ���B����k���?�f�ګ�9�.ϋ4�j]�0F�u�_}���?<�_O���?��m�E[$�t��<��ɡ��ʯ[|oI��	N�lf[�x�ۥ"_��_4��g32���<���Y/_cQN;��|�s�j�['����f���a�WN�ӛ�M�=���=��_�G��}?�H
T�K�.@*��=���צZ���W�=�����o�տ?}�����Ѯ��ݷ׹{<�6_~����囖�<)������Ģ B��캞�I"�ރ�@�L�2���W�hCk׾w��闟~t������/�I뽚Yx�U���ѕ��v���Կ}%p7]{c�u\jjP�	0����~�
̯됙����t5�p��#�����i�t���3;7�(}�7#k˽��~�<o֏��D:$�p��h��i��*�����5��(�}�^�L�
نY� G
Ԋ���1�!:�kS�d����_)o��nq�l6��3�X��
�}�Ï)��)��w?e Z�\i�QH��F��zp�d��b �H�s��{�B(֋Q�4�>8~/k���{�7�<c������5u��Y�G���H^�̏N��×�2
�������+�2/*�p���\�
��y�ُ}���M;�����h���Ӝ�y�a���� �{q\'�u��rN�+'���\��o��!(8���>\�RH����/9���!�16�h�{��FSo�ڔ�2�Q��'<�����ܞ7ϟ!.���88tpF�9	E���)3c��������~�CVj�1-P5�,B�|ɉ��� ���W���}�Y�U���Lѣ��ӭ>C��[��}�a�A~���y�ͯu��t�{�f��x����M���o��s@�|ux�	��5u�Ou�]�+���/��l�?XzάS'�m��H;~�408~���]ǎ���v(��N�M�e�(:�i�mN�F�ٓxUy��w�)w�����޴��)���8��.ϧ�ā: ���˓�G}SF��Ӝ��^H�w4������CGʧG��4{?��������:��O}�)�C�tN�����u,�3/�s��\�]v��BM���;��R�.tʌ���gs����Gup��mj�3(�p��u����߭|v���^����U�"�Y߉��ќ����z�������*�f/ʉ�[��E����
</zuQ&�_>x2m����?sTl�iP=4|�|��Ū�m&�S���c�̢��wZ�5g�#��X���3X�h��?��4ʳ
��HN����z7-+�1��ؓ��:�����ݸu��\��Cَg9(@�,R�O2�4�@P�f�E�`_����>~�`������.���������ѝ��d�����v���ZO���Wp�Dt�v������c)Q��Y�]������~lx��z����ik�.��߽y�7��Y6�g����}r�)�6���u��3u?�����R|g�虈<ۥ��n�O�V�����M��CH	��7p��brM� S�F��v5Zyv� ����v�}еu~<ݺㅠt��e�{J&�� Ps緋z����!߂�������YP%�����F#:�_SS�0��F�Z'x��ʵN��$�a��Gc�C��Q���dJ"��*�e�<�Μ�XE9��x�J9)���	ׇ��yCiP�g."g�Wkrz����*/k�/jԳGI�,Do����/�E�A��8F�Å�=f�g!�?}�Mk�͚�_��[H8#�pZ'nxx��n�|�H���_zm���w�x5yٴ����paxL&�g�3ru�#��/�S��0���v�n��Ykd�A�Q����сD���ˣx�a��A~�UR�P�7��}�'��������?���'��~�g�9��1a�k^?O��~(��(g��/����2�<�����0u����:��7W%�;���Lg�<~O4�g���H�҇��Uŷ�s����N��7�,��,r}���7�\FT�p�ţ7J��1���ҶޠB$F��q�Rz2R��W��y������q�ݏ<�7\������!��ن����/i��e[�#v�\�3oz_�eZ��4��a��W�Zz�Im����ͼ޻���È��V���}�#AAI��B�
v�F	F�̽n�_�$
2x��w�O�p�o��)��vW8��WG�Ce�!�2v��ʏ���/u~)�L�?<�}_a��i��g߁���v���&��|�g�v��i.XxN=8�AX�:�����u�A�'�6i
�|�N:xૉ_��=Q���A�(gKNWV����	oH�~�|Ye�p��w�ҧl�^��^%�|Eg��(g�]�ܖ5Wo&/+�s?�l}���S�X�FI��j�y,g�_x[�b�[zp�;C/o����I�|u�Ƴ���+������U���_jю�6J[y�gBK]�Z���g|}��֯�F����+.����k�4:����ʀ�5��!���h���|�w颽�=KV>Y��]�<N��k��-�%>9�M�w/�������$+��}p������_�m����JQ��ߖp��+=3�_���W�d�����+en�'l�'�E�&��N>�-��u9�͹,TY2֨	�H�F�u���X��1�Ç��rԮ;/�߳���}����������w����l_$̌��s�C�_�V�\��j)ʕS|͏q6H�]֩@3n����Y2rE�*�������N��)�:���4��`,Z�>�v�wf̎�\e\���m�|����E���Z�Y^�ʄ�@b��y�
���SfbV�+���gv���sE���	�X�aS{g�
RXuS�D
��T��� �`z[~����W_�Pw3؄!1����C�1���[x�(ͽ	/R0F�����mB��E��{�8�\�K�vk����D�3m/��6��Zf�6CZ=y��������G����ѻ$�e���K�{����/Of���NcY�p��	_"�ɢ�K���9�W=�gY�f����
?�tL��������zQ{�C�ݽJ�dޟ�ʤ V�$����9{/n���_���aa�$�u?Ӹzp�G�����x@�_�}��©h�~��rс_��!	��@Q|�#�)�����S�?��2P'��u1�'9R�����ngh�o#��>K��&�
�W=5���sv\��o�h��ǟ>��Q�8ޯ^֪����5tq��h�7vzp��c~�aW�U���:�|�AX�:K��4Cy��Gބ?Z8�{�`����u�S�#he[�u��p��ȡ^on�4�B�a�~>E�@�d�R)*�c�����M�)c�Tx���l]�/�rb�����[��x��g��m��u���E�].g�J�luL�e;���WH-݈1���G����޻��b���ؠ�S�0#��&y��R��r5�s�ɐ �
���~���=�;�Y��J��{����{��\��F���4������� �<��,|�,`y���\k�i|�Y]z3�t�����������9���L�:���
N��4yK	��5��[&��o����t!C ���BȒEk��p�:��,-�cc�qdJ�����Z4���O 4�,Z/zS��ᴆ��M�����;ɑ[����Y�UV�G��~����_Gv��QՏ[3K5d��&YR_�zEA�����d!��mu�b�L����d9JE���}$�9�f�����af�%�F�{7ﻪ+���#Z�˜⒤��I�NK5e��I?>\nR�{��w_~|�۶��W�>����^Kp<39':Q��8<ii'k�q{R�M��@�����˸��Y~ѶE�ZߔL��Y�d��_���7���� ���כ�W��S)�����>F'�Y�ہ�^h�~
�e�aá7�4�8��j���G�?�(f�,HV~=���+ε��ə-HN�X��� ����`����٠�,�3���]�~�{=Ű
9���5��I�bh�5!�aSM͖���+7�����bg-�7A�P����G)_�~�M��?��'J�C�t!������T^��Jw�A�U�̉����bx.�h;ǆ�|�mX�� �7��>מsT�,�L �J�R�j5�G�/�������;�?}w���o�G�Ԉ�)�,g��L�X�1�����*f`��ps��[�0JV�z�k��Xh�ڴ��O�At>��]��*��	��h�$��M(�У�;��W�g����'N��L�d�{�o�o�<l��O�.}�c�^�ۂ��4V��G��_��������zC���Ţ���s!Aïc֬	��ҝ��f
j�S|�T�FuWZ�8k��<�sx�E
��5\)�˲Q٤t�Oa���ow~�y����:O�n)���-ț��A9:��wz�S;��x���7C5�N�2:����ڇ&wr8����7�P>�c�V祷.(��|)��v=)�`�\΢��1�e�~y�k �ԢU�*��I��M�L�E*�WZ��(m=S��]Z�X\��F�M�l/��:ໄ���K-'Y���O+��;��w��u�ZN���^κ.Z,�(��d�$ͭ�I������� ���G-7S���R��v��]��U���M8�?;KJ���~�_9Ȟ��->M��믫,���T����x��k&��V�b�nx�~��42V�T�٫79ι�B����n�|.d� [k�O�2|YH+s�"wCz��Q��|��d0�0�Mk3�R���?.y�lz��|�]�O�����)%���)�L2Z�ѱ��tl�Q���d�4�Ay�.��!�͗G�ep�6}W0E0x`�)��X�|`)�V�����Ѹҋ @��������3����6��O�x��C"`�#C�[c͈�4�P�3���S}'��^ʹ�X�rLa��I��X�[Y��$���Wʮ�Ӣ�:R�gu R��)9�R��X��oQ�x�1nh�/(�V%x��a�k�(�!���?8���������h�����%e���R���Ȫ2��	�Qjn�zg�I�C�ƗY�W��ĉ׆O�%7����+F�Q	Agu��=���t*&H�*�U����BqZ��0�)���|P�5㖂x)E��u��&�6����b��yV�w�͔Y�k쭥�T*��3�nf��)��kEV�P��h�𓏐Qx��x	Ǚ����~*JYb*?�L��i1��-^OY� g��!YB8G~���a��������\nh�Z�f>����'h�|<��:Q)r�]�F����V �)*���vF���Q��cMI#tXPb�h��k�>Lc��3'<�/��8Y�}08c9��I(c VK̌��E�֑�Z���#��1 >���K�GSl�{a�U	9�S�^=o��&��b?�3�� �iV:K��
��u��Px!�n��zn�R��
9�𞼦��m���}�8�~��T�kU�"u?Pނ%mʴ^[�-�+A��d�p�t��W(�zx��6��R����0F�+�pE?k�=|����?$L^~�	�Ze�J71�E��]
����Ya�4e��!;��><�� Ȅ^��s��	������Y0�CHvJg���y�O��}Ხ�Cޕ>�Ari��X#z���ş*�&c�"�Y$J;�ŷҸ00�R"���Wx�	��Wa��5�Ki(m��xxu���úG�Eӭ����0�>�;�[�K=������[q(�+�Jo�q��]���Pmx��p�Gǎ?�ga��Q�������B#P���0̄�}�݋��?p��܏s�U�p�P���̭9���xZ��ތ/�돒�w��[lZ�'�u� ��K�����H=Ҧ�o��)5�R5≮#7W]�o�K���v�6�-�0!��i�:��52hJ�0�/�QV]ݐ�h��Y��\��7]�����F�4��D���v8m�)7��1��+�	0<!��ܱC�9z5�7��e�N|]�����pΐv����aE4Dg�ʎ5������Y��x`dvI��S�! ��Yo_G��z.�����1�)<w��/l�F�Wb)���Wy���L��W"�:������ڒ�s�y����,_��_e�ʑoa�^6:_�Q&�OYuI%y��wɮ�&�jٔ�2=�����ܫ�˥���(�H�\��`\l�(�!��`o�!�됝ɳ�s:��i�������*��J�+�S���y� ��7�Y��0�h�!S[5x�����RT~b7Z��9Y�Ci�����	���)M��	����tx5��q������7�t��4����>������ׇ��|\W9�,?�.���<KA�lz���K������䔙��nL�u�J6ؿ�����SK\<��#�Rӭ�4%L�MhP��0��)+#�6�Te�`�e�	��C���|�Tv��5֡Y4� GQ�QN.1G�T��*�K9O)���\�X<����Fm�����P�"��P�q�7�k�m��lKU�=BB��P�w��2}���QA�x�G�� �W��J~�yx���>=��4���j���2y��T|x��]o���*hH�\���8ol��Z�Y 7:\L ]��-�7��؋*%?���e|P]�%�bA���V#��S�{�*l*p�%�=>�)?ΣV�6cMϊ"���l�'��������K!�kiv���c7�"QL<�[���� �vF�	��GkX~ŠL���hY�j^��A�op^GG���px���}i���°~4�̐�� Qx#����\�Y�;��ua<����5N��ຆ��v�@4T�=�ȑ7�n�=w������ яg�F��γz	_�����n�Պ��;O��4�ۊ�8;�P^����Уp��}�Y�6<q<��Q�{��� ��ɔ�2��p�����dm`:R��R��p6������ͺ����Ѳ�P�o�d�0���2Bh^�|�4��W�!����c�b�)^H��k-�x����²0�*z	ςe�Ays�g���7�aK�鼗��4�␃u�z��F�q�Nv������s�Q:BF��g����b�k�ڣ1��q��fP5ޡ�1ä�M�V}S��js�	�� s��?�z�E��+\��4u�U
X�Lz��'+Y$��_����YR.�l4�-��9�W`Jפ����Qc��o�|�i'�4�r5����H�M��]���8VV��;y��V�������|������N�cF �����xY����{��\k'��<?^���SG�1�2SOR^7�I4����24�֪��r��h{V;(~a�1<�c�N:����ž:-�mh���w��0\kR�.�,�>�F+����j����iL��fMj!W]� z�?3[�<�4*\C$��[耥P�>���v�^�}�D+;�~k8���[d��o3��k���F���[�]���Ŝ�d���X��k����Q�0�(`����.�H*�񇟦����p��g	��A����RL�8/�XAa�N�S.%'�4ZR|SE�Fd�`:%[�upgz{�MȄ3�}�U���	�YX�<���S��-�Ğ��1������*k�B�����y�o���㭫�P�xmL0��X�Rz��^�#�G�5�x]G��2�"�9�_��7�Q��,�	ﮢ!r1�*}�|���z�1v�T����J�\��?���_o������*�T���|	��U3�o�F� !:��գ���.
t���^[fV�����ʏ�.��w��V�Q��PC��~~�������ƪ�JX��;ue^}�o�[�=z�����|��+Z��4�2��$nt�\(Ք+�t	0���w��\���o��`�7�h�v����J�����4R�f%�F��b5d5�#D��������O���1�x������q�+pr����@�����bʅ�s��J��>�Q��\�'��V��*`M.OJam|Ye��w���,��MӍ��?I�I�F�l]�u�E�
�X����kX^���If-Y�۷�������J1�I����xI�:�  @ IDATp ��й��4���-��M|Y���lQ֭�T��T٨�Ȫd�<��s�F��-��G����V�޽j��Ң� ��Y�6��;6C|��5�Y~+��FɌ����G�R��],N�$+�h8�����Q>6�]���H�V��_�=�-�4��J��=}h�إF�L`i����mo�ܷ�3<��ɠho�﷣�.��6Ỗ�'T���	Kr>^)t����~�L�%Xsj�/a0� ]��i�ϵS���|����k�����j܋�0:��+���t����2���^�6{P�z�R����GiI��+��֘�Ž�q��E�a~������^X�z�*޺�`�\��ת'x�r�p���X�}��1��zr�ɺ�c���{H�ۮo0-k$�4�����i��]oO�,`�qh�Y�JaS@�$�������HC#.d�a���OL��V��:�<yp�����y�G�Bd���c��՘���3I~x�����9��zǬ�c�
���J���/,b��s�/Ċ�1����nK���;����s�������|�p��u��Ѭ�l���%aBQ-gz��/4��Y��]/o��r��O�� ��1�ZB��L����*ؽ�O�AB��sQϤ��+.%�"��/]��U)�!]���sܼz<�{mO�1/����¾I ¥����Y�%(+�۲z�ֵ�Hʪ�t�4G�g%��J�C�b��p א���y�3��&?����,�=e�4��&;�A�B�%C�8~ȓ@��?�4���ɣ����]C0<�,��Ś{�+���H���e�UZ���\�m�+�=��l.���̧��9��*$��V��uufz� F7|H�m~]���:���ΐ�x�
=tD��w�X�(,��-�A�N�V����;�����5.pY
�x��y�U���?����tn(��
��ݨ�jgJ�<j��?�®�R�4�c�P'*c��n��7)pr.X��=�u����ʋw�]W9�[ԁ�oߜ�BV����O�GiZ��t}���~�ӧ|�	g��,���s���ϓ�#\��:Xӥ�rN9N��Ą�ߔE|KT���r�ǖ�B3nx��:0� |W^���Eg?<�\�D*Kk{]Ih�gq�dG��aO1*��\I�7&v�Ru�|��"��^�s�<ϵ��N��r1z��Y�w�����h�[y�����?r�F�1\{!y��ס#��T㱦�A����8
-�DG�D#�eލ��^���rʗ$+��,��Áf�Z���E��?Ds�7|������\h�4��B���skp�n1қN����/Fl4�SЮ�/�M_�/
0yQ��\e3��S��'�(�(��T�T��W݋FGޜӕOD����C�g��uY���,��ǵ����������o�q{{��Y���Mt m��^C���ʉ=E���C��E_�Zj'i�&��Zq�A��ɣ����c��4�O�;V��,���.��'� �����<�l4���LL�l�i�`�W�1z���e4���!)Х��$i5�2b��� @!_fт �Z���}zTN,��ڳ��.&��~�Ne9w���̟������03���>�������u+�~2[��B{�!�g�!��\"R��N�'E�F�ŕ+1'f!���z����i�)��<}t�_�?r��.	����g4��ǂg��w��¢0v|�>�Dz+x�=��M@�guz����y����ۆ �rn`~o��/'wP
(Y��W�-<��z!�X���w�};����lâ#�J����)NU��56
�Ț4�tb��D�B��o��x?�3߾�y�g�߄*eOP����S�p����70ä���v��࿄�
%�N$�(xevx)�{��4G��֬��1$J�����$�G���ɨ���@�z�$�f4�� ��܋��v�ŉJ:���(�xa�X��-�K�.�Q�&��E�x��2�Ka;��	�#�]�	��)� ��ۢ�YH��G�E[��@uW�	>!S������VD�k��`ǨwYF~J9�\9��"��6��z�4�=�j~p~(�����+���^�8��:*��nu� �/Xh��Fg��G0]<��z̨�=4:���vv�{�ߊ�;p9��o��L�.�y����X��JU�����SZৄ9�X����-�h,e�[�Ճd�\���XvãCw�"WX�8ᦤ�v�������L11<IN!�2U�!M��hhmup*��WoɕT񑝣6��{���b(���O6��
J���o=��"[t�����Y�W��5yR�����T@����ߴ�ACc�Δ���ʫ�VY����7�a_aCY$ˣ�Ny�}����&@\Ȃu��K�h���ڪ[�o��gW�����n�{9�,�_T>���G��5�F.�M@�mFm���Ɨ�Y����׆��yx��,��s��ɧ�7yxY��_���sqI�I�����Z�����W_�_�][�����z��A��hۡ,e0ʪ�{�`p]'�������OF��+o��%L=��<*���P䝇	����Y.���x���Y<��E��knƣ�Y���U�S�@�9ĜH��A����L��R�Ű�7,	^��u�Ƃfva��_��x����i�|�h��;?�p���o��x�M+?�������|��˯f�~JCD��AD12o�p�
���F7��zG*���4,5.�L��͘�ݶ��ǯ��Y�n ��2���a��/�m���d
����?��������û�k��{����'��ܬB����cb&T�5��Z1b�/OKH���,�F��71�a��v>A|���'�?<|�Ż-�`�h�����
�7+�e#fI����)�>(^�����o�_�/�Aֶ��b�ZV�_FV���Hؗ�5C����;��Ɣ_W
���xx��JR¥�n��T�3~�)C�,O��(�jHǮh��ྰ}U��kz����w�%��G����v��FT�:Y�ш��P�K�a�(��������7�����?�d0���^�-ó�g��8s?<�y�:Oу���rthlWCUz�ZPC�k͉��4��)�¬���
�a��s==}֎u��܁!w盍<�-���l�����X�S4M���ʤpc���>�E=��݄�U��mZ��xM�#��N~���Z�a����o,cC��P��=�⸔�n�3����<�s���\EX�>�~���9��n'�`��%��_�`yZ�����;�k�r���{)S��^0H�$N��e����ͺ�Ko�L��;�J��c��^�P�(�Sx��E�\=^6K6��gX,��v�:�ر�Rc����,T�V^�L���ʯ����"�¯ӽz��)+�;b��eh�<�M��x�(��(#�}���\�K����X<�@���Ƚ�f�����ޏ�q�R�d�۬;����+�bX��f7+؍ç��v��w
Ut������&CX�2��,8�|��/N��-�)Y��*H��hx�1�܈`0Ôt�^�Lt�����Uf��XG����g2� ���/]�r����s�����V��$���5m3��U��j����э�˒;�U@�}�<��巄/W�W���t�_�.~���(�B��P~�_��s�5>���k�eWge�^m����У��L��n�B��&�qN�M=�}m�F9� ���]Ĉp��~�Z�f�����4Zd��f��)�t_�Y�9��_�G�3V�2�띟F��U�7_���x��~?k,�enFO��q�ED�G��)�q,�_�@�1d'!�*�jY�K^�aJӭ��o�_��Ь1��(h���q��)ORy�����-]΍
���o���>�H�z��Q��;�'[t���jţ�5�����)O�F(���$��d�=��7�f�JB�i�k�ɰKY�.N��%%�����]8|����Ƿ�>����;�-�4�2�՘�9�brϻa~Q~^]d�v~���8ܾ���QK�5���-�x�H��C9���/#
�ߔ�R4'~S�g�S��Lz۬F&h�ʌ;
_R��MP�$�Y�"��%)�A	ש@�9+%����FK4M�V��P���rY�Q�`�υ��U��ëꥨC�~փ'�D�2�����O���;Ǣ(�uo}����xқD]:�9�wLw`���QV jF���m���?��
;�v/�R�i��R�ltO)0l-����az��/.�=�&�Ļ|�$�KaJu���vx�2\f�k�8���N�\���1q˗+<�p[���*4Z�ʓ|�N��,en+J;.�N�pxm�ܳ��wu��֮��0��W�N����������;�X�+d(x)�'�s��m��Q����N��s�S��y������;9�GW��(��k��}-@��u�-���ث���3:DY�/e�9���ۂ�|������"o�ꀣ9
M�~����~�ZNo�]�Z�Ec袳_�+_�����NL{W���B�\24���0�5.��<C3���{y���op+<T�.�K,�Yћ����e�j�b�O��}��<�24����2͕h(R������\,L�x[�C9�&�R$�<t���3c*����	�E�x.�o��7�q�M`o�,�*����Q�p�%�z�z�hZe�N��;�k��/�L�q]��\��-]r�Z�K4B7����_27�-z��J�C��]��x��n�^�a�gaU�ޣ��$k���"aAO�6y����{�F�׬���(�~�_�´ax��� ��z��c�h'�*81�G�w=s!A������J�
w��V�z����eKC<l	��Y�ndA��Ï�������ߵ�^��Ye��m�.3�G�b�Ic[�0�@8�ϓ�8)z��`v	�U��}������Q�^����5�NLV :K׫�{�t�������徿�_�������������?}���ΏߏRU�x6������U����f�@����S���zQwM<h������Z)3�aR��M3��NK�T��	+�ہ;����,V�t��ƲR	��,�*�a���>�;����
���=j4zߤ�l޼�����m�z����򔐰<�[��`C�ZID�c�wݽ���� ����>e����u�Q���W� �j
^V�f.�l2Ƽ�-N�ȇ㹙��Й"_�n�c=4�i���h�ҍ����wd�<��#~�.�*�^��U�u�g?����U��1���Y�\�����Y���Y�5��΁g׵�
O5]�� �Qr�f����vA����A��7�3�1���t�R$�����Z��a�hRR�`P�,��">1^�W�մ�-Í%�ʫ�[�5|@����2�]����y^#{��K��;�`���>�c�N�Es���a��n[ռw�#:-�c���躏���ȫ��m�����	�8	�ؖ4q��qv=�8jB�@gJ��������b��w�X���|����]W����釶�P?F4M��/ř�X��HO�p,�:uc!��W��_2��깎Sۈ@!�8T���J2K�b�qf��ԥ`���Y��,Z�k�(HC~;��Ka�Vf�����G�(�y��⒢����ڏ���x��C������D�$��i�a�}��&�@��y��g`�.�;�7�$��0��/u�G^�/�O�%���[j�^���V�c��>�@��^ɶ�ReN��~�$䈦���K3��k�Ss˶@���)�� �7C���V��LnN�iH��c,��]Nf�m� >������j8��5vK9��B�UuDuqt�W�#����ɄY���I5ί_���Y���M;(^�-���� 3�Pff�Y��Ě��a���r���׸�(�#�C�>��$Y�r^��2֛q
����Õo��ո(P�)�O�n���cކō]����&��`AXc|���z����X�r"B�	�iP����1�{�L�`��q�'�)�[BO��o���i3׾��!�ϟ��d�U��A�Qb�k�[/�9��y�fK��ޯ?~��χǭ\L��|3٭
'KN��@��u�Q+�~��K�{�=�n^j��L�MBPQC.3��[-��0����Z󝒔����2��=�\���BL��-;TN�����\	�׽{���K -(|�T9V��n#��oT�!LE��2�"h��EP��K�@/���U�UO��Ϛ���}ݞY�8�����V�b1��>Oixf6��@��?�ܼm��9����.����ryf�Z���,�x�`Ň?>�m�ߌ��5x�ʛk�����Q F�����������
��%.��G�ޯo}�yKht?��Ѝs�U��Q{��C����b��(��w��!+��5����c��%gp�~Sg��}6�n��i�=SQ�0a�-��)����B�S�
����c�XB	O)�]��s��g�����"&�e�\<�t�SJ���������Z�(��X��g�(���!�u{�!��EW�!�pV�*���)��#�ʼrЈ�_�\
�ă/��!���X�w2��I|�?��i���z���b7Dh$yr�p;�OQ�Ή��`�kڈ^W�d%|���g���o�rZ�J~�)�gib�uN�F���+K���uʢ�*����� [���^�5y;{��{lj�[�P�}�$�X����x�vp/s1yQ>)a&�P���;I���2#G�/zw�3�<�Dk;��?�4��Uc�+>:�f���e�խ�V��Ћ����O4Rߖ܇��r�s��а'kM�ЍB��N�-� ��a�^��I;z92��w�);�;(~��k��`���#��ڪK�VY��)5�Pgߔ�������*���d(*���C���ď�M����ڬ���B����rFV�L��׻�q���P�(�SG�&4�H*��Y�®8��-�1-�i^p��aw�3���+�')	0+�=9i��i��7��G����V�O�5y����>�pzr�߄��5�L3:� ���0T'�1�U�F�R8�A!hX���h
��N3!?N��	 �~j���~���R�����o��`�́�|���Ɣ/U�?j��w�}�=��J-^�4��⮯�����3	��z���\O�>lT:��G��mgۇ*X��r�u�Z��ULQ1�׸�x5
����r̮���w�M#ŧb,��4+�O�hN(V!�Ǥ�
�2]�x"�UoXc9���]3}мt��d�o�xk5&�`Ze�@�Hք7Y��������o?�i(�E�ԗ���Vx����-O��P0i���T��I��y��LM�YJ�4Kh��QӸ����:�D��teQGb���W�~��S�1]�͌�� ���,�xaY2�E�ȵhr�[��O�p����P��1qL���4��]���A�t",��6+�U��7Y���ߐ�
8���V �i�|�l<m�M3}>�Z��Yzh�Ooh�����!,i't�Q4�Ƃ���K���l(�[١ ɧ�2�k֊K(�=d�����p�k�|[8�w�z��9(M'ep�++�g�B�)�>w�"�N�u�߂�z��%��Y ;z\�V,HEr��;�].�������p_u_u�µ��42h:q����mL:d���,�&dY��|��"��a���fĤ�r��/%�^$�l���Po�J�{S�K����>��~� �zv/�$��He1K3G����[]��\�zӚT�~�-��7�]X��֬Y�\V��T���\4,-φ��LO�
9?R��&9���(HB�0Rg��B�<�h�X���������,50��2��,��$zn*���Ⱥђ7uZ��^�]DS��d���cE@�/����X�u�Ս��8�^��\M����X��r&�o�.޾}+>Y������z`V��s��-�W�+�]�C��z��\��ڟ0�n�9�FU�cud�G��8~8��J�/^��)����֑_/������A���Ba�gp�垯�z��MȢ��3��m��Al��1!�L��-V�]�+L�B��:\TܫYUn7�����T�R�,�?=�!%x� �����^l1W�Vp(�p���y�"�"��˒`3ԫ-uqk�o���7?��i!��b�Hf��֓zUc{��fY�Q�0C�ر^��-�a�K`��Gf��9��Խ��_=of��u���<ߩ�S��D�a��f�/�¢�����^�ߥ�_WLC���T�p7;��X
�����^@i�I�NM1�P<�A�d� |�����pz�]z�)��/S&���_`�`(3�'l��Gq�y\��P+
�����o�6���n��^�7z��2:Z����E+�/�b�	JgJ!C;��ߘ�U�0����
߬��
r*�Jm(FIC�kxZ�v�^��J�u��SQ�="٪K��A
��+ܷ�p���	 P� p���#�`hY�c�(%[��1D�2E!j4���c���®�|Xܭԍ#z
�,��O5��~+#�C�`�E7|�E7+aoh�50�1'���Q�ܱ�<�s?�=N>JW�����V��;�z�����V�4*�wx߄��M�����0[1��L8���ݽC���w�o��x�_�;a�бn��://�{���2�E�Z�Vz�|�s{��foݏ%-^� ��O���9�S�W��z+ٕ2N�?��c��R)'Q�	�r<��^(M���&��^nV��N�/�;��f��6di����(�eS�?d�[.k+%9�g)��y,�)��űM�~q��>��l�wn\l�KV��pዏ��ً�����!��Ǘ�����_]5ɧ�K�r�� �O��oa:�*/�?~0��In/"G�!Vy3Ԋt$���<w�x��@}�\&��u�_�\)>�>��]m��u��Y��y#��7��~Q)j���`D�C�ua�"�dӆ�$��$����ob��5
�6�P;u���pcp�ed��#Ȓ8���T.�\�B1�Ni)����S�1�:�OCh��9��s�m�t)�㿩��$?�	-Bg��ގW��;v]�+<\�W�'x-h+�^w\�+�lY��d��G�]�Q��1�I�7��­Q��#ھ|�hA;Fޙ�O�/!X���z�'졊����S�&���@6�%���|@�ՀEĞ}'S��	P�6��i�㗓ՆB2�'m7�}���xwt��������;9F��%��	�P&n7m�����R�Xj��)i�R�l�a�v��b[�����T�[ͪ Mg]�a(e�
s)�۵f�ب��k�,�G��
145<��@a�*��r���Lb�)�U���9�2�;6����!�2��R�GK�	!�b�m�:a���z�T��ӳ�#x�e*���Y�����۷/������om���h�8���y�.�)}����"�W�%���7tCC	�-��@�R�I�N9�w���z�b����E]z�0P������eΣ����#7*�b��)����w���,��>ܻww�$��]7���f��;֭�EB!����9,��G�u�t���Ց8�Q�f�Q����ʷi��f	�:R�#��l�mw��_���z,W������@�5���.�z������:C�)p�Á�䏕 ������Fa��xƮ�ܹ��u+S`�#Kޜ��7��X����/�]�UF�7�l�2&��S%U8��4�l+v����,K��ͷ����Y��^>ܓ9���H�����ZF_�Y���V������Ф2�\�pd��z���w���a��cY����󃇏�'��}:��YF/_n���%��Z�͇���Qr�"|�UV�癍^ש��2!�1���t5>��(������*�<��:9�U;��G���G��%_(%��uT���k�+����E4+%2Z��ד��\ˏ9���K�,���}��[6�FC�����o�V�H�݆�6�*ou�U����5��衞�����/��~����Ky��G�Hy��bX�F�Vg���:��|�l�~5ڶR��o)*��J�V���!�}/3o^6����i��{��Wmɹ�P�'�P>!����JqgT��#ȇ`�'���> �r�3|�mX�9zV����ZD1R@V��3X���ҝ]
#�/�4��Z�\D=���:·oRw�~���G���7m�8�݅���YSN�p�t߳מd@���ҩx�A�Sm政��!�S6���1x�O��?s���/������x��* +���L��f*ؤ�sZ�4�y�]� ���L��K
RZi�C?�m������:��x�Њ0N�����1��z�C�P�0�
���q<�����?V�����ʽ���./�FS��ur>}��^�E
A�'&�x���k�3y�CmJ�,49���~�
s�e�/�V�z]�j���Мn6O��zO9����,�#{F>`M�̚3	@�G`�C'��#��*��ʖ#�?T��N(ǝ,�&����Ð0Z�*HaL<X����	�K-\�(,	��?�]h�埀S��XN�P�����q�ݙ�P/Vc�lU��|�r���?I �5&ڑ�^烶��d�{��;�>�)uJ��۷�;�{��S�um(_�$�M"1�⽔0��� ���k	�')M�)�vF�����bhzSw�jꃠ[)�q��FNxu{	C�Q��NC�����gED�,� �ƛ҅'V���(]�J�JXA>��yT��uuhuv6�R�4���(}�LYHOu�Ӿ_����,�MQ��	���m�C���m��m�t��Li��}��V�,:�hp�Y���ʛo�:��u��6 ����?�|�l��q]k�������^<�$�~�����{���hBҭx�B���?���>�g �:��������dy�zC�!P}d�T�n�h��Ω�O)�Z
�3\�M�tM ��si��7
rtKy�K��O��:�t,���C"�߉*d6���偅��O�NȤ�A��AiT��_[��j�`�=e����<L�˧�Q2����4k.~���ѥ%Yu!y[c.�!�X��	��}]�)G
�N�7�_�`�~\��R5L����&�w���,〞:?#���]ꉖ�����x� �'CS�-�B��k�%�r�7��tN^��Ս /}�uL{�1���%'�@�D�q)�řL�rb�- ʖA��t�ф�i�^(5c����)�`�g W�Zẟ�h �>�ߊ�NY���>�4��An�l�]!~�������AI+������1�bl�z<���B�$և��1�"ܿ�5_E]yG���t��L�m�,��q�����8=�2 S��юb�� yM�%-�0BY�8�����X�z��s��xMXמ;(!����
5&����y��|�;�2|4~2UN�2���y����7���`8��I%y�;���Y��V������K`ގu�VC�NÍZ�iqP]�S*�!��Z௪��j�|$ޘ
]~��y����C�[�y�C�)NV��p�O��%:�)�U��SP�i?Z(��-��|6f����L](ok�G�R֟z[|������<z�4z��g�5_�}[��7}p3Z>?��@^$)��u�X�X�����'��4����]�%��W���\�෷���9�nW|��b�5dcV׃f�~��O�?��������f��s9�E X��O��O��w�efz�͊o>���Q�(b��zy�����`���wm�ug�BStp	�nvn��QhJG��슪ή�����S�^6�
�1��hX�%,L��m>�z��;�W�v���7H���<Y�&}��x-ݱ86���"�p��P�,�a��U�t�NW��\4�m�k�]�n��U��u+:�a�w�#��>��|�����������q\7Ly��놻�U�6
;|�s.%m��T��U�+.:P&V]H���xuLr������	X�Y������)aדO& �ey���U�r�~J%u~�Ӳ;-:mY
��{>���o���NH#ё�`-"�ϧ�B�Ϝ�+���P=� [������~������RJ��}��>	��@��^M1������o�z������f�2)L{�2F�sgF?���t��q��_��O���9|S}y�Qؒ��s�S��8���?X3�Y uZ;G	����3<���1�c9�u��g�a��~�<���m�Bg��f5�����������O?��-��,u0��i�U:Ao�g��&7�`��Φ��s��o�}������I���
CI
�pT8���1�&%c^S�*8e��Lvߓ�QQ�*��9�^yW�¡�#��{|�h4��Â-}i��:֛ �G�ߎo�}��ر�S��A9c)�t0�S�(B�����1p|a�>�v� ��<���Vh�'�|Φ��P�.s�M�c�#�uY�~&��� ��"Q)C�\�GgWV>T�]����x9"?ְ�?�y� w�����+�0�<���Í���i��'�%rv�����|f���s���s
���ځc���7�q^�m��
>~��S��͔/CQWk�_�]T	^E���r�54&lUg�4����;A�|K� ��/ݣ�ƿ��Kb7�FA��*�p���G�Q
+u���<�NE"G���$_����I�hcIB�q���L<������	��<���T�&0FK��{OB�MАp+d�e�ʇ�z�WK|��f��Z��?���E����Q�o�c�(��ߵ���_���f������Yp��z�ر4�Fx��h?TW��!{��aE6�����]��c�(�s��_���A3y~��ߤt}��d�����z߷�*�d(��XlZ�,y�K{�࿫w���w�ޯ�:A�|��(�xOJj�ы�����A�r�ձK۩'�g�ǄP�ESW}_�v���oFPv��|�Y>�0��.e��g�V�C7xኮ�Q��l>'o���	|�czΥ� &@ٿ���Hy�s��������NW2�~_��=6���Ci���CyL���9��:�ܝ �����������m��t����,�U��X�&�C�(<y�����=%���)^�ƞ�9U�Rʬ�d����S�,#4r2K�唉��e|��G��>��M>i��{�<,7��rp��c���B�0qp�!��ᒲ�=e�=!]���HJH�\�{���������ǹ�ċ�>k,���(����IQ'�ܪ���8�'�|)9q����r�p�a��OR��Qz:��v?����ɚ��R�X�]�Q��~�?�绘�U���:��37t\���c�'{�P�*����_�����@y�{:y*�H۔x�3(��B���q��ۄ����ï�~~�4ך��k��o<A�ƨ��VYh�����P/�΅����: K[r�J�fu��l_�!<:�;=@S�כ��F���x��1�_^&�Iw�]GO�}�� ٣�Uw�=к��wV֕�i�+�����_��Y�1(��w�����O��`�OT0Cr�#,��n�����5P)<S"8�Gi�`6!h�8�:Fh�dd�ۿu?�*�(�|��W���{T������2��Cw��$��͔�[�<hHq]����نea�nf�IJś���ԙ�x+GÎ}����?H���Z��,}���a�p��ح�!��B�`1�����]H��wh_�G+Y!+��_�����S�E!�A��@S��\���p?�9&-��X�s���(g�ԗ�!��.X��|�)`皽9��wf椖�]�F:e�Y^�x#]8���^ή��y�w�S�R��	v�滇�>�<����3�	OH:,���Ͳ�U.kh5aP�7
4>�6����4k���͆�����|��|}&��l�ː�S��e�~�/^؄{�H�H0S�A�� ��;ӓW>��Es
��cʮ��ϱz�G��	(ܱ4��\|���T�ޠg��Gc�{�3,[��`yY�z�JQ���	_���O�$��s�ՀD�wY��~��c�,�9V��� PL6�`�m����#`��!����h������I��E�vx��Mg�@߄��N�,\�'���9��"^�p��R���ʣ����$�Ҩ���g�%�N�`�����v~J�2_Cj,���[t��3IKo)?���� Nѹ�
g�#V0�~�����O�0��ۃ�Ω�*�p�+�a�N�����8o��|	u�~�Oi��±Pb���ҠZ�>32s�(����������>����Ϛ�n֯�z�1
$��,�A^�B���J`����&�����O��X�+^&�=:Ξ/��W��El�8�JΨ+dڬH/��w飻td|\fbs�:�H�!y���d���^�����]oʫW��dc�,�C<��݇��3�[ۥ��R�Cn�<~�뇇���&�}���n�Ϸ|�|�x����y�|���=|3�+ܖ'�.���!����	E�XO�۴���rE�ű��E�:V)�����+�HĐL��t����wC��+xo{��(�/� �|h�}�VV�s.�n�l��C\�γ<��W�8��/��+��.�w?�֛������V/mՐsH�@�歸���,t�������8RMv'�E�?�;֯�#N�ֵl�v����~�ax�@����|�i 2�&��hH�uLak�4J��7��x���̌F3o$<���"�ShXJ�T4�=F� U�)h��U��"N���"t�V�O�*��Ih�g�^�d��>q]�|�-��NB�z7���b�%4�����4]��j&
GK |Y��͚]���@��%�/ue��N��vx���5"��(�W�C�؛�/�(ٵ����x����o>��!�������L���ĳz�����i������� ��p0LG�қ�\|�!�+	���+g�3��6̢~���~����Wxe�zw����tش��:�����{/��ӏ��o���f���H�!������/ʸ�������2>�����0N��A�m����Kw���w);�Zƕ�$��ߖ�S�
��5��3�1�q�bJ�=攆�c�x��9^��_����$��p$,W�����b�&�����i���w��ǹ�����|y�^p�l���CZ�h�V��0��V�w��JF?嵆Дkx�����y5ޔ����J�4}�Ѡ߾yZ��j|�ДY����g��������B��;����خ����YÃd��'���t�5;�e:YKNZ����tl������T�Q^��Sk:+�}l�KIgu�J=v�����ͧ-�a���*7�'��L�g����$*�kd@C�O�{�)��~8�,?��ԡ~Z}�����!�XqX�u�xXZb0���&ϑ�Ƃh�f�w�����c�Jv<K=h3kKi)�'n)`��X�E��w����ګ��[[2�w!e2����yu����Φ�J"^[���sh_���X�~xp.��s���ە��i\�[�ȑڦ�3=�pxS,u�$��]�8^Vrǀ��}��NO�O��c���\?(�?��n�~��:;fQ�B�}�^��4�|�k���9�ٍ���y�3�1x�@x�I�q�֊ݵ�^�}��_�5�'?+���I�,����q��ڀڰȝ;?��*֋�T���N�T.=0=Ĭ�ö�F������_���W/����f{�I9�[���U��U#j�ڰ;�쒕w���4	��U̥�A��FD̾i�)�	W��5CoY����o�A�`M�ߓ4����k��n
+�u���L^��|��r�f��e��ҍ�R8���7MᦔQ��ऀ]�.�.�٪�/��3�Vk���H�c6+.k�3�_��OJ�_7���'_���pC�z�˷���������]3����z������q�64��d9���h|��֧�~6�_>N��>d�yu���[`�a��#������a
N�7�1?H���c��������?�����?ܻ{?���GA�h�i��E�9�^���D�)�^h���O�=A�LΆf�X�Zt�j�	d
��K�Y5�3�@8~1�b��`����V̈k[x��c+%��FI����#�w�>�8;��t&Y�����,�����7su��\)2�	�  @ IDATx~+��ga�� gp:��������(����'�>=�46NA;�Aa�^\�,_N�೦�'����~:P�5$:!g�[i��Yڟ呕�����Q�K�V��F$̴����?&�3��r���N�D��q��^�4�
��Y{.���SY�^	���1OO�j�2y�z��݇՝�s՛���f'V�c�ExP<���0����j�Ү �f|Q=��c���M�f����a����,.��2�6���߼Y݈/Ə��6���������$���12PVm�cc����R/�l7����.VmJŞ<z��Ǉ�~����?�?f�©w�5�T�叔��D�������x+���46�hr�B~^��,s��It��J���/��w}�ū�x߾����һg=�����+�f�����;��p˧4�}�HKm˼�H�����N�݉�|�&���A4�L����-Z��4�"�����w�}$${۹@����*�qɕ�d���H�������~_�[a�6��/PZ���߳�Nn�g���q�Iʜ���c#�q�ӱ~�Zw�r�����|���g�ۻ���jr��۩���m�Ú�E�/㮄�8~��½ԫ�N��8�|=kW{��)�EVjwr:�ζ�)Aq���e�X�&�-8�/HU�#8�Q�Љ�u`�R���M�0�	G����e���/
���*�.sx��u��sY���Le�i��D9a	�|q��\��()X�&��bC��˗�'4��	{V�&Ew� �f��Or��,'T�F	O�y���]?����O���_��n����𭰄BTJ���欱�����Q����?K�t�_L�FV��kY�D���v>�7|�8��̴�(8�F�d��y?ڳ�x��p���ǽ��M��wa�����ǂ8)�^��{������:Y�X�j���:e ��x|2�
7Xq�S�Td���������������x^B���`����\W<wy�}?���y��~�Э%V�țoN�l%p��3�s�6�g+����!mpۖ�����{0]Ͼ��~/��,7��p|>�hɚ��ݠd��R��%�ao2�Pk��N��u~�d��@w�T���8�m G٢@<�"�U�^��)DfS�f�ǔ�+��J���=liiP�;Y������~[ϑ��_�,E�r8C��0�C��Q���㔗�Yd~��~��D�᷍$��Hfi�8ߤ�U�zՂ�o����%~^>>����h�q���dI���+�Cwe2K`��\���$��ri�^�@F��	��ӧM:(��Æ�fM[���j��EX�`Ѱ%;�����6�k:�a`���d��7���\�Lr9E����ʋ¢͡�~��Oc5�:~���NmC�)��$C��ް��@F��.�����?8�̺ym֩l��;������W���y�p��jY؜ʤ�����t.�G'y���1|��W���|���b�7�&|�"��2C��}q-���;i�<o�[e���
��e.��R�꿀p���pǰ]��:��p'NnV�w�����ެ�$u����L��À,@�
4�[��zo3&��0=}qzw�/j�t����n��yܒ_}�E��a�x~������A�RAP�*�Y6�gu��U6�`��
G�L��Xu���nt�؏齵cR.�5^_-8,5j�b1ԉfKC��y�b�U���1�o���;<7Pb��w�ߏ�@��	�7�Wa:7�hT�� ��Sq�L��H�g�F�T�{�5���Q+(A�!��J<��B�i�b��!��[�ҕ6s/�j��v�i4[
�5{,�fR65�L�~������M�}�r�)E�B�/�-����b������?;w��Ǉ%�<|�͝�/��w��_k�,`����dk����gŽx�BÝ/?|��*/�Zk���B����'94��пm�¥�8C߭���:������ޔ���V|ȳX�G9�-76��yV��=��Q��k 9��R �R3��0�'�3��_D_H��((;��y^�oKp-�;fgRϱ��y�0s;�(���eѪ��8j�v~����	β&����F��C��;7.󡔅��5y�Wҧ��R���5�q0�GX��wpΞ�-+ҳ�(��j�t&�Ͳ|]&W&����Zy����j���HgY�����N
��;?߭��|���NP��²�'��$���Ck�u��T�,:�ӝ_��0��-�z)���c,W� z�n`��b_�b��0������[�b����ƅ�u<k�SB�&n�<2)�l�NvǷ!�c�0N��
�^}���8��c�G��u�,i�^����_����]��iuh������?����yC�WS�X��Q&l+�l�	^Z��AR"Y�w>��������Z�	�);2vjzy ��5E��ݻ)�f,6�l ��� $�X�HE��w�Ͽ��m��:��o�>�*���f�lR�6�,}��%�h����ﰩ�3#^�C	���ԏ���쐶�lc�#"��vZ@=�S�G��\�k��"�u@�v<������$�E�#����$�_<OH�W�ɧ��<���HK�Q&C�B���P܄_���/��xl�������N�|
d2ч��j$�P�`z��h[@�LIp�ۓ�'Cǜl�x��+|%�_�,(s�܄�� ߞ��&��m��b�8���|t����*���M�}�%K�c�����|�9�U���W�����hih$X���#t9Q�RM�X*Zy!���Na���}�hs��<{��0_�E���Ꭹ��K O�Z �A���礴�^�y���Ύ��k��b�9T����_�0ed*Q�cm��ht���g54f:����P�_��|)��zB�e��������囆I����
?3����4�b&������-?�9ߔ��ǿ9��$�*aʴ�n����:���%�Ƈ ��[�m)a	���i� �%�EVjx�y�Ʊ����}�����������e���Ɖ'\�y��M1Q��(,e��ې�~e|*�c+�7RN�	�8A�f5�G���y�h��0]�s/W�c�Yy\�T�N�ࠎ:�r���#��}_��X�g��I!�n�G+��u과��J��
�S��C���l蕷[���
	��:g��:3��8���g��qR������93k~��,:Ū����p�k���G�¸�A�N>���c�SX��,F�V]�:�5&K�t@���z� ?I���7
�((xt�&l�%xO�e�+��(C�R���-�W>(&=@����9\
�桡M��j�yb���&�_~�Y֡����H��_Gy0��6Ys'϶���n&��L�w�MrV����s�Bn���]�X{�)�08꥘ڝgmv���{,������Y�>au@��Ɩ��ܠ/Z)������7�y��k�Ģ�-�{�0M�U0���B��;�ߞ�_�\��i�n�8����T�aY5�馍������N^hy��;�?�Ky�,x�1��~?!��p��7��?���wP���8�� �|Bk�l�����j���n[ {������)�sW��8*`E�������x��~�,M�s4�P�[䋱J�|��p�.���f�섽Bu��K|��v��5HG!9	���c�~Z|�~��c(��Z�vDO�Ƭ1+��z_�ĭ��6�M�cs�|�J��u���w��Ai_Ih�+`�>
wM�f�W)0�*�Q�k/9w��>�B�"�]��
���#Ay>����+0朆>�#��*�No^�{���}���)�ҙ�S|��T��wl���~	�.��|�b[]���6�p�i�	v�N\���
��'���I���?����Z��׆;2�?m�A�2�`��ψ$g]�P��ֈ�̔�Ӽ-�F�I��r�%��z*��+��	6� 1�,!B�����k������w�L�Gi�|�hh8jFY@�!�������og0e��_N�y�y����/�+��B�ȼ�ǣ`u	z|v6]�Rk�� �~����g���l����w����r������!�]
zV��V'������b�ő��������p��t����E�B��m�^9��3��
����Z��6�gӖ�M#��o��o�&�T[��1ez[��+))��s|yP����g�ps��#��_9){��da��=�v�?Hެ�a�fmfy�۰�?eQ�5kMÊ`��V����l]��uJ-�����rh���8���eig	��W�/��s��G���ׅsF��Ŝ)'͚�o�\���_~f��+�_Z�����٧7Y��Ѣ����:[83��a��y�0���l�lS|(Ĭ��A�e�J���4ܒU�� ]{�J���W���Q�<�uX_��`�r��!h|�R5�}�~ei���!lx�hx�b
��������ډNm3��i_Nޮ����M�L����2�d�{xz��=��m*�,��i˹����������c�N-C�}.@K����X7Qr�Y�<~��I���_=Kkt�d�,�֒<ڷ�ǆSYU�^hg��s'P9M�}�2^��c�.��}y���������\��уĴ�B�#Y0��uz%��y��(lMzR��YP
0����de�g
q�D��-���/}�a3��ұ��R�4��)`�����H�/Ĩ�b�E�>C4	�q�,�X����YCmǄ�ĸQ���pl�RC�^��p����a��'�\^��o���V��g�Ne!x����0�{_�*�"�Q�Nz�Iñ��n���Fѭ�%�}Ch�v]���As���D�r%5��Ʒ�B�ӫ��%%�����TB�a�ҷ�};����0���ǘ%{�I�`���=��2C�7)vа'����E�����Zok��*��]�H�}zކ��TY�K�x�d��	���(��ʭ�
1<,��4�B���2�ǲ�#�O�>+��/��N��8�V�`v�u@N����=`���2�?,lƂ^��t�n�O�'�ga-�4v����'�ql.�p�_�)?f�f���z���N�����1t��9���|x�<i�φ�"ܷ%]���{4=�r!����wx�.|��݁:�t�.pذw�<����pGYk���Q}�B]����X�B+�_���k-+����ʷa"Y�œ{Zn����bO'������f}��1�0�-\��k�x�j���fcÐF�޻)k��bu��`�&W))���:0�E�t�/�x�_=S���w�{��W�M��X��6V������Eio�lQ��BΔK�1Lg�1��u��8���#y�-�JZ`�hK;��E��#��[Z.�9���x@-Yg�<~;?�k��X8J��F�7�c�]�}�)�����hl��\��������5q��;Z,�b��х̊充sq͒�������U�VvCpߢ�B�U�[M���: �fDC�߽��O�/�&`EcW��!����J`�R�v�;�z;���`ւ��X�*���ԙ��[u��>�Z��n~� 4ҁ?�V�̲\����໏ӻ]��~����������O��rP\L#�����n�~ˌ�C�߼���Kux
�d���<�*�)�{^��+#���0ֵ����g1�*�Ys7��5��Y3�B(+�7�َ�n�-���e��E�X��S���zp���('�KA�k���[�J��)TJ��M�U�%�(�zN
g��d�7��c���}V-ȴ���90��l�0��$ ��rh&��W���J��.��z~܄ �W��gذ[I�q9V�^@t��򳾏/`��3d��x|`��A%iG�A5C�f��g���!�k+t>���rv&�qG�n�	އDQ�D�=^����������%Q�O @�Ǿ��M��}f���<"######����؊پ��e��հ�[c�H���0!�iD66S
��΋�*���PĜ'�m�R�QX�LO*�y/z���r����^�c�RA%ϸ����
���`$�	�|�& �C�Udy!��\����l��
� ����˂0����y����w���/���K'�m8�P����o+tQ��ǔFac�Q.nZG����U���W罕re�y�w/a���.�	�AA���ǔ�n��aMS�Ʊڙ"h�.�~7������qm|��r��Kt���Y�OÈ�O��7�o�.���J��s���noj�^�́w�l��n�m-��<ZʭZ<������~�%����݂º�r��?<b�}�Kt�y�"q�Q~���ɓ'OY1���z�0%��� ׬�,�̤x�'�_��N���ir�$����k�.e��b�3V�B���9?1}�E9�d�u����TT$7&�L�_C1>��o�Q(��}ϢLP--�������{�m@#8嗼aLcq��Λ�WeV�y$O�=��t�����=�s���ef��F����Z)N��O�<��ϰL��,"�o����oA�=����4�b�&gs~�Kۆ��,�����˜ϫ%/� �7�g��.�����ʦX�����
��~�T�݌(�ϐ�DL\�;c��f�
+%[�z�Mӫ ����(D��)߼��4}WO���K�����%�� \�D0`X�r>��/P+#?A�ߤF<�+Z��իj�^��W�}ű�(�H}�LZajҒ=�+"�aLw�E��9��3��ɤ��j2Ҩ����5��Üo|�!��䷸��_%�=�����5�_�n�y̐�+��8�{�6�j���^DWXm���*+�N�j-K�� 2�ơ+VB��K%9@ �@0�[��Vb�K�)∺����i�xI��e��*���o��Ϟ�h��6 ��d��[�k��g�����g"��l�R��)��<t�]��;�r�Χ!�C5�H\�'&�E%�!����^����N���8N,��"�s*�1��⨥̊X��*@�;Ŏ�|6���Ort�穙n5��
�e��%(a�a��9q-:H�MǰUV/����P���)˂��	�{]��_�k��L��b�_�!&QYx���dJ��;��o\�F>�ϓ�S�:�W��]��Kru�"M��u�--/��	�=���k߽�����_��Nɫ���~��j+F���4�"Wʙn��|>T�z�RԄ+;0_�a��OG����3�ˤ�΃���$���Ά5^+`����e#��t.�+��#lu}7�]����|΍����l���=��[�{@I^>1Y�x	R��%����d�mQ��
�҅zf��������N���%&�_����@y�F�*�*i�w%V6 '@���
��`�|�C�2�^���*eʡ����W�i�C�kn��.�7��$�;&��.���D������ji;y�X��^Z��2�ft��1�4�B2���஛�B��׃��K�i�s�q�E��]�����I�w���9s��'��vr����y���n��!Ɔ�}F	�Yǫ����=�?� vՁ�7�Lt�-��Яb%�ݍV�Y�����Pu�G��,lA	Z@W��9�$�T����}��O�U�š0�%�ʷ�*q�ڸ����Q�u��m�i��XO(<�ow���&:)�1$@����h�;�����P��+�I�:@ې��̢&�X�{|�@e;�Ή;��
S���('��~T��;����]>�d&a	<ʔh�h���މ{�ܸy�N*�.˨O��d��`���𴨬b9Q�s^,�2Ǣp��� c�b�w�ǻ0�K�u�O%2�oi�}����V�D�	�%N�\/��d�7L�0�����0�9v�3�Qp�h|�eέ�����Ь�V�zN�[	��T�(_%G���L����B[�k�l(a��U��..V`��J�[�x�=Fw�.*�w��YW���q���ޫ�Xi �	gզ
�K�]��p���j�J&�7Nɜ��V0�/��w/,3��2s�N	Y�
6�ƣH4��M��wo˘�^ҡ�~�9�N�q���-���?�ۧ���Oᖢ.�sD����Gi��4����`�����J�>�KNa��0l�.Vg���`�#�xY�s��?��[7���V�,��e^��v*U�i���V^��ҹC���i$���歴�o<oyM��|ɭ��P�Щ|���J���g�)��GL�Έ{���Ƚ�T:<6�Xv��?��<���kQ���a�*�-',�]
�iQ�P,ߥS����~����U� �g���쓧���+6+���M���&8�UZ7�W��`1Z�"��킣��<Y�&�<�^;m �|IS�ܯ�c͔��*x�e��t̐�
�4�<̣�uz��H�=�G��H�X�HOٓ�Iك�P��=;�Ν�B�toH���y�tU����$t�v7�{�=$u�a�T�驜��s�<��&�����I�đN��C��b�?b;��=F	�Z��KL�Yg��G�O�[��?��n��.�;g�1FlL���������1e�²��j��Gg�N,O�Snhk��S��*�P��c5�yA;���Ǧ��u�{�zy���yg��煦�y�xBf���3�X��k����++:��ԩl�8���E����D\�Φo���X
	��}}6`%U��eJ�>�%���}�Y]�z���3������_��x�p���O
���3
�����|�� g?!I>�1~�]i�8�������{,q2��N�_��H*T
 +��]�R��9'��G�h��`����������¹'*|jil���H��;�BϢc�ʄ���R2+Ct!s�rf���� ��;O雹k�@����B{R�r�6�i�|��3��U�Lx�l�Q��_�yZ %��%�fOIuRrP�	,-4��|�P����>�_,a*b�!2���p��=C��� �Ga�
�d���0�(R��_�Nhp,?79t�Q��"z �xJ<w�>��!�]%� �U�5�~s�f��J�'����W�PJ��O�!��:��?0��0��o��nx��y�l��|ŭ�G��g �w��m9��Q�����[�JE���'�΁�gxP����4�țy��f�>��mt��H�r�����_�˧���W�+� �7�a���~O������t��{�A$�aw��k>�7���g܎R�~wW�Y��0���p�1����5ia6�BH}�q�8^�R��'|i�<`��'k���ιו�ccȳQl���]��������*0n&j���r�*�ȾS�(˷~��.�t��zb��On����i��wglb���]�rCl�p6^%?5Y�F\�����u:�S>�w�� �+���:��c�j�+,Z�U���c���_؉t!�y8`(��4�#o���2���YM�Ӆ+�,.��ǣP�ΦηQ:�4zSEH#�Rȸc�B�5�<,�锇(��d�%m�x�(O��U��������"�I��U,K�Q9hZ*k��?�j�J�CĞb��c�U�G0�[�|N'�{�"�P�m��l�nd����hP�6� \m!��;<B| � ��C`��3l`�f|�\�Gc,��-�0�e)yP_VO�5�hy򓧮^]��������0"Su�V�:ʩA�kCH�
�x H�d����6�p�H,;	���o�7�8����Mџ��O�;�|�BnL&j�'���[f2O�%�Q���
��0��*A����#ٯ�^���8�w�J�+����ó��t�o+����b�� 8����#a�i��^����~��/��r�h�q�]��H�������E�F��T*�N�]�O�I_�ap�r�8���s���/��B����?��ϡ���$oZƇ���j%��p���� S=yOck8ER�$"�è�T�x������(�&'9HՇ?*�4;��9�	���*t���tmJ��_˿/�D�R����w'���f��-,�j�o�eLE(G!ll8v>��<}�t��{��E:�"����=�=�����#����6u�#�o���F@y����^;*dG�2����gy��r`vN��ѕ&%�����B5����'oZ┫,2��B<A/W���=��hX+�L�`�4�B��3��u�FY��69p��+G�t��Pg�#&��*|��I���'n ��Λ��U!3�5���/&���ˢh8~%m�W�BT�~>]��{6v^��ͷaJ�]7�n�xF'ԫq갆��C���2p�p>$q-��R"~^²���t�-�·�U�p�w=��"6P��A]Y�p��:��hy����]�OQ�ܻ���,�_id'�n�	��s䨓����ON>�Nv߿�|d.�yY��B]�{�}�W������4�nea�m���]eu4)h�q���_�H+{�ԑ�X�\���󮬛f]ˣ�Xy�Ʀ�����3\E�!��l
��{DjM����(� BDx���rfxtV�q6,�w�nT�σ�7�!���ByRђ���Nk�" ����89��0����\fQ��3�du��n9K����o�в�ێ)|h~s��*|N̷�*��	9����6;���c�B���&���\W�l�)���D)�6�hV�R��b{�	h�� �<*�=|�h�ʸ�v�{�nr��
k�8��N�J�r\V�Ŗ�N�{nyl�<[�m�_�L�˦&O=x�����'�G�����8T2��!�
���D����-��%ec���o�\���C�|'��}�2<��Bb�@6#a
XF�d�4�0;e9�dޓ�2�B
�h�`�Jk���$�}'��|`�4wE �=𵠻 �� �T&}�" �04�ۧ��ׯ_�>��nE���C�r.�L��h`͐&٘�ɳ{���a"� ����$~�7	b�`p��
+�ᢙTt/�� ���,��>��R��]�'do��2�C�K�f,�z�O$�Ƃ�J�Q��8׍R Ut�Ţ���S �M��s�Yp���4��6��c��ζ읋E����GWL���x����Ә�����^�bӀ�"t�{�H�1L� ��t��|;�OK�k�@Z>���` �}� �a���:�)n�f��onO�� �����[����{�F�l��l�w�PEh�P�!CTs����4C	��+t5x�)���p���5�V��K �?Jv��g��4�FVA�yx��3�
3٪t�k����P����ǗO�J�T�T8Pʅ�������
P�J&9���5.>����633����p���޾�?>[�R�w�+u�p6��k8��4T�Z	�4R/�DS'[��y�ȶ����I@�r�W������t\~��'V�ߦ�î�lŢ�
���6��J�1Է�m��0RX��!�sW)��Px���?��]��١�
��v�';tt�>�D9r���k�K�9��I���F\J�f�U}�l�`u�c��q��v,�[X�����ؠ���*O�(UF<
�wzK]��egi���ޱy�	v�_>�z��)�2�:���2yJ�������q�!G-r6�*%˔����W�S\��D�@?Ş�K1�K�"���8��gZ��K泂������y������\e����2�����z
_&��9w�w˝�D�N��,��ic�Ë�=8�	8%���:_
�bOI�H�K�P����י�a�v�m'r�|a�0,%勍	P$�C �&�p,�؀R����$�}&�;��!�(`�eS1�vNe2y�(��h� h�$��P�%��/eU�#)'/��s����!�/��lt��ixS�p@<������s�*c�E���f�$Ñft�jj�426�����"�$3�g M����W��VS��T�(�!s`XO�/�}*�'�?�ܿ���%�-rt�)�q���]��&P�rkU��n�+0��6/��/%�\J8+a5)+44�'���i��1O��+0��� J�$nl�x�1x��ɹL`>yZ����V�SY�/I|v5�`V���T�,Ky�+��t�z�M���*]���y�9��)}t���'��I�$�<��*Dy�?���]��
�_�g#(�-�<�'�|��/�d��s3��=d-����	�Lf�I�_����L4�S`*`i\�WH��W�\g�����'
���j=C�ѣ�ˤb`*�ȹ��g��%��T��U-y�I?ʛ�Po:�X��{��AڔO���ԩ+���o��5��w�?�c&����VX��/�Bk��0�W�3�v�H6�2�^~#=#����g�3�	��L0ˍ�M�L|�<{�}�"�����W�6ĥ ����jZ��|Z˿���+S�-�]�So�(�U���o����u\����̯,fZ�׆����C�)f*r��F�\l֩�b�ۗ�����F7���<�;(_?�����#�w
wpp�a����-�����R?���66�¡�B+�%|��2������_0~}�|��m�O�y�!>�s!Խ{��[�Y��
Ie�5�-U,VQ��L^�"�>M󔣉�}�I�w�c�3�S�y�',ߟ>�a�����`!�Q���	C{�����=���o2��������s󖍷JL�r�=�*ݶ��[Γ����>���`h���oװ�����5L���K�r�$�zeCI�\x_�fG4xP��;�QЪ�^�J���:�29���a{�\yx�)2M��Z
F���Kq$�o��܆������He �f�������H��S~�+�f����VC�,dz��5
ބE��	��o8�����׮?N;By��/��D%��П���<���Ė�1�C�,�� _�ީ������4���
ڼ���$��7E[,�g%kJaC�!]u�$n��EZ�*��[)`�ʇq��f@�ZӍ�?[� s9�-��Ũj�C�Ԥ	i��0Ӕ
����?#�N$]��=�f�{)��*Q���Гt�xV&�W��7�+�Uk��*�J���٫�=<��yG�{�f{�e�'���N�g�����M�����j��m�,l�R)Y^k�=�G�+�wށ�?��U*$+�����^�T��� fE^� 0y���w���/+�� S�;�4�1�(��gv%�0�N��7��{��� @��J��!�O��V��o������� ����twѡ9'冁�B�|V7��f�#'���s7e炸����8�a�[�mr�/�R(�({b����i�w��>�no_��b�
�����J�p�i�L+��en2�y�t�ܻ��{�[ehұ�e�=���ΙA�C��K:Il�n�"���x�g9̮*}䯟U7g������oާ\3��N�i:v�K(��������G��A�����}�%�d����n~���T� r�%�BΨ��Q�a#���_��������n��dC��h uk��^�?��E��2�8{��O����5k�`8iSq+�ٻ߳�$��[x���h��37��6��`�:�#��g��@������	��ʜQ��n�Zz�����M&��+��g_�),eh��ЕͭX�D��숡1:ӳn:�㜉��L�wҺs�<��yAZ�0o�:�^��t��yh�]�鈹X��7$̿���	�P9�����l��p�f���@Y�F�E��
/���5�8e�sͮЙ��'���P�B���s.keh)�%_G��I'�0u��=��/yD����� �V(i��(�JU�Ǻ�lޤ+�8TA(�.�B�M�LE� ���y඲�x�9t���ǭ�2��2w�~ɜ��҈���㠠�e��m=��x���m��y�Lb��P�[�%Z���+�����,x�b���?D��v��zNݰ�D�P^y�(�|"�U,W��'ϫ�$M	#nMK`��&*�*_'�y�m�|���
m
��T�����]U/�	����R^�VPv��QO�;��I�_��MH�z��2�����WY�ی�$��X���;�[G�H�R9W�����"�q��%{�8��
x�:+3��f"�Y:�0��P(�ʧ�!���^��*2ɚgV2��;�ڠ{2�3wTg%��3�9e�2-`?.�^�����ke�9�9���v�?~� "��\�V�X�b�H��j|�J�u!�D�
A9)͚��+�_�:
���ˤV2�s0�V0����x��4:³r	���[�Hi�b����뻌l`�I��t�|�'|+�_Z��2�t:>Oa�
f�$L��p���k�
i����.�&[\۟l�C��a�4J�g(ǻ�ֵ�}�������Ϊ��P9ܬ��/��A�>��Ƅ�� ��P�<���M��t��@�=�bM�X���pɺ{I�s�ÊQ�76�'�ԏ���(d�7�� V1�A�2��VRR�^���JE�<����f�_e�24�>����S6zX��?�Jڤk�ʗ�0HM!n�&�Ʊ܀G��kZ#�O.S�i���0=_�˴�g��R���;P��i���k#�啺2�*,�U��c/��\,ݍc�Vr:L�i�I��u���^d�,E���iY+]���{%c�O��,X�<*��#`��eL%�p�W�W����� +k��|'�6.��\Y�l,�HЏ2a\�h>Tl����KW����j6'����v>�� [\Xw������{��ɪ
�h?���\�bC�P��ə���z�=:>�鈕��1Re'�;�g9��Q� >>�p^��`�k�.V�#d`ؑ��k���`�g���]8S+�:�
u֡�(�`'�ao��r�0�Q�hKj[D�ʘ�"��"��
����ߠ�ék�#������!�)[&K'�@�IQ�`9���6��
��D� �
��1�yb��)v /����8����R�}|�c�b��@�1T�z.�%/�r)�*�n�M{	%p�U��4��:�t:E~/��������~j�?��w�����nd~��Y�{�� ��
���� �*״��[?��pn�s�Bv�U�(`��2u�`�q �تc�le�L�O}��$p�\�E�3�DO��i'���a��a���]��5VX�o'�X�
�  p�L��]������h߄7ƍ�)�B��0B��b�?���,� �$��A����A� �C��'��X�~V�j~ q�X�O:� e�M���;p���c���@��c�S�p���4������^@0�(��V&PҠ.c�>� �}�Jf��dn�&
�>�kES1��JV��<���"�Ai,x�a>>Z�93�����2�W��O��q�Tz{q+�3aV���$܀m�m1�e&3V�	�q[敔��yB���=뷞�{`��`�ږ�R��M�"�(�cfOr�UVN�ux`���n�7�H�����!��!+�8k�t��o)WC	۳�vP��2���Uz���t��An��"��
�b/O�0�����p���%a��4��z�c��	��?dU���|o���MC������(y��O��<}��������UPfdv�.�^]��%�*o��^F?W|69�@�ɻx�\�����q=�o���t�Oi�v&����`J��#^���8N��\Z3�zk+��m�m>�YܦU)����ز��[��p��L�j�JX��������`ަ�Rz�G]�f��Ȃx���s�~3�xU�TŦ��W[[7���*���`a�3���A�*-�0Tj�������q�:��$� ]ȩSw>�/TE��[�G澋J:-Q�.�f�
D�Wo���fg���H<+3gy������MV�;�6@,Th�u�lq��w�w�{���<���T�A{�>Q���Gޡ�>y�$���a�2Ľ=�h9v�:{q�Y��g����8�X�Tu��4�"�f�D\���XF*��R�(w\��P��Wr��>��
��uѐJGtH�`�.�|;b8P�k�w���(�o�ud��?�2����A�ǲ�z!-�w6���|!2
��3�GɃ�����-������R�Ik�����S���EV��t�(/g���Yfw�R��q�K������z�M���� +�l�+���<��Z6�@t#|:��q�V��3�Ȍ������
핆��UWn� f��x��v
E��.&�6��l︶����ڣS�qҧ���q�7���`$[`�F]�`U�L¨�8Zo�F�<�b:b�^3���9-bN�\E����1��I�Nk°�YP��yƎ��f�Z�xf8��1u�܊|�I�ݻ��ߞ<c��p(  @ IDAT^�[�Ƅ��a�+�w�\�*�y>�熻sP<]^�˒�/*��H� R�
�n�K�D�)�1��}�jo[���'�L��.��Ĳ&�;�h���Mz��F��'j��� @.܀)#�3�z��ec ��K�w�������_
��{_�3�K�ڛg+����p�v�ؕ�H��*s��|�Ս?>b���ە�aa��
���q-�(aTD����;^3���ǿM^�e?"z���6�&W��Ln�=�����*��Zv5,�P@`�"��Tq��C����E�{�nޏ?FadcJh뜴VQ:_ ��
��Y��^�&��/q�'��S Ўr�2�'n����R/���v��܏eڗ8�#��w��iZ���s~
��:^租�F�w�����;��2�����s珧�xVYÓ�v�(�eUh�Ip/��}��[�U�Ώ�p�e�h6����F�Ռm��Ҥ�K��W��i4,��Kw�~H�;nhI�+k�s��/��Y�-By�&h�Ǳ����<��kC�������["sh�A���{&��o1��s��qy���:%^*:��;wJ�ҁ16R�(�]C��=6���r!�m��4�:O-��В,��E%�s�p0sɻx����(�DrA�e��?���?�Fg�C䶖�k[��ġ��){�g{�2dw/�OZ�~x6���Y����r����۷��~�9ُ�!W�͑J�G��1>�6Z�,Sٖ�o� r��� �u�Ӽ|$�J���>2��|�k}���槱eٸץG�c�i6s�a�c��0:\�R(��/^L~{���
�Y)c�M�$�E~�pd�2�5m�
��n�������F�h�R��By:�8�a���9��)�<e!�F��M �d���{�_�K;$ϻǻ���+�G.2�&��af�G^��dV뗼�tG]"K)��YZs�l�e岰����u��&��,�����������9z��y����qJ��!���#DV9�1yAӱrF�JL�ΙBaS��|hY��F
V�������^ y��<5��,J�®� �D��Q���V>͈��$fDS��`N�s��ֹ�gv����RVGR���S�J[�p���7�w9K����ѻX,.�v]��:���P��֨P�X�V�-���gV�P1�`��Sѣ�<_�-E��6�ش;ܹ��[]Ā���aI:ٵX���H2���aA��)� ��|҈S���!N�����2�bP�`eN��O�m�e�A�|+���jF�k��7 �^u�-�����d������ �:�m
n Vڼ����phR˧
�x��Ff������� m��heL������iun����0��>G`EA �'4
��=ZE����6��_���bFA%�E���'�|��+��LW}e@*JC���N}��L�V�Y�
_�ipH�6I���(J8]f���t柺{u�����\��t(C�R�A�N:�8��J�	���W��qh���x�^W�y��)m�F�����V�����ʗi(wT(:�~������*^���c4&�����.�XBҨ��Y<<���*Q
��
���&
�&S@���Z��#��ƕ����E�Պ�p�v}���C�40X�D�S'����=�(���0{��PpN��w#&�����*����;>e����ƗR���:�yf.�Q1���!�R�'3��p*G~�����M~��	���$�I7��v5<�I�/� ���'펖�X�1��K�������#������-Gi�<�]�O��lǰ���U�-Wk����2]���	�y��o-/��W�X���"�3�_��W,��p��w�U*J�(���c�4l8�*������=0�JSҘ[��wR�dS
�O�"Yn�%��l�|�� �2sd�Q�_p<����}��:ܨٓ;��O�m��s�j�#1����Sٗu������n�.;���p��"���
c�ɹ!��ω�H���c� /��� Yb)pѠ�a���m���2zs�E]�{�<��$;�`�1#�'*� ���uij&�[IRQD���/�L�K� �-1$����(a}����($^Wa�c�35�:���3���� �*f�!���� �
�̞M�̗�׆]�Z�X����P������o��/�M>!ղ�!a8�jݞ��z�X�����h�B7A*�V	���e��Y����7�w_*��x1}���K�,�r���⻔ 5�-9���m����D�Ø��
i%�� !��N�bd��^��b!��)����*�������M�)*6 ��P��z}�ǩ�<���0��L��� �
�dY�OcL�W���a�gj���aP�S�:B-��(i��9�yʖ~��/�)�v��W���p��V�s)Z
o{����Fr˷^�Y�<s�4��򐬌K841��oiHn� �)|K�*���������([>�����פl]���>��W��4�{�THp����-o�<�M��+��7LgXm��q�F	A.��W+>~��y�~�����^��<,�̈́�e�S�M�������V;㉏~�d�R�����g�n�ѧ��
�����ehޫ����_�i���z���]u�IG�r?�p.�i���U�w���G"�d�m������Ml�
�)��r�<��`Ag�$_ԧS�&�tK���d�]��9_7�8��I�����i;�ί�	����L=����	�z�ܷndB7B{����xx�1�~]�W�[>q�@��)�	����6U��T����;eW�X�����g�5��W�˘|p
�߼I�ʳC��]����^��ڍ*(J��C���(n��0n��o���,�x��c(,/�N��>��v��Qڎ���5��U��}����l�a��U�3)U�ͷm��Ϥ���޵s)ye4�<�W��0�i���X�.hcl�	�����P�KF"�P��0geSE�p�N��38�lys9��^�.D�R"��1�	�����q̶]QʬN�Q�2��V&�F~�7�&eۤ����؄�҆جg���:��1��liD��)��&��YB��`�T&+�h��.J$b/RB�G�,bj[RЃ��he��bFf���Ț?�-���W���	�F*N�!�k2���G��f|N��.�2�	S��ǧ�5߽Ĵ�#�3%A&�����關���ɳ�㧯��Ȝ/�/�ã�#<9~a�I~�"�E)(���,����2�)
J�|y�*���d�h)���3�D��w�=|�k%�r0����4?��h�/�8����x��峅zz0J�8�`I�
5��4d��o��h�<�$x�:/Č�O��=�|�ŗ�S�<k�:O� ,L�h�<����۠p_BߢUѬ��8�7I��ĥ���-����[N�w�UW���C�o�r�-�K���eނg�=}�|�ɿ�tbN��·+�]��F5M��� ZA%��TY�t���{��0�7�B%���y�i��.�r+8��t���I�4c�����?Ҵ�e_:��`�{�ӽ�~���8�7M���<n���÷<���RVh�3�P�K�sM&�����.�|z�`4���i���5>��_~��袿���*�V�ڽ㚮����3�v���a',/�{5���J��a��
礋���;��k��\����o�x$�J��"��xR�C�@L��� �3�����T)�f���-,J7���Y%N_e�0[�c:9;Է�__�fn��g%�3,�;XeT�,��P�5�ΒC�',��{�)6������ϞM޼}E�)"�W�)-:Z�=��y��(te%e��!���u�4�;3U뗊�a������;�X2��ѭ/l�U�̃i(w,��7��é�(�Խ�TU�c�V�)cK	��^c~��0�5O�MB�0p��C�* �W�S2���J��P�gn3���1{�iQ;G�/9�L����Ox@��r�[�m�m�����6�*Iy�G���j	%���J*���j/�/<�B7�%��v^��s��na���ܞ.��h��y��ŧ|�Hک��L؎���|����߅��{�D�P>ó?RF�@��'9T0T�4\(����Gxe7#+�����.+痝'�H%^`i�
��@� �����T�炐�d�P�Î�Q 5-_A��&�)�zӁ�䎲��l:*ZV�̉�4Y��8\T󫍭�Z�'#�Z٦U�����7����R��S�)#ib�G������_�:y�{&\Ҩ��;����4KĊG/���4����	C���%Ҭ�I4�P��Qq�.2�����N2C�A�Hb�K�K�z�ɞ#�a����6+�W �x_�9���O��ƅ�>�T�J[�C����-��R�(�f^G8�7.�TÔc�-���:O�QAC�Y1�}��U���@���'�׿��g'Tm�A���rۛ�ؿB|���s?�;�8O�z㐶�"��Q^.��W+�����$�4|F`�c�3si�
��U����7`�2(�y���U��k��E�aSX��aX�'=�@���uQ���T�/��9f����ٴ��%��4��w��/^�}7?T�R�<?3|f8N��5N�Æ��n�*V�Re�2��v**}u]�ؕy��S���~{��m8>�|�����-�V����J�0[���k��G@��86�i�����m��1��꫞���m��v�T���M�za�pJ_��
[���嬊�s��6"���<�4���M�-w׷ZO]y����[Z�_�|��Kq��U�X�~_e���V('�ߤ#t�yj�RdUp��WNWPArh,ǅ%�<?3�ǎ��V/yJ���������9�L?��Z��n`��H���p ���2�;�� ���9D*����b[V��le��2�I����<7J�`ME��R�L�Z%�:0���/���4V(�*眓�N���AN�gԹ��ͩL�{�6y{4��������4���.�+�h`8'i�js���o9(�0Q�����<8��0P�N���9�s,����*v��O�J=�&��8'���K������?�?�������{�Fx^CH,�Z���"Ǧ�NF���rLJ�qֲ*=͒�b�dZ�yV��V.B�=�2��R7����θ�_��<9ԫ�-��w�h�~���;K�ߣ;,��{�p����bD�a<�����ahM�*"K$lAY�u�_�$��i��5�E����CbS���J���6K�a*ͅVJY�%�nLWK]��U1+�{&��((���������-�]�>{9����A�R)`&�o���aò~�F���6�T.�Sa�B�����S�
6�zYYLW���$Y>�-A���&����u ��Z`�3N����4��#����s�	-�Dˏ�eJ>�X%���j��cQ�a��L:��x��%���nJ�>�*��\J�|Hy�|T���ۯ�{ ���Q)s�K��*V6H��Ge�孛eb�+�� a�2m�/{�5���^��ثV	;b����'(�;�%U��g���?��A�<�̬��V%�z��y��I��6B�W�j]���r^4�?)�|��U�.}ķ��9݄M�Jl��\� ^��n�ICO��,�����ɏ|m�.���n��Z���+:�����г��|�l�M�����\	U]*Ư��PD����5|c�j��?|6>�r�wZ��z���߭X�#��F�a>�7l�4.�\ʸ�Ư:z�tP��&�MIU^,R�q�'y���O�SF�O,�«�_��"�����y4�a�r �W8)��o�����l=S>�;νT�n�������U��7�nt��N�W���c�������T0ٛ����#�3�����#(=<+M����.�-��/�Y}��l��-�}7���L�wT��Q��Eǽ{4��]k��d`�ԁ�k�ISփ��̡`���`Z�TX����y	k�2���_�;Fny;m�*'\c��M�e%�a<�۬(ߴ�{�s�.QR�ky�C��aA�6����M������Mn�	�	�:�>a`p1��n渒Wq�I���,u�R_�-��i�����)�!��H�se1m�y��_ܘwm{D��j�c��O�G�:��p�M
�,nnع�mX�̫e��٤ ��f޴I�h���^,򑧏Ѫ�<�V��/y�V3��ߊ��@ k�~e�O���϶E�e���F��8��Wr���ׯ���� �!�!��;C�֭{�t/��Uz��7T�A��3jahf�2�K
�ރ�&�;.j��k$kࢰ�/��^@t?,:*��o!f>��H;�*.�.������m��_�|;y����9CKoP�>|t�-�Ι��j+���Qk�	���n4�*���<�)4�t�S`��౽�-^
�g\y���צRi�
נ�7�?_���{}��Jb�T6�w�*(E�����r'��8�$ 0m0�
X���_3o���c�J [����op�C��c����5pN+��"�4���S�(�(V������O� ��{3Փ&��`�? �f��\"ބ]xN�K���7o�s��d�f
|��`t�0��~��#��1�_��L�|ˋ������#�SpWSXF�aEտ�l/��"r��﹄#M�5O���}vh'�*�I2�޴�k�
�)̤� �'����W�5	�K��U��2������0L���Э�J��o7����t>�U��@7��#ʊVv����_�WڕH�ğKy��Yx�i	��J�4�0?�^C�_�T��ڿ�Ge�a��Bb�糧�y5��+/��߱�G��/���i�����6�
�S��C����q���H�4�g�RN���1p�s�=�*Y?�8�Q��G;5������*�2ꡬquS�q��Y�X9��Ў/�ЎH(�<��Uh���[��^[�����(n�a���� �@���<�
'=L�!�Cb�ʦ�	'#3�-W��|��{�S����O>��V��k�AkTћr!ҷFN�W�e�-�Ӟ<{J<&f#�<�1rya�;��}�E�-� o2�y�=�\D �3,O��ͩ�R�2���`�n�y�ese�j�o�?���K:���S�(Mb��|DNC���\�NQ��4���@���1u<��/*�.иd��6cò��K :�x,!k�d�=;۞	�ϩ����ٓW����{��c�ݛ7�b�t3l��.` �?@eǺX@� �OVX�!w���}�u˝'}�^Y?���dc�]]T�̡��GF�J�`�|��#�ې8?��1�(e��[��g���k��^����� �+L���JC ²��Qo�N�
?�7���T0�6��W�ʕՀxh�~geyy�/ʊ�K
�cY��$<��W+>�XX%�X��h�X����F�Pd���o�c�r���.����E�0X�,K�E,~.��x�Ƙc�IQ�+��W&u���g�ٚ���0��oV�feiS8Q�bۥ˻��׏/\8U���-s	�s��	z����8F�U�*S
��߂_�K$#J_�I�~q�R>_,��\��n�������������Ȧ P��VHe�~�+o�c�'\�o$�k%-����pr��ޞ�#+�LS'��O�:X��@��=ϰ_0t}�nߔ��l����o��X���i��a�8-{i`D��&��ĭ��KoNy7O)k����栍o\���j��]�7@E�	<Ǵwp��!�}Ϳ��y�]5n)�ԥ�|�����`�yP0^)�����[�[F��E������}/x�i�ÙF|	�����_��g��a�m��k�W�'@m���(e��W��*�y#�A���4�~��<���N�uY�+��!H��L�i�=[�Ȱ�tB��~ZO�>���������	h�Ȇ_� o�U �]����8g�a����4▍=Q�̃{-ma!������Q ��E���e���PT��:;%ALk�
��:/J�ICi��M�س�̟��]�-��X�\q]�hw�̍��Mn����5d���ӧ(�X�����[Љ�*wI4�|"�N�����I*iQ�p�>V��V!��Nr$ Z8Lɔ�UV�k1\pu$tvj�{F�<}�Ԝ�(�(���4��K�b��e������6Że�_xCz���K�Pjc��U7��ft!
�Dſ�S�tg�/(�.�p����t-��M6Ig���0��"��'�΂�^B4���~�+�+��.Xv���5:9���3f��u�;8�rq��Ա3^&���|�hP��'���DGA}�iMNm��,&�4|qbO p�
��&(���T�MYbnS��@`�?D58�S��:��Rs[w�]��;��p�YP�6���xbe�'o�矉����a��",(2j�5Q;���ܩY�ƫ��Y��!�X��I��C�*^3�|Qq�f]��+�g��X�X�G+�^���F{~��'�������w6'xxsre�Z�N
P��BSFm��:,!<i=ƕ<�} t+�ٻ����O�� �M*Zx�v|��HN&�r����"IU��?+��dx�;�`�Ц���05�;�(T�[?�;X9LWӱl�b�5�x68���ݯ1�/\��q�L��.n��h@|%$4I�RO���Z��0�;�ZFZR��2�o͇s�6�(eN�M�G%0C�/���a7C<��%���!��B�IY5��
^p 6�
o_���A�E��]����F8�*6~D��1���O��F_�:����܌g�^�^�|7��S�	4Ż��_
��o�g��s�7�v�~v���e�"���a}��%�v�A��;�C�3��G�e��򚺄�������cƫ���Ѹ��eܾگ��[҃
陏��Ȥ��=&�~��$���`��x-�xH7��6����3�i�h�3ٚ�+Okr��![ dc�kU��ZFI��������eK��Ǵ�#|눲�����V��-�h�o�yO¦�3Uf)+�<�ᵟ=��`�O����=7��D�ve�Uꔸ���\,�m��А�$��߭��GJ��TRh�T
��W��m���^h-ӗo=oVe�FZK��!�m��U��b�o�.�s�++��oq���w:��v��2c��@�4Sv���bO����ߒ}8��<U�Qi��P܄��o�'/0P����*#^�(YZ�����=u�|8��X������j	;c�t��k,n@A���:�r����:��E:�o�]�X�y� �X&Xd	�d����W�����Ï�#�;�D9T�!�/��mX�/�pY{�*��E.
��=�n�S��GYe4Hb���wyeu� �l�'�����y��g[� �&4Wn3ُպ,���0�@bj�rb���S`�d�N6�ي7�"2C�v�����aA9a����D�2(a�g�p%,�4��;Q����8�~�>���|�i��D#��IS�[N,16���iv�9o2�1�;����|��RdVV҇Y<���i�1�.�^�<�͞Q�[e�x��X��Z���P9�W�-�W�we��& P�a��5�]i	�⎆玡���_� 3z&d�^���2<�p�@/�A��s?�4�D>S���w$�>-}n?M?�!��>����D*�$o���3�i�c����S�U@Xړ��}sgcO@�9Y��19��|<���Ҫ�X������H��iH���y���O����1.��,6�۷R�����2=^�C��w�����e�]e�PE�����~�G�0>�ֿ�}7^�z�-�Bs�(к���hX��1F�����׫a�����t�eg�����@�8U��W��*�\�7�W���p�*yJ z���U৳d�`}L)�T#�ʙH��¯�W
�2�sR�\P�h�1�F��f�o�<����!wb|�����K�<e�-�Zgx(�2��H�Ќ�rҶ�5��7���PF�@�����-�r<q��2=!-�� �ݬ[��UFk�PJ^Sz;TKO���O뎍W�>�l�R�zT�UY|H�l�Eu˹7n4�	]6�$��L�
�,T��K��;i+b�m'�r9g� V<Z�}�<��yl�k��B�A�⾎�̹f{�.ݝ�Q�d���͊s�o��%��⴯��J�h�4J��}|��A�ٷl�=�(w7I�D�:OX�EvBC<�6I�h4���8|�{�)�$�}��Ӆ���u	�E�P�U/��ʿ*����Z�ՊȤ�6�}°Н�c��y��oĩ�M���#&��jQGN@�i��ֵ�F�\�&�S�&����.��
Y�*E��J�����
W�x�Q6n�a�����BZT�-8ӓZ�����O�[��ZqĈ��%�=�[xTݖ�ͪ�q�+C�bn�B$pz:�a������fZ��`d�t��\�Z%j�������	��oD�e�=_��R�M�j��
���Q0�rJ��r&W*�=4����T�/Q`h�V�
K��%Ll%����=(�o�rWhͮ���MP�����2�B`�����b:^���FF��']�{��2����B����e�ēYɛe  n�rS[V��=�d-�$g���^��}�	;~�Vf��?��ި�hG�4�� ���T�A>aW=]�U����r��U��sr�q�/]��0c7OD����N�^���G?<�ˤP�2���jLWf�)czt�i�)�/��^�x+�@��J�z�r���ZE/I�e�e`�*Ǌk}J>���o��&�I'_F����ea$L��K]�F7���F և�0�W�����&^����[�!�	G�/0�u8�~7,a��nZ���o�{ux�ۯ��[9�-����G'����V��d�n�����-��޸��9*�����Ze+����r��+�m��3J�B��9^|�mD<.����F�LH��/�8OI��V;I��e���Z�O�Ç�ɣG�T�Fg��'�X*��1��vv��rW�!o�ogڡ1i���'Up�+s�����_V��̰�T`\���:bՅQ��?p�|2�'�J7��7s����S+�A�	���?�̜a�T�M����>e79|��;�Ca��v�����PF9_��2��m����*���7�s����9���(����=oVY%y��F����{e���
eR�5}V(Y'_�fd˥��]:a����1;��q@��ݚ,���&����GQ�;��vB9�T
.1�\:�r[�;)Io�I�����m@�I�O�r��U�Q�� B��$m.lc	O`MN�3,� h����"��PI�!n)��%+��i�c�X���;ʎ��N�;b%^�iE�8�o���P�I1�� k,ZFv޵��SZ�����Z��ڹ����	��"��2"PQ4�jˇL2>�r���;�0S� � �9]������O)��nΩ)�e�!�BnZL� �b�#�2�M(�h A������Y��C��QKC�9:��g]��\B�rr��r�!��a�T`�����CM��G>4�Zq͛w$Ѣ�x��Z�'�k\ޱ�ʫ��X*Rx>�4�R¦��
2A ���L�a�M�R+��0�t0�Ἄ_0J�����I�ʆ�,�(p̏~��t��/LÄ�|�{�	ůhPU<���|��U̪�� U|݅U�bѠ�(�D��*�j)�u>����HYZ�,�%�ޗ�a(��
����ۻ7)R�R���͐�;�7;���3*iTܜ\�Er�Ϡ� ߍ!`)+xh&�ӛJ��cY�ws���(�.(�[�J�xE���H�h^t����7l_Ӳj��s��@d޽���������O��{Z�)�9_����^<l�~χխ/�;N?�kw�uo?q��`�Y��i��8�խ,�ǳ�6��w�u\{��uq�y��ƣ抡����:@�1�q��怂e��3�$�R�B������u%�I��{0�n3_ȕ�쟅���ݍ��]|�.ei)����D�M��XEZgD;Xn������f;���8����W,��x ��X/<���XZخ��r�y@��l-���o�M�g�!=&n��"r��7�Ñ�i���?�:��+�̦��7,x���\���������E(gW�V��~)�LV:؞e��I�N��(��%��JOw��Ӷ�6HeU��:Dy/��_B0��r����9���t����1��w�_���[#�ƕ�(��{�]�m��w�,J��(��Q�C~x��*���6��Q�r�_���%b�|��hX��@���C �Ӗ"Kq�=���S~$�m�`��|U�>�g�B����´n��c�D�+�m����:�C��-�"����ᫎ�`��<H�o~�+\�?Ƴ[��xR�rʓwr�|w�SA������F
=�@�
��P�$��c��
~�����n�> �Vb)��ef��L��n�	�
�"�c��|�w
��i�l	��R��0��U��%�Qq�#=٥B/����ͭ�%8�|/w�_��,�Â�ͬt<��O2��a%�ְ�0�� ��U�<x����$����)P�և�U�V�3��W2�w�������;fI<�-Z�^�V* ��fx/�e�����k����{3eдl�q7 V��|4��g�Z�����H�3�U��E���ޤt�QB����|�BRy���%��<��)����;��F� !��pw�sV�,#�Uj<���L�Xc%�����9��v
�
#x�~i�=�����Q��L�1�NzJ)���W�vӱh�b��<�0�<x�kf�!���tWq�:���~�+<a{��0�޳���p�p}G>/���{�_���0��;�gx��|�_��S��U��k8�޸X�"��>\�m>�v�Ooi�e����NG�����{[_;|��qS�r��4�/�V�M_�e.f���*4v\U`R�M2�(OKŸ���T��#�*_��W�ׯ_��f��� @��dbO�p�]�{�X�i#P�h ҩK=��>��rt��C��3�)��RssU�Uk�
�\�bi�YTA�MPQ���]�>��m$@?��Kl1��:C��9�3Cso���y�O��,d'��wnL~��a��V	9x�b��91�������g":q^�[�]H��y���-����*jT�dY7��m���͞m���X1x�<����8��X~�!�����uFm<ڈ���"�?���x���d?K;uZ����m<����s5!�2}����u���㐰\R���|�#���w+��z��96*c� s(��]�R����T����Fƣ�J�t@�H�gD���w�=�qM-��o����V��״�K�T%�p���a[,K���,:� �t���qS_U����k�nHe�X�Ι��ǃ��m�.��!�?��vF�S��=V?�U5p{�wtޗ���2�0���-R��jc(A�2$LgO������X���+HY� T�(_0_���p���~��Hl/�f\�4¸

��=�F0<��\Ǎu���׆�4�0�?��m㍕ޅ�5L�N���.�B�3\�wb_8-^<�_ �~�< L���M���`e��w�o��H����;�u��(���0��m����CG3��*�x�w�7�+,i�m+8�q��a�z�/�X�eO�����n��0��+~�I��_P*��H��)Pt�L��N�J��%������a��ƥ�P8�H7�=q0y��Q����i�.�v�F�p����wƉ�;1d��f�[X��)(z���qI�(`���R�i��E�r��
/qB���I�m=��X۸Y��׆�xQ4Nؔ��s	��5=�Ǥ����5�oZ�g����U���K�}���4��p����B��Ȏ،[(��O˶�7�^`�ѝ
c|yux��.���i?y�� !��[��-|�[����p��2n%��Q�Ϝ���T�J	�����pM�-N<�,�Fs~�Ő�]6!U�z�����٘�m�C�טc�5�	Ӯ"�=iPg��J������� �����L�^�~�m��`w��F�9g�P�Zo�P�T.m���ez�,��i���X<f���3�6ω�H�Ϙ�,�iR?��\ö*��/:,<~�C���٩+QbU(C-J��i4��ў�K&Ż�{lE�A�_%��%�BH��Z���N���5U��X0r��,����S�q��8>���%啓˕�Z����E�ds�>�I6�ժ��|(�N2�U,�lT{�i���1����	�OΘ���&|F@2ej��
�v�w�:�zSz����u�
��jd<�:�OlcɼC�*�Z�l��T��,��"���FhJ�������� �Vx�+��O�<��5����r�R���{�~��pj\K�㛲0�`���A �6�w�K���@/�n��g-;�~�Y̭!N)0����>I�@��1C�c�T�V0U
�BT�6S����63u���\�D������|�A!���hl"&n����d�Vb�0dփ�U�djͯQ2(�4�V�K���%C܂�f{��4��.I�g�1�W!���{��H�5}l{� 9p
��f��$L�.�rx��!]�s���?��,4�+ص�I��>C�>eDa7�H8��x�a`�]�s1�x�@���+t��]a}�>
�����/:�Q�md�xǿ`������yu��C<)�@�J#ƻad�����[=6
����~B��=�gI#i���K�7'�=�a���c���H��o��NJ����\�8���P��/���&`y�˯��L/��_���0�@P��<�����4+�S�E�(�����M��k���k�e�eztK+qE��a>�L����Ċ����2!���������A|y���`gh��ͫ��%h�G���fPp祟�/8�-�O^�q# �r���p�o���
F�uS�0�)�^U~W�O㏴:M�^�f��:�����?b]HGx�1�e �F�i�����z�.9T�����!G'߻U�:礮o��R�������r�}Ҡ���P,r8�3N�2��K���I�i'X��VcUGގ�ʒV&-P����ʑ-LZ�b��o-�n�|L�\ m�</�����p�p�Lngn3C~{X}��U���w4*�U�<�BH����3┡a;�$U���x<��n����6�ho�_ [�:(:̻�3]�rx�Y��2�s���F^(g<�֓^6(�Zˑ4Q��B�Tҗ��gpQ�/�lA�kX`�� �cd��|��CF�L_�W�2�r��9�ȗ�d{(��'T�#��(/��9���`*M����8��r	H��d[	,]�SC�f5�ε���B��_�7��E��(���� ���u���3��K��#���[F�ˇ4quh���U�Tͦ�˷2Ȑ	�p�]�ҹ�.���e�/�r���8R����,�_`��?��:f�"vJ���=9<+��k��
e�-�3��I����-L�"�*�f&����\A���K�CW� D�"#fӌ�MR2�\&�H
rU�VƜU��bc�ݷ�V3�!��B��Uh�Q�b
P�[Šz����7�40A0����c�j��A�Ѵ��������4��0��Т�6����RM������z��Q�s�²��2=)���ʖD�x�<4Zj	�M�)"����4?����<Ki�4�g����]&�>x�pr�9W��K96�\�i~�{����h������/qi0yC�:!�,kPw(�eӷ���������p��l5�4ۓGE�v���u����}iz6tN�e�k*���_Qx�~j�X/�]+�MG�N�0�q�Ǐt�g�m�篂��5k�K�c8���A���a�iX�囧q���U��;w������{�ǉߜ�|�Ns�.��m4��,����58���r��;L����]X�/2��z�<��������抬E��;nw�@a�K���/<Μ�������O�W�7��_�#�G+�G��(��h�p�b�o����W�(ױ��W�8���t.� �v��%�Ǯ6W	�B}  @ IDAT�4�f1+��H^��*><��3Zۘ����֭K�+ߡ@�Ѿ���}�m�V0;��G*@�}i�ȇ���m�ӝ�����>��<�υ�5�xi��VMIh'�p�:�;��d	�$h}y��C(HU�|�2c ��¨,X��2,�:y*a�)����.b.�:Z���SX�/-힪aU�ᐴḘ�������~I��f|������s'������b�n����M����(x��e�|������(ܪE�Đ��c���o��6���gm�h!KY�D���L�t��Y��$n}��xW�s�@���ԓ0��/�(V�O�x#�8U$����I+Z!n�=��x|@w(��z�`�ىw�#�s�bt����b�L ����p��H��^�&[L�g�J`+}�L�f6j O3�7���(�W�A��Q
���H�5U��[�����@�R�(\�{�o�e�ꉀ�Y �<G�J��*X�0ə��|�ਹ/3���(,2|+cѐ��|�}�9�+�A�N���"f�
K���Y�d"+���TX�驲�s�+�U>)��'<q\]�{U�@ڜУ��^��<=^��3n��哜�6�f�����JZ�F���W�Y)M+���45������O�&��e��-{u�_�݊7h�-��fæ�z�y/�����vҖW�y�	��?| �+Ƀ�>���~N&6O���<����<w=.z1w����;�a{���?{���"�`{ʕ����0B�SXL~$��P%�!Oz���~���� 3��Dc���x�T��?�@�zVY%�W~��,/�3��O����|��a�����\@�Գ|���kp#�����g>���O���a��;����}~���"]/���*�} �a��g��]��8UO_q�[?�ޞ���&��,l�Oi�������w�A���a�u(��/����=gH͎�[x���>x���w����G��s�>������M'�F�F��N�2q(_�lӐ'bJg0)JH衸�'J��������W��s:��|����{.)�X�P��oL��|ݹy|�{�F���.v~��|��R��j��:gF������(i�e�E���f���״F�,]��d��ƍ��߅5ϟ� _OB�;g૕E�S��v�T��rSZ�͟~5H�@E�7D�s5��R��]A���7��&J�{"���f�
e�UN9��r��V�qh�Q,�h�Kz{Ǵы��a�P��	����]XX�c�"YUvI�:���]8[r����kt3G��L{K٩e�L`�r:J6�a�%<��l=�B)��=�w¦]��R�wȤ�	z�o���o=ڽ��ّ���쑼̻��i2~�?���$}yݲ�ϫ���v���O���^�O;Y)�0�/�� M�P T�r� ��s]@ ��B���u�ô@�`*S
y�7T�*`SA�Y�I*��ďh(k�+i�f4���g\|'3Z�l�J	#��U �~y͕J]և"�xqO���W,q����@�|�ԭQ����E�>*^����_��k��$I�ݐ	$�Dʪʬ�]�3���"/x��	ι9�3�TB����{Wus�Ď�f����Z���WK����&��<mū �[�6�eC!�5��z#}�h��+X�&a+��'T��Vn�����{1�m�W��8	�+�3����A��=O��S���8�4�~�ȧ��<z���Q�I8����an� ����5Lxw��e�n�;(����q�����v�\j�Q����&�+���D�TDq����:T���~����a��������y����aN^>b���]�~���I�r�!4���7����ʔ=�]�+3͗�]��QE�.�(I$��H�L��-C����S�����	d<g�[���n��[���2���o�o��7���?����q�m ���U��6��mz���ģiδ-G�C�Ӏ�"Q�ԀR���[ ���F��}�������yL��	B8ʅ�E;�a�|�in�648�-�;��"�����@�'���5�پG󐎫/�A����s�Jc����re#�\�d�ҹE��h���r���F��G΀��/f��5u��-36œ��o�Z����9��`iys�%�˯�J����(p�C���ֆ��l�%){ �n�^L�{�~�)����6^����ܣ���7_=��cp�>b��=Un�jD{ׯ��+�MoNu��̨I#�#�����y�1QÃ�d5�����g_<�~�s��ㆎ2lvʷg>
���5\#m8�^^�McE&Ȥw)F ��NYN���ҙ/�*�x��G��W\�S�`y5�QB�ֽ�`�q�f\eM/Ì��y����t��&?��P�J]�[Ă��d��}o�Lo�~��h����H y�⅏IM��Oe&�dF����\����tڐ��sx����5�8`|�U�Z�t[���ݕ&�FE�U�9n"h�	Xt Q�&ؔ�X����7���
»�k��F��-��]�`�@:�D6�#|�$�M�B��4F��z�OQ6К�G ��a"8H�H�$L#ݎĕ9$��I�Jv���b��j�]������W͌��ӊ��pk�%[EI^\�F��L��C��tWQ�\�lL�%-�y��xyG�.?�����4�>�)�*tG�.�e(����o2l��ɷN2�No��2���k���mMj<���-��W�D�*�V��u��/xa-�Y�Z��;B�d���L\=�*�w}�0��P�=[�ae��a%���Ҋ{�	�T(ۏX���9^��th�={��`�]0����{����T\GL&Va���§b��ɲ��ѫOiI�&�#���5�g�o�-#e~�d��#�=u����F�,i�'~�����GWd����&���TFӥ��p�oCHN��5�*��x���{
&�¯B�L��7�1ބ��L������t�^��tťʴ�v�i�Sf��s�O�Ό3�ϧ�-�}j��_|�{�y62�]:�%�,g�7�f����r5�<��B�+:�-Ñ��z�����^T���;�9e����A�FL�P�cnv�Yg�X���O�D�*]���4*쁶a�Vu��7#�T8�!9���ix���/��l�Oy�A]����`�y��{��)2�ޡ{�m���rk��s����!�ڐQI*�B�Cm��'�|�T�����?���?<"�zV.v��O��!��yn~h�Z������K��鈅:�S>�X#o�h�/�������U�|Bg�e߯co�#U��bգ�o<��nmT>|���,�aя;�W6��0��5�$�����U��2D^��H>Y�X��Q�[O'�!�?�"#�7�#��a�������y6�0���U���N��o4�2���"Q�12m���'-�k!����ƋX�=��?q�Oo�L����5�� LC��Wb���o|�0�.�ى�ni��n���6��J������L��`�G���8k_�UZչ&ej�I�������0�l�J�� ɗ��pPX�3���+�RA�Y��!��C�۸}�P�7�������B�2s�ӌ0��kl2?n��/<�I���E�5���D �'����/{}�t�LqD5���d㋧"5֤#J�|S ���^ƛJ�ol�[���HX��4���{z���AH��5`ZH�7�I�!�-8�D���C
���J�6�챚F�ĹI���Wo��߲��!HØ���B�SL�l�i1D!�����t
�������^�爐暹�Q�V�~�ਫWw17ƽ����3+�ޓ&�l(�#�q�ҡ[�]!ۊXT��	�ȹ��
sL*7�yZi���ӹ.�3c��R��h~��U|�G�\�U=����u4��2L�\�b<��
n�����}4Lӽu/�;�N���|�r��[��'*�1Q�{Ӛ~����*��������5NC��<����5`�o4�u3��]MOٶFy����ʘ�Uވ�����eJ]`��lhi�/�i�^�	��$���t"
�rO��n�H��C��@o��ڭQެ��s������v򺧉Xd�x
�� p�|W�_�+��4�!tq��w�*��ϩ�f�HBu��B���>e�F�FX�T~b>+5i�<��0e�.���f���cO1��[/6(wY�qN�81�:���Or��K��y�r4��2�����ޥW�r���C��j��mq������)������QkN9�+�"���yNAH&�R�<<��n�1�{�����#K�H	?`�U�� s1�&��ܼ;�w�S�eG�H�Ud.�&�Ե����ǥ,�����KZg�i��3?��\�g���X	�I� ���r��_/{��U6�P a7n�����g�pr�'64� k�G5\��q�|/��UϠȗT�;ˏX�P��k����%F�9�?����%C�5O�	ބ��|I���t�c!c� �^/M�FL�� �?��J�JS�
Y0��)�(a�A&�Ό�6���ި�dZI4��<y�!�I����dB��=ё�c��8�\��Vs�f�5��o��oӎ#m�8?��|��<�M>�o�P�iz��n�(g� �m�%�I���2��<+���O�h���Oy�Y����2�嚕��0�P
�Ɖ�]�&"~��&��KGi��|57���h� W��A�s+���U��W��7mt��:�ѽ(��z��}Z�.i��g4����_],�E��I���`�>k���0D��m!@�p�Iŀ�&?���0v��,��,����+Z�:qٍ_<���H�@�T�Jq�(�%Z�"�d����RT!nI��4�K�]r�a�9�U���7_m	��.b�w�M�����4#��<F6����xL���	Ty�LJӼVÚ���f5l�����3������{XEU�g�>'~�ƙ��U�՘ţqf����/2���a&i��y���*?W��.�%���V�ܸR�����a�<F^�����C�3_�|���!O�Y�����L8��|����O9��p<�����z���Q�艶�`_�t�Ӗ��l���o���;�:�-{��b�|��L�*���&e��.�;��c&�x�!��g������8ϐa6�=w� {�>YWa|`�q���3Gr#�[{l���{�gO�İ;=����􂱝�%������=�؎Ek`�� z�>��>w���)���	_[g:�j�Yg�/����^�l`��n�0VQ���)�\p��	 i|a���N"�6�L�p.��Wؠ�v��xo6�E�Z�G��}2��ow�R��P���Y/uP�@�=} <Z~h���1 4��`,J�����ʹ��D��9t���c�<���z`J��pt1D�5G��_^�a�&��2������Y>r�q��gCD�ȫW�	�U�F�n~�c���I?d�
z��(��Bf��*�1�"M��MV�W3����Ó`�LZ>y�������K�N!~DAH�����-5qK:'?$6�o$�`c���I8�z���Hz�;����O ��+�I8����XNxVhSQ�r���(�m��C���/J�N��]�&�/�
��承��w����س���a|�k���ۻ���\�2�Y/��?��Ƶ8�(�Y�GLw��]�����wK#���;"��k�s�h�m	�bI�d��=6l��JCȉ���z���\�d�/UX�n% U����0��J'^���#7����/Wm�c#H�	��t�
�Ù�8�e��'VJ^��M=<*o������5������������3��g�4�����#���ౄ2���]��PV�*�A�
j�k��ʷ�����l ��m��j��6���3e��f���H�G��㸄��3��[�̃	[�f��/q�q�S�g��e��{�W.�1���u�~����Ca���ʏ�B>����O�1uk���oRƲ�"�s��]�7�i�7������t'�~�\p���-_��t1#ď홦�e�V&�3��3A�a�������,�9�>:�>f���`�W�W��7)c���K/��?�ǋ^3V	�Q�F���[.�Q�3s�^s�Vd߯S?z�b�c�E�vu�glB{x��8��D�h��+��ιr���p�.�P2<{����in���t~%��!���$�e |+|M���W��嵍;{�l�ً�|�S�L�?n��x�yk)0t���B�!*�W����oR!�������O��^��l�iy�k]ᖙ���^@� �2«h�/b(<��N�!ˑi1�"�bhj�ޖ�>b�|0��dLQZ�߰^��(=�w��қk�_+��Y��mK��W��)7n�r�H�`Ty �a%b�M+ƄCw�=�Ғ#d(�&��m*t{vle[�8�7G�%�&3�����_) ��d��/G��Y�	~���� u@���B�g�q��"Ӓ9|6Ôx�!ޒ��P蠿/x���gķJEC�`�6M��d�7e�����D�gұ�"�^^�4�A��q*v�g�8dYx���{�|Up<r���#��/y���B+ύ*�U�9U`���5Y:����/�۽�p���ځ�ud�~��x:`��&��{w�aG{�֝�A�C:�ջ1|���=��I����x�0�@e����˕yu(K��fŗ�EY%�wa���C�ޮ,r�y��&���}A+������,|p��8>����]>.��'�n�> ,�:+��v}M�f�Gy���aJ�
L%�;y>��<A0��/q�V>oe��U��_��#?j�oB���m#��u�eh�O�a1q�߆���	'�*��*��^��	�p��Lg�������8�r黽��q}_��zͰ>'/������m��W��3l� �M7i�.��˲���e���[������}��(�����jjY	�~�J~#��b��m��G�]sue�{�ql��)�-gE��e�v8�hB�q������i�X���C��t$���!=a�0��hp�o�K�Ḥsv}ϫlBzJy�`>Z<i!'�Y�v�k��s٨�v1wH�M�>�|��7��5t��+�(�w�0ꆰ�N)�6��@\�=�>go��i���Wʵ�]�:�x�&H{DN�{��S�'g���N0��OѺ2uo��G��a�VW�{uj>�!��$���l6���]ʍw����u<�� �&�7|�C�pʀ�ȇ��O��6���������W0�8�wװIӹ�-7�'�κ��H����tM�2_|�2��g�%��'�!"0ŋ��-��^�v�F�y��v ���8M��W�)�i��(RA���2�fe����.׵�f>�B��nq�=�@ZF�����鍸�z���13� 2��ZU8+��o��$���_��+L�U ^�'j�D��6�X~���#fF��NB(��! U�d~A�Ci�8a��|*{� <%��a� o��BRX�#����3oS�hϼ4��,��X����a�K�� ���1�+�]�o>)Z��@�q\>t)��&a'���=��D]Y���e�̤{*	W�nm1�w�_?z��=����Y�}b��N��0�p��`�K���9q^^[�Sq��0ɮ���ixu��{6�W�>����-�b��`l�?xp���}ʑ�|灹��ϔ'�R-ؼ7�ˣ>�O��o�e��u1���2�4�OD�Z���gU"
$Ň��X?q0��L#,#�OC��qX��ܭ8���t��L��A�Fz>�G��.�wӜ������U��=�Ű�n˧0�i-��f���Ø~�>'�ާ�j��������2l�e9[�c�?E?�Y����OyC�w����m'v�3�G���'VC��a(ϡ�44�Z�ָ�eAٳ'V��5I�Bdk��`�8����_�#��b#Vה[�Y�b��e�iv�Q�����\O�C-�v |�0�H����ao<7�vYW�ih�cX�9_ǧmO�=�a��k��#�%z2{cѐ���E8��n�53�\$7��0>n��D�Opq��!�&�{�@����^6˪z�$_H)|ǑK���5�bl1���v��B���oN?�@��eY���|��-+�eީ;�7/�'-��zs��N)S9�}��֯����fX�Ы�u�+p����I׈��ȼW=�_�N�q�Z�j�)փ��-3���I�0��R��x���-x�$L�?��L�[��t��*K��<8Ʒo���-���x��HU�R��#�2Py���Gf�E�1�a|�V�\U�I���^��D���|�-!/N�I���D]���ʿ�/��&���t
u�+�x�ݦ���8�M����s<��+%����G����KX~oiq\~��l*G��/"Y8ZY,i�{�_�\��
^�V��ij�����BG�	ch�Px3�@�vv�ǭ�]1� K��O8)�n�*J�hja��͖	�
qc � %�?�1V��
_W��r����,=�@�r����x{dS1P!�����}&�j�y@�-�S�3W������;f�/cX�|��+<[������qD������a�e�_��kZ����;�EY�0��a����g������Y�(p����|���o�`VE�;?���+
�\�*�t�[%��1����e���Ȼ�����׌/�P=�W߇ӌA܆U��{q���]���^�4&.��n}W~U��G���>iҚ_���Wq����z#S�x��3^i�-L�����~�k��v>�$��ބa�yMx�i\�yMw��GƟ�|V.��nؙ_�*i���p�Y��K������ӧ��O>_<|��愞���/�^G��k�1]�"�yU���F�5��]7���A�b�N�'}��7�8��`����Y���z���E�<^ݥܱ���1�;�yj��۾��Xl�L���fH��/�s�1jaqʾ�鱶�G�d����P]����yRg�'�	���
#~�Kh]�A7¦�Z� 3�`��[�o��aZ=�捽�nMa���)���gC:EA��C�V��o�VC���|C��1��^�7�o��/,N��#������"0'SL3�=��@�%�4P�n� �l�i(Ӌ�oH	��;y�LJ\��q�JGF��UCiD�K��f�L^�{�L�:ι�k�d�G}���<C����<X~�'ߒ�0��Uf�c�7��3T�n����{H������vp7&��|�4+#q��pH?A�ho|B�AЬ��)t�9��
���"���5�|r��ϼ�`w˖�g^���0܅P@CD��X�C��P���K���7s���߿�H���@G2�"�U�L���r.V�)@U��'��P0��O#~�p7%�5tz'��ý���&�0��ě�,Z����3��<�s�&>�K�)��=�2�K/�Sc[��g̰�Sf���=�?��W�+NĐ����݇`�J+J[���r/"w��0�]�v��^�(V*V��!��������r��C�۱��J��-"+�Yʁ����U����s����2�����y���?�å�������W��t>G{*+�_Z�����_EV)�V��H�sލ��&@,�w�h\S)�o��#�5meo��Db�he}��?�V�����[�ȤiLx���֤^�}>������m�H��]3����x3��jٓd����.ˌS��3���l j��m��.�m|,�F�N)�e^6}}��0��B�'�=e[C̡{w�w��/�}�\�����k�@C��0U��Y�W�n-�2��A��e"�&����75x��3ı��-{��ۡL?����/O?g�-L����g!�K�9=Bn�`/�G�wi�=�`|��[8�*�M==��:�r��AT�9�By64����)nv��B�oǄ��P/D�_f��a�� ;=a����dx3�4�Ҙ�kT��i�p'A W��9�]���@��#a�SÛ�/������9~J����.됔i�u���a|�����,C���.����[7��<_��B�x.�����_ox�x��p�4ѹIK�oM�B^����w��@�H3�'�I�r%��M6iJ��}d#�w����3�����g�<n�
#�zP�ge��~��(A:˝y�|�&�k�I�f*v�m��1����� Vf�V��h�����aV9T$0�Kx�����V�*��ӄ�;�G,^{���f�D<�xkZ�BOt��4��N��	p'��O42��eN0��b�LI��-�%��#�g ����"*��%G�tK�'�����RQ&|�%?�73���";5���>{���J6-�j��g��S����x�/]�B��c�ҙ�C��0C��� »�Օ��?20i��R���W1й�qx�䙭cy:�S�D�قf5"C{�����W+9鱅��m��3��
+DitX@c�#G���!g��ƚ�^}�>X8�3r�aI��X�_�V?xC6��U7
�t[��{x�!�{�y)�Q�����˙�O9$��+)�u�/м&��,�O�z�+�|�o�p�����;�}�S��F������/�vU���8�W��ϧ��9��m'�¬�ֿyl�?a*�f��Y>���[��s^���tk�eXy�e*5�[9jX��P���0ꟴ���8��%8�^�K}�tf�����T��o�:IjX�@]g�5�a�[�����2fϊ�H�C좖�M��o����CCYޅ=$�X����x9uDz��ObI��T{d��樘=e�
�<#���Q^���ş��>���ހvn#��[d�а��~�L�j�#C�/^�Z�퇟���ū��ؐ�
����+u�@P��nP�:�U���;I��o�Z|��3�<���T©[�4���t�2��p���;oӃ�D�K/x������f���Ј����w��[[<ek�����K/!a܊"G��4���C����ݡ���?���kI]�>m9ZI��mO��L�@5�-����G��/B���F�N�W=c�^����r�*p�[ҕ�|V���Z2�7dq�j�@��R�9E��=bֺȹb �\�x��U����>�w:�j^�;�5�-g���e� C���=ˠi�|ק�Ip櫅vk\�ߗr÷E ��!��h��6*"g�������J{6N�)i'�ĻX%��
q����;�|��	� �9���IC�p��iŐ�m���Z��̦%�^�#�	�����:�q�$H:Aٟ�ϑ��M<�S��K�(�Qb(ڵZ�9	�a�o���M�!�f*x�;Y�HCzEi���A^T���ISP��'|"M�:����������~�����Ƥ/o�|ȟ �a�8�.�j��G>EnL�7���^��!���r���^0#�yVT�D�(��S9���U���јtn؅�����_<}��ϞB��`E����K�t��.����s��$�]��<V�{���"�`R�C�7���ሯΎ�h�T�"��
��+�}���u<&o�_�p�0���0Fس�F'����p�E��	�#F8�>��e%���2�3�9���,N�FY�"3�	c��sOH,�\+[������jz�i����'}���O�u��~�G�IwIUc^�ch������ϙ��f�<�7�;���}3�?�+#si�d���N/��֟!�D��^H�w��lx�aB�[A?��p�x �H~5o�.���Dh U��cSk��=6F~��A�!) ��bˑFD�/{D�Xn���n��z�x�\�~�q�����Wv�g���J�����琹�ҡ@W9�������8�5^.Y��}��p�u�(�: ��^3Ϧt����g$��S_B��9��'M�~�����OO�6��Ɠ���O�1�5�ڢ�x���u::p�ƩN�g�xg��_�Ҫ��W�|x@������o�b�e�D���Iػ�ig����'�x���J�Ӽ5��4,##���/�d\���k�:1�d1�`�h� �2�F�+�5��X�4��{3c�'&�D�o������ܿ6���9P�H>�~ZU����ҏ^��`f��~k$@�aU����ɼ�-��o�NsFt�<e�-a�	տ��MhNB�6H���'��ZƓ�֭�1L����m��]\�@�3�����[��+��ΰ^s<[��`�
�-�v�ꯠ��6��/0���-oH=�|�!lV8U6�1�39��W���3U>��yR��7���]�Q^���y��3�p��>'n�_��e,�-�%!-/����~�h���+�&�ȷ� "V�*D[�(
��dHOC�}�SE_ȀVY���u�!�*&���������s6R<�'���Y��c������(U���6���ӳuD�����L;���,mढtC^^�i�I�(����&��p5�p����].���SN��T��?e�|�a-��I
�
@6�-������a�(τ7�6�	7��K�"��ʲ^~�{��s�'����O83=���
P���
lq�������L��-�p��-�q�m�'��K�Y���<�w�İ�sWa��W��2͙������P}0+45��)��8�~�+`�Ox����)������I~
��p*?*GW!����u�	F���k	.M叩r�r�Cnu��bEf���0pO��h�q^ ⾀.\�t�~&�?�[���
ٺ��_~��'α����`|�Q<=��J� �K/����=�{����;(��|���}����p����Y��[�zA7ez�o ��uʐ�#�O}b�\�!{�1v��8�C_ x��|t��"[n�B��jS�$[�(,�'{�7��-6�� :���>`�D{��'L�V��>�������9'$��v��O�+�� @�H:s�|	m�Zj�/�[4��/^�E/Go���}$$̷���$���i#<r-��y6 YZ���ʡ�e8]xƱ���P7#�D6d�������Q�V����u��,>�=�i@ !��[PbDHa�H��X��	�Ba"���/\B(K�w�HP��_�0���k�J fF"7[�&����z'-� QE	L���Yѹ��8"�[���^�QEk3=�b�.ϡ�,�Fj��� [��_\�ސ�{Ӯ��*��R)w�E�\��?�W�)�H�$P��7ᥑ��?�߷p�߸���$;|���i�U�#,7�򠊶�l>�ӓE�چʲ]�
�s'�_�-���wQ�SN�5nrdT*ft7{˴��ޯV@���w=�ު6&�rT���Gq��me������ �a�����^Tn漓��1�ز���J����bex�%��'�Fn�#�9����.�k`/�52�{���(�Y%��ͻ�ǲ*�^y
ۏ<�v*��)��͇6�H��q���7���	0}�����`��t��V��|�2᳴	g �s���׌�{+I�ʋކ��*��e��[�L�&Pnb�y[����'�)+n�7��0$p�r�zM�"�o�G.<�{5f߅oJC-oA�����l� X���M^��h�AYx���˘e0�J��}>u������o8#�v�MP�Dߘ7uy�X��g#�Jy���Ǻ����Y�| ǷPv1��{���ȯwl�����U�3��kzo�����;��H%鶧%:���:����
^ஞ_G�WX��~g��V��ۆZ7��K�䕟˸~�o	6�'q���!�~	L�*6,m�	��N�HFW�&a�|4������w{�1/��[x�
�}��r��Q�Us>���>��0����R�J��$�����������Mb1^�\�  ���n6��ɴa��Y�U�ԗ\�,|$�g� Vo��ԧ���S\tM��"�'~�q�e�!֧u�6ʫ�%��T�~(T�����Z�pR��/Q�v7�?��*�� �@sb0�o�L�bY���Gt1�O����2p�a&�y�"��c(��1�@�6S��4��
��9��4H��̄%܁�C��y
����`8�3=�I~e�5�U�u�O2I���IcK�$(�Ʃ��� Ş��,�U���a��m��o��,^������w�����&�@\~����w�/�N����r!24pkp���&�!7��G9���
d��s��aR`#5Z� �<��Ъ|Uvʂ-w��;�ӭ~��\���s��q�7j�gN�;c���v�?Z�gO�W�^Di{���>���^+qr[���`s�Il����J�9��^@�A�g���b�dA4?4�>i�b�>�D6�_��r>k$�q�H��<�-p��+�T����!2<�T0B.3��FK4�j%D8�"Ӭ,B�I�n��0w�V<�2/�,J\���7�yϟx�8�a���tMB�Sf��eJ���i����~L����:!�a�jZ���(�	lu��r	[~�`��^ ˼8I�jB����.�%�b��W���}�����^8�����x�_��r�ߍ��+��5ЅP]1!��J�h7�2"�"'D��vt�c�@0P\Ģl�0̡�ʐsne�������h,Ey�I(�򑷔ax�i�G�Qp�A�&��u�2L������"݂��z�����N[�%?�k�Q����X �.I)�9x�w�� ���px��>W9#0�#gvy+��\�gv5Ky��|���=�!g�φ��~	wp����9L�ﻫ��<Ò4/���0�ԇ�O~�\���ss��s�yT(��=���d�N��-��A�e��s�������\<s��w0�v�Sf͏�=V�2O���y�����[zGϲ��36c<��[�i +��&=��zx�aF*.��:�/G\�kd4�0yA��#��K��tR%I�� ��^�I��|J~��?�2���WF�	☆��;/a�Q�(�~�>�!>�I>��Z���1uT��i� 4sQ�kH�B�V�dc>aqY�6~E������!B�K�����
QF�!KhC���᫃q�i��7 5����/]up����Z�>�.�1��h�:�4���X�#4��h�.r��7���QX�W�j$�"�B�p��U)ʤi���}��+W݉U��i����,��V�=yc���P`��:Ro~]}��LCG+�i�2J�\��V���_�gX|���0�"W�*��Q�˜��8	��=_w]�u�0�~RQS��O��v��礱M@9�����ᇟ�E�bn�B����z������8�y *x�H%$>΁Ȑ�3$�CX��G��Pr���̠Ɋ9[������s`����[���/o��]��aw����Y���|F�>MY(�&��{��\��)���JJ�L�&��}O��^ʂ��N�J�&����iv������c<�1<�6��3�lM�s�A�MKG���M��C�%�CO`�[�R`Sn�.�I缍�%i���M���k���w���6D۸��o�&��D�[�RJ�i=⩿����zH�CW��v�;�1�ps��i���,?o�{zzp��D�	�P�!���!�2H�)����u�'\����SN����e�+�Ȅ�|u2p����lV�
r;�Qzd��h����A�ċ\8� �:Ԫ�F��?�0�.S��|�%�ܭ02L�Q!���>m�'M\���"{�	WQnwc#1p�%�N��tLp'���QF�M}�崇��dZMI}R�3��!��(Z1F��}��kO�� �sψC�CJ=%��)i1rp��Go�+$��>�m����쿨�#��S�M���8�wÚ����n
��zӴ���<�_��昞�4.���O%�|J��;�U@�fj~�q��03HB�b��An�^fNH3��Ij��Sf�mʆq����m|�1�2�߼��2Q�>e�i�Q����x�X~�l?)���kQ14[w��_X
�1�J�X�*���!MZ�.�\����)􎬔���  @ IDAT���5��f:"=�+�*�(
(���@�-M���ݞC74�!��s,,-�� G��:Pʢ���Be&�EE���|rrْB# �OP�_����-4�<|��h:�ۊ���R��Y�W����V��:FL����4�+�����B�(*��yl3���I ��m��T����;��U�m+�M.tW�o������{��x�9�.CW�����e>��6�����������n�z��}?z�x��3V!}�v�����f��ت��[���D����>w�V�k�k�s��Nnx�^:�B���4�5�B���m�V����UX䃽5��u�$d�{��r�y��6��fRn���ee������"C�	�
Q�(l��Ω����)�3a5��Ï��柲��y�gp1��Y�_�7\dLo��!etaEQ�!aaj,릜Z��|�����%_����,�Tq���k>�lp��k�D�K�|�#��j>xԎ���ebj�u��8Ϳ�I�,Q��r��qUe��'1~�=D��{��o�oY��r#A]b��aK�%�M?ޝs���̋��.�lK��=cҚ����_��c�.n��"Q��Xʞe�3�s���ׯhT���r˴�{6� lq������)�}�c�/vz�y�{�cU?�{P ]��M/{�\n����ǜ��>~����kd��6/{D����'̉:ff����X��.�4y^��o��r!��]�l�������,�\g���/Zֲ8	Xl����s&�1ƫƤB%��e�������+O!`����=^|����Ê�e^DM��$����<ᝲ�9����w��qy���i G>~"l��*8������W�&�}f�����e�2iĕk���ƐzI�]÷t(�#ܓ���0���W��qu�v�>�]}�O����E�7�bg��<E�XG(����?�S� ƹ�����!-
"��w�s�ng9��廑y� ��f��i$'?e^�y��e��Hl�7���K$&#⯒�f�Ad�f�$���&ў{���7��f��ç�����e��n��U�#�����M�Uy�K�.�O�J���$���EC&n
�>�:I��*U �7�)������W����ҿ���L��m���/�c�=�����~8).���ŋ�K�콲��K�Y�`O��f�]�vyk$�K(�� ��8Uy^��4���B䆐��,���zq�!�_oPB/9#�=G�:@חEҊ��ty���&�LF�o/>�����/��|�a�OX
��wjC���N0pN�$�\r���OR
t*(=�˼3�%g����#�iG J�Y6���U�P�z����R�4$U��Z�G��0�������Jag�*�S�&�k�c� Y���̸���O>��)�C�����^6�L���1�.�)��)� V`�F��vA�3�Ө*-���LOb~
c��9h�M���ß��'8[�(��_�r7=��YƩ�%� I�IK���\Z��d���?�Mü�r����d��S��c��Af�4��\��w�E=�)�P����(K�{�n�x>(�ʔ��(��-�%".��_�
�ߏ�K��7���e��4./��<b�ի�Lg���Y�,8q�/�c�:�{�����w��W�_�J\'����I���I�t�i최��WL�1���[t��%s>���k5�t)��-F�eꌞ���6�?C��� �W�Y���������{�~����,+s˳ñ�U�����濂��`���V��p��$�'�V~<��sr?g��'��r4@9@��p ���J�� `;�=�N������rR^��2���Op�5�f��I�J�>��7�<Pm�&�AKd;@_���b$֢ x��9o��pǨB��o�i/�y7d�&�p���>q⧂�.̢��oު#M#�0����2 ������4L�9+7��Ej�y+"d�$�.-R�r�$$0n�@(�y�%���]���d/��H��-�N�'��0y@D��?ҍ 8�e��
�Г��7�Q�ͷ�x�a`�&Vv��#���a�ўZ(N�vb�
3�\d���q�M�̤o2g[��Z�|	w�IM+R���/ O�Of#��X	+�b�o�WZB+����
g�\�VnP��H�FZL��_�0]���k#/�T"�� �L$�b��%Dsɑ<��B�I���a葕�[����e)`VR�]ޤ{Ƽ�3��p��R�[����?t�?������H/ث7�ٹ���ǟ~^�A����xV�ں�^��۾�㷋�������7������ �x��ܺw(��i"����rX"s�4Q����?at;	��ɪ;*&�uH���%��
۳
)G��%��)��|kl���i�828��O��e������] �O�`Ȁ=o�8�("ȎF����{�){�h�d� �:����:)�\e]�T��L��a��
�|����G�� ��J|���(��P~/0���r���xI%p����񦩜N��8!i�^`X��Wi�gB�.4��+='�}E�Z���a|/��w�N�-�L�~pP�	A�;���8��x��/pt�a��ei���&����S�-��	��c���2F92�8�2์ɕ�<�5���Y��ғl���V��yx,.�%NJ����H�Oy=�k\�e��\O`�C|�g��W�9��U�/R����)���:��C���O�z���G�i�`ϯw 9������i�8���:5�A�[(mιJ9s�Y�����_c ��٠��>yq�'=F�7������J�C�/1�~�]��v�tfGGl�Sg6D����H�e��a��T�Ѐ{��9�lm�f��,���L3աO�W�H|�\�cξ��߼��5u�zU��|
C��������O0�����0�7������C��eG7�wp'?1��H�yY!B^���nz�kC��W��.�� R^��9�X�?��p�?qR�Ut,D��>'�}R%$A����� �P!�Z5�[�����&�!r�iY3.��TV���H��Ȳ�Eއ"��D�b�ٻ�NUՊ-=`"
�Kn�)2��o�i��� �1Zo�� 1����i�*b$�K�33G���D㦕]:�!F�! �7�)��^�R��'�aR؟�$O<�̷j�"�\�� �:�+���d4�� �HvP��/
=#��\Qɫ �?�#�Oʹ-�s
Q'��@�����-�)`U
J!w��!8(���I�U0�C��2����TJm���^�G�-) ����RHǲ���*���|�^q0B칲�_�9�C����]x�ٍ�p۹ (��s����!�G�ޱ3�;����"���=V����B���{	����G,ci5k���'2A��������}�����/�`;
�]���R�X��+����j/^����dY�}geJ��,:�C����la���J~�+������[��W��?�!//=��c7��P�2�������UPDy
����Bg�6yȻ{$Ik�^2F9q��"b�PBM�0I|#qQ(�/����*�2l�M�6:`��p�R%��i����K�҂�5���|��/	�K!�_Nbp���������y��·��0��
�@�!	\�*��_�= L��Ѱ7i�S�K80�X����\��/yR�xb��nx��ޖ�R'���_z(��ʑC~�iZ����o/��/�����Nᇻ+��<K�H����H�-�G4��0��Z+:͊9� �`�������ۛ�0�4>�'K���|Բ7-��=��~��w���?0���	���i4�q��s4�4��4�^���#����oρ�(����ik��
?�8��n�A���9e���7��P�G��YZ�5�@�$n�Ue�]��!X��J�i����×��t&��U����ГՎ�������Y�e�
?���������M^9i=fO�tzE�̇C��:�pBV=�S,3��"� �y�Ӻ� ZA�w�2OB��L^[~�ox��X��`0>##��,>>�P`ʿ8;B��8����J4~S���u�v��
�ɵ!}��EL�/�RBȦW�$�!�[�k����]�GH�#���l~���H���ƫn�M+@Bl�Q�ЃlHTh <TrUt~������	�TAZ�-p�@e�����$��f(1�T�|�3`�0^�K���*n��U��zt���xw}qtw�ؿ�~Pf<�q��f����w�Bz�����D�`�§��$���K��D(��U��q	�UƟĒ�\�������N[�!�8p���ĳ��"d�L���$�?=|�s���Y�G� �0�z���/��s���N)q��N��;�j�O�'����h�EKw��g�[[������8Ű�e�{�}���[#1�ɐ��Q�{3>��w�f�ʣ
�y'(�W(�������?<_�~s��q&�
�F8����@��rn��x2o�p��l���`t�^`�d���N��<�Wy!mV��=Y�J���9��Q�fAz��0U���NV����ar.B3��-��{_� U`�'�ଌ[��|�pk���=�b\��B���\3�W���Ҳq⩜{ٰPV텷h�~2'��a���`�U����;/�*z�<�;4������mzN<_��H%�L<���,o��m:T�^��R�.y(\���K���y�N�f�4��NϚ ��ƍ�ʋ0��r~{��OS�=M~'�@Y˒΁�G������԰7��Y�]�����[�wp�Mvτe�t:�Ն��֐���&�K�8!F��o�0�T�O�!�%�(�i�:u���R'�7�:�������3܍-|������^慆�<���q?�3�;�B5z4���^!yG`eG>9x���^�utgh�����OH�e� �g1A�4�0�K����؃�^<9
�f�����Ve+��g�>}ʭ�)+w����F �W�c�0�\��,��B����	���_Ƞ щ<c�����{oя�G�k蠔&�x)s���'����\#�4o�'���i�VGZ�WfH�zԼKk]����y�<(K�fb�CK����t~6hR�BWt3��"��̈+��zɇ�0�dʛ��`��rzG ���oC[[g��:���	m)��ɪ %�;���c�#��T��r}΁Ǘ�t�q<���_�3oE�V8_�}Vq�&"6�"3
�*�*3J�`�J%�f�L^`ja�G癡�]ex������7��wS�x� ��w=�Gߢ(P
�1��?���	V����ps��KälX��K����),��+����4>��������?k��˿�����iȄ��pȷ)x�L�J��jV<3|�N�œ
N"��m�f��Ŀ�E�o��V�Gv������WH5&0T�7k�[��b�����z�M�^�g�U&�bx��[x�v�>^T�?���ޥ�eq}A������V���:�ʦ�F�����\P]��_z�Q�n2�g���_�ắ�`��굻�SIx�YW�Hs����;��0����S��%�\s��
�<QfѶ`߉��/U�V�r�
ݗ�������\�����]w��.o���0�r��f�CȒ,�&-�?3XE��3 ���S/����c�@�͐2"�JNz���WeH�ۥb�R��RAA��1Iؼ�����|+��ȯC;�n@����^��u���8��c�S�S�IY�Q�g7ohQ�5\\\��2=a�]�Gjϭt�o��$DҲǎ��N��@�F����Wd�z�#_�SJ/ ���V�ʸ�T����h2�Og�ieM�_��S���iw��mvg���ϻ~�M�=��O�N�3��Q��._����У��-�^[�Ũ����\O��'�w��hd��9�vͰ�+�c�Ǣ��W���@��{/���G����{�^�N}o����wc{��_Xͥ�c#���ꜜ����W�Sq#5�%���e�������O��:z;�o�ApL`��ĩ�d�$��<UN�_-����r��70�jԸ��8R.>}�ۑM�#�m ��Y��%�p�"�?l|u����!�c��"�Q�����{���o/`���'�|ʬ	q3���\r�8��\�����@�N�(\[?�t�F U ;�6�`C���C�S�c/Q1��ˆ�SWLZ9A��p����,�!�#e[FR6A_�N0�,�̀�w��a��w@��5�2��P�?x�=��Q��eޞQ/4&𬓴�+�WٳH�fX=Zt�eU]�D�3����ad����>� 6���aK�L����6���=(6�O�<(h��h�F-�|�BR�(�*$w��P2}$���i
����Af]�����Sa�̂��-��kUR�L�ʂ��mFY�p\#�-[��wG�OǴ�ޯ->��^=��f����&�v��,�E~ �
\��$(��q��/s+<�b@�WnV�C���*RçJ���g�c�# ��Pq�/Y o6�4���N*D4��`�8F��X
���k�Q�'(@���������
��m%����u&�2����n"�N��闗��/>,^�>�|7zڥ������{�ܫ&�c6d�f�аk����J:��C�R�J0��1x�Ѱ8Uy�|	����?����ū�/�XYt���u����|�T�T��U�jc��5
����}�u�A����t�d�G�R�ާB�g��� {R5t�	�`a���0�S���՝����5�v؟��G���	6�]{�\�/;�^�̥P�������u��TdHG`����/9�-C �o�����{�9�q�,^6 �'�/@)�{,fp.�}&��e�i�^B��s�����_�8�U�N��AIy_Èy�C�=�8�����,^rx�K��z��~W䋆��~��8�d\�V#������]�@���A@�oQ�ҳ!-Vj�b>v,�k��؈����Z��OJ�Gza��Wġ�O�?->�g���Q�4^4F�y�G�K�eS��,S��^S9h�R�� ����ߡ6d��<���,y{Ȟ�ω�a��5s���0����L���C���(����g��GW�p�q���>w08�qؽxJ�����#����h����JP�x	�;<�k�!��
_��gT�ȡƅ�n��O���҅Li�-���u�i��0�����m�yjo�gA���u�~�X�Vנ��0 ��Y }�i���蔈�����ػwi(��M߫=-掠��~�k/�e��&m�I[$�R.=�_��2��g}ku�_0lO��	�m�r�A9'�|��%�i}Bo(�f!ð��X78��.��5�H�Fŉ�5������9�\�hŐ�Q�k���"�knu�dD��+�]���z�
8�~�߸x�x��P��S���Adz��7��K��u>�����E~� �B�>����6�9�-2�j�w׋������(�W�R������_3gL��O��ȏ�(����X���E�ߔ7���М�	x��-�+5.4�п������F4������P8���	��|��QI���P���(��i�Y�!J��q��Z-�2��7m���Sf�fA�`VJN��g�/L>D�m�^-�&��Vԉ�+�	��4|���k��M`� Mjf
�o&i� �Cqc��2�^��/魹:��^P�	���Q�m�(����b8_@>��O ƍ�V�o+3щ��(�*'�g~� T��X� �,��/��i��4��f�2D��ɯ�޼5�a�k_
����4��z�*{4.�S���4n�MZ*�j���(�+z^��~s�x������p���Ұh�j��2���.���S��]��Y��I����GV$�n�g����1N�N�!���1=j�g��L��P����M���x^j�Dޣ��5e�<�[g�o���u[9��T�_~�%y��%�����&���y+;+h�S䣻x[\����[�����2�B�&�ȿ�x�!��g����! 0�y0�<����74�/ʖ��(��r���'w��p�}��z<X����1$�Cb��,7+G��42:�������ٳ/3��^�m*[�/0�^�~Go&�`��� 7R�.��X����9|Y����5�0y&�Ι�'G��
����!-�_g.�2��Ӟ9pð�(�fsd���T�q�J��J2s��c�:��<ý���������-4�%�/�D�a�21�(���!�w�J\>xL�'��+�kcl�4HN���@K&�LyB����Q�[d�=�g�r��b���ǭ�[):���:�{�|����=H��F�9�W��ߤh�� ҵ��_�z��	xR1P���1�+G���2$��[�$�L�_��QrVP�D@��W�\[�R��H��YCD�}�^|O������#ʚ��4���a}�6:�^ � -����L|�,������H��A�5��)O���=���{�g)�^����=`���MW;(�AJO�yԟ A���4p50�W�
N�A�|1}{�cT�N�0��/�5ڙg~i�S�\��ch�����9x�E�"� w�����.�{��ۡ��:�F_GW*���zO�;� �K��^v���@�r�)h�^o��}J.:��Y� �z�) �m� �Y s��#ȍ��'���]]/�l������O��؍,k8�����ͫ��k?�:����M-�Q[B�]�9����dT�#��%�D����m�ln0|LCt˭��3p�9��䛦44��{qF�¶��6�sh@"�2K������9�a%�c�VRX�ɰ�
� 	�^��I�>�~H���E���@2
 �hM&�<�NѦ`�%;|b6��CH����K5!���\���Ui��2ؑ�Z(�^���U��7pjK��9���-�0Pd��{0V����;n�%߮d�-2V��!T*��GH�`��;Wg��.�Ǖ7��7҃��b��K�es>��j@Yz)��&�*/�nR9�q*Q�unF^�0�Y�@ �`���X��y���P��"&���kz��R�Yu�
��LK�����c�����PIi�&�1dy��[6{T^c�e�,�}�P�Ǐ�1��῵x���w1|�X�r8�pg���)�\`��@�l�
h����9%�uM�fK���d�:GѹՈ�B�� �,l���̐�	�88�h�{l����8{�m.�h�k|��K��/��S���mZ��{�~�����/1B�>�P4�G3�>~�$��)G�h�Z�kx�Pag���H���+��C���6;dR�}�cW��y����j{b.����p��Z��4�X-�9�>d?�ﲝ�b�ܙg�o���]��S��`�ĥ=��
��g+���{,���᲏�s��|���c���(<�o��fQ�$
᪈A�)�VV�]���Az����Ċ�[cW���F95�ݱ�i4y(�=A���{�]�����(���Y)E���0�>�v������3<��F�����2d�|3��Tmf<��+x�������6+o_�/�s��7��R	�<|����S����-=�ۈ�q�p�Oa�Lp����G6w�~{�]�w��c��Y��!�ֶb���{"[�H�;���i�N�b��.`Z�B�z�	໛ ��?��⛯�LΆ��٤�A
�7��ϲ.ߎ~N�Ɇ���6N�c6~� <մ�|.�1�\��%����oH������l>v8Z�{��1
K9����%�<�3�d��_�Y���1AYB�8�f��{������L�)o��olm����2m9U�jʓ����ke����^n{�6il"+���9�h]&��/�7�+��W�X�Q��}��cu�˗���}�$�������*,h��8
S<U�v���<�e."�	iR>g�F����� �D/v��<{Do�7��=�E�p��m,~����x�(�� �EQ�W�=Z����h����UO�h�)�řwҠ�*����bu��U�!�pȘ���l#�gw�"�؞�uz��6��f�n<����- �Y4pHS�1n.�
��j&/*1��mE&Z����NKVcI��5��J(�{Z��w$ӧa����q�K��!��d��\�x�y2&8�#,�$.�Iq��$~!nN�#�kJ�0��ܭ>PAX��0�J�J�ʧ��X	ZA�W�ML�7���P���ӈ���u�o�DΥ-��0䛷�q�MH;��T�����il��!@Z���Sn������<�CLxw�x��0�(�m�^�\A܆W�k�2�(�-�IGG�(R�BV��3+�k
�7QD���s�c������կ�.ޱ�㇏0*82���Z�w(���*��Xe��p'�����'����x�p�Z�.�>����aAWa�[PJ^c��#�����AZ�#��-s��}<cx�nq{�Θ|�(
ޝ�?1td��
;ʙt�y�\+{�4�����1:��n�a��t��h|�q6��5�=���m9*�{wl��r�#L��R�<e�*G{�=^I�ǡ���}�����G5Z�U$��S����Q�#[����s2�<�|��ӧУaѼ?e��޵�}z�0����QN��J���^��h�a�ػ��z��Q���2�|���5O�
�p��a@{�Y�u�Oq��lR��N{cQ�5x���F��O����bR�e��r�Qd��z/���`ʖ)!�n�&����WϨ�0��]P�?f��m���--�-�#�	�R"E�~y*�3*c��{{̜U�����;y���o؃*��0���'�s:�!�|86���� �?F'I���kl���٨����向
6��P�yoX�UJ��Z�M��<��e�$���|�+��:ņgz����B�8]�\�a�>�p�OO�]=��Xtȟ�"��o��vc�^���_�{���zX��1D�Z*wd�r��B��F��hok^d��_ӱFu�4��K:O)�������q��\+{f�	o�p��6�$�S��@Ƹ��>=����"�':/=�`����F>(�u@^;%!��
��X��o��ߒ��0:>vC�l�O�=;�pN8�"y���Ij�d-Z}�\�~��޿n	b#E�:�d�{KOt��4��F�8"�G���/�]3\j��B�&l�N'����#�o�3������Q6?��C�٢����������k�y��i���"4���[S<�QyQ��Fc��p��q����_^��l$6q�?�ޱ	�����e����5.p*h��������䯮�46�����L��AX!��w�ۭyE�|���J-pG��%�5v��7�X�$�G��)`rm��B|,�oP����q$�$A���g`����|��c8����%^���Z6ܵ&Sq2=����1��iU���7���(�iX���cp���g��B^�P�!�!ʹ,�`L��f��$ݶ��ki�r�SAP�i��Ǹ�8,��|����/aF42R�P�|��_�\C&�^���$���f���C�(߄��ch$q�E� r��0��;��ďa!�Q!Z�g� :L�A�a�T�w�9z�f��J��������za0���?ݏ�p�AE}B���!}�w�ȹ`�t���wxw���,{���5+y�I�ʌ�dޗF�&wE�+7�3�v�y	��H�+g�M:�zG���m&�g>@�#Hdv�׶4]T�\�z{4"홰��ՀcN��Ç!�-�%+���H�c����g�1�1���H�9\��N��?��y��k�>m>[�\�gϞ-���������o�p�G�0$�E��3�B��1�p��Þ4��n^zM�t�R�ǋ�o/�;LDy�q[���(C�0�Ϧ1�-��"ֈ����/_�/A�8��J��*�F��~������F�����\]�����t{�=�D�z���F>OX���${F���C7�����E�o���I���=�nz���?���ſ��B���9��	�w�5Ce? ���59snF�����|@��=<V�����?��?1/�aAz'�(��{�� �y�ea��F��?w
;fH�|�Đ�;`NFخ����WE�En!����4&�`�9�g3���e�ѳ�/=�Vp�]6Vv�N]�������+��G�no�������k�tn�JNܜ'i�[A����h{%�m��BTȹ|���`7߭D���2c �����'�՚�c\8j�[�9��y��S$t�Je�S>��9	k�U�m �츍,�)pIQf��qa��G��T�8�"G>�R���p��q]``0;/���2Mu��	bB��ʣ�YK^g"��ޡ,R?���Y�8%�O��x�Ec;Yn/p�"psn"E,�[�U^�x�c$}��.��[W)Y�"��<�`o~���u��wV���t��s`�s�o�\axQ#�f�
����	)~_��Q��E�#gSK��� �z�E=�T�ȑ���J�rhXt,��:K��5�I���] ��&v�zTH��y�x'��NTGEO�r��S��7�j�-�af0�F��N�Wv��`T'܇2�2|�B�R��n���5�*(� (0��b1���
9��q�m.���a���+YpM��gE�YmL+M�J���r+L\m���������H��<-)\�H�������)�9�ъ���2h��C��:�b�-�uR��0�<����-�N��`����ɸ��W��<؛��̃T�D���5��L$J�5����=�pg�Q�6��POLK!���������9;g�Cz�T��ƒ�`^��F�Q���[��A��K�h0�-W+1�r�~2��zi>�Z�Gp��xhqs��b���J�>}�G�����^��xO�]�+�j���m @��`��� n����i�G����B�p��M��}�H�՚L��?���X�I�Ռ����� @�F���<2`�Gf�U���������G���rr9�/Ӫt�Z��m�x���YU���5� ��8*�W	�G�v?f�G��PXCY���T�"�L�y� �}h#�ֻ���$��m�<�؄�N�)�0�<�GG&�A/���)�Y��b9���p�ʄ	�~5�l�qs����o7t�NÁ�՗�.&���n>O�G|@��*�[��aJA �k���o�������W�p��l6< ����L�^K�s�����-�Sm�������G��p.��4�N��G�G}��#�n8��a���j_����P�fK�<	�e��+�a_�������@V9C|7õ!�3=�h~�h-�R^V�O�{��,�	um�7����(`��y�u*L����,�ޮ����&Սv��g���J?e����M�x�E�?��Q�����8F���F�g���-&_
��d4�}��%X���)��G��+����M����o{��^^���.���9X��xrT�C���vX?�[�_�*�WG�0����EmcEp��¤^Ym���	�`B��j�X=�^�rﳶ��|˦�Y��uL��'�:��[>Yɐ��AR*��<,]z=>"<\�����m������R�ɻ���:.s��j���)���eK��Qw���Q��}�O�
_�P��������;�.N}\�m-lM�x�����^�տn���(<K8'|;�͢�0N���QX����[@���0joF�.�۔��(N�X�sW��W3]�O_iׇu�n�9I�.)a�4��&#}���vL)���D&ތ��ؔ���^�=�?˽��,�+B�e�፥+�_��@O��0��ALDkb�[�.=<ydz�Z�L��i����W*���6d%��C�`\�k�3g5�W4�3�0�ҷ!�d�,�� /M��!�d״�.J8��Qw��<Hp;�4"�@i��P!Ȓ��}��z��y~Zc�5t�t������+̍�$��(\�бp��
3ļ*pt��OC�/"���@�b��������~���l([,Uk�-X
��e��4�ʎ��#�)ץ%)x<�}�YTө�F�<�#���pz�!x��A?�Y]5�)b?�8" 8A`k���;�"?��N���~��_�8��6J,gM�����,=�	�/D�-\�6D��R�z�-\#�i��q�;iaU3���~e�񎂜��q-Fq����ҟ�p����efՠ"�Ë�FA�>/^	@��Y�N�MqBC��q�N�ʖy�pp�g�*��R�mՂN��`�-r��0���U�`y�NJR�w%��R��ZJ�{�@��b��,�I��5~�׏������֖�h���5`��૲+A�r��b��f�cd&�z�EÁ�.1�g-���D�`L#����t��{C����z
̓���P,�����ЬN�ȍvk��
S�TǄ%�R2˃�;�G[Z���X�QJ)���Q�R�œ?�s�s�7e�-]�q[I}��e�����r�m虶v=�ޕ�W��?�sCw)aK�2�n	&x1�k8�u�:�6��Rf�.%�����[��lf�^+���r���o}Ck���W�{	J�!b�^�� �����ǇX!X2	�����|���)�w�b��O��u�������r0�Wt���C+��(-��hF�`Q�E��QT�b�m"}�mG�����D{vj���}��6j��5��[9���!���Y�,|f5.�n�g�n��,X����q5�����+�T�o�(��AoV;e7��eS��Vu0��}������U�¢ɡ��t�u��)�����<db	�±a����o�v��	�pp����ӟ��̂�Ë+���p����d(��or����oGq�Tɓ<����0:�:.K9UG�}Ј|Rf�k���W��ۇtt<��.W�:v�G͌�)�G�X����a�D^�1�]N �<C��s���ذ^�wT�,]&0Q��3��I��0�M��7eY��8|�p?�Q��}FH����of2��f���L�B���Po�
>�~�2<�l����5Iɻe�J���N�U�c�'��2�Zi[z:I��(��x��6�4cy��nbE�K9a��7��<r�*j�`�SI	[{�%d#�WgC���U�%X=S�j�%���|�`�󼟦 x5��un��TqiL4GM'x���!�(a�1C��3yQ\j`�\g/)�j���=5M�ж7fW\>�`+@ï
Z�=V���.�u���N`�g���VK��U���m��qೈ��|1�L7�oN��Jˆ2�4!0e�`�x�^<Tԉ;�ר8>�h؈C���b�v5�2���R��g1�Y@QQ#(=�^n���h�'L��QN
���9)��ܶ����5>����RxEC���u6Ci�[tP�0C/�ӱ3re����o�P�^��Q^U���1�.3��R��Qw��0^����3��XyR<k0W��_*=K�Lg���v��rbS�Ü���*G/OQ�7X��*ȫ��.,�!5�Xa�#���Ou���o�Chj{E1+��6~'�K��������=m���|�6ŋ������\~-�M�b!�H�JyV=5�/am�����r���x�k�J�j,��	[[9�p�bC�Ж��C��g�v������:�OJ,oL�6,��\Kㄒ)[�(��fDa�uJ�ӡ�+��͚l)�|��e�nʊ%T��m�,Q��m���sz
��hD�4�5!A'��KI��ә�#��^"s����6�s��XJ��ưyJII�������Z���^��o�y�����ŀ����GښSGC��-���<hh��o��W'|$��}�m�x�xuf��e����Q�`�����O���K8LQ�� ���}������í�5�U�R9�y�"yTa��G߇g�2����/�Ȅ�o����7Ѫ��Ix�U:����G;�x=ȍ�/�KB��A���?䡜��,T)`�*��}��WC
Cbd�o�������i���Y���}���u�)4_O�.��]	S�=Yz  @ IDAT`���xҷm}fy���Y{/��0L�ʮ68�?Y/����-���?��?T�ߗ�R��udl�_~u���r�}w־od�z�+�%��˾��,��m�G�Y���tЉ�?囶��[��GuXWY���Lg���Z�M�`/�����6S��5�W��:���:�M����+���i�O��Y�S��˝���~����5x�'
x��[fշ�,���P�O�Sr>/���d���f���vLG�W��aB����+m���R�/�S����j�u�I��Vr� )&�"��J�	c�M��Kװ�V��0G�����Ӵ���Y��!w5>(#B)j��vKp��1�I�k6�8�b`i���?��4��7��x��i�F���Ĕ�����a�F�[��$K�I�[%S�e��i�"�Zv>̱��ٯ��[�4�iH}��x_i�Є�;-�������/r��`�Bd��X��i���c�
�0�P�#L�j����j��_~Ջ������y��i�w�0c�*�B�b4�����e��2\�H�&��~a6�1j�����e�e��|P��z|�Nkv�+��>��W�V׿�����R:����T���ʄռ50�kVr�)P��@��!�������+�ѵ��b�N�	/m�
��~�̶+-��$Nc������c��������'�^3!�����F;+ó*�acȲ�������x���V��7L%��x���i��D����q3r����fv>i��*�y�޹y|��Æ�p�5|���ɢ�3X���bt��^��`xvQ��l,��0C�(��RXU����*fs������c��uJ��&Ȓ�2
�SJ̚��0Kأ�V�����f��T�����m�;.��l?�a�����naZ�t�"������NZK�rP`5���r%�Џzy�R'W���᫿|�E�Q(8�����T7|U����Fq{]|kB=J��������3;	��ӗ	�`x43OR��k
e��ޱ���oQ��Z����7�~3��R����G ����r0<nF���{�kk����ۄ�_����X����N1�a��Qcy�ǚq��[>iX���aF�7�ݫ������ʚ~�`q��6���
�(a]-�=��!��NG ��}��l;�%�r|��$)���7p�
3��A�t��ף'�I����(�ҋ��Yϩ\�� ���n����)a����0J�tF	�T��{���Gp�R��1�1��ju�	��N�FQ�y�:��=X���
���9eж�L;+����-=p�]m/ʁ-G�ZuY�io:��C$:���*�d�b1��Yˋ�Իr���7��W���U�"���
)_+�xr�i��8ٍƮ��E�W��L���t-��S퇻Ï�ϥL�k瓸��u��i��� ����=��9�����*wm�u��*�@_��W�-����έk%~x���w���a�� +�E�Y��N	?��?����Ȳ����I�-D��09��;v'��ь�ņq��^}��_Y��3�]�L�Y
���с�L�9�sk�,^~~�pC�]�ʞD%X"235�.��̐��7|�Y�B�zʔ*�l���;Ș���O �h�[�q�h��q��0;�c��S�i�M�\q�E+��Mi���L�5"�
��J�B��|`���8��$�d��k� �)b����Ҫ2�L�����C���AB��V�^�2}?͢v;d���������}���텫����w)E_����@2��MD�1a+P�xb�/��=[�i��,ƹ�u6��n>e�R�͔1�v������a�Ű��~y}�㟿s�5�lʋ��P��.�1A�%��n�f-1`���¿�Z�N3�>Ȑx�p�ɫ�ó����	���8���01��˔�sC������@8��oj���ŕ�R��B��0�ՠE�D8?���]/ܕ�37��;����٦֛y�Yu�k�/�1̳�z{�#��
��b��X����5/�k�,m����*Sl��_È�j^�^,Er���WL�]�%$	�_G ���ĩ�f���5x����X�ף�|���3��vg��4ef��1�')`R�!��~�H��)����Yy�a�oս�d}=�R;3L��Ű��;�4_~�p��q�X�Jx��aC1mQ��h��5���0�|�Ѿ4��m<�Zªa]�@�8��"Y^W|���:�ҋoX��}���͊�^�eM��+�j��Cb��{)���srk�MG����q��ݬ_ߥ\=��0X</|�u>��j��`6hΚӬM�!��S��w)_w��z��"�SҬ!�z`f��N�J���˿�)Z�WY�Qf�F~^�py+���|�2��Ѭ�6�ٔ5������U��{	'�(�1�úD������%��0�N��β��e��ɠ\;�ՃHQw?�1��>�}��?4�<}��p��4$��p�����%^�Y�Y[~c�Q�>���gȨ��6�σ$~�0�N�-����	��:��I�ţz%�(J[�KZ�V�~~�$�u�@׃m�(`ҙ!��`��R���Sؽ-RD�*�ᤞ�˩����e|����I��J��X�������ڧr9Jv�Un��"T;M��Z�:�E��r�+��~,����|O�)�W)`�ɇcC��-�Yj��$�o�����k�x��ן6��֨kˣ\X�8ͯu�Um�+}yN>�;y���S�������u輜����*���ĕ���N'ϕ�$��Q�*�:R?\N���T����'��-�Dnu.�c���A~^��J�4�	���o�����eJ�y�kL�A��v�i2qx��y�w9D��� �~���
�Qp0�1�n~�F6$/}���i������Ǳ�A3x!v�aη�̣'zb	�4��|=R�fx�Yw���[σ����b�k�����|�fx���ݺy�|�J޿>|�INǑ�Ŕ�mR����_����a��T�"VV(>.�6%�hͬ{qژn��gV+6n�꥘���a	�R��AXf�����?���y��Ə#|�Mi@f�YO�Ņ}Ť\ϑ��L$�aAz�x�����&LGP�a�VJ�F�`<��zK��-�;3���j[��W����㮗PY1s�Jo�J0��*<�R/��UӤ�e�H��p~��f��˕����G�=����aF,$7�UgX������@8?�z@�ڬ�ի��廓"w����4�(V�W��P�4ɩ�`�|���Cݖ�Mh);Ƅa�ԥ@_ɯ�f��α��J&-�
_�j&\�9�g�|���M=��_��u�8�`��UH�)*:-��',BeO���L�a\����d��L�����u-A��RKvD?e=�k���H+��:`y��!�Q��MZ����x�(�dV�/�;�Ͱl�d>�[��y֡�u����I�U3���u�^|�B��]�֯�N�:j]Bk�M/���l�h�r�����nV`4,c��g8k H�X��_�����%��]OR,��pv0�)^c�&m^;��W��5�M�3p)c���}w7K��Z��X{���
�'lw���,��b4S�ݔ^8�n(P+��SO^�Xz^��(�|��������e�����ry�%Y�R*�{]����?ԉ��!�W��ه˃x���v	vjh�`����9m	Q?ÿ}�MO����%ʂ�V�y'�q���/_4�l,�����ƴ�ł��N���IC���\������8�!gO��m������1�M����|w��t9��z�`��S7���>q�6���4��z�����\KhJ�E�щ�T��8���O�eZQ���-���0�4ؿ�j�.��ϔW�:���	]��X�({:;+/H��Ѯ4�;�����)�T��:����u��]N.p�����#���@��/>;|�!㣏�K�j��H�5�H�`ؖ ^�X��,��#��<�j�zt�w�o�󺟍���"�)��Gx��o�Ng�B6�U� z���:k��?K����_�|?���1hiGǆ�4tD���2G[��[7L�(�g�����k�1hT�^d�NC]�^PB �}������)J� �4���
�U�,��ק���SdfHn�R�ʟr �3����AIBo�a����>jX��n'Ԯ�}oz�?5��<�fY��1(V��G����`w��j��J~Х��Gx'��?|w��6(eyQ���h,`M���˯���(Z<�1����a���^�1.=��z	O�64Uo޾v�Iq#�/����+��Y����e�Ð,FKȌ�z�� ܝ���U�&(���5���F8}?K����P���Ƌ����r�e�y��+����/t9&{l����C�Z|�.
�L�gg$��L��k�bͬ��q��`���Q C/ךn|�p�͛Y�3΍��W�7�D��ᇶ�!X녰��o$ ���h��zq3$�U%�t�w�=��\9S=��T��+ ���,L�R͠c���:L�V�����ÏR�j�E�F���ִ7
��cQ�w�����q���e9�e��w��t<i;'3�X�VG)��=�.��eJ� P:�<�������Sk��i�U��7�1lq3�Q~���YfA:�+���C�v}W���f��E;2��
�a�k����k+��~�0=��穣����Y�B�v��Y �?��E�ږe.f�3��˰��s
y�����X8�&��Y��E/Y�Z[��c�6~<��a���C;4�aO����xá��-��0�[à|f���<Jh�e�c���~CS:��ͰK�ϑ���)�,k�H�XC��Z[�x�'ʘ"Z2��?�T|m�B�v�b-x�og��[�n�0\1�q�-����Ě8�B��XiBaU�ĉ��f�Ӌ�7�"2���|�x�O����]<v�Q������Ӽ��$�bl�S��8�cבgR��\�(�����N �>a$����4oV���	~8��O��������u�[���ۋ�Qxz9C�>�p�n"��φ��m��%����5F���1מ�e_�Vi�u��C��hD��#�>��EK�(=�O�h�/'@KH�g�I���#���|v�ͯ?;|�_�`_'�َ�,G�	�Y��y!����+�)��Sx�[F/�-�W�� ��+�⪚��J���^XXp�#t�hO�Rp�;ް���F�G��םJ�Zb��Ad����׳��xV��L�ҥ��^��N+l� �����$���>�����<*�bA�IO�&ˀx��U��3�Uo]!�
��}i��3��E�3O:��C��qb�[�o�6c���?H	�S�~��{�/2e�i�s���?���Ãm+��3����,~�,D�<��r�.���C��4��Q��E*�K�2F}j(�Z5-թaP:�L���W�i��IO%��a��4��:�Yo�B�$����ƼQ�r]x��Gw,|�K�4�5?O�`:�;JN��L�2l7[��1���	R�ȎS�͸_q0)�Y[�"7K3�#�J�{�EWr(��2]���I`T�+�(�k��cK��z�5��ʣt��yJ�9��
ܮ~O3]�b�M�j��6�h�mX�a�C�Si`B�6|���i[+4�k֐5���ywTڳqv4`�8y[��3q!Ƴ�Y���S�9k���pgi'����Y[�W�eM�����_6��������:��gx����c������ȴ��R���S����s5֖��X�?4_o��E�����orB�����C�xX>���r��QJ��rN�U��Q̮6�غY�e�E�V������L!�#��b��A��XMY�ia�~��?���Ì��-��Y��K�/���!��@���IQ<;|��w3q�r�=���A�j[�F�
���]-���X�sU`ţt?����j�K�Ǥ��9�p�x���vG����ݳ,=X��c����~?�t�j'�"j�Me	��	�jC'(�w�?k�B��[*����ꨎ$Z�TWu\�{���)ϡ���gŋ�:�y����#_3�_[�;Jps�0:QN��5
��aTY�<�$����>�� .m7�L�'[���A[(���۝��Џ`s�.�8���_qߏ�/0<8��y�q-~/G0�8+<���N�[��"�����	�%�L&�ɵHsݲ�p�/� �}n�3Z�au���.����T��@��F�{�z�<Jc������[J	�Pf���]H��qxf�9�m ���WP|j�1��:X����}#���z���������Y���g�=K�Na[{���ε(ިce��@Z����Sr�m������Ⱦ1ؚ@>@���B]�U��Ϻ�Z�.�  ?^8Y��W!�-=��rVgR������?�o~��xi� K_���`��ެ[�ar���n1����$��N���mȆf�wEe��@{�)�����!�gL:!�e�cU�"ة`�3ģ�'�	�5��]%���_0g��?�^��'�`�-�yl���w)cwZl/K�͛���/��`�OǓ̡�9�M�F0&�3!�h/W�����|`Xi��7�fS �,3uLq>J�&�Qi[�1�9�Y_�Y��^C17Eƥ�����9�<ke`�����,��Im}x[���8���y�Qј[��!�������}7��$��pVo/Z�¹�	!8F�ˑ��'(kvE��Y��|.z�Fr����(�`wu>�`$�0K �i�XØ��g�TSL�{��ꆜ_g%��NU0�#��Acv,/�Z��2���A��^���/@0���I�xgH�e{&d^C�p�Q�X�40
~�_9��:��)V�׏,��
��j3�tTzϢ�����Dx[�c2}�Ys	�Y��f�����:�I�o��R �j��5�������R���~��o�w�w��?������K��뜬M=��E�P\p�^�{~���c~�w�g}J����<���Vڎ�f؟��A�E)��4_ԥ2W�Gu _|�c0姗��y���ȫ)��u�f�������e�x`h�������cB�� ��HY:�i�	���R�AꈰJx�a~t�3��"��$�ᡕz�,��⛔յq/8C�zDf_Os.N�1�0D��S� {e{^B��޻p��F'p�닱R�ݐ����W �6�,M�^ �_��QС��p�90�e=-zYʠs|!�N{ՀL�ͤ	���*n��^e8u,=�Is���f�[��̭GwϜ�ۻ��ܯ��mR[)�}{��y���Q{>{�	8��oBh?��n���P����'�ͫ	�'�6`|s�����w`���F],X�͞�k��G�X���8C@�j�d�(��r��~�&n���>l0/UN�=^pW�
:���)��O����%D���l�E'�fA�+1�;OS����������۝h�徑�x��г\qf�ڤ��萲�:�x*���L2BF1��7��}�Hkؾ&'YF�kB�����c4���hpS=o��U�Pe�F������-����=�=����j#��A���27o��Y�o� `�Z=K�a�[��Q=i�#ZC+k�=X�{(�Xy�1-�+� 5���*~'8� ����^0�.^̺�ӷ^լ؜�ƽt��,@��6<��2Fx���d�2�x�����~��yc�����_����ËV�VA�,�U�ᰗ-������e�"�4m,� �L�Z��1����L�Gi���1��`勢7�0�����~y����"��܋ ����}d����GK1�P( ӛ�^>�����1�"�|}�ů������M��B��fd�d�m����F�.�a6ۮ7S��
=�axhh��UV��U�Ը*	��W�p-�8��zh�{xI1Erӈj #t
�cl�d4*D��-ͺ甬��"����|Iq~U{�<4���d��Ͳ����J���&���ߗ%N�Q�&Q�j��S1V��ҳ��%x
��kRСu5���{M����L���b��@�ce�����&�a�$0o9�痖r�\m��e���S�e48V?��c]�׆{=%��e�Ni�E"�m�5�㩇J�������󇬀�̐�a7{>jw/^6��t�O����ʤ��l]�?�]
ړ��G3I�]5����W����v$H{��Ұ]y��0�!�~��ˬGv%XC�aϰ��pS�y
(e��WZp, ���5���Qtg��)���Oi��+K���>��ү�f���}h�$u�~�ϛ�^�5�����R4u�\�j��{��,��Iz�՞^ס���g	��I&e� 3�,�(��-��%nd0k��(z�&��Zِ�rPPuL3�gOP�(�r�@��lx�.�+<��kkˮ`�M��<:Q�S��*���t�E)��\�eT9Ѿ��}�z)���|R9��:�. �V���c�/���h�WT���u�^!����	"�`ld˛�WZ�IC����g��/���Ľ��t�tV�ׇo�,���OX(z�$gr�T�7**-f�	�y�:V{�v�S���U{�K_�'{��'�����ċ=�<�+�drcW�\'��u�n�$��'�����~�v�ET��l��"�Rb��>_NV�-�lI����r5�!�h/LV.��,'���2Hp_�ö�+��GOf׀��-���*�pԫ.�Z�*9�*k��(���=&����iF��n0�u�SFi���;���:Cx����� ηֳ�އ��1!Lӌ�+�!���0��h��T|���)�*q����R����̌k���HC?�bp�`�2z^o�v[>�g���(!� ��p�%OS�l���0W>3��s��� [;`3~#�U� ���`*��U3��"t�=O��P�A�}5,`4dr+��VV9
�=��E��;���A���z�|���i��=�(wH�i�X��)M��aη̟��"�-_�y�w�G�" w���-B���r�"8���L��<e�����H؞z�Z�f��|��Lk�`"ᤗ���'�-x�4g�%�
ݳ�v��z[/�z-����nk��(?#L�~���Z6�g��|J����`�.e'hF^�vB��^�ӫ�\N���`�cR΢?a��ҁ��e�R<����$xį����i,�Qzz��e;뛽J	y��%�m�t�a�rՂ������q~)��)B��+�r<�J��7?����ɰv�fiQ����4�zš��T���T�Qb����usp�!�:Ӯ×���5�\ڵ!�� ��������e��O�̄��Q�Rn�j�[Kہ��b"�`F�)j��#�ae$Fy�5J��O�(k�d�5.�a�j"��9������l-8(J9Z�u�/�L�n�dT��V`�xE�7�Iw�`)��$�(�Ewt�Ԝ¬����G_{��\g�bKPb���){m#������NV���Cm�����ݼ�n�����p,Ǫ�-�Ii%�RXmw�ҟ���-� W	��-���&��JQ�˄�f�m�S��K�[����e�p���{s���4��p��_�������"L�}�yZ��W��-i��v��}�:�׷ށm�$�l��B�ԣ�i��� �^E���u{��5\x�m!&�X��r����pJW~��8bl|��T���g�����~v�UW�T/20J�0���}Vg�/��ڴ"�83i�ޒ���)`c�*_��kq�J/���ih�4,�Fo��E+�F��S�OnWy��׹e�&%qa���l�<;H� w:���g̸5�r��>i�l���J�9��~xz�Ch��̸���6�g����l2ʇ��a4� ]�C 3��.F��S%�Ф�ɓ������d�鎃��0�ِ���4�0���ڂ��i�I+ǌ������>�|nNۆ�?�״��S�B��-�����Y�ꤷɊ�	8�1!�\JC�FA��<�#�@+�#�tT"�N�|��+%�O����ه,�iΟ���"ja�'1�wr�6<4C����w2�Ά���L2�9�`?h%����Z���M���T�����C=�0ŗB%-
7����!�ٳ.|�h��俆HSqM�/��$�Wq�9"_��%��;=n�׫އ�tM�J_6�9[/Q���@�%�L]LZ՗<�c�c���uq(��f[��<ZG�R��K_��fsU��]��>��lxWp3��zSɊ�v7x��UC����Y�G��QxM�����U��r�$߰^���s���aA���j2[��GX����l�E2��u���x|�R*jsS��?L�6�.���S2^��W/R��X��}�������~\�V�|��D��nh�ڀ��4ZdS{�k�Q[Ѯ_�71�zGᕾ£2�(����]\��2�)��m�5�:/��@Z��@4y����j�1�!}���r�8���g'7�l|�nch��|*P��V�k� �Vy4�iYra%z�3�[Y�ze��bxgضD����Q[���la�<Jq(
�ȫx�X(_,lcp��-�+���t��gñ�Y�����(���rR�K	Zý+Ԏ7��?§pmݟc��ܕ�b)�:.��)��W�l�u�j9;l赬�z�t�S0�n� �$*�C�]����q'�2^�C���4)�������d1�{���%���s��9|½\��\�����a�b�YIm����U��'���`uV��?<�v99T��pp�~�R��v�8���'PF���Wٔ1�M/���E���*��}��2�_�S���z}9>����������os�i�ňFퟜ|��+��z��ӟ~���VK;���hRdL����\���So���>�����-fF32-~�
�ʇ3��U~ߔ��v���3օ��{#�CR�hurۄ�]��Nuɣ7H�vo��������F�3�5>{����F<\�|ȫ5�n~I/k�cԉ��#���J6���J��Izg�Ti���+��㨱_N�9!8�&g��x����R�^T�R���9&��c��pY�0|�ȧd�2�z�S`\>����u�Ժ$��j$�+���z�U4D�o.��Y%L��l���K��֭�4�� �	����￨�N�i%毬��h�����)NmP���iL���l�%�G1)}�����ӫ�ϳ�XTP��aڸ5n���i!H+>[�ق�V����:�^������P̖gFqFX7t��	UK0pbWËOG�-vu�r��KG�{8��^�J>-�a!��8��B���WD�֊4,��ʷ�G��OQI܆���(��ZV�Q�k̆4/�|Sg��\tZ���4
N��*��M	���t,WBh<�1���Y��-��ge'��i�J0����HƂ�?��y����9YW�]
�9�=)f�������l[�5(��D�=���|Xg,LL���Y��o�S���_�3?0Cgz�pM9�w�ߥ|ќ�����gH��I(������j���R�]�S:w>Q�<�:/�Y�L��ݢ�U�+�Q뫇o}��Խzh�r�^�;���2����(SwpF���`Yu%guڿ�'��
ͤ��i,E˰rJ����{C�6%��k�hA-�b�a��K�g��,�5.�Y��C:�\SP9����t���΢'âӆ�
܃�A�*l��ٺ�����(���#�Dq���XA��� 8\q�Ȟ�����TL����]���ވ�}��Ôc�{�`����#�>58A���q���v�&���3%��ҙc�[�����n��(�]糟U�y�Y������l��)0z�����E��%`��k�ʡ7ݏZ?�6+N���;��n���𸌧�JZ�wթ��*S9o<s�">:��A���D��uB?|���׿�E���GQ��D���p���n��|���[�q�`<Z�r�J��agk�K�E��+L�G�\m�].7\oX�F�)(}�R5�\�z�N�/m-@X#+���0��<-�s-�$����X쇿/Y4���$ƀ1Ʉ�I9B�+�^����̰ŦYE���S�x%f	Z�^�8�؋��4�����h90����,�Bc,Ef�q^=MȘ�x�����t�hc�+��Ę���J����g	��!���hhϊ���n֟�h���;J�y�_���_}�26�_��Y�����&l0�0Q>	��n2΁�A��Ǥuˮ&��o��]/��?������.^����O1�K������f26>�S��=��Ō��y�襎_ǤK� ���$�^QWKM���y��?�a,`�\EJ�x8_:�/{�Qg(�t�m���m�#�뭘~3��OYH/E+�a�uB֐�U~Y����B��زnf�lX�p�`��L\s�z:�N4`v%e�u*�����N�r�:�Dk�f�
��Otj�M0� �t���5��Gx����*t��)����pO8�ϰQxJ�� �ה�5����WنDȪc`�x�:`�)�f���E3�El�t@�J�DP�'Õ|�(S���_Q������`���߲���77�l��dzپj� q���Na�L��,�p������:*X�/K��IPP	K�<�L"�o0Rz�zD�Q\x�e����=��N*|,KJ��������ed�ѷ�۞,3��=kU�y���<�m�e-\([�l4%���	��Oꆂ�2��,I�M;7V�Y�:(�^̤��`:��-�9
Q0�8�z�z����xi���+���.L�Wt���ǳmŏ�6>�Y��� �%m�3?-���A�^pS~����N����T���ʷ0�
��|���2Ǽ/\e�%e�:��N��c��H���ۍt %���;�~���[ܟ}*�|�?/��g�<��|�/[���o��� ��1�.����w���"��ۛ��M�����㽴���!��i?��z��i/���'e'�ZNh���o��ޢ>a�x�Y�M�!�X�W�x��0ɂSY�O��U��j�j�����i4�a�k�e}Q��k:˭ك~��ÝW�7:dB��͕�z^P���ֵ&;xZ4\���	7
�2��%��5C����b����d��ԍ���U,��b�|�53��5K+�N��eE�k{xYz���H��&���La�>���	�4��0���L��f[��
� @�8fB��	����n��2�	����p��p$�L/��1�[̈́������}0J�F_ĢJ���{��v!>��AX.% i�3�5.�:/V���0��;w�Jha���_�����֎�'��<M�7[�vF���Lō�J!��3��Q��2��+B���Z).��\
��A.5�ex�d��y�jV��U��#�sq�C���)�B�&?�k�N�c�w��-][n�Ќ�fW�?~��А ��E��sC^�ﲀ%��@ �$]�r��az���,�X�U���p[�1���oj
Bg=�pYĵ�\3� uDC�P�ip�}fA�E�U��(��o�P\��P��Ux�:KX��=zPC��L���k�jCs�[_�J��cˑ@�&��+�E{���l�0��rƼ�C�O?���-|�5��y�0ц�{���׷M��M�}���ܐ�e.��(+�K4Y��S��1�Ro������y�������m8Ń��)6���N(!�R�I��F	S�J�7m�GHY��R����{�ٻp��t^
�f�#V�w�0�=/��j����(�y�L���(��ye����zN��e7��(���%�h���I	.
�8�� ���]�-|!��|Ǌ7������K����h���/c�~�S޽�q�?,A2���|ɣx�/N���k��z����Ȕ�t��u��^d�ز�{��-W�E��aY6�B����*�yY�n&���|�gqa���(g��S�bm�\��O��븸��G����}"��N/�_�؃��Nq��c���,HW9mHf���R��2��J~=���2��d�Q�W}���z���z�wo�/j�\;��`O]�k����]�c��o��Cyr݋����VW�$G�yW���YzX��f���)/U/���U�OO�����٧Ƌ�c�8ف�F��j����Cz�N�T��*c����r�vA��W����x�o;7Nq��xG-�>N���&\�ZZ�D:{�[�b�/m���z����jג�\�`�P��DЊ�7Jk�c.?��e��1T�L!�����H�3+��o�*)_#b�	o���+��1=q��
��8�;�+P�8����G!����3�-�F�� [Ew5���!S7�x-��J`�{����䓫ƟC�����c�)}��f���_�O����G��Sii��,�o�O#�J�%�4��Y3:# ��� ��o���!�ogY�ڿۢ�@2��e��.S9� ݣ�eAH��`S����7�:ʖ		`�����w,���=��m��
6���XC��ߕsz��@�`�Nt1�D'��)��O�~����Q�Rߒ��f�S6��η�%�j
��:=)ኙz��"�5\�Вo3��D�1���"S�����2=����;�`��Z���)�j���X���U������O)�w�Nn�6�����A���m�t������H����7�R�2�˷$���L8�I]���öm����~r�w������h��k�1����"}��^o��ZTԦ޳�{~cW���>�aC�&� Y��ɡ�YX7_�/��݇+`�>��k�������M�͠V���9�8F0�ɺ,��G�,_J��G�XM2_2�z�ۂ�~V����G�K� LuS����Z��[��F/�(��¹���Q֓��]��h���E�]�O�@u3m3��U��E[[F�Ъc��^�f/)�c��~9JfyN����>Lh�����Ϩ¬�(�i[.�2���y/�̀n�$��r�@g�G�Ў���e���-���D����?[����N~ʱެ���V�Qtuccf��|i_?x����,�Io�ᕀ�1%�\W�9E����s-D��C�-Λ�z�J�v��EY�D`_Vo����T�'y�'���+�	;觇��+ޛ��<��(?K�G0��{Ǜ���&��,�{��*|_���jZ��|�iFV~z���R"����!��[��Z��'�W���z��5ș^a���uH��V�r~����>��7���x����6ry|��%����ڲ(�G�2yӁ�b`NI�ȣ�s��f�0��,�-|�`D����4gG�-���B�E�7u:@����j�u�n��M:�R�p��3r���~�o���u�p=x1V���BC�4�4DaAL
k�%�%&&~Vx�,CD��S�#��,�Ҙ��榗S��R�u2*�q�4\O��~V�C-�\��$D(WC�5�h��n�#��,ajvS?��s<�&%̶�B�Y����Y�^F	������"�ɬ0nO{T^g������tٝ���,���a,6����.±ЫM�_��N�ba��m��<m���(�g�
��!i�l���?oCb����|�¯C5��͚b8f���a�����Պre�'f�{@��f�4)�fx�z���U�,0�8	�L�6\�(R̏��7�r��ᷲ�eɩ4O+�v�ѐ��v�(�2��͔�����A�^��K
pp���gm\>5�j�����M����H�e�q?Oѹ����o�
LJP���z?h��y��/,�Y��V�Pap�9X�%aX��(�����w!�n?d��o��ml�n�y�)��:���	'V����V��y�߷�W��V�?�!�Ѫ�2�ki�x�L������ig���sZ���]rC;�e	�X��i�V��T�Bg��L։�.��M�[�~Y��Qx�Č��r�S��+@�cm{�y>��wNlћ�h��it�����]�:�����"	�"�0<�4d�!��]�*�K�!���)1�wy~>�5�I!d�U�M�L��j�[jh��Z|��)����C��R'��k�|)�X<w��(`���ٕ�QyZ`�L��e"��O��AS��Zf;���V�`���	�2d�d8�[�XuO�|���Iѹ���)��2�\�=��`⮰~���F"��8�t���T��o�/�����Q�_$�ś��仙��4��V1B��p?��i�4I���}�i�0��8x�@֤��k�|�,��+�UY*�>�[�0+�2��������ao��N
筶�|C��-C  @ IDAT{{���Q�N'���:G�=L��3p���_f���y~_g�	|��uԒ|J�\��>�7����d<ЬҨK�����{a���c9��&���������`�;��l�ʯ�t�+�T������m���W��/ �H}��P0Ǭ���/�R/�꜈���8j��BX�l�9�<Dܻי8�.�m���"��䏕2��ۀ������	w�-[<��-3�'��tx�����t���P\����kV�J�2�#���q�:+�1`_���4��׿���D���?��p���h��3����+x�p�2Wf��/���L���@��`�G^'aw��2���*��cF�O?]:�����-6��4Í�!c�Z�YV,R����S���U��c�6��_��Nf�X�8��G#a)���,͐��jf͙
\���ef�S��P�������s��JCx�G��������iG��3i�f�~��O>m�A=��9��c��r�
��,`��T�V��Dd��3%��D��Y���D�x�n�_�����Yݒ��o�%���dK1{nE�����׺3��x��~���Z���᷿���7��6��b:�7����B�ij?��-���Y��w�s�Ǐ��9�w�+Yj���f�<�|��X���@��j�ך0s|z�a�:.�,C�6ǲR:�5-F����q5��)�+}݈�P+ߣ�{f��bP�b|���ơj�&ɤ6x;֮'����SN�5�V�6�z�17�
!ł%x	` .���(*���-�sE��L��Ҁ����@�E��8y�"4�N��c^� mG�hh���N@p+v�����ԛ/,��&�K��I�p��1�V�+@�$��ꧼ�u/3�%#1�\�w4����DUf���TR�F�	��{r���?O�yi�!x����q�9{?$1��L�=����f�����g�z��:u��S���R���	ϣ�/���F��N���BnjdpP�
��
~�w��e~��3t]/Gq��l�
8�=�e?V�Q�����|K��k}������+���O�S�Ҝ:ݳ�u˫�@�da���%�~�������p�>嘿s,B�;�F9L`�k���^��T.��]iM��9�z���+�A�'G������91�a��	�=X���+�ш;�3���Ǉ�\�"Ռ<Y�u���#}%�~P*;�����f��+��}�����<�)�f�_z��~���������i�9�`t|҄�Q�j��}�
����|'k?% u�;$��S�o���^���h�_�;�(1!�c�O4�^�J����A*k��O`���*��7����fף
�[�V8����ݓ���9z�����aV�L�T�����.��[����z����{���G�P���wm䝊�ظ;�M"[(�(A�B�u�J�l?M�u�����s�z����xY��P�Q�uQ�����4=�Yѷ��d 0VBJ��.J�~Z��Ptb�D8�6����W��%ӊ��3	BB���ȡ�����(cZA� `9�!��Y�zc�z�{�T�jP(�]Ϗ�Ӑ_#��@�,,
eC��+m˒ ^�f����4��igMs𧬯�����o�VYV=kd��� Q�i|��au��,�+}��%R�7��e���,������~�LT�Y��/���(v�?J�E[`� ��¤;��:XD)�9��F�]���҆�)ۆÕ�#�gՓ8�l^�VB�0��1n����5��z[�mx[�e�(�L�\>7�����p$�����R��	X��`�[]9	~�]�)]:/�0po�TR��6��|N�s/]�n>N/u��yY�1H�)#e2���I0�4%��E!���2���~��o�5Ac�(��:�|=Y���/�~�3L'S��bɕ�v�*ޗr�D��~��H���΢�:���[
�!@�ા�_�9��g)_f8�j��l�U��װ���X�KO��Fw��u��8C�c������(~X-�]VwK��%���\n����R��ܺ���-l��^<eW/�~�zZ�O]Gq��/��W��������Tb5"�:����`����yWb�y�ZQ�'\i�������me���.��wW�]Ź8V�+!�)�ű"���=�7�M�+��Ƥ=F;���J�����S=�]<O��pTٌEzb���s_�X)L�����R^�(M!k��?��ˋ��;� J��)��^�܍�M�'�))]�G����W���TZ_�(~��N|�GE?���r}�g�[9P�����Z�c�;��SWC84��уq�z�܋�`L�z�P���|�P}SA��ΖpW�<�뫥��g�*�ҍ�м�«�UV�5��ƭ֭괶�Q�i��%ua��V��*\�t��^�!̽�"�!�t�k���&`�&��1`��~�.�?<����Y/�G�~��|N��P&)`Ȯ�*?3MK1��g�� כ�*>eGo�i�����~++%�0���m�NN�1݇Y-��<ςc8O���j�5�X�(�'
6���4_B�����g��,qQO�7A`Y��a�˞u�@L64~l�{��RJ=^c��OP���Wu�}y4�8�[sk��������M����`*��aD��5%�~d�RT�E�5C}����GB��$��-��(�GshY����`���q��F�_%��h�}kf���|�l�X�Z�,; ;��a<Y�2u����Q���܀)V�Y�t3S���|y���ހ��-8�A�G�:�\�P��ې�{g:��,Y�"�����o�o�>V
��n�;�S�����	.�74�΢����J�z�p0�pD�W:��K��w�l�t��Q�[�?F�S�uF�̾��2�U;^�;|eP?H�I1)Le7��Ce���ˊ^V:�|`DUk.�Sp�efZ{H!�t(NGQ+L�V;�ڐ�P������:}���f��';8����u=F羕֫�(�޴���=�k=!
����}��َ-��BD�3Q ��d��v����(a�1�rX�͞��1E��*���u���M^��e�3�N��(fQ�Ck届+�����P7��w)`�G���N]Ǫ����N�_�_%�U}Oˢ�:
>�u?7�R<
Ǌ������]���`�}ְڊ/�y��`���V鄿P��U���=�r�M; �@�L.�Xd�U�dԄF����tx)_T}�-�����F�ï0�B�rh��Mo
���l��&� t\A�Y�Қ<{F/��,>�C�t���5\�_ŗ��d̒3a�̴YH�ʜ\^�6���|�O��)�#%�hƑ��X�o�ݛϋn���eW��Y4ȭJ=�E��0����E�]`���H���q�Q��G?P���*�Ńw� j�&����dם��~�{@�B�\���aI����1c�c�*6s���޹=����[	�M����#/i]�{����0���^������qr���x���"]��z3�>�
�����nʊ��q�$�_0��H,]�,��)߶*���ȟ�q�M�עo1�*�JBְ�a��o��#V���Pbv��E
����/s �O-&�ে��=L��:R
O6��¸�w����J>��b���ë���M+�6�h�%XТ��Z+���ޫѝ^�8�̆��~9�|-47��@u0Jf�_k(y��w��b����e*��|P����S��'D���8��
կ���\`*c1������^��G�n�P�ǌ|�Vѡ���\�'��_� ~_�	)��W1\�����w ���i�?�|�Ԫ;��PUkY�wt�0�y��c���c��%ت�f�Q�Ks��s�&%̒�7+��𩼎�w{4��[o�1�Wh����s{�1�ʐ����b�1�-�����-���N�onB�9�m�MJ��٪4�I�"d5�ax��.xF��$m�!<���N@0Fp�Zmʹk��($):�7��}A��fV��lE��t���;V�|��hS��%�\����R�r ��hA�/�C�(E�G畆j����Ix�W6���c����Y;w����E����(�-��#�C1�v�E�n=[���H�v�2:��x��ٗO��S[�שS�Ҟ�!��c�My�Ǫ��	�(��P'�`
<P�x��0ނ}�[��;i���َ	_�	���,��{�|Dz�ߕ�����-�.N)K|��x�7�z-��o=�:p/�ee��ޮC,+E��X)�ub-��덎��>V��fb�.�ds��
�s�3ч{G�=h_��d=yNp	HY,\mJP�]��y��ֈR��@ɞ�Y�6��O�ՑM��Q�t�J7K�>�Є�!���ܕ�����z���w慯+�z�>����X�_��=Kr�|��2L�Ǩ����N@��<���Y�A*����x���{�Z�[/��vO���WF�j͔�����/�̒hf�V4A���L������̀4H��jS�-��.��S�-�^|�f Y�݈��W�t��#/�Q���9ș�YEB�{M}�����lY�f�B�I�6��iJ���d��)A�f9�lb���}k��m����C{̒��F}��զ��GM_Mſ|�^B�O)3$Ec���㶍9+sZ��J���u۰�y��~<��/���ӆ=�j�fT6����� �k ��0@��- G)9+C��>jc�?���~���4��$����|B*�L�if�G�����u��|NY��=!l���,`')`��d�9u����z
��Z?�g3�*~�35V��SNO�ޙ�A����|��(�c��&y\o/��,:G-x�<�����N����*�-E�a`L����E��ey�0�f��(��V�KQ��>V��ynX�`�����	�Wm���e㧕O=�o�@�Q�X�Ϊg
�;�XE�aj��9F��SJ��-����Y���Oz_0NKgY�JB�l�Mo\��wp���W+ǮxYvd����9�wJ�Z�	~N�Q���,��`�5�i꡺��3�'�a)!��/�Ҙ���9��p�ЄD� e<O+_�����L}�5�I�Ճ)��h
1��b��9K7D_��t5$o,h\���5�L���n�-���Q��'�_o�:u��eG����&��\>_Y���j<>Y�	�_����/57%p��#r��<M���k7�M��v��_+��jh��}���'ڝ��Y�(iv|0���zf}�T�ҳ�z͓�U�1.L�W��!�p�ꐢ�v���V�|���	��s�>澄ĝ�����~�	*�w��=L�ni�L:�o�].	�u�i�:���:����:����eBx��=��c�p
�
$dgy��qg�������"�����$ɘ2����~��W��qRW�t��ׇ�UttK�s)4Z[�1�i���,d��g6פٻo2�tr����������]���N��No
����;F��vO�/48��Y��#<;�hsd��߽�:�נ����<؛���[!�d�u��+א���̌��n�6�xDC�����YC
�ҟW�{��������`G���\Kb����G�3ԓU	�&�
JPu����R�޻Fc�N��E��v��`���-:�� !������K-kp-��i=����W_�Ԅ��|r�h��
�٬KSr�Y!�/��Ys-?�,z�/������p�����{1�����$�g9��j(�6x��칯���Yv�ZH0$E��qq����{�aP�pV�a`,��?��{0J[�/��uѾKq����r&H(�O)���a+�����T������P��~S�OM˭��_���iP
/��VC_s��cj���{1����4z)�|t��(b�	K"+�^�q�^��Zs�R߬�9�g|���+��v�����-����f�F8_�+ey� �+G�.�O�6tc�7�ސ�a+��b1�n(�zUk��|�G���M.��`��X�&%0)r�����a�(R���w�~0�a2�e�L*��eC篮F#)�S?SW���YrB�M=���_���U��et!�hp%B���b�HN[@]K!w.k�d���W6��I�b��C��r�*�Qf�~�8�b D'����߫�������� � �C�
�]S6���Ktz�}W��S���p�Q��Q�am�����){���<]iͺ��0+�똥N�>yϺ6�P��%+��s�}�<����כ$s��)`���/�F�OZOy�ޥ��8ܨm;YV���u6�����
}l�7k�3�NK��Y���,11H����_� ����`�R�s���c�=��[�=�%%��G����ݞ�
#	u&�u?7o��i����N�k��0{�� g���߄ߋ�v�r��:��g8|A���NZt3;h���c���%��q� �Jr�����
����7�������6�����~��95׊,�
3���:��"g���8��n:�-oJێi�/�l��.o}�ob�)���0{�&�_�;����D�=xfgȰ@,���� � ����8�2�
�σ��=͟�Hkk\��a�����І&���t�MB�����)A�7���~;É���Q��j��"xOn{Ყ�_��jhq��
�U�%�[LS�i�E�ޝS��<[/�<���+1���8�Q���Y����W_}�l�Ŵ^��j��G-%�4�ΫǮgr�֭�-2g5`ӝ�ʗ#�3��"�Y5=�9�Ճp�8�8Lg�j}��Ԋ������ru=�s�OYz�̾G9ϋ|�rt��p�G�6�w���ӌK���	-�2z#k�]�呂�4�`K��Y[�K�zv�w���Y+*�U�`�(4��&��pɒ	5�ݭ���>ɐg9����J��]ؙ0�JQ8�B��ޕ6����hh�x�*Ryg�}�p߅R�LHIە5Eg��w��D���>����|�i�(K@Bö�m%�侩?��>n/�.+m1$�B�t���'Sp�xk�3#k�'���D+�Ugiכ��0qJ _[Z*Ǆ(M�g��ɕ���Y��Q�����a�4��U��?��dؔ6��{�K`m�*��5�k?��eN�ô���(�,bƗR�`g���]i�zWޔ������A������H�*��41�k���h�%:�,d��:�GA:�(�< �{��9f؆Bc���ڗ�8�6-�{C4�%Z���V��Jp�_��?!�:6r4T=�{7B�[���Ȣʡ���Ű���bv�`��=���:f`7�i�%��O뢸�4�8xu0�r7ֻ֞lf������4�+��ً,��P���o����x/��nT��W��"e�ř��Y��U�fx�	H�f�F�Ã���5
X����?OC�f��|��sƆE�@1s��x�nT�����ە��L�������m%f��U�{����a��Cy��o��nO����%�-X�N߽x�U\������l$X���C0-�"��(&���Wfd�e|���f�zm\{�p�T�s}٢��L���Ѩ�1��&XQ�����.y�c��,^ƀ\<�y0�Hߎ"��h���u�Uz�*�]��j^����"�ǺE�u����"����x��[Y�L�IgI�<@���\��y�[w��o���sE���*��U��]�d��*@_6LIˡ��6i��ü�[9���!�=�����(�n~'�n��Гvw�yG�ƨ�qC��xL�(Xi��t�zo&�)`S8F�i^3�jX3�XC�����a�S��=]�,�KP-�2k�Bp5�R0�) ��5��3�(<��I��e֨��k�����e�@�T�#(,��
6�׃��­�7θ�%��rVe���Q��K��$�����:�~�ʎu=��.e1;�V��l�R�����u�R{�5���"<���Qj�$�hwx��ZO�c�E]ͪEIRUʲ���blhLP?�he���_ߦ���Ь���dc-�+���Ǫ5g��i96�̧/8[��EJ��fkR�� 3�_Cz����(i�������0��5�z`nqY�j�z���3D����?w�b|1<S��\���aR�(_W�'�zuwf͙�s��p}�0%q`ZӦ�b�R�шm�Xlp?��*��t,��0�w]�p4��.��
�5<����c���a)'f��MP�}i+�dO��Z|cB��£���n�4m�\���[8�ꈠ���]�R��/�@�~��~Ĭ �ƙ�9�N��^��ʙ2�~T�f�>f�S��Jۮ���ә��,�|b��N��i�{���Ż6��v�D��4��^�2�����#%ʚs�R�����uȲ�������Wu֮�'�,�R9�bf�/�Q��G�jN��F(�,7ꐽ{���>��]vi�S���t����1�6>���:�;9��|Jc���=���p�҃6��K���&��������a�[��:��
��{;���j��'0�N_vY;az��P���:b�|���97����9?�}�������E�|%5�2�Y*�2��Z�o�cxP�7>���So�:��tR���l�SVc٬`����{+EIH˛�u��s��_��=�P��� �,��{�%�Q���pn�O�}�X�	��c�����>�_�z����ۿ����!�w� ���b5~�ˁQ%�z)_,L̎[<��q�FEZ�_���v\�Yp]|�����[�b��z�'Y�.eq�;�8��f���j�1q�1"=��VY���������W�w�>iP��"���y6��S�^e�z��~�-qe��->�$���e=_�ޝ�34�q(i)h0���������k�g�{d{������t�U���sp?x����X:�^ˋyOS��))
�gʚe�L�!
�YRWR�n�t����i���[�bf�ys��c�O/�d:E�i~m�&�>V9��~7M������c�\�V��X��=���7�W>��B��}�J����H;��Jr�L'��}/�^]���X#yf���_�s��ز,K���Z����6��F���Z�5I��L$�@ ��HbZ <��A��%$��.	���0-��Y���n(��Ո
<Ym���ʩ�0i�����[�n�z�) �[r�WA}H%�-T >����Q�P�͕��Wu*t��;
�U{6�6v8�%-/1
�j��I?岌hZ��G�7���K��y:�H�fY��פ<⁪�����M�v9N���k��Q�誼	��Y��j���w�?���4y��Q1��vQ�v��9U�m@���9���U���_Q.�I�Q�i�ĳZ!z�dڸ��w����Y��N41��`����.���4���Jl��H���\���T�.�8�i���z0bf����)��SV<�.m߅S��ҥB;���[ʐ���h��ww��E�v*������C��'\�cD��<��Qi�(��&D=�,i3f�:U������qf���#��Y����=����(8U��&)XY�!�G��}��,�-Z�G��=�b�H��j���ZW���	~��?�7H�g���y�����>�H훖���4���]��߸7_��a�c���jto�Ц� ���ӣ�����wh=7��8�^�~��V�;'�i[��
�O�����y�;^ܢ`�1����z�~ �б~�,��M5H����Oy�6U+f���6S��-}W�{Y&D���}
�c-�pط�ap���|�p����z��Op��<�?U_|>8:��(���b,n��B|�>����,���J�7�L<~@��Jk�;;/�\+�_�g��]
j����#�R:GF3� (9�RȻ����q�OxM��X	V�&��O��,L��f�)����}p:~��L���P�N�H�Ϗƶ`X0?򶣛�%�w�w���r]~�ƝAul�!u��(���]����ӓS�	��-o�"��q��^�'1�G�cW@X��T�������-�hj�������<ĳ��H.�(���L"�)�M2z��E ӫ�އ��t�i���1�=�P�	�+qĤx���2İ���C�(�0q�X�k��� �]���No����-v�Y)�+��'�x����?����U�)$:ym�`<i�5�y0�sĢaR[�p�2�i|n�[�W;Ҷ��U��)#�(��S�rOK�/5`2P;�ơ߇ ��)4z��!P!#��k�[HN����:=�p�h5S�6Dh��o��w���a��Z�=1��;�Y���j$�����L��g��,l��}uA�2N�goU��	�[Z�^�$��#�pkQ<�?����zWR��tg�rI��NS���b��iA��08}+�
�.ƈ{qI�����iz�{�/A����;���W �`]wN��ZXRkm'g�Fk$s��\Ь]i?9!� K�Ҁ��۪;�`]���tm}ă���!N��[T�Qa�x�!\�p7���c����x q�OI��y[w�x��޽|�4B���!6����m6[v���q��~��&�}6ܰ��ZO����x� _~r4�p״��:�Pd�0��7���O�ߍ�/8�Ҿ�?z��~��||��x��֫u��W�k��>���;C϶#y�S�h(���m�����7CK:��lC�O�f�q%p��t�qD��D�����@i�T-��;xG�}$�L7�B�m/톫r!ɻ:��Um��U�����������^�jY��H}^��L���a1�,����W��ҭ�*��%�$�zho۫�3��l��^���~���3�5�t�wD ��#h��p��*Ȫ*�+��J���'BG=\}���K}�Q�Tȭ���ʶ�E��� QB�ߵw�W���4m�XQ���7#`3��#x��j�Y'�:�(6�i�T/�T��»���ެu�Z�-L2�7EG����]�ftZQK n�r*���<m�ā�mG�h4ݽ�=V3�!P�Ãm�j�b��J��c���%��n3L�i�k��=�4^w����<�b�`A[rҐ�m �e��: ��>LT��<��֐|���V��6p��H\�K����M� q��%���MƂ�-o�3�8�_��KA+-;��xŢ�(�'pgjK���̊_�$o�W��`t�f"�/�� �}4�Bj<�Lu��{�9������ ��T�IԖAm��(Җ��e�e`��@�t�x�_��pu��"��n.R��;qH���p��V��0�5�Ԧ�"(��S��^�G;C[�8�K�ȟ�B���\��L\�'�P��t�^�SJH0a�8�D�XD`
j��vZܸ����-Q���3�9�\�G���bĪVk+<q���S�>�����Zc�4�s:�JJ �ۗB�4�蘒.��zP�P��0��@��OAFtN-$����C�ދ�.�,a�����U�,�Y^a���S�W���,��4?��n��2H�'�:K��= "�m�K�D�T�cZzV�z2SPʉ�kxUj1�CЂ��6^�;|��|�~�x�^X��M`��j1�_���.�c �f_�2xI�{xgh&mR�#�p��?<�/��K��5j;�/���y��z��o����������<>����q�?���1����}˻�=��&P�?1)M��_L�'Oۦ��W����@��9F2k�>@ [a{�E�0W�g���A����!��Je�~+o���[�AY�V<��D­�L7�&�����%�IC�.Ap�M�G�Qn9 �rxf��k�V%$}��4F������J�i�K�����	����3�K~�@����`��$B&�����(1s�!(j�%b4�>9#�
4�7��4DzOD}�(���p�ڒȵE���9�	9�_�����'{�mM�V�Y��ӵ�D�őTɏw�U��%��h�1�!]ᨑ�)����)'m�����h�T��G8)T�0:ͧpV�]˛o�e�1;��2$b�����D`$�$|�Q��(���k���8�^,(h�A5}5�L�e��F�?I�@'���NC��Њ(vJ�iς��pA���H�|��o��Ӯ���l1�'�<n`�.�(m��Ee�I�;���t,�r�f�I�j�	OyI�`LR�Trj���t�:�*#P�!eJ� .�n�ؾ�/"��0a����T)ੱ�]��w�1i!��"�9}n�S�R[�p���Y��2O!|��Q0���&핔���ţ9�Kю |�|���6$x7�bG�R�d/̄#v%��U�@�<��t�� .<����tN�����]$p��&m51��M^jV���0i*#uS��A`㚝,�&��.��R��� �j
��4�9��=W�Cl"ϐ��4�i*DZU�G(,g���Yx�,�������g�%�%��Q�����*�8�F�]`?zvԝ�E�;6�JM��)��+���@35��$�JJ%�� L� �<�^��>�"F�:n]d�(<�7���+	S�� 2%}�#�Q�Уi/2u�L�Ρ��}Rh/aA��&�F�t�b���"Fxu���k�O��O{׮-��N���w��-���[�hN{>��y�{㶣�k������KqS��G�9yTv�S�8)Z�.u���ө��T�c�̠���:�ʛ�oi)�D}�d�eԷm�>�*v���̆���	�H����I�� uO��Q���^�ǁ{x��r�2�#?<��w���}��b��|�hX�鏞sc��/��S�X4���/F�kl�ӎ�s�n�8��iq�]�Z��W\ۇ�y���0�1f�?���N�)c58	H��VlI���WD"��\e&���A�v���¼�ϓN�2�z�>Q(�����&�X6�Nƚ���w$���J��6|%0��S�S�DL�Q��RP�"�C��,F�j����%�w?,�K`>�N"s�b0(#�L�.�Q�� m��ȝ�!x��<+����I_B��������� �ܬ��k�O!��NHZƵn(EV�.2���# @�P���W5F�-Qd�1}��e�Y��D<�c�r�>�QN�$b˒��Hg���ip"��x�F�R��`����.���Մ� ��PW�<�L�O��`(��f|�Ь -��PB�i*X�X��`Ж�}"������a~tF�z��aEK��g�h&t��#K R���:TX�'��~����%�H[Љ��4��CkӔ�>��[5r�T�)-��m+��F�������Aja��NK�:H���Nhm�+5��^�$���A�Ep�U��j2m�]]����2j�4x���~���(��S0�����b� 6@u��j��� �&�{��ZXB�/��y��i_��[�25?�:?�ތro��"�ؚ�W�{�e���%j�l�Һ�G�Sh*ܸ�G�d�6b�l�p����d\���<��:��X�v�p��+6fG���Fkoo���Y�C���2��_`��^�.�I�j]����;?m�0qG�tv�8�Mr�^� W�h]?�L=n|G�!S��������Гu1da�ۉ]���kzү��h#��|_M�u��k��\o�j�����=fmG��=��R�`V��1�XB?�I+%���C�{�3��FZ�(]����6h�׽�?�� �G{ni�����8���=�k{׾�[��k�ϋ{?�ky޽����ᥝBW�J1��EY��S!X;KO릝3�5b҅�V�%�;t��h�հgp�`�A}v^Aӥ�GW�ߢ�ϑ�:<c� }�(Wco;;:8�6ڸ�9zʯY�50>=�wj7/�������'��/�6���}���"\۶R�|�`��}x�������oh��'�4>�iɷ�]!���p$~W�h�� Ȉ�(!�@n^	�oK�eX�h		��O"sӰ� _�N��xzwoD$������+��F���YH�6lG`<�G���Z)s���J��b�0S����[�)i81����ŝ�!{jN^)���hi|`)H�����$N��~$C,:�����;�����:M�r��˴��#��b�K���Y5�����v�����C���E	^#|ZxUd�򙪲�5i �`�G�Y�rĨ������r�������	3��4yk0?�+�MP���4 �TH����C�x.�Q�ʅ_��%#�k�oݹ�֕��$(x�u�R��G�u�E2 5%�V6��'h0u ���K�Ϋ��_�/�D[�y\̺r�z*�j	`֏4%.�W�H��C��_�>b#S��\'x��T�%�(�-e��a���@ٴ[��كP��6K8I_���)΄�b?bJ�\���'�QȨ]q�Qq:hZ�xI^��I^��]���	��k5�-;Z'���b7O���*�����C��OI�B�|��Y��b�e������#�w������O]?�6tG�@�zsA
RxP�e� xd�2X�},����b�]XPQ���i+v`ְ�j�VY�JcV"Yl=.bT�� �0�՟���	A:RHDлD0r��>��ɦ���8�$��=�Y�q�
��@��n���=͓Ǜ��Lu��SS�Ȇ�{��yv'���
�_��tH�=q�o:�SN�L�d�1�H|�I�,��Ua,`����{o��)��7L*�{����^���ЛG�Pӭw���O˫?�[<Ϝ���0n{�}����<�;.إ��y�;�-���(-���k�}N�N�&+j��!�I:""$?y�� }�.p�Qu��eRM�V����߁8�)�f���&�+˸N�O-��T;�P��fgN�;��x�ٝ�!�uU5sC�e�����L��<^m;�a�/���;�[�C)^=�ڞ*���m��R���gx0��ωc���蛔đ<т�C������rW
#�����}_�������#�� P��a��R�f��#�&��\�2�B�8l (���FQڍW�������� ���0��-��)�!"7���(�ؙF˅�����/�'%>�YnN�v S���k��!|�p���w0)g:b�T�\d�
`Tq��~��hԀ�2��c2J�;~�]äj�Bģ���+���$8j�!�r��آ��i��Id�\����=�ЈMcx=�
��D��O6�����D���3�N"���J��ޫ0{
�18���N���o���l*6�ī{���{_Ի�t͜r��S_�4#�GnaFvtN����t�vv�Q��Y~>��dX60�)�Et��4�<�F�qibGi���B�:u~�!wr�1B�t�j�\�X���%|���tS�ӎ�L�~�}q�]�J+v�����<���M�u�ܭ��.@�� \ �v"��j9r�c^V�>~���k�*�2=F��J�_��<e���^���������N�AJ�{ZaW��C`e��~r��`����@_C�����NG��K��:�C1I	:���O��<��=<�v��p��]����"B�
Ya�G�ݫo���k���C�>�k�����r�1��[�0h�)��$��؆�ߜ"�th�V�h�o>ĸy��-�S�j
Ĭ�T���@[��o}�����Y��S
^n�B�8� q�L�x��4�@�i�	ڥ&'�	���jn�-��#�
@v���wg�}��E�4�6f��O����W��yӛ����J0]�x*8ȯ/���z{����!�-N���);k�'3�ʮ,S�6Z�G�l��=�$pyJs������ЄAՙ�@���|k��G��L@�cXu�v� �?,������jX��Ñ@~�w�Q\�i�V�7�ܾii��8��7~�oW� �w�	���4�h�D�|~V��4��O���A��)>$�k�#��~��U���
�¿��e��ٳ����:��hw��Ϭ;���?�U�1��cYI��W���M��V�0�]� [�ako�̓�	�E~!���@૬�p)ķ�����_�1�����:��*\�L���<��� :v`<E�0��vꥁA�Ҵ�����p<U�0m+�F���_
�����
7N�����o:�(��?���s�4},�U2����w���zc��A����,�!����  @ IDAT(�p>[ǩgt��H�}�\&[~L\:΢l�̀ ��m(�8�=Ezکh��j�hS��Q���S�νG&�4�"SU�a|��e�4�f.Zt�C�\��oO��Q��@s��s����@�Ax
@�����ԦH������X\�Ku��Hz�����UWN��Ƀ>i�p�|�MA����H�U��5r�*��EV�d���h��a*:���t�J�E��9�y1?���%]�#W��|�����4���B�ځ����:_渜DX�Q���'$�Вn.�^����E�0/�xR���$�Y?W0����a^i�L85�m�Hj��'P#~钗08|o��i՘��ޢ�i�I�eN�D(؁�T�����,��1AZq�	>�:]��vc���vϞ>D �dˮu�U:_�е���%p@㧸�8�X���F�(H� ����Yᇮ���7#i@�������;��@�77���wO=����0q�2`5bG�J��9d�w��}ܙE�a�n^`�:"]��}	��Y����h�Cw�Gx�-<9G_'n+��[��A��q����ҙ�=|�=A�z���V2����Zc����e�"V�C�k}��ڽ��~�Սn�l MYo
�qG5��0���)<A�#�e�-.y�������{�N���������.#0j� i��&�&\��udN]�#^p"m��q��Q����E�hI��I���>���iZ�I��GIwދ/�ضY���_�G�{{��#�q6᧽�4.Y�Ż��3�|ǿ�-�m�|ǿ��o.����t����=l=�|	��.��[۸����<
�"�ڤ�]�VJ�.��o�/�����5Խ�ecs�լ�h�ϻ���Uڜ;*��w�!�j;|r�p�[~���9��hpO�k��8F�����Auq�4w�s�"�*S��ާD��~ÒQ�>$ן�1�O��I��W�B��^�тS��#R�w��ixդ^�!}��<ڽ������^��:�<� �L6�s�P��2��}�G5�B����г$��.	�p��t
�ѻ���f�{��v
����Eo�:d�A��L�����<Fp��]�=Y�ZB R��a!�� v���VGvt2NA�Aq�y���E�INǘggv�JA�ߓi��tJF)\�EʙS����c4�gG'�D�%��Fӷ���S���x/�.]�x�+s)2Y��}J'�j8m6t����'8�c��g����.����`z1�d+j�2�Ε�n�k�˚�>C���1em��⽰)lF S�`4醛��4D9�Ӱd������!)?����� 2�+0�`{%5��D�idq]�f�z�t���"��s9���Q����e�$��H�Hi��v��t���K��w��<��꒩)]�h��9A��nb�����(
_h�t]���^S�E�5�	e
y�0a`H�O�����1d���0��4��X�����W���{�4�W.j<!�z �v��CN��D�2�ߡ���W? �Mi��
<�p�%2�5��G���G��Q��S���N#b�=���C�#�i�C^��݃�|�!�m ,|@�c��*ӟq �Gxm�P�a����`�ڥC:c����[���x��N}j-������ѽx����d�ԍ8�nl�<�v�8+9�{Ys |m!���3���U��46�뀇 |���S��M�:�	p�r��T�.�d�-E;�44K*E����`���l����n9+����Cxw`H�F�T�R{��4�*�=��]����<��ڻ�P�-�¸F�j� �p�����+h�	�p��rZ�����K��Gkk^�4`�]�QT�>�w��4}���i_�X��oy��]�����ӾO{�����ڗ�ų�œ�g�A�iG�Vp]��ڠɴ۳r���W��@�n�G�ĕOZ�6X2O�3��>��T�׼������K�[�6��� m��>#/���L��WpQ��>����i�+@r�}s�"c�ay�����SH>��p�u���`�
a����*q�wۉ3<�C]������#��8I����|�������Xw𴸾�4�(vk "IB�ډ�=��Ř6	H���'�}M���/�������-C�>I��MO�\�@���Q+�>�ߙ���.�8��8��
�<����>�9�ma~� �m�$Ҿ�O����<�ga�>�a�@�9f���Ѹ��Su�N?�h��8��ʬ	zW[9�TS� �7e�&���}4W�:�c0���S�ɹ��1ƽ@ ������T3�\��h\�F�=�50+��yΐ�S
�N�
��=�d�i�+���ػS�%oma�sZF��B	�P�Οp�U	вz��{�Z׿T�?���m"4F��|��&㗔���J
u$ߒ$�F@�g3�]")��S/�K��� |.�itjg^�"s(�t�e|�Q*=j}���W9��H�W���f<�Uvr�P�VG���q+�E�z���)��M�czj��<�k���B#e��u��|5_�:DTK���yZ��E�[<dS[���Gx4~��	�� t@4�
�sL9,�.t��D�+ݓGh��?���{����o�W�ܼ㜑�5H@T$M�u���ٍ��2��Ԃ�7���N�v������4���Q�
ӏ+0��\�-g�9������w�L�.�k�S/j�d��@3�W;�ͬ��g;;�2)�E�MM� �m�y4��׺��9@/�<�=���p�_|N��mb���YQ�C�"U`������h�� 0$�9GRAK|��i�ֹ����x�M�:\�w��ZgzT!����*N��!�E���d��l5n��\(7K�M ���b�r.����6=�iH�kk�c���\�
ϣ^��{ʧ �^��>8��4e~�hu��zI��q���^����*-����qZX���}������<�ߵo���^�Ñ��XyLg�(\IM���<y&� 3m�n-x�����֓Wx<���>^��q��E��
຃�6e���y��apYmB�~�e�쓨p�����B�-���!���Π�t�1��e�&1��_�Mƾ
���۲Q�*���O�O�ѯ!����X*�IhT���eL�c�ʼ�}�����vm;��)��,]�$�RT�O���7Ja�U7u���3Ҁ���5���F2�E�ֿ������h�g�J�X�WIS���G��
�,+�.!�C�r�+�d̖����=H�wy�O�h���E���N7A�������ná�����k{w���n�)�i���Kw*t��XAM��i�����)���imz'0�wl�����?��;F�+�h���r�%:8����/��o.���i��{�c�ߩ���M����v���QKӎ�k3��ӿw����o�o/�a��F�%\1eC!<���V(�z�NJ:�յ�����M���/�U:���O2ճ�{�����~|���A�x~�qN1Im�b$�A~�X��ď�[]W�I�f�r���`q�/L��H��I[:�4�4�-�B}���Qi	�P'�ϰg��7�4��&+�<L����M�ΈzP��kh��� �]�����փ��|���$����I{;�y�]���~DxG��~ړ�4nU�/��q�#��+�>e��� f�U~��F)�W!��?�#F�t���Bɴ����#�>Z��g���WO�'��*NB�:*δ�X�-Y˔{�1�H��Y����E���xJ�8_��Շ�lX���*�T/��\�C��>M;y�L�fTJ����j��Xpd���LC����fc�h+��{�G��\C�ۂֳ�A�e*D�}���Z[\z��(�]�B�E��ɍ���`�9�H�Y|Z��|�^��[C�u�F�b���i�7W�]2�:@h��&G_K�;7ԷS>�O�Պ�1uׅ؄A�Ҷ��&i����������cD�Q��F��Y(t5�j����� }:��,���<I:�AhH����@7�e��G♎m�����/^TmA1i�n��k�_��8�3W�
/��q"V����h���w-�>�w\�1}�ܾ��x-���hq>�����{5�L�s5N�.8l��{�c<-q�~�ױ���2�˴��ȩA��]�i�
��j%�g�M.�8�o�dP��g�/� �B��T���+�A���xƒ��[�������!�^gh��=I����(!pM1Uy���>+��0z~�Uƴ�k�8��d���AL����������<��OBePI@��a2��U2
wlq �;pd�2�r%�u��a2��#~�7�����1S��U��O�ly�?���$rM�]���.)�x�,=l�k�G��@��R�������`a!]2���ǧ�a>��F]^�I�̯�e�����!����MaZ���do��L� =vL*�W�s�h��?f~�݇�؏�d�Si����(� �t�I��S��=����=~�}���|��p�[�P�Lx��_���NB{�u�
gk�}N��3�\�iKl��i(�	�oS�t(t_�|�}��_o9g��(~��Uw���ea䑥�thv�(8�c�\�cnm����۾[$9��Vd�^ P~� ����<#^7O����޾Q@=�NP%3\�S�)*T�Hģ���^���
*4���{��E�����ع��6�Ə�������|苂����^��@�4�25��	K��o��򦾀D��ɢ�%I��b�;�PzPq��mP�LĖ��V>��4M��Pb8~���������e;��7��f"�EB���V�����U���[�Ɏz�7U։F��T�b�!i��>\_���)��G���WU6̖^�!a
�|M6�g�U�>�Ʉʦ������+�L����I4ZGh�#��"�T@Y�B�A���g؎y�1�%$-����	�wd�C?G���E��aS�������;@��eZGH����^As����x	͑� V� �8��J�b��W��b}H��M|�th��-Ӧh�s
�U�g��m�S�|�A*8c���LM� D���4�XO��~���o~�M��œ�ᴢ�-05�P�s��S�0b;`�	��`���I-��$+�yH�W��֓WVLڕe��1�D��ՎJb��y�	���֥�����ٟ��׼�{An�8�G��;�z����7�ǰG8�}�~�j�vn)�>{��޷����ϲ�F��b}�ײN\�zl�3(��"N�>͖�y
�3!1c��Lg�I_�P댏���E�޼�\���3K4��LK�|�X�H2@wK���=�B7|F��@O�u m3E�a��h��Q�����i���Y!Y���%U�/����S�={���{mg�WQ8��B;�����3<�A�������i��T�mW!͕�W�H6Wd���7Z�1��i�`�<�-����Q�����"�-���<���L�F�t�Q&�i!#�Qd��8��nl������-���J1�פ=d�h}A}�����wF��_��}> �t8�yvö����d��̛����08���9%V��I����`��k��:�!��ZY�����B��sqt�5O�@eZ��L	l��B�C;����l!�E+�[�Ht���0'�.�w��+RV9;��Ԯc�iB����3���F���`L�4y���a!���$�~�ʱC��sd������`�N瘷5?vj��Z	�:���SMŊ��*�ZA^q���V�[��V������t�\�ܭ?�CM�S���!\Mo��.3	 ����(0�0%��+'ߩ����g���D��M�-�bD�J ��S' *��O� 5����	�����YZx@'|ֽ~�c�F���z�:BH��^��h�$n����]�}�F����ى6D��m:��������ѓG�/�z����L���ϻ��v��c��ZN4;f"���p8Z>S��Uf��UW���4��:Z.��0��>d�:��۹;�g�:�$v�Y�p��ֱ��>��?�¤#t�Z���Y�'���G�u�I>F[��I���o�����ʾ���gؠة��ӭ���/��M���.k{k�A�v4�Ǵ5hg� ���ũ:�8�0ykB���I�$lfps�|����x����<y=~��z��n3������`�"��*L�X��bo��բL��Y�W5~���_���ݷ���ՙ.�g����qz�Ц w.O4]@�?� ��(P���=��x��* �V��+���m��^���Ԃg�W���C���:y��Ix��u��m��l�~?}���>���.|�<�H���w���ƿm�Ҍ�ѧaX[������ȥ��a<�g��l
G܋�m�ҳ��ҕ3�!;���0��ʤr�6�mQ@ҙ���������)?��?�雞}J4�����}�hr̞�^�,i�����RW%�@&�`�j������0�3���/�Ou�c\`��-��{w�w�q��J(�Fi��r7.	HG"�ғu.���r$O)��eߦ6W��d�{&�>S���N�;u�(�"���_���K���+	�hr��MA��@@n�X
�>���FV*T2��ދ�g�a��L�h�Vp	�̎������uNU)R�b7N��Z�5�a� 4ާ0'�q9���
�l�lr��X��.Y����B@���e�j}n!���e�p�4�B�etՏ[ph?4��n(�ڭMtn7�~��9�wԨ�E���4 �O�U{荺Q�V�+Û�#XfŒ��4�:���`�o�:o(�@5W¬�xs��%�`d�A��f�"�I�)^2�iGjG�=�4�Х��+���͓^l�1�}��DnȺ�	jS� ���Z7��xo�?�r���{��)�އhM�?�3�����b�e��c!p�J?L���>�0�i�`y�`��<��]���z׉<.I��4�Lݤ��;#�VR��g���}K���PTiOa'7���C���>^�s?��N�iy��*\C?2,?MgF���
 ���I��\�wO`r*��׏ �LB�Ti�w���/w�~�{��AV$����C����#��(�]�D�`�M.#YW9�w�S$2m}b��Sj��1���8�uJ�i�kh�C�ϡ�#4c����V�4�i�g�z�V����A��ח{�f��^hp%���G�O�i<�JM�Lg�����د�0MrB�1� 6����5E� b���6^�8������o����h�h�(�i?'���4����u>��Y��������l3^�%j�h{����.ܠp�%���~<d?�Y��R�T�p/M�>B ���ݗ/��씡�a5�?�>�#�m�M���u^Ol�IGw!�eY�����R�G�c���$l�J��#V"�N�{��k�u(����P�
&BE��~�M=��d:�%Hxڎ1��?�+l�<�}V"y}������q�j�}�oR�?�O��8�����_[�[����۵��8��SQ�'��+��;<��ie�R&��U�[W?O����3ؗFv�p#�tlkR|�E�1��S�,����w���������)�1h��b��R�M��!oq��TL^�,�ob�Sh�Z�k4a�EX�������h4b�x�
��\�I^�=�Q��Ϫ�g�Z���jҦ���Q�U��#�vL����$���*i4U*!L�?��>-pz��n�äE:�aa�(
PD�
 1L	2��a&����� P�n[�e��D�ţ ���0O���J������>�*�����G�2�"'���ϭzD��%S�?��^�y�p6
_���2�� �hA��|ʰ�	���4}�#ˌr�t���pe{�p�0���۽Er���K�+!���^�T�N�S��hVM�g`�j�T�{ 
��Tbm5�h���2�Q�Y����d�zOX��5�'���2Ƽ�Ď��a�� ���H]+ R<5d�,I�e��,�v ��16��#
��g={���o�����l�)D:�`yP��A��w�ק�J:В����������ۿ<d�؃+�h���v�(���2*pf��ܥ\=A!p��f�@�4��B�>A�26�2+"�z����#:��1�X?����Pe�e�AXB��_2��,uh[է��M�����^�gW�g/�w�����w�y�}�l�#Z4%���K����3B�&? ,�- 4���B��*�#�H�M���C%��ܶ��bt���E�ii�_٧�k_B߿����?�{�+���E�E�NZ��O�0VW���q S��+]w_0��#\IƩ>0
�jg&�t�X6В�P!����s��=I�)�v�;ݟ��}�������#�թK��X7ؿ�ta�wj���h0����Nش7�\G{��o�
�bϩ�C��L�\�bx��>L����. ��V���vkj�Ԫ���6%F(8�b�O��؄��K�֗V��m��k���6�ѸP�0�l2(�/�����~I�sHZ�</+���6Z�f�Kq4�'Q��m���]�%N=J�?/8.��wI�>��G��ƶ��5���%�MK�:~����7��\����k���E�}�Sރ.1��9��y�H7�����L�����P��Ȕ~�8�.������v���/ͿiCȄ�B����C�.���'*x%�%��\4[6 [�xu:� -���>�DaN����m�iu1�"�]"��ԡx��ȳx}
�W�l;%'�:l{�<ч�s]آrC�����2EVIßm�t��Qr M���Ҕ%�~�Pvy��(�f�`f�P��'6~�-�h�f�a!rS�yh^}O-$�U�URd�F��̣�UPq���aW
@Ņظz�/X�.��&��F��P���Sx �0�e�c�WpI��r��K/��0C���	�����Bt�;�MC�S���}���#jp6`sQ0F��T�NI���sSH�t�(�ה�l�C�|�����dF�<e�Nc��7�:@=^����P~�܍�e���P��l*"�n�(�Q0R+e�)m�D�04�9C�u������2��!ґS^�e��SKG��
��
�F��AYwU\�;OR���U]Y3uX��!~yo�&^��
��ӯ�W�9*����X�֫��Ѹ	���!�?e�F=Is�'5��Fe�7z�o��@���q�y��GU�1;�>�Yg�E!X2?g��BB��s��Վ+`Ҡ�2ū{ w�����U������������sZVmȪJ(1��dQ���2���{����ў��tvz�cՉL�!�O/ah�*G[C��j�kh�is�v��-�ƻxf�-�����,�[� ������M�������C: ���6; �}X��-��w�A[����Lj_Bc��i��]Bu��?�lj��� #tp(���?D�V��W/��S��͸�\�m{���{eG��m�\AU�v��k��(;;���Q8b�ir�ۺ���t)|dO�h�b%�=�u� L�@�mo�S����d`AJ���b��5��c�=� �8@�]e�St#o�k��,'l 4�`P���޿������<���6J�!tQE���v���!��0�E���l�����g���ԼyYU�&)����!U�� X
���������%8����Q0ԣ��]�����+����w>���k�z�v������u<~�3���}{�7���G�]���%oWp��	.QKߓ���p9а� >�uJ�� %}�����DA�x��<u�3b���b˕c�A��h+j��b�3��GO0�������%t
w`�H]x5�L�0���2)XpO>i�ɯ�gG����FL��<VN)�Ps3�o�#i��-U^��4�$�� A�<��i.1y ��:�̅x_ԅӿZ�	HH=1�9�O�? :E�x6�^�q#N�ƺ\:�%���� =�<;�R�Y0Ӱ�&s[6�ZW5��R�R:�a{����hP��X��I?�|_�#Sx<)�Y(��Jɖ�����x慎Q����p��x�a�{��i:��	�lr���ʳ�:�� /�"�S����d%
���a�X�1�=/JkC��ѩv7h��~)|�0U�H��t�G&{�t��M�i(�uj �)���ьf�D��w:D�Z*�e�+��Hlj�ʷS��t%p��e�360ƼD��2C�	!DFY-�1��B��::�Z]9�"�3f���u�:��p����_"\'1�  ��f�z.���xMyč��� �h�"��}\mP4=W��ʆm�f��N����}�a{7B��_���n�� �J����rG{��nF�m�)�Q��-ׯ���*��lN�h��r�|���M�VInl����k�b�C]e�C4jW�h�Z�#�Z�Yڥ��tW0`�@iV[�I�*�{BK.O�m��5�x�'�g� %芟^#�[
^�H�-���z%0��Y��]|c�b����y�7��bK�W:H^2d��Q���;�����?�۟��%��j�vd�*tN����OMP����Z0�jɧu�*?��|�!��;>��"��&T�Kڲ��iE��r�)E@R���A���C���fe�ww��y�fj	�e�����d�zŗ��u�����uuu��y�[���fԖNڎ@�Y��_�6,�	����UR�4�S�Nכoh쐡���%��#/���!���U'�+���u_�qَ�p�����V[D`#������c�����7�k;o����]۷�����[X�;~my�����n<������A��C��$H!������L�pM���R>$�D�V8���#��	���s�f���ndt_�Y�g�����{��rH��a�][�� o$��y���L3н�{�]���?3�aG��o��Ǹ�q���m�UR V4�C�mk3��f@���c�A��HH�ȩ*�vfN��X�f��;h��l��ӎ��;:��|���G�E��fF� _�C��$p�&����V�q��c�̓Y#42�M�J���$#�+5�����#i��*;c�P��[�Ќ +Sj��vtbL����8�`f\���I�Z�/~DBK;�"�Q��r�t�-L
�ڦ),�"�M��>d��W?~�{����seyb_5��Y�	�k��g�j!�p��
_��)E��k���)S�p�BB��@���_�&A��ܩGWEEc�+�q	c?î�8�Z��:}��(��V3�t;�0�ĪV���x�q�҆b'�"�$0�F��2F�ȩY�Y�*�Eq���L��T҇�@W?����QDn}�/)w($ϩg�'O㤮D������M���S})��T�r�P�
U�2i�����!v0
W��Gh�= �鴜�+�E3�������"�iDm����C2+���d���5hwq�4��32 �f��1�[|h�M�fu�N>I'��
���Y�u9d��� ��,N��&���J�v�QXi�p.
N2M�-�5qU��h8L�d4f���](e���y��U�c+�i�l�%��0�q�#�jP��ԯ.n(�Z*2	S�2��\�'���yv�i�ĕ���x��=TG��ʯ�L�m�6��K�YɗN� ܒ�²�X�2��'��Ew�(��!�==w�Dr����䅶��c�>c�4݀�lգ�HW�k��m���BL��[���&$�Oӄ��GlKJ����W;W���P��y�G�FC��+�oҷ5Y�"Ϸ)@B3^�,�6}f�4t�+���t�b�b=f�"5��W�8@b	a�3�.R1�}�1�g���#!�������w
��o���0�+��7M��4��ޏ�m��}������ߴx&���������v�q�g�N�<,ֻ}�L���)�J+�\�ޟ��5l��9�Ѐ�z_����Tn� 5��du�%��:A�M[r0$�Ќeͬ��<u�L[q��mLT���>�&x��3�����&��qk6�GU�R���� D�H��* O��A�J� -��d�HO�d�{#�7q+>���m���u��(�L��+��6��7�\�I��`�����L�h��
"�<��l^�CbTF��S2���"��dRf�~����qG�>@F���rm�@�c��Źh�����;yG�X��~VH;Ʊf��T;�*x��x��o�G=O�j��FԮ] 0��*}#\�>lv��ǿv}��;b÷	:��i���g�e�nu��&L�U��@H؈.A�!�U#C|%����+�8��8����Q>��[�Yx�&�dG$0�I:�+6=�a����#m;�h(4�w����27�g=j�k��C��cT�f�LI��*�R�i'�((���݆d������\��c�M�]�d�����)�ʤ����[�
�%DB,�d<^���?p2jd��~skb�q��;pFB���C_���A֑�6@j�r������y(��1T|��f�::����V}9�`�}�v���<�	S�j%i�aG?��-�)��[�Z��y	�
�j�\�p���E���7؞a�������c��4$�����W�
��Pj�d�b$���җ�"$+x��0it�ЕQ˾g�95����}�V�l��άsӡ�I//��4�>�E�˗�P��hWJ��H���Vv����1���b�(��+��tVZ��2_Tg������t'��ԥ#,��@&�
r�d(W��eF��)tK����Eީ�Y����*(Fˉ��>F�
42mT��<��2y�Y�~��+Ʈ�R�lT5}������[��.��փ��k�4���C�t540�(,?�Y+�v9�4�">�����r��/��DT��]$;[`�y��eԵ���)�-��;;��%��N;��4^�/3(k-����ݫWYW���3w�Y�
�:�7��N&5��Ǜ�ml-?�hGZ��:t�K�E*?=F<������#oτ�X9�9�]�3?-���-���	.-O�3���a
9��<��iߴ4�_���,f�U�/ @뿃�Qq?%t�^
�
(����K�����h�ԓ�`���wW�~���ݗL�/1x��Kk�����m�����^y���?v����O/ :�ͯE_<ٽz�W4����U��)/w`��?G_<� V�l� ~l[���PT�`�v�-����[�RA�4��'ЦZ?��+y&�3��U[C��l�3?ZRH�M���
��xl�g��ݍNڼ�AƔog ��$�˯��Ѐ��|q�mF�����1�� >v3b���pec�`0nnD�LEfSs�6%X� 8Ҡ�$(x)�iSLԎC$4�@,�v*.��w�}�͊���'~���:�fF�
����y�{��Z���9�^[����M��چ(�im� �i�0՜h'N��$s�Z�$E����c:��g�U���V;/=ٟ2�D?M�2�YT�׮B$]�kJ�$��e����zҎ��!{�����,��N�|3�j�ڑ"�����c�%LOphǯ�	�ө
#e�!�9���YL;�<RV��~�J��8y�����S`�s�B��i<B�($�]�UXK�:g��0�vj��K�:�o�J��IJ|�]�3��*�Ԉ�A�,�����-͆�-��$�"�j��R�a�v
�;�<�<G��K�`�x�,U��-� %�h��3p��$�\[�2��.�|�%�xo%�N� $��+���Z@=������s�Gx07ywU��}7]�&���u2.aXB�����/��FB�w��:�f���]�.Nq�{];B���~i@T�I0��)��u>�AK"La�ѥS(%n�����Qgi�i+ЦXu���p�ʎp�*��A���U���G7'�N�k�z��
6N�h�B���IY��e4��ؚG�ҕ��9�):�hͩ��U:���J� /�sL1��L�it<��`�_8��]�gA����U@"�f�v�;���p ���A��Zn�X�!I �>��4��b��
����-�%q�����	+|]�Wq@����
xv���]���{�іI�I�*�n��X�=�DbH��5m�Nཟ�^�g[\�MPj���o�����������)�]�8�������QG�.��Q�u�"�Z��d��vƷM�(�Zz%�YzЌ%Z0f�Tt��s����2�'��:�U���g��g�Md�=O_~�4+�q���g�c�G*p!�Gڞ}�<�ٺ_�E�+�q&��M����۷�����3��!+�5�e�	Y�풅8���?���?�^S����7r,j'�@��rq��E��N~��:�M���ƶ���o��S����S"Y!���N)��2��2I� Ty"�"�Жea(��������_�7�!6�E��@�r�6�N@��#�E*R5��~� O�u%]��301�@�"�,��!�GKg�v��%�H�d�_��Ʋo�mu����!��}��n
�Z\j�n&�i@��!�,~�40V���h�a딬�=��:�9B;�JP3��*��լ1sF���r���U:H��0R��/�܎��)�]G�t�j��őo��$W���,Ԓ�3�Q��.�j��&Q�V��� ;(�������b��ܤ�%�

����i�Es�sz�*�ecr肤��4�s%H"V��t������7�ߕ�|�w��mU"s�Ѡ�������F���*G�Z6T�l��a�3h3��s��<#��_���t@Yތ����.Р\8��}# 2)W�����SvB���|51(��iArB\� �e�� C߀���h@(Z�	�4�T�Zh�W��ug*��j u��t�Ǥ3Y���v�K�hx���L�����I�0�#��m�eꙶ�M���憫�بW�	�ntu�������.'���h�1���&m?Z��`����C@�m�iA�Sah����圞rJ���OC`�m�f��w.�|��2U \�.A�)W4QԯU�>lE���r����-Fꫦ���� O���|��u�7�^fʵt ��m*�(�|�=�������T(tE��h)�d�� X�ỳҶ��$h[am��9��T@��N�����&ֲx�T;v�Q�^�ÓV���,Q���M;E|�4��A��98���e`��L�غQ�4C���C���߳Zt��&��x
CSj�J��[;9��aX^y��ȳq$��;�۽�zO��q�\�ޮ&�}W�����������~.�������C����]��Ĩ'�X�։��W����P���}��_]azQ[*h��$�oT&P{��]��5g^�=0o6�-�D��D�U�sU���v�*Xt3@ [aaї8F��k�(��Sg��Tc���ݻ����kv�xL_ACD�qWy�3�A%�~3��D�+�fym�%P^x���]`��|8}�ǧ�E�$����q��4k%�(��24�ʚ�;��\m1%�_�W��T�ͧ�P��8������B7e�c��Dd����d����@��֫�a��{y��#����a!�me+��d�,��_�#�PᎾ��S�8*�Z����pI5y�S�Z���6:!�F�=܇������߽����m�~��%���`�c7���)�i�1�'���a.�ŕ$sd$��)<��"�H�����{|Y�U$`#Q]����;A�z�4Wl,l82+�/���U�!�|U�z�f���yة�C˭�c�%37��.@�rT�LC�Ɛ��>]� ^h��q3����9ժ�+!5W��ڸ��[���ا4:��u��Z�O`4a��9DTq�JP�K���z0����Wz��С&Ɲ 9b�V���VJ�`��D|������g+�&S��v1�mr�tf-'�7�DF��1�,ª�vC�B!�4�����!N/7��f��¤Z��? �h�C�|�m�;2#���X��7CEoDڄq�Grj!n�+B�	�=��lqi�\�+��v�&���bI���t{C��P ��6\N�` ?ƥ ��Ro�2�3� \�66��Z]�_�ڙ�#���+�u]���|o�h_UZ�zs  @ IDAT%!��R�
`�XS���c�C'���	����9i�‸���SsS��,܇�%:gJ��/(S8��oϻd��h��Q�:����#��O�+a96�ң�&��1k�XUx�7��bl2-���4g]H;һ�w1'P+���4jJ��T��x�?BP4L�yq(4Y��)xB��(�%4�+���UM��2>g+��jI��0;+���� ��=:�w�c\��w*�m�n����`G�M߹*�Z_�Y�ǒ��[��ۜ[t�,^�h뀣:5��Ҧ���Yz��;0�W@�B�q�����5i���Uk׻�k�����c���v��������x:����dM=9T���w��v����C�SW��
)�L��C2Og�p����b�3n��v_�������B�p�i��s������9���"|qj������Wd0 n����fY$���:��]���{�ж]��^�F��������4T�HQ�����J����他K�4���M�������Ն�>�q�c	u$K�{���!1` .���^3 �`����?�rim��rt��d �2|�IRB����I��5f��2���!���x,tr��-�S��:n�!�٨zQ i�F|���n2�m)\}!"�q��'!6H4�J~"DCl����<�#����	�1���?�����	S2LNh�s�d�IS�	"�>�\��H\D��"�k�AG�vAﾪb��Iy�#

����YE#�՞T�MG��;H�t2�nګ��#�L���|��F�����0�����)��0m�Ǹp�m%iQV�ذ�Y夶";P�z����{�������fcwm�y4 1����G#]ImM���E�G����3
�ddM���_��Z��亂� �����*ՊH
�������#�%����W5&i�NH-��
��#y��^���:�]�k��^�W�0���#��ى0E�h7gY}'��	9ʜ���`B����+ݩ�p4xJ+K�Am~ˈ��Ey�F����Ǌ�N��d�w� p ���h�ċ'B���QS��iR<�����\��V����`c�ȅyҐFy2]H{B0΍�+j���W[BuzaQ<0���ˈ5�)��v!�`ii_S�_�����C�|���]A'�µH�u�z=\�Nqn|���s�]�\Zu�B^�RP^hO��I>�fz�Ln���&NU�i������t�XI��ց�$S�L���~�v�{�O�7����D/�
��,2�P[���2�����g��t:�����Ll`�5:�.\�5��C�o��7��U3vt�αi��i��r�G�ήX���4'�$��/����<{�m�ꂂڽ����\q6��@!!_m��|L��}Nk6<w+�£������8(ap4_�|�?�ԡ�o.���L12�!�y6�s*I�
�G��Ȍ �J۶&)�!d�`��t���C�gN"�+Ҧ�����Ȱz&��=�ǽ����[�c��;~�]oi��[x���������g�o��3i�si�o[�D��>خAl�`�GJ� Zē<��E�05ȘbP?j8��'\��<��j���.��i���}���/_d����u4c�� 0�MCH�g�?�\�2�f}_����^�/+���~t����>������;?d���l\P������q��=�ٽx��>�klܽ�\*�S���(�i��ҏ;Wj��k�!�
c���p�̵�e=X�4'�G]�߼�'���������~�>*���%\�v����]�.eVε�=�a��n�;6�1�rs�|Pp��O�(j�`A IG*D^zi+�6�w|Y����������.�ڈ��bR �n����H���{�d~lx5�[m5p"I�������.�u߽z��G�{���ѭ���b��U]\��S�nM��i�a~
VJ��ޏ��{>��0:F���a���d(��jW:1�TF4���Ǐ��v^�c�>#�%��	+/����4B$6F$ _������,6;
�2�h4e)�&qG98��a��Sr�`1K�
K����WV�)�Y��x�:���ش��S !
_6R�� �o{� ]���+�>�G�%��Z����]\( 8, �-;��4��=�پ%B��)i�pC�=7`�F������hK��|������/yvT�V-�0D{I����M2��!(��6����Y�^gd�!��\ӱ�)�@?�E��`��@�\]e�6�N/�O:�n�u��Q�X��r�$��>�\u�h��ݗ�:�tD�� ��M�+���(���1e�(��C���Nܩi�7i�f��F�/Gׇ|w�f'�'ZX5?��n
2iAo�'�K�e�_)@Ux+���W�O&���i��r���EG�Gt�`���4x�k'>����f����!e�����%`sCia��kۜ�f��B��Vs���5�#�g�Hj�t�<˩������%��BRH9�� ����Fl�)h�:��&8�����fzN��o�
\Li�i����I�zbҕ�5��E	�f��'Y$'L�:�������r��9��ߜ�g���Q�;[�"?�{۶�^f�c����Ή��A>]�U�����OOy	 ʫ�ލ����~< V����?���r��I
l�(\8ēa�j�uS_��nH�g��9�}Ks�����O�!��7׺�c��|SNi�,���-�h�ƨv�>�6f^���`�?��0����J��cr���RS�	 t`U'_h����U��Z�,"�y�v��P���	�?��X���p(�O�)rQ�	B�%��|x�C��V5-RPre���a	X�_r� ���$�K8+�TVM���mP�)��+��S�V-�mB�[�~k���7�NhK�ch>�헶w�X��齝���c{�F�Z�
�㩗s�:��입VF�ը�[;�].h���}��z�+�{���H� f�_M8������2��k�MG���j��̄�,c�q�q���G�p^���?���ﺉt�V�����-#�I�gؔz�_SLG�od�Y
.RG	av(�Ua	�\����QWQ���+xA��E���mm�$}�d􎟕yV�h�~�v��7o���`��ۘ��_)[&�شIrS]����qUA������6ސ�P�[i�������D7��t�J��
�W!����5�ڒi�딉��l�*�(O6XV��j��,��<�V��J\*`H�9*�NȖwb�?*�'̋H����QxO�����S�����Z��]��D~����!�[�V|�y��}w��%��Eo2�u��j`��[�"DC0���o�C�vz�>W���������AUa��]�?|���8&�f<j�ՆJ����Y�x7�xZ��0�V?�^xW�/��V܈s�]F3M	���#B��3jj�T��o��wo߽�vp�
\�ha�<|�*�M�7V�h�$�O�O++���uV�:R>`Z� ��F{��?N��C^|�E��&x�h_��K{��������~��2-#|9e
�15���ļ`���mA��ضL�!���![����O~�q˕���L�(��U����HrttWsD���ɪiڛ�i�s;m������F(�����G8>����
�P9��K�pV)�Ӿ�l��;�UR�2p��Z�I����!'�;>���P$X�-�,��5�p�b��q����Im���=�,0<�C��Rl
YP��S��*DyH;�-P(����YWi/P��#;hy��xH��/���0n"$b:�|�����h}�/�n�o$���g6Ó��+h�۾$~{���u��4���� �i<�}��~����3?_��I����|��� AAܲ^�I�vX�uDcı*�xJw�dZ�j�,�ڥa�c*�zkk+���㇇ъ=ʀ��oF{E[*wLj��[�jj�t"�Q#��Է����M��>8#�w
m+��M�{l�>tkL�?�p�m<ъ�V�>WcW�}1@p�*z�$Oʭ!?pV���)Wz�x_qD}�l�Ү��e!�A���4p��RFޫVӞ���� +��JJ���=M��K�/�ΰ���ŋ�B�͗Z�	:�l�bE���a*��W�[$���\,����!�9(� [9��é��H��W�!+����$~��e̦�Ujz��p�LO`\�G�� r���[�L�a��0^��za�R��nu��}9�(#v����z���h���u��6!D%H�NQa�� ��="%K��#>�0�r�omeT[���L�����r瘮���E��������䣡�,�&��Z�iG8@nj�޼����Q�`@�@0��)��R�U
Vͦ�� ��+�f:C|�k��ik�f�d
�/k��t�=�\/�Vl��	��E%�)��W��Vy����"4�R~W *�E}Ng31��(p���\�F�V�3F�$W�	$�%u3"��@�V2e�Q;L���Dǹ��2YQl�fhL��IM�ً��w���7h>@$m³��$[v
v ➼��W�V��L'K@�!����a�*��l�DbL��fhYhvi�q�h0X8�|����2�+��F����q�j���0MRߙ�i���S�{h�N�rt���°�S�~����E!!�[�+�bYsN�7�]R������4���8=�
�|�|l����v��	��܉ee��y�Р�厮3�]�%L�� J~2�)ԫv|
��Rf�jGm�L����\���g���t��q��Q�8A���ʌ���ll�u��	vq�J�)CO3y��VAۊ��.�CL;f)�2k�!�4�3�r1kz.D��]�,�di�)_�
���6�N.�pu�#,��#���lb5���ږ7�g�L<��~#  =�gc��E��IBoKI�ߘ�4���ʙ4�8u�W<KG��4�M�Pt�?������k4�k�wx���4̫OP��58�cw�m׍$�����G��HM������v������*5�RJM$%R�g����RY��������"�  xdZ|m��n�Q��ﱘ��.�E}Y{�V�O�� �����,�::�$݋�w����$DL�26����'wf��t������N�YAo�4AƳJ�!��`m�~��B9
��0����n��I�c��d�h�a*?Ⱥ��}T��Wx������j��' ��(M4aV��m#h�=��_�W������/��0�,����J�nW��o}�|�q2%�E��y�<'oT�����|�����or~;��O�Ѿ�Ǵ7@A�f��(����K"� J�� ��"�=,��k���[�e��0��i��fR��c�UvZ���꿒s�Nf���$�����s�U8v�v���V�<̹�i~/bԯ;ne|R���3��5&}ӎ��9+
Ӡ�Q��+�5
`@�l�=�6���l'Ql���VJ�N!�#���4L�f�߈�1FVL�����]r�J 5��u�F�|ql���{���ϥ0~^�;�]���#c�����(a��!��5���xY�^�`=�S�L�J�=�f�1�"��/$8��YZ>x5a�Cp�6F��ځ�p.k���rVs���a���"8)(��lo#Ĺ�r���Z߄
Z0]DG=S9��)��������Y"��=OQ�&�h}%��^-F�x�@~�<fΎ*{-�@�]=���1BVQ6��oR
���I��YI���������ײ|�Za���|U���V�=ɡ���"�L�Sl)���h��3�˲g��l�Lp�����$[�ѝ0Y8f^�(�[���bG1�:m�[���X�;�Z2+��X�k����|Y�i�m�p4��bh���}�X�,��Ot���ެd�M/^�S�ދ� �|U�q��V�kgx1n�Z�U��͛,5/S�m��v��(�T/ڿ�py���/
&n5��_�1�b�@R��[�'��)�Y\Q;A��d8v�&�TN=q��kSu�m�����g�}dj������m��?�@2y�?ܻg�s4�2�%a.}l)���<��Y��Se���L��ϳ�ܾ��!VN�h�uO[<9Z���J��G0����dxx*7� >E���d``�5R�}��:�%�M�L��|����3~����IQ�uʞ6�SQN��f�8J�����3�V��O/�^��n��	Щ[�=S�q�M�t��{�R%�?��^эҁG�E���x�(f�+����6Ͻ��w���hb�jE�V`c��棘�[�)Ń�e0�Q���i����BY����M}��G�P�|��ʠz�����$Sm[��r�I��X�	��S����S�~��Rm��fx�B�E���g6	.Q�]�r�D��L{W�1FDk�!�������oR����Sե�kX�w<kk�	`p	�?K�������~������lq��F����Zy��Lh��,�um�'b(x��]VHuG'��p�W���	L�B�2aF{�T��8�V�L&���H	�8���[�4��hI%'^_{Šhi�F\�{��0��L��]��ʥ��ӈ�ٔ��� !w��G9�˒�n�%#��4��鄳�F�*}��MVG�q�L1q6Z<�z��ʥL�U�i؞�{c��t(�/�{����jg@�kh�H-6���M��7cZѹyv?�h�tJ�Qw�N���Y	j
����������zԙ���A�:W�i�[��s�.�'�-�7���V;7��'���>�F�p)��⇫-�g50%2�d�xT����:!-��Ǽ N�q���ɽ���U#����k)-�>8\�ߨ�,�J�n	��آ������y&x�Z	�y�݊9N�:;�z��U#�����Z�}&�vS<�z��`!�Y}�u�b��g�l���-�x��e�O+!���V��|��p�*��K>a�艂�#���<�W
МW8u�w�`�s��M��"��|�c�������P1p�����$H��S�.Ep��>��tac�
��İ���e1e��1�^?�s;K,�ש��f�����B��V݆;�m.8	�}l�;g�,�y��󍂵��mP��+l�B�`u����˔�y8`1��e܂��dM?�������d"P�'wV2󓊶���W[�p�r��@�dRQ�����Z�Q:�m����ܙi�(`�pS�f�j��ʧ�c�	�h�v�L��)H��R^ؐ���m�l!R�������ژհ2�杛���,��4�V���+�mҼ|u�� ����|��j?���Rp�L��ږO��߲�R���G�������Sߥ���X���۝0�6<�]/�~8������xG���A#�[0���j���~UF��V%��\��׀\2c)`���u���{j�2E�H'�Q�.�,`"�=�O�aW����)�k��B{胶�R5pM�J��)�������!���-2���|i���G��h�[�E�l��>��{������Q=�o�OṬ��|B�d��:�A�ZA6��ԯ��];�FPk�����*<?�x�2��3�E�qiC���<C�{�>��/�%(lW���q��!��Ooo�O�����4Ztm@��Y��{[6���6���I����6R}ԴރǦM2�Ձg)u�La�� ��梒�	ٵ+`����F�O'Z�}��*�ʮ����":��v$k�Μ5Ƶ��X�>1�VW9��tU~k�˜�UD��J�b�:����"�:��������zN��JYm�����W�>������^\
����C��%�Y������q��R������;wm,<��sr���~���Y�Jͧ�I
�N�۹y߼u�y��Y��)��~�䛏
� Ng��1\h���ZnXu�/������~�H[Ey�N�<���|Y�]k���x�у�o�����tW���]�Ͼ��p��OZYu!�|��ݙ\�2�}���!,@��w�ՙ�X#�F1�L�-%e?i*�^D��k[����W4��D7;M�!�	.�E�Ír�3�b�FXt)�YJ��,cW�K0}w��g��D;NK�%��#�0�s��7-�O�0ܞ����ę6�0�Q�����7��*C�b ���̧���{� �[x~{i�0)X��Q&����l����w�[��ܓ�Dm��`΃1�#��^϶����X&(�Ng��qNMa{Qβ��!g�v5e=>j
�a�S��C�gs����G7:�1��C�� &Y��F���8j�rb'��?���}�<l�a�+�N���?�v�Ŵ&��(T����!���=���0�Sۥ@��n���on��匁S��	DD��?~��w�n�9���<ܾ�s�ڴ|��D�a��h���d:ի\����2�e'��A�b��ӦhX�m�j|u|���ـ��xu������^��S�kW~����M�?�EQJ��'|���0�%EW�o����.��τ�x�4}���g�&m�i��N�;�:�{�Z��b�q�#�G�]#��l�u���Ѝ���/2]��X�ɹ6~>JV0�>�Eʋ�R^g;��W7�ǒO�DiG����~W�/�\�:-+�
�/�Ǵ��L�Œ�S�dR�`C��,��>������`8-���W�2�G������ߕ:��|� q���V"����p�i�_{?|)|P.XΟFg��k�rSrZ�h��J0�r*�>�|���f�d�p�W�z~����{N�Q OG'�zCi����~�a~~���^;���h+���[��X���6D�[���U<|�:Ր.ֱ`\L`�|i
��u��l�ٞ#���P������N1�@g5z�4á���:i�5i bJF[K�EDc��NH~�h�x1��3f���N��8x���4L?K��zW�G�myҬ)�E՚�hY�X�?O##OL�m��+�j
��2N�����x��:`Z�\S�!���[sM����d��>��J�1q���>��p�J+6�:J�7��]S�b��U������d�N�3���0gEg�Q�*cj:炙)B)?W#���+�ڻ�������/�l�؍q��(�FN,��Z��gdY���Y*ߝ��Bӆ|Vi��Y����6�������O?�Ҏ@)K1�Y�[Oe�{|���1j��>��5��7�7n~�u����==���03�	�'�j'8>�� �p��^������A�f10-��{2�:}Ã-BN��oZg��cpx����3J�9��}��aamc2�;��x��٬�D/k���Qt5S�e��z.�w�F3	���$�d��Dӑ�QYς�N�T?���tuu��<����~�o��D���3��=����l��$���o��[��o}\�(e��WSً@��5��G) ΅��?���mJ��.�B��e){4�y��1.�0۞̦H���d�&�P�˜�?���M��:�����]l��Na��t�m6�~��|M��0�8F���8��3����[�/
O귦����P�����t�����:�1(�Xo\��EK���E���ahY]����᫿v\K>-�}ޅ3��N�Կ.�$`�߳�T����_��р�<�x��4��i
qS7�w<̽����X�ǂ�ϛ�
��.�(k�SX��e���;���m#���,i/��j|�m�s��9�#��/�C�-� G�AË�F�<�0�
B���)�
mU*kj���i�!�Bahy^��ޣ��4Jӳ�O��X��oԻmyQ j��Q(`���!
$�fs���>��K!����t�n���yʘ�6[�ӓ��z 8�_	vJ���Sذ�)�>�]�i�r�i�d5�d_̑�▏��$��utrf�_���Ԭ�}�̻�2��O9.5}���>�u�p�ƍYUL��7���	9��yF�'�^�Eb$��=y1����A
�GA���8�%[�R!��_��y�	K�wi��q]��,�)8\�H�?�J���3:�w����������GVk 0U�R�ƨ�agxs������ �ǟ��/���E���[���ʚ�@(=��͞1:M:�
�ϟ�I�0�& ��p�p��Q#���u3u-D�<!?�n��+0k����
ѹ����WcO�T*�� R��6����@�!{�nȝ�M��p�.���м� �Wȑf��ꌔ:��hc_��Ѧa�Bd�2B�p���U��z�ӝ[1��9��i��'9s����g��Ǜ	�<��ȡF�I�f�W���ԋY}�v�|ɳY��1��u1�s��EQ�pd�o9���8\�b0Lt�\��c>�]v��Չ��N4���T֡W���V��_����Sq+)rO)-u�1�������#���YS4'�ҶYߌ��Ͻ�����ph���ɧ�G��;Zxopլ�����F��Q�kC��	���c����������/�����*fП����D�M1��092�xF���D4�4��㘇O�bC�p�BA���(��-�hےs����)�'�`V��1�W?��%Y���<���!�,�GY�ޥhP$=i�������ՏR�v��ʻ?W��������#�$k� ��&� 5�~mS�ڤdpG�j�!A��^SGՍ?歍(�|�8�^,ޭ�?j�����wa�k1��EB�h��������ϳ��)K�)�g���J�v�k�Z��#^�+��7�F֖כ>��A� �NT�ҕ��P��A'�X�{n���w�B��{m?�Kmz�������p���/X��#��T_�h#��S��0s{���ٿ��2
8�լ��?��Ӵ�Ub,�`셕��bP�͂��D^�Oݦڜ�A��dy�*]>t$+����r}�l<N������W?���ng������&vg���)gx<���a:�i����ÍkW���/e
X��Z���o��O�������&ZK���,z�e�_�ՠ��,nf���H�.?0�����{���|�Km���'r�
]�%:�3}�<�՚cş���7M��7瑆 >vE�|��r��'�L�B�/b�p��$��
@
8�4+��-B��?�0M����0��,C]`\�
�������O��_he��y>�N~1<������W�Ň�᫔�{�\!X˰ꬾC����l�a>IOs%���N��|<I;ʳ��)��v��Ǉ��_������3�^�5�+_���iۢ8k�x���/N�1CҠ'�����|Ƈ��E9�w��ժ|>h�$�k[���?�*q��gz�𚠋\����t�����~y�9V�+t�=��n�f��e M��?m+���=#��rt`�B^�I���6Ɵ?�v]x�N0�T,�jS��Ջ���lE��(d���6b_�Q�M���b�e6,�E���V� ���=����|��~>1����Fp{r��0> ��̷ʷ7Cl=�V�i�:��J�P<�:'�)`}(e�S1i������r^�� ��N���ߡ�x�ۙVH�����0Fs1�r���cF�[�ȩ2�E�/:>&��G�܌�R&i�6���0�!`R������ّ<�Ϫb��#�ߍ�[,3T��?=|���Ͽ|}�9߯�9'9��pq�a3-W�pFXY(��	E|oL��cb�6�ub Fs*nl�dN�m;֯�p�=���~�˭�p����>�+'�!eZ�(!�a�	f+MY�XX�^�����s���g='S�l�'���}��{1�a��+�Nw�����v�=�,@8�5�t#(Ϸ)���z��i�SB�0�x�O8�H�mx�$��? D����KXv�����y��Un�/�>��:���5������)�/�q��i)5s�W���$\YJM����Șb�~Ts9%�Ƶ����A� �6&hF��~A8��yJ9�u>J�X��V��N1�*��8lm��<���1k'C���]�{?E� �O�[��ht���$�����K1��-¡��������xG)_��b�>1d���O���������/9��/_��p����S��l�ܑ;V~Y�9x�&|�`Ã ױG�63е1�cb(`�:��qm�F�Ó���FW���W�g�wOS��o�d�.��	�o�Y�}ӂ}}�`~��K�ͦ��C�������SJ9�g�?��e�oˍh�T�ݔW£����bf�#�1<�����c5X�o�F{�}&��-L�~�ig�O*�D��M���Ƀbh���)�_j�WݗrT;nx��|��W\b�{���8S���bԯ䏗�ì�X��x ��a�n
�^8�1���	)�>��jp�%�:R�o4���c���k�F�Yg�*�@S��U;��u�z� �����������S������9GinZ7Q�y�`���7sRk}�������O_�Y����>o�� ]M���^��t��ٚ��+� ��/�<𗯿O&��I�Ϧ�����1ᴺ,c�^X����ʧ_��n����mq&�߮����j��~�V���}�y�G������)m����I��e6�[���x!��9g$�{5�5�jisK�_��E��<FFH��Uo����1;H}كiAH ?aD9Xs��&ҙ��:���k�/�Iߧ��@[�b��'�Ja@6��w:X�	D=���[
�=E���L;&g�t�N�:#�P<�r`)ܟ��\V=�V�K)���7+�bB��+{Z����z����v�v`q�����ӏ�����ѵ�ex���2�1"�P�<���O��WSt'�o}�؊�ۍ@����/����x���s1%�ϙ^���0B���W��\]Q�~���,^_��Xg�&jds���t�v�O�H{w�����X<�/�����p4Uu%%�b�c��U^-W�f�>��k��a~�q�=��ocVE")�(�L	ӫ97�43fU��d��x+�^G�F�i�#|�g5`�z�h�b�;��SDMYU�_RFg��4>���z+o�s�����?�.�n#�p��������:i){O«�g-�f��.\?>ugRН��$�ܓV�=zf*��E������COm�Mh��{��_h���]BeY����~8s @鿟I��w'��6��q�#l�hϟ��=K��
Ǆ�Cn��[�%����N_�OU�r�5���=����~n����1�_�=<܉��5�O_�M���s������A�|�s��]�\þ�MR��6�У�R���鬫/ko�����
,�G�;?VJ΃��8V�Qi4���p«sg~���]:�ۢ�Y�����ܾ��(�7۩�Y���մ���~�,�BJ?�՝���w�e�b10�zY���~�G_� �y��7
�|f����sy'>˽�־���Ý�i�d�r~)�U}�<M1N)�� _Y�!,�uX��j�T���M�0�Zq]1)���D����� <�J���������,��_V�ZY��_����̾q���,�>ScL��&���˿��o�=����������}�ot�&pO�)����V�	O�.3�7p��蜢:
`��Ū�n��e����-6\�?=�8x�V��hj|m�Tfðȯ8p�]����O>9���������|��k��R�k��|l��.������!�4���3�K{�-u7Xz�%���(a�k0@�?M�:Y[��?k���o�
����XT�BJ_�՞b��gk#�\���}����e'�4xӿw�J
5�e:KH�S�1�OY�b�T���Rl{����/�
��oW���ma�Q7��k�b�m:oe��D3�v�0	J�B���c�\�8�G�%j� ��� ���T�Ç�^g�⯋k�)�p�,�ʛ:Izw
�Z�3֯����Q9�& hlSYd}��KQ[q�~ o7m�z���k>"[x/f`4xg�1��)B"x��<G��	B�`��,R�Y����KЗ���Hb{�f[��;̯bC�Q��=��։��M/$���z�&G��4�u9�s����o��"�����͙��F�ά|�2�'��Y��a�0�T����7���hW�a_J���qN⚿���H_�W�=�;S?d���;�X�7-�ȷ�T�p2��t��w}�6~��v[��3��b���'�������+M!aF✋A2m��<X@����0��
�f�,b@�))6N��m�ʱs,\:zS�4�Y42�m�}���Z�'�_���#�Nm�s��������, �`�Z>�呂�	!N��8�O���>�asA47��]�P���,k�N��":���q�M;�J��Mۤ���$���X�9��Bʆ�`�j�i���Y}#&����<��=�}�(3kH�&���Ӎ�k����i)R���ӥ�4w�3��i'���T��F`�r����BD�<Sg���Mo=�|��vg	���y��]Vڙ֢�5�2��&��6�^Q:g������-��zОd��z<�G�?���� ����N���V���w��RR9�'��)�2rV$?&Њ�c%|R9� PY/����S����E�=q��r�L=N1�����ˢ"ֳW�FU�~�S0��:�����KW�)���jԿ���l�a�+��fV�����9��ʰ����q����m<�J����Qm<֮���5B0XXb(Fc�	fp��_6�<��vDJ��ŋ�}hL�Z�x>��������|zk�1]eŝ��'h�g@!�G5x�Й��;�o94o)�)A���%��$�k!k��j\4���3�Q!��R����7�C� `gB,qJ;�*����L�V�����^��s�OS�����~�Q�R.� �B�u�c�fF��޸q���^�s/x�zQF��Tw�md�fU7��	A�f"p��*|����m*ݨl���q�Z>O��c�3&�U��9��`��E}���.hz)��ύIx_��o�Qc���j�-�ޯ8b�D��&�-/��7w޹ߕ"���~�y9y�n��i��{�r<�E{�س��:��-
�b���zV!&�EG�Y�fJ.�왹��fa�:f�y�Y˽�:M �g�� >u*��}�t-�����0�U�����J�o} ���4Ԫ�BG�UL�N�X�zo�@�FM�͘�u�IJ��|:���2k����C��v����v�� ��p�5��u�~�>�z�*9��E{�<m�ȗ��̈��F�7?� ��M[�°0����yk`�g�M��2S�cv���í3M{%��(1�}�Χ����N�2�)!s�Q�28V�n8C5ZRyfv��ʹ��Yپ��Ct��K9�=݊�L�5�t����QY>q�r�m>�8�o_��W>|��&r)�Ͼ8\��Q�E��eǵ�^
�(�!x,<am:|�o݁�������6��"ڤ�D�kX�OD;�YB7Z�rBa.b-��׷	��)?'��]
����I̞q����t~�)���r ��'Y�*�mx��w�}����R�l�0A���I�E�g���fӷ(��|��3ϩr[�;FU%j/B������K�ӈ���Ch�M���١Y��/��R�	����p��).�ףǭ(M� ��Yw�������j���;����o��6,�de�g���M�����M?6uc7�J����~�7&̟K�_�P�!�2^j9����C��Y�B`Cէ=��j �se�og~V7J1�>������ F��?�B�"�d�֦����y�t�ijKFΤ8���� �P�]+ �A�&�����>kP0֫�g��/�4M�<xǗ���"�Ņ /[���4�٨ror5��O���UK�&�WSoR��;:�Ό��s@kY|�����;M��������j� �n4jݐ1SUw�f9�����X�A9S��D�ƪ!�sH��F� ��2���M��
�p���g���QJ���ơe+����Ž�k���t[�|����Y4@�,8�*�k��\
��:���?^�f�²�7���(��c���6�����س�K��	���i�چr[���z�_m���Y�z��ׇ멵%^�����c%}t�G���C�6<Mc�`0�3�	�,�`Y%7�;��׼Ii�-��X�ӹp��N*aY��x��U���6��o�Z��<���a3PS�)T�u��\4/^��y~��/9�5Fl�  @ IDAT�C�.�[��}�`R&�̆����آ!�y)����b�S,T;��Yσo�𿽘��e7�}y��V�__Z�;�[�����MHpDtH��8�o9�|&q�>�ő�6S�y����כ2^H Z0�>�R�q��:�G!+<�=¨���h�,AJ�t*���q!ݮ���P�Z���1D+[��Z����L�޷Zx?
X#d
ؘ�G��*3��@_�N6�BY}�{���,��{ܥ����$Tl�h��^4_[H�{� g�?'�;(�����?��I
��f�b��a�Ѧ���<��`�c�.%�ݾ�w�xV	�t�W\��,F�*K��'7�̼_8��1��}�b�c&�*)K�g�#�|F��ھOwv�w|�XGO&�4���/j��,h�q1g/\Iٺ9�RY?s�����Q������qD)�+��f�6w8��5G���
����E�$xZ��~G��m)t�DM�ݵ�6g�٧k���y�3��Q��(�u��U�T�ڙ�9��|���	�-ſN	��;c)bY;�5�ʵ�����	
�x�Z1'J�-P��"��"�"6����Eco����� B=��]_�1��(�;{��%D^;�y���ՏS&��`_DGϟ���R��!�c�ڂ�-7��B���G3�����_w��M�_S��S����Y=N�sH��:c�+����B�Ť�������~5��SjY�Lѿ	>#t���J���@����r�g���ń"�+�_h{��L�8�҂����g�m֣�c�� ^��c�k��
c��W�qdG�F[o�wp���ƚL��j�����6R.)��8t�Y��d��,+�9��b����Vwa�1�J������>�j��_@��p~����A�������(����;�̀�J`��X�(2ng��pp
�W��mm�iS�A�_V{¼�>�ˆsr�+�)�K sȯ��g��25�Q>.�omc#X�5g��z
t2�ϔD��e2۽0<L��/]��Wc�S6��J�����N+E��o9��L�aPGAVVO�%a���QȢ5u[�kla�((��'Yk��9�'|����(qɄ��ף{S�|��{Y�l�LY���b����J���J?��h*k��Iu�$�N��).U�@���A�s7�:fc����f��gCo����~�͵h���c�/~H>N&,����&��)�ڇ�S�.�����.lfK����и?�����$^y��5�x^M?��bl׏��<�{ģ�&VT�
�-�VDU
dڰ?{�O�
�14ak�y)�T�"�b�tӎgS��w؄�|#̖e`L ��t�ɽ�ǂ�}:Lq�$P{��S�AL2����B{�-I��Ƥ\�S�jiܹ�!�2⧴I�u-���S�O�V�l�&Y�չǌ�^!�s��.���1��x�)�o����l#�s�:8�тKG#�q8�j+(0��Y �!�kt\ÿ�-T�E�B��2�g���Y���s(�X�ڲ�Q���8��s��cU����,
���ߗ����\�W.m�3m�q&u#I��E���_����.,�8RCZ�t֡�A,��l �l{^�vpK '�N&��N{����X<z�*N�S�d����0�����l#WL&�<�Y=d�X�9YW_~n�|��ᛯ�/n�:K��wC���!��W�L�3��<��tg��/Xܹ��V�7�����^̅�%`�% ����7!l�j�`�݉G���TH|�(�Mv���7%��"��~	xm��[u5����^��)K�% �C�~��j�n=�-�;�~xG@�#p�ь��+����� NM�88!Qm_K�2�U7+����z[�ߧ|K9ʗ-*t�s.e��pA;�W[�)]h ��l�Oo���脉�kф�}�tx)>Z�����}�7=$T�¤L��Δ��hZ����@���9����,!�}ʩ�|]����>���i+��䩄�>~��Z�W����,���l��f�,�`�����a
�T֋��.���C�k �g�־`��wG)1,aV�W��^8����y�X��CSW�:;�o�4�,�(R�|��h���4�ۿ~;���;���:|<�,�tUu�fa�(�Pt�r�4�~xʑ��.���و$����l�;���r��W�r�����o�����/�m��^��C2-P���#>���^ŋB���/w�5˄~2:R�t��q��sNA9��h/��5��trڠ�U�Q�f�S;i#%�&�4�cKn|�lV�"�d[f��6a͡в�ٷ�ĉ��b��۬�A��+%�%�>P=��S}�gP��A��5A��Եdho0���#��}���t47�a�j�Qz�O)��o�O[�����������s�]��oO�us�-^gc\ʻ��oyT���aRn2Qd���u�vkĚ80�R��Ciy"�o_���ZvC��b�E����J�SA��h��3����5��q)_ū��),�/�w��g�m�s���=����B�� {��ŕ`OTF��C�^״@q#r���
�"��
�N��E�gB'�B�'	ZS$'#v���a��Qg�N����yO���Ɯ�,�?VL%�W��v"�T0�j*�����������{oT���G������S��W	,y�Z���7D�CTW
���La�'n^�=���,ᅱ�	C
�8ï���wp��o�=mM2��F~�鞫ڔ,���/\�=9�@=�I���c��l�S̉*^��ōi�J��f]�+��~����0v<F�Ց0��ʂ�+��Y���Õv���Z�g�O����.�&�ڤ�C���D�@xU����}�3ʓ��/a9SG)a�X�08�+��'���#��b��(@�Lŀg��A��S���8ڿ{�XE�_��8���c��V�N�Yq�͑���T��n���
S�]ɷ���a��l]S�Rm���~ݣw|J�&��n��PT�\Ԏ�U�˦8��,�W�O���Z��Δ�:�\��Rf��������-��C+F�;.�fI�
WH����]a�Cx�r�(�Sܪ�j�	�xS�>)'1n&���g|r�C�:���۬�e�U�l�qϨ����go���YS����K����_Ӡ�[� �a����M.�`�B���?��Q&ݨ)^�?s)`�@lEmG{�"��N��ld��Ӷ��M9����4�Q~�G�9d�����w��(���N2�Z`��TV0ӹ�Lϲ�?���u����B�G��w�ڒ$���5���"~R��$E�3�,�\�Z}nqzt���Tv����n����\F>����)�� V��
���Ĵ�>pA�/J0��M���ǟ�>��AC�[�JƐ����)�%��(uŮA�?p��"l=�����o�myo�T�v�!��;Y�b�,%���7�V[n�B�����2����sXO�o���A<c�7t��߅���B+�z7�z�O��O�f�'b�O��CA���0BV�w9�ˠ�>�Lz���q�wSJLJG3�t�B���Lg%��7-�d!n�J�⭆�}A�w���Ёa�W��z.n����Z��+p��dVJ_�*gK�����!��AVU�a�g�-|���m*�1Z�爝�qdJK�4��9���$0%�O�7V�F���m�pu�E�yQ0��q�A� i���WF���jY^�� c��NA�AR`*�rF�0.��c��`C`�B9�3��~Ϟ/p^�5m��7��,���Xy"Z�#�
�-'�]�B�1�,�+��4�Ⱥ�f_���p]�^�9�i��i���0J�:ңv [8vb��r(ƵW�#*6��e5`���@5���TʫM��A1�D ,�L������G�L�Y(b���D���(���Xݠ���o}k�2�S�z9Em_�C�/�4�<��`u�W,�8]�0%�O�������&�ˊj�c���Z��}��ʧ��&<`F��#����A3������Fu�#԰4jj�E�3t�����(,O��K)��XKi`ٳ=̫��Zq�&|YemH|��}^%X�����eS�����JN��Ʋ��)�ߊ�$��g!���ҕr^C�#b0�E���	�U/�����w7�+^a�b��t*�V��O��^T�p7�+t��5Q� ����\3��	L��C�z�Ry���f��œ�zX�q���_���a�µ�
�,�PY��a>�L�%+�0�ϔ�z����T{Rjb(��gmA�3*�Zim:��o�T~��}�>bd!�~3~��k�=4�쵲�S��)�Z���������ύU�:��f)|h��(\Nu�u#ژ�b���>�2��g��וg#f��g~��^�/_�h0F.���p?0��`��3����ٟ���)Ȼ�mm�Q�N�!+�;�)�取2U������H쯥n{��]~�X����k'��]�*�J"����/���5"Gj���.��#�1
�@��|L���{��W�xr��>�,۫�=n�S��~�[�#�ު�+'z	�H���8ݼ�.|o����L��+�B�{��/?}M&�lqz���@7xܪ�D�O��PZ���U���?�Kǧ��H�F�Na}�^�t�8��:� ��BHCd��8!��K�Q��� ��2��Q�ri�j-��w��t0��%F$��$����2{�p	
9o�8]�m�˪k�}�ؠX���+��W�%rVr06�se�A8���x?�T�o�,'�\D�%X$Xy):/�p����D�k��`��.�Z�X:~\��V�пi5�\c��>�H1����l�Wv��`�Xn�Z`�v�״����6SI�!@y,���Y��4���0����`a2���*l���;���9�ho`���Ɯc����"Q�uw
�R*����b�����C��	���	�,���j�
^����е�|V;����dm�8����1���|T]��2����]1��3��U4p�k���0)Yl�Y�,���8�&�	�Q`���NT���3fc_��0%���ʫ�����6XV�E�T��X[Px������	���B�>|�5�&��i�~�Sy�ߟ~0|E/���m�1�3����s2�pu1�du0���Yc�6�c%��_w��Q�e�1��x�܃�;\��X �=� ��iB�>��W_�d�V���ch�Óôg`P>��C���ѵ�4~+�����V���>C�Eb՛4�',(q��V�R��p偤LY���3��;�?Wܳg�T`B������%�j_�O�c� ���Ϛ�V@��o������=&��M��'�GQ�_Za
?ܔ�1�����P�v����J�]½��cC�)`c��w�N�I}�r�G�.'[8Z�l+����,ާO�<َ!XֶQ�Wc�o�h��;��z��ҌP�������
'�d'O�i��i��������b<��Ԯ��9�e�����՟%��o�55Y]N4s�m´�1��P�j4�
X0�����C�j�5��&z٥ľ���l�a�[�>B�[����� '�Ff�~�+7`V�p����Poq��X�OL� ��N��&���Z���~+�gi&L�	p>���?�59l����P|�"nuE�{5����bb��h@��� N%�)`�f2YÝ�1d}����隈g����p/�>�����5���0x!�vi���{� [~����M\��������_������/�Á�Vw���#�J)�|`���&��<0y�g��~1;��^��R�|1?4�*�zŪ����۴�JP˛������;&�>
�ș:f��w�7�B����ރ,W]�e�� |f˅^bj�OV{K��9՟)��ø�$tu��rZ���>L1*�|&���)`�Py@*����^�$-�Eث�5J�*L�}����N&Mp���T?S!R���K��^��8�d��{����jg�y"3��d	�W,AyLw`�h�;>?'[ql>{meg�1׾	�l`+q���*��+~`TL͵����;��^O[F���LzN�ډ�����r&�m��:p��0O(�p�\Q��a,�A&�Q\�v����On,	�5�o�E,��-��ۤ��ڞ���o*��*#�S�ԥ�Pӭ����ń��e�# %�)R�v��X�i+��,:0�xU;=�����V�^k�Y4�9(�k�Y�G���^}��M]� �T�X4�:�'�?h����\.�H#'mY2n	 ��?Y�E
�!/ūgڳ4�m@J��t%�oq��+�+ %�mS��]#��r���ͱ�/�	3���~`F���t�5�VM���s�\�x-J预Q�X�N�GgaL(v�k�E�H#�Ok�^���^��Ee��p�_�E}�"�lգ:p��bOW����y7��ن� �����?��#���'�Q�X�:�<�뱅 );�8��vZ�a�ӼN�`��U����i���R;���{f�!�;�~�����^"��w9�]_}�g���^���.C��5��耼��̖��Xue�֧���vChR^������×�c�dЊ��6�rí�
�)�ǳ�9�H�`X��f��|4��런�Nh�߄y+g\^���H��6����`��o_����w���������x7q��~,z�Rmt�.��K���K{ӫf Y�z^�vt�pR�W�*����>*-�) �M���ʬ.��zY'ާ�����M���C���@<�X��߼�|����U�����b�Q��_q5҂Y�w��W&�l�o��K��7�I�a}�������B���D:�ZY�àQ�<��g��L��H�>�T�Ө�LZ������WQ	>�F���N��	.���Gf�ޡ� ���G:8sQ��
�3JS�
���W悦����L�y(�S�������ض� _�z����͡��~-:�vL@/�*upԭW��W��*3�C#PY.Җ��o��`�ߤ�� ��V�eY��W���M����r�?��}Nc>�!`M]N�m�M�t��)��4��;F��Oc�c�#�w�L��h��Ђ2]S�-ւc��:��}�m�i�B�kXW������&\?� �<tM�apнf�O����A��aɫ�([��G��j��f�<e����購*s:��"�]��~di;�g�ʙ~>��c�.���Qz}e��������4��]g�����󹔼WY�X�^��������瘥-(��j�w,�Y2����EuWG8d�>!�wV't�0N�F5��F���S����W.�o_J%���fꭸ��&-\�Ԛ��5؄�)��)�'�}�Rt\,2����U?���D#(�?��xR�2�5��*�@�\��,.7w�3oϦ��a|�o�����ڵm^FfD=䐯e�tZ���
��K;����p��oK?�t�JS��~�Y�L{���6:J������L��,EUU�w�˩8�����G\<��H({�9Ks��QUi)K��~/K}J>����<��»U����x���%>�s���͆�h��i^�hH~Q�R�z��tJ�,�V|�6*O�̙��ƕ�B������oС����sW�aH�Ki4���/��mY��ą?m3m(��:�t�Z��0Mn�wSA�20w+\�B݄	c~l���7_�%��W�y?�n�Џ=�)p`��-������-c�{C��r}�o��
VM��4j�?F0s�	ɪا�M�^�a���0�u�i�E�4̦��\N�ƛR�����w;���M���Pbi���Bb+�z-�T8��X�K�05��As_����B\]��&����o��`�`��_��w�Ѐ.q�s/N������6Z_�B;`�����N��|J��I����Y?zW����u���9W�{���V�����+m�y�U�I?u)>��J�]VN�z\0��p��Zʏ� ���̅��D�������`[��@-�U�>
���I���s�?
��r���9�~W���}�7L���]���!ia��Q��Ì6�^0.�ʅ�)�_�����%��E��im;��
1q�[>��jw��F h��Tn���ޗ֥ݴ�p8�B͏���º��^�e��߶�DC�`h�M0�ϲ��`	p���0�7�[˹��8d�#�l�9SD�"$
=@lQF��曕8�����`1kϴ[�(q�](0(�C��q��;(�⓷�\%��S��n����Ꝡ���ǈ!�v0����e�h��)���i��^�=�8c?��S~+����G��^mg^�e5K�o�iϦ�8�gZ��m���y'Y�*�ReO�smG�������2�����yL��ih��*����5���AG�ܻ����W���!�v�*ъj�>˲�T�?� ���~�M�Y9�j;��
�ɬ]/]>|����Z�k��ٴ��3��W�p}�?��dx���]����PU����>v��+���賺��~|�#�A~e��շ��]}��?�����'j� ���?׉,|Y�(�e�w��;G��D���-�s�.���6(����J�Q}Ѱ~�=�"�p��Ct1��F�6:>�te�������_K~vP`�W{����� �;����G������_�ڨ�M���(����pRp)�a�\�fi��G�	�r)�.³�Kɟ�U�g(d��R����=�2Ur�'v�S>�k�i��Q���p7����^�ߛqQ��01���\�����Wv�ε�Zrc+V/���z��zX���'XL'�I�=�3޳ޞ���{��rh[���|6��V�2��W̛�ӏ3�1c�?XI皊y�B&���g�@��	�~��)~ş����xV�q�)y[���{���{A}~���8�� ��������:�����;�w8'ǉ\�-p��X���7{~D\�ˈ�[i��rv�z�oK,��N��;��]��y��¶�N��=H�c9�'�D��$�<="�zT�k�iǞ� f0��
"K+�-bO�E�s'x�D�}���fG�O��.Vغ��,�<)~͡�)c�+k�Fga��S\,��Ji�ؖ7�e��9����{kivl�z�����!�(Y�f,!V\%�N��
6^���4�c�	���
��~�4hؾ�^�Ya"������X>�������!;}0�����b[e��)�z�ߟ�ٛ��Np�ؾs��^>\�l����\z�^A	�U\���"E�l�ގ;9q�ޛv������rs���ӭ4[+���ʶ���(�a���F��Yن��+��(�Tp��gΦ�
J�̆��U6c����c�>����)�O�����2b���)ĳ	d�_��7:؞���n@ݽlU���}������ݙ�hvm������ڟ#�+���Ca<Y���o^�z�򳛇p�<�o��(�?�4N�U�%����?���?�H�,�p���`h#�h�f�J~�bͲ�bw}��~[\n����^\�/3��k03te}w�� U�JC;��<��/�H؞�Õ_�yZ���+x) ���΅�h���^��vY-S�C_��������/8�|�*��X�����O5���EV�S�K0�)��2�g�Tb�@/l�aʿG=w*	�⏅�U�A8�~[M�mceS���~���,���U��z��b���������G)yVN�b}�|�L�^�T
/A}�ϫp�`sJ�(��G���� �R�����]\4B�Z�X�S]�;��Rgnڤ۴���2u �r��Z�T=PiuӚ�	I�8
�ߕV�E���MKᅧ+W��t#ߺ��I�}��|��}��N��z��|v���W���X��o�urm�������_���!�<e�Y�#�_i&�y��x�c�w���5e�c�3�[pϥ�Uף%˺ɉF�����g��H�Д�4#(T��g��2?�X��Sex^Q=Oh1��^a�.a{�[���b *���Λ���{��	_w)&�O��o�Z��qV	[\���nUd��h��Z��<�N��w��4�ـ����½@�v���c��q%���As���y~�P	��_a�}u=��lo�`��_ǐN�⭔[�mu��j �#ejM�UBiw���+��MHa�>o�7A1�
�k�(ʞ�z��M��,���DN#� ����d�ږ�p)`��޽z�%�S?�!���o1+Sm	�~<F�gj�"��7���,h'R欆Z{U%�:GM^g�)V� ����jv�	Gޫ�j�������=�P*e�+\�q�r������y���k�/?���;ۃ*�������]�;v(<]ho��7������9���J�.;��@��$c���_�=Ӵ�=/��?�������?>��a��5��qXw���t���(_V@��ֱA����O�c\ �'g���O����#��?k�MY�b��[�n>����o:���_�6ʯ]ﵛ���~�f�,7�B}���D�����OR�RN���:�<v�zV�K	��ׯ>���>V�zၲ΂8��F�QX��&E�z����n�����çr�C���o�8|n��]h��v��ҩ�Mw�Q8�b�_�I�7�pȯ��N����>9\��n���?�x���?�����6�9V�����y������͎���� ���V��y���?v^l'dy��'�n>��o_~��Z/���&_�:A[1�@�@� eH{��.�z�2[��Jy�n��;��볕æ�L}Z1l�e	EԦ������*�lQ�-�c�*��J�
뿸�'�0�S��w��O#���>F��})z9��؆�u8�X�.����H�r�Z�O/������=ȏ	�-�OY�Y7V��ۑB7�_��|S���m3��r4y��}���l�Km�������xD@�WO4<��u��G7�>�jy����_���?G�N�(�p�=Q�X٠i�ʋ1��e�����M>``���\�X�Q���᏿KQ�\��������u����ׇ흦��A�۪�_0p-�[�(�\ӯR?����a�����G(F�ǯ6�t�N/��`���`,��[����@F��j�!/��׾\���d���F6��t�؀�����u1�64}�� ���ـ����R���$�F� ü�ۋ~��y�#nwo�}q�I��&ӹ��G0NО����[��/����^(Ԭ���?�)8�N�g���[�{!S�qC�SqJ)�@��D6yN��	W���]+?D!��rŘh}�3�m�����D�b=���=��PX�yǩ�i(�U�����n�M^�7Q��q�4OS���O_��=K+|�}"ͻ�~��]���c�}@}Ҹ����"b��͆�C�h)<q�)V�%L����4'��6aC�t)��v�?q"kCJ�MY,��@�@�� d�4J��X�ް��&7�=��V�\��.�ۢ�ӆ��M�&l�u�c.�5�<o�����`A�3���t��On���O��������)�1�n���voj��H9���%� Q���hM������$����d-�rp.kх�[@\�$�������_|Z+΄k���������:T>!����u-e�,ƫ�o0l��T<��]��,a���e��iGn��ow:xΧ0|�r��nn~�A�/-H���?��G�O[�g�¹��O>�y���%�n>LX����hR��Kx���ne�)#u��f���\��CE�xEqO!��`X<!�
���Au��Bh�p*����FG��|>�%i�~���H��k�]N�	��RRX�.D��?�t��on>��|���V�����~��M4�ΑS���V���n�퍏>l��2��򣄍 WB���3,/���ܵ�����|�8�]��t~���M[	� �������]����f~3y7o}M]���4����:����?��F�cP,(T�[h��ɻ���;o��\�q��E,~��Q�J�C�,��Ŀ�[C�u)�V��������?J+I��5Qq�t���۠�����,F���M)6�ejk�.-����߼Y9`G5Mw�&����!�'�����z����N�����||(�����p?F�`fE��ݪ/|��'����o�r��������֗��]��y��O3��MU�P���s�"u5���>�[5���������W�~�q�͎Żw���	ngy���"���.e����E-
Ze���n=��D�\�w�x���	�ߋ��w��G�������ٙQҵ�qǨ�5`���_�ߋVyh,�AD�3N�M�0�:u���z���B(`�ō`�d��]h$�����_X-�����}��O;ބ�N�<�,�cUH�{8`��W�̵ ��o�~m�x;x���Kܐ~�>ř�V>[n�d��}���Ҭ"e�*Q�k������ȫ��<�|v\l�<{>�iW���A��xQM/W��Ѫ�N���A�v�@N�>�tҮ�n]��rGQ�[�+���RJ� ��>�m�m�t��.$a
.=@��~Y���*g�o�N�E���*�i)���&��w�;�3��p�UB��V~x=�j��\7�������/��*��wꨧ��ý��i��[>���[[���MA4�²뜶�{G�3
V
�(b���]�콚L;N��r]��S�����{���I!+?����q�JJR�*ۙ���~�J���yVxeͰB� a�;���F��}��:V	�M�c����(G�}�.��x��a��K����gu �L�Qx4���)���:��bmlUX�]���w�U�h_��qhe��0�O��{���ۭ�>Jyi���br���M��X®4�h:S>�����2~�U{!�����t�Hݖ�A��L�u:�Ƣw������>ِR�#b:~X���O���~���}�$�;J�����:o��b�i�w��K�9JI���z!�B��8�U��YJ���0U��S����8�y�ii.P��g:�T{a1���{E��dJ�`/S�������s#ɟ�����b�l
>����OYE�P?I	c�6]g��:X�uy��k�-�r���3���*A�l��
ӕ>|bz��3ܠ�_�&���6u��YQ�5�n�΂�Zl��	�V��5}���2%(�"8YGg3�(�q��\��h;�nJ�f}����7�����"_���);��sx]}3YV�߿ױ`Y}��c=*� @��#���v?|�.6`��ʕ5��r;�}��N��;W�ƍ+_~��7G�_�Y���R�P����;��`�qۗ?�\^��$�9e��^��L�o�=�o3�<E[C�e�l����{�B�����;8�/?�����߿/ږ~ޕn��>ټ�D�)�IfhX}�)����7#���G��o�̂5Т-l**�+�3Y�"*:�@��\pQ!�����@��\(O�=��C����<&d2�U���͏R�����v\�J�7��l�#/��:I/����w_@���ĵ�gZЀ"n� 
��y)��U�	W�+�^���5��h+�=�%����g��c����o��)k�fH�/�.TXD��I.�<a��{^�ŭ��Wx9V
�hf�k�߳>ה�ނa����E�>�#�����d���i�5�x�Þ?��e"E�(Sc���/���3�'��x#��4M�e%���>k��C�SX^������t����Q��_er�$�o��fg�|1>����2���6�}��m�7�}��I�,�5aR�*|��~j����p|�8���!b�g4+�0�W�\��1I�6�4�Q�J�.�?j�˦N9���o�o�!ۦ�f���Y�nT���G#L�5��Hq����5�)�s�*5V��9��/�gd?��M�s��a��7~|	J�F�b�bE��K�Ք���fN��s)VY�&����wy�u��[���L���.+�=�d�����5����O�: 	)N����w�޽�&j�=j�N����}X�(`������vZ}�~��[�3�|��{4|)gvrb����]��q򾚥M{R�(�;����>uX����X�l�ڻw�D�o�v�'Hυ��yM�����S(z�ZD��b�U�΢;SP�����:��Kw������ڏ�G�xwxz�)�t�i�gf�ά��R�.\��~���]��*���Qt��X�(�dZ46\ ��la�?8�ʖ3@I�%,]38�a%7}9��"���5mfB��؈�X�>�;EIߛm��di��F���;#����~x����G7?7��X�(bh����-R.m���E�j����]S�Y�*]����?��ߦQM�R�m"̏q�!�iO
�լ�7��R�_�h����x��Xw�q���'Y���^���vR����p)k�l�����A�)'�|<+.��HFǗ���S����u/��'���޺���%�\�(!��$��M�畻�{���;%���&z���UN1��Q�������[��!�a�2�#�E@����F�.�H�U�-p��d�����R��{�/*�+�~�A� ��>e��������o��*�d5_+le�թ�U��9-PvH�4��b+őV��L�3������
��	���6��<+��}~�ǔ��n������ޯ�&����R�*jW�-��Rm�U2!��@�� T�*��D?���,S�8+�I>o�+�=���V����Rނu�oB���+�q~`�L{��&��I�ʅ���^=�O���6���>Nq�s���_���Ó�g���f6��q�`����������$�!_��ֿx�{t`��Ǎ޿����W1�u�য়||������?�����q&��|��)7�R`�cK�w(0�2�S�i�A�L��6�������L�����|`���L ���)[2p@~�4�����W�~�����ty�r�*q%��^��`И������(���/�M�a���M�=guL P�XY�޽��H�����g�4%��'�ԝ��q�����|b��)K���1V��?�D8չ�/���v��Ʀ�.��P��/�BAsh7�!��������m�/}�2L�w����e��SH�����Q�kN�	��J�YtQ�R����j��� 7<�E08��l{o�(]D�1�M��L�6��,�����9�_H�����7���}�b��>Y��J�G�ՠ�<��,'��/�Lk'J���5�?�}Ѫv�T~�����w
����U�b�H%��愂���U�~|�0U��*���(�s��U����)'�hl�����dm<ۃ�<�b+�}jt��^���C��*��pS��K�Uek�{5��l�]�=�x������>�O�_k7�;y����/L�q���/�j����ch�O[��V���]�Or��w�_��h��z���rf��Y.�y���{}�r��k�>����g+_����;4��#��s,�*�#C��k�-���=0Gc|�X�}.\p����"m�0w�e�FA�~����^E��&ޗ>P�y9uG1�5r����U������~a��������'夙6݊��o�>��2wQ�}�UJ��䫗�����]��N�[+C�h1J��<�wϮU����ƚ<��8�����Tpubl� ^�{%WZ�ۋ�������_�N�ۻ���c
(�^Ъ�q.���r٣�%��d�BV���˫	�{�p���qW��w�
�
Y�!����5	w�$��)���o���B��D�0тa�q�+�(i�D����.0(g~���	���KuR��p������O;���k����r��m��.I���h	����X|.K���']9|��sp�,P[f�8�t\�t���#�cf�	��a������ʋ	�aF�Ü*�t��@��3��G�+󣜯�f�j�̋����1�BcQ���M�R�yT���.k���qEN�*�3�*�ܦ�^e�;jZ��ֲ�@`�˿��U~jMѾ�������M�g��p��;������~�S�pF����D�lZ����Ȍ�[ui����ݟ�������'f�Bq��6N�ǳ�����YC��J�9t6鬠dqK����:���"q���X>�k�]LR[���u�c�
�6�$�Od�8����v������бU��?"�������$�MI�˚��T���ǚ�դ�	��@^=e���W�C�h�-�v����7����R֕��7�ž��O�<��ʆǬ�	JSShX>h����<wVJ�Q�  @ IDAT!}:P���p�'B⺲����|s�쪏��z�s�8:b�SW����!�0�
ؑ��NX�()c-�#��/�+m<>C��^4���~�!{ɖ �y���[�ڗ@:�����Z3X��='w�|�T�4a8�a��c��X���b��a�fz�Z��M�^�z����h ����.^�)�+���_~�9?��-`��*��0���Z�O��l��u�iC4-O�P��q�Ȣ7��?e��n/R�v:�N��J[��� 闬���Ac�^c������ր��G�1��^���(�R��a[`w��k������@�|�_�W�L}ig�h�ra�]��8��?���E�Hܿjy,�����&劷z�dXD��>pWq�([���D�Q�Rܮ@�x.w�q!B؞�C*0�ھK���z{zy�LB4P�<O�U�D���5����7X�{����+x/~@�t��@= y�}���q�^���Ȋ���	�FK�yջ-��๼��=	W��D��*p�t��R,8V�����=}�d[��;�Ni{N{���������@5:�k��y������Pw`�d�>��1�|��ߊ�h��m�`�	~�3/�I�0�[�f2�v1au���S���1�31��m�F������1��Oڶ���ºfY�*�d�O�w'!�"����h�Y����'�l�6'����6���y~;�/cw�]W�$��� Ip߫XU�����#�|���9������uz��Z�⾂ @��O�{`�H�}���KdddDdddf����>�D��BX�Z�@��
\@�JIj���0
���>LNϹ�(b1z־z/rJ�t�a��^a6��1=UÎo��΢u)�=��uR�����W+E��Fb5�հĽ/���?���3�k���d�;e�Kbuq��;�r%?Cq�����'y���ì\,��}�l�a)`��󦀽L�x��qt�q&�峆Ƀ�^fhFUq0��k�
�!y!k E�⒈�Ug��L�:0̗p�`����2�6%L�*� �2Y���~8pG�)���X�� SG���$��5���Iu�G�b���0c����{?˞T@me����.��0�W�Á��q[�l}�P��Je�c�3DEPn"��1�?�>�F�F(e�a$���Ǵ��K�������̒�gSV'�p��^e�-�J�� �^����4�!r�_�AW]��`kL�,���N_�ñ������~�/~:��]U��Z�숞�Ic>M�?��<�[0y�Ur��^�(ͺfh"i�H�
���%�;׮u$��Q����)���3���eX,����d�.�bi���S��k�^���6
:��~z������SG���?���pE���ZV��cE���o[��q�P�ʡ4���ñ�F�p�D[��(ǽQd�l!�:(c@��]@C=��F^w�v8V)C����z�+ທ�|�g}/�n�G�o���X��6T�護+�ԩ��]��}8����D��]��!e���7��� Lh8beȓ�!~�6���D�K#�Jwފh��:
Ť����Ig�!~ާ�9�p��JûI��)�������`�/%�ʹ�Z�eW�ݗ]��ڽ�o^��+u��@����Ľ���*����(`�0�W-L��%N$��c� ��,�4���R�{��>o?�_=�s��~�0�ܥ���w��@��s'������/�8V���X��!m{��٦�{Y��.���j�P�t�~Y��ể�؀��`�C�d�:�PHr3�A��y�'�	���°���z@�k3dci�˗^6t�0ƹ�`|���*��+�ےf�%�1��n�c*�ˮl���A?J/O%�LSy����71�̫�)4N�̀��Q 5Y�Y$|�&9�R(�c��'��0�1��&4L���ŏD
��?���'���X�����C�T�e�>^c��a
��N��Gy��I�t/K��v���<	1E�?��B@��%��d���wc���%�}>f��e�3dJ������B#l��ɇ�<tE���E?x$��m �$w�"�^��a�I�� $P/7�w�2��]�h�)S������T���:���c�DW��cf�%
(N���!���!UC�fd��L���f���(`�!�r�),z[B�B+�S����V7Br��
��ߖb(<eA��á~(ÆEa���*4
X��h���i��U��7gEih��G��z�:V����=�����
�=�M�-�W8�W��o�.�򱭗��)��)�:8�&6��dk�Y�K=£�ɓ:#����N�Hʑ�f�Ni��k� ��a,�q��<?�
�,����9�[�f^���U�U'lQk7�tS��[����M@�f?��X���m͐<�Y�-;���8v��~=/ڙ�}E��k����"�D��p�o�����K?�Ϟ�0�>�tZ����gU�����z�Ғ׺��"̣WN]�	�S�����r9H��E��YZ��p��f�m\�"�u�<�.�a�o�W�E��G�A��Q�_ѕ�
�����9N#2ٞ�8��o_/A��b�1�v�m��w/��#�m��X��z�����9/~�E>�$�,�T���qb#a%�\=���U�m�����T˄۾����ӷ����y�!8�Ƿi��6䊻�R��<v魔{�ݧ�v�}�S���C�0��"a�	i��as�t�}W'+;����ug���bWZ,����)1
G���P̬���94�*�R�Ӭ���������9�1!
X+N����ޗ�+��Q�6��?�b�-e�I�^ʺ` ���R��Y����$��:)��w�h;��h1�0۟���w:�2K�EL����|;�)y���B۷��Na	�1X��l���U޼x���[���54&)���y%?~`�1���a>E�T����P
�Y�Em�{C���.4㍕��E�.\���X~hY0)}�U<y��Rp��e��zi���˗�sxZCh�[%�O��&ҕ�����!�*�(bk�au�B�9� X��U�d4��6C�/�ao�f}Z'�p7���������oF�����?�0���X�X'P7�2�t��=�G���0���ѽ���/.e�/"Ï��F����(q��\oIa9�[�`Y��
|�m\%��8'pߦt����Km�vB����~Q�w�3%���X��={G�7��!p�~,�vZkd����|��8)��ь$�)�g�ʹ�+�g�qėo�{�o���E�Ƃ�u:f�Xm&���H�x?��ᛔ������ڌvc��4���8ʗ�&�T��13�@�?��nVI�i �h�4ojký�/^<���O�|�͟�
uڎ���.��U��>�D���_�0ql�d]2��ZT�RO�J{=y�j͝�S��?�j{G-�{��e��k�`V;�p�!~8�t��|�7+�A��(�� *<�=�����ڢr��7�rx�X#�
��!��M\�u���쮻�^���v1������H�Ed##����SY ;��D��Jʽ�V�j�<��E	M�c�gZ%!��BF�����vZ�S(K��[e��m��~W�y @`j�t�f����C�����z��4ƞ��D��J�ۜ��J��?��g�'�����S���)�6��𦠻�?��$<(��kU�)�z*��d�;w����>L8/<�4'����䱾�]p�W����D�Icy}E��XE�=m_��;���/���8w�$]?������߯4�w'�%��P�S��L�F���%ƣ��U�МbC������B�/�l'�&~i�@��6+_��M�%;L%�l�E�z�B��o��,��B��W��d�2��bk?�f���aiZ44���=��´�t��%*�>�2���9�v�o3�.�}^�}YWt O}:($�A�{=���"�he
:��0����7B�0��*�cɋ�>{��e��0��mY�?K�����_Q� ���T����(�#Sd.]�o>g�fm����V�����J~fCh��n���ݶ���'-G�a���M1��~��'��0��$�)_�|V�e�l���8i���B��aʔ;X���c�}CW˟�Z�@������)�{��I��,Q�I��@x?��v�6t�}��(a�P��0�^U:x��z���딬W�������Zc��X)S3l�Jf)��p�z�`G	�D�+J�t�'�;�t�G� S6d����ӣ������y霫sp���dk�;y�ҥ3T�������6ڢ�ɉ)xq�"X�����`:�T���>zuz��B���
�׈�k��VJ��]�)nK�P)�I�@Ie	5�L�|��Z/��O����Z)2_��{ְ��`�������&��hrГǏZ$���O-&l�Z�x'#��]ǂ��G�н!���נ�y��[J�3\/����*f�Pe���V�纡ެ�8傯<�U���Q�&�Xְ��,ޣc����x9�^�	ڈ�;]W�u�ʚX�W�o�]�.jS��c[o����ےu?/�O�uxᜯ��Q-����k�\�	|����u�	�}�S�bM)׹�Sb���9�W�?6�����;]�G��)`; �7��2��7!v~����oUV���Sc��E�*E/G��4y���U9"��w�SGdˡOeB��
v�u����!�9�]�*�.n�K�Na�����y�l���o`,�?����nEY��|X�`���6����'�9������aܯ4��;<M�-��ij��Dܥ�q�S�Ή)�-�ַ����v@�����U�+�]:�H?��>M�q_>>O���?�GG�� oR��4�Op����U�nN4����8������z	�/��r��y����y�|�Ϸf���6Rv��8�t�W�^��{�z��Zɜ�K�`nTe�6k����q�q���u���<��\{�����Ö�nĞ�{���41�Y��?��iW&4dA1�@�r�R��_|�Zw6������}��w����0�)���l(��%�h(����mCd1S�X����U����3˫ن)^��s��f��'ܿ1=�e	.޾8C��{�E����K�U��є����Ϻb�˥E���c䫮O"�������3N����Gy1L}�fӶߡ<نfާ�^��2�l}H�L�{�ऌ���h#T�#v�"�A���ϖ9�l���LH\��Ke5T�b��)]C��;�x�.�~�V�3�Xy�Q=\����2M�����7)�?�X�*�����ʊ8�Ce9!X�ZWul�_$��*�z�]	�_kf�����͹�"e�_i�x����O�|��	�����kY<1S_ֆ=}8>~V���u����e1T����N͊�L��@dwN|�ѵ�P]��E� 	�	��
������4�W�Ȧ���"/���"�e���[+X��<��qt����}2K}�kr�&�|�g$�u@�7��QC~?���z�nf���ς}DQ�O�!��[K���_�r8�ḡ����:R�ZJ�v:�u�
��eV�?f�:���*?K�����#�������ɡL�/:l�8+0E��xg����)D�$�Ks�sW��4��լT��KN�Ts�������y�f���z�����O�%#�1��=x:N3�>�/��	�)��΄�pz��i��{��w�Ixm�1Ō�p�l�J+T�be��A<����È7�?�1<#��ů���k��-D��~��આ���W�zM�z��#�Q���f(�9��ve6Fb} �4��DGp�������SV��r�tc+�6��Md�'e��4���A��n&�ݧ���N�zZF�*�G�Ŝ��넚<���(֧���-\�X߽Ā��w�M&���{�f��i���.΄g>���n@��ӏ=Iˡ^���W���O@<���l��󤕧g�bb=Ztw?.J�	��5�c=�hq�I�4;����Z���#e!�w�v���m���R����U�O�+�����]2ܬ9��a�M�ƺ��n�캅��)�&W��	S]�0��D�������
ob��KYbD�"�l��b�ڨ��D ��şI��B���%�Y��m73�b�x��9b��0V��.�ڭ�q�:���?7���1d��w-H�m��)/̛b�B��0����ἝBs�z���9�3\�9$��(|_|O��o���`�+�]˺]��{3�c_��@m�5��r���Oh�>RF�#�2��X? Z��_�:=o�Re�|ŢY[|�O�`If����=V/C��3xe{G� ZJ������k��(}`&T)��T��qM�%(q07m��['|����A���yO�L	<���w��b�#���I��t��,uO����պzoZL�i��8uk����u: ���W �|u�0'��J!�� _��3�쾳u��L֮Mm?
б�K�d�6�dG;n��͒��I;�. M��83�J�E
,ƲpD	<�Pe����Z|uW\t���[=�,,��7�	�f�P�54bHq��&��<�Kx�YD��gY�����[$���_<21��h;K	OA�pV�����d���C E�j���f0�r��uŃgϮ0��P����L-��C�Ƣ��n~r/�
ꬾ(a3+?H�l[8_�`d�5�kB�o!�͇��L�+�z)_���IM�!+��}~RE�����aL���]E�Ȗ��QbV��+�p;lz\*6.B(Lc�%4�АI+�Б�ۧuFl̥�׌w�֐�j�"�5�r�~�:�ʰ`�4���~����g:�̧/J��Y9쾬\��]���h��E|w���~�f�0���� g���+�
ׇ�O��wH���W��u����~�T'��y�Ğ�JV������������7?S���}j��*�ͥ����[�aD�����"%J:A�����=��P�������H�I��,KP��W�?¶�Q0|۠`
��hǁ���l	����_n�����K���u����L�ț��r�i��~����JGd��];��]H�T�S�옺\�w肷��B�Tm�c--���0��˭t�n��s�ٰ��x񼭁�%\��(CB�0!lbR���LwR�.϶<g�Gl�!;
��I��%�@�ey�9�W���D�@�Q���6'���W����c�fU����������<�x�A/�($ Y�
0�d:
X�zg+�"�a$��
xc�W�k.����ٿ��[p�^I;�������J@�6'(�p����W�G3��^�k3�k�?�ʝǔ2J���W�e7���g�!���Vf��F�%ؖ� @�x��*��'�P�LjpR��0~���,sO[Y�]�W�{�fk�e]d����.�ai=�G{Q��(���u2d��ю�&��w]��5��`��w�d�.�f�EN;|���뚭l���g�j[-��~6���,����|�޴v���n`m0��A@��2`��k�m�j�E��7<�~�i���̭v7w��N�@W8����N�W����PV(S�+;SY�U0��аFݼyk�n�K�ŝ��^f���y�o�����k��w�����|��,�����4��%�Ϝ�)~���r3Ͱ���R��̶�Wd7
4�J^f1�p��x��<j����:\��\
��_1�^}W����򠍚�bk6÷���
g�4־PxiA�䫵ҢD�}�%���?ex[{������G2�w�~�|��W�S��I�4%�<���*����n��4Cl��p7�+P�)�?Ƚ�qx8�$�p�٘��zGU|����X~҂�z���VZ�)8طE�bH�pp1��UH���G�N�ՇR�[����W(�nE�
_�*GA+T��(��2�m��}�����@9��4��� C��y�&Bw+�|PwA�1R�ջ]�x�t���uq�vIKg��{'��۸=MB��G~�}��:�)���6�y�~ ����~��o�\�,��p��kC)���VGQ��4i���.x��~�vZ�I-(�ӱ��s������i����xc�4��#[��Ĺ��]�o/Y6t�6
&T1�-��a��̣�$&��B�h�)�yCa��m<�W#A1��L��E��?��k
���M9ԃs�UN�|��Y��g}�9�W�%��E�(��"��eW�YCXY�!�e��Ug�Y,JA@���);��^_`)y�a�>i9�7�g)7ÂVT[�Z��f��lQ��f�H8[��+xaE!��	�'�k��d��0l'�Of�I~>��L)IA��o�P�P�[Y�j�/�6&��y�=�8ƻz�Gi��F|����;\,�QS�@�8�ř}�7�Xt�]�c<�Raɒ�)J�:���rz�=+�3k���&!p��!Yå)�]u��PR����K=�u���HH�"��B�&�+��"� ��u�|�ۄ��ָ{��eR~lف���Q�ɫ�E��5�._M���0���B3�͔�]^|%-�B��L"�3��#����,��w�wS`ӽF�B6\����ͽ�x����"z�4���z)E��[{���|�kK�<	�f7S/�������F���[ �/����~��v��f�C���}U�xV�.�����y?I��r)������J��ꨭ������T~eG���X�0�nK_�3�_����&Y��m��OR����Yj(�{� ,`�%{S������v���j`}B��������AXr�w�>,11N�,��y���aZ���%���� �{���p�	�㴫���i9���j���U���xR�,<oU�k!�g�<��ԩi��5�3D����������h�u���A��W�e�K�����S�m���l�sf��Rn���u�g�k(�*��rJ=6N�x�(oj�o�ԓ��p��4�K��"!�/���\��d�	��8Z���\^%	���b^���ƥv�3U0qݹ�cI%�	�4���iC�1�(�3��+�����L�li!K��k5P5�\`�q*M�z[ۼ'ت�	\���
�1�]�C��]�v��-����<��:T�Jm1o+��)dA'��f�M���1�*T���1���Ճr/
L� S.��,nB�^�ꁧ��^O��pƧH�=�{ֺ�E�B#�m�q�\��D������u��[iH�]�V���ml��DO�,z[�4Lu��Ζ ���>v�z��L��-��kG�W��׹z�mC�b���g_Gf��H>$L�tf���I
�9��1���=�zSf ������c`쵚�Y1A�S�>l�X<��8�D#�����Z&@+Z^�7�ߧ�8���
�h��9�waz�W+���x0h��8�x&%�0�����A3�m���$�!��}ݹ{�}$YS^��=���k�e}i�U��$�n��f9ܳ674��E&�06ԉ�D[{YѮ��m�mI��"r�.���o���s�n�\���'CϪ 9.'�6�.ޥf2*1_�K)L��tኯˁ�}�m�c>9O�S�1�W�l�+��]3^��u�\�	+
����k
7�+�dfK*>b�SZݬՐ��P������V����e;,�$l�"�|���ײ��~Zud!XC�gR	�o��a6]?������఍S�ݢ�W�x�" 4�R�o�����\�֬�x}.��$��vV�/�Y��Q�H0{^~�<>�|���,m�o��xP]�D��[��X��g������ffF�֫:��Yk��R�XU����z"#����_�������/h��v�Wu�R��0cT+��3�ޱ�/��^J�X��rxv�┧���)��W��l_�0_.����k���G�>�S=����/7?=~�E���#��w��9_�d�ÌfC�H�Z�\�z�	!_�%���[��i|�U�:��q�Km���L���?�T����"'ѓ��N������<w���%E���	��Z�Gm�l�{��}�h��m���V�4��QO&8�C�2�l��]rr:{��s����+��Z_K���E�k�~#*FI�D��{*h���6��8%�q�3�x�0���:����H�
�1lfݏ�����g7{5�s��ʨ�T	���)�J� ��@���/�yr������~�\�ɞ�]�X֦��F0���RBz���P�I(d���}���h���E����*Ly�]Et��J���iZ��ޟ\�V�p�]���y�s��`���Sxw�V��G�Ѽܬ�y�}��l3ƁB&�W�����p���z=����W)�8�A	,��i���u/�	(�X��%8��!Ȉ�|�ܣ|�7��z����t���Ð�RS�#6s��)lx>�\�B�sт<D�=�34H��4D[g-�`�c�${�Q�S�Y���6֏��:D1E��ٮqr¦���^��>�GըЇ�Y�^6}���8cͤ��q�И<���u���cu����:� Z�Teq�x�w��J_���ۄ#K�g��tr�*�Wsz��$�8�=,x��r	)��x;��;���%�vD����_��]�������'��+fB$&���*���M<{ږBy#f9�	cD/;j�����^)8�;�`Ǚ�^��Ǐ��_�~��̼�㜥���w��g�P�_L�ڒ'���l�����J�$� �P������0�38��6���
�jdx��HV%q(d��gX.ED-<��k�ڛm�}k��Q�_�f�e|n����0ka����{��!=5j��U��|����G�)Ѕ��;�xo��	 ��Q���岁�?����,�\P�bYj�^uh�ٹ��}�N�F�+���ƕϬ.u{��	��l�L�������ʡ����|����v���\�v�K�/3 �n��f��:/�>��a�����kB��Ouu�]�^�0a��G�;k����|�62�>��P� \���smYɂl�
�`Klml�Х��*��2%�
�i�"�#�˓��-��S��4q�����ro���@�uz^e]ɏ�\=\�G�/��W�~��p����Wt��U�c�O��C84�\�Χ$�z^�]���ձ���E�/�LS'ɂ���a�kf$�d��S��Ʃ��>B����b&��g����_g��£Y��T$��.���^C���=�Mp���,���ϟC�ƚ��}0�Ί��Qw��7�f��je�	�<��x'%>�J��'�t�}��� � >����ޙ�5��Him����8�zA��Jd�?D�#d	ZL����}�v1��*���ښ���ć,o�i�(d!}�8�Cd�D��e��d���zl3�&x)a� J{���c�Ì8��g,H�;�Ѕ$��Ǆ���n������Oqܟ��9=Ds�箥���� ��~�DL���
ٯ7�u�|���.oW������ޭ|��SZקm��1���l�<�f2�;oC��)=��A�|�a��[`fƸ�/F5���>`BSh$���ϻ� ���j�ދ��˹��:]���S}�%0�/rM@\i��Yl<^d�]k�ԨjD�]גK�T�	�r�>.��X'�z��/J� %;����fp-�a��K�*���rl��0ʔ-O�����&]x{�����Ǳ�/������F^���b]Ѭ��6�
m@=��w1S�8>��(&��n֌�z�	��ȅ��쵠jm/�U+�O�o˓�F|�,k�^#G۵`j~s��AB�p���ݻ;���;�RB�$�d�9	.V7{ENϳ4ߥ�!����)7����8�mHm��{L���Ҭ��߲�5�Ca�q���&�t%�xG(�o��=M�|ym�Ň�L�5
����0��f<��������,a*�A{B�u���>.�x߼y}�W�����/��6R0�7=��?�\���bR�W:|Vٔ@@���>���.�N�h:���a8�n�HV�G�$V/	@�g�y�UVIJ�G��o��!�iǒv��m?k-���ͯ7���ެ6�
��֋4��^oj�g��߼y�R�n��/��w�5��*�z$X?d�Bs7���Q��2��	�axfe0t�����㧯�e�V�my�f�E����ﺥ���\�p�^^�5u��Q���HE��_�1$t3�>	�z�ϺV�E+�tխs��/���N��-�(��D	�)��װ}iV��d��,\����Ney��.Ǳ��_���S�xg(.�C��-W[=��s �����g�����Sjj��X��(��6������w�w�a�%����l�u���(��X���=E帵Y�,|�מ�M�%��S�2iCSй���[;!W�U<��+�����aCuݷ���R��+.YW8�6v!���LHLL�#2JUkm`�
�=;���[e���6{�Y�R�.\(�2�¬7Bfp��?�@�]�'%��Uc�m���o��0�:h���F�Zz ��I½F����-~�c
��W���,�j�	!�JNoIȾk2cK��Ͷ01��r/�o�D�t��	��i�����wE���HK�(�m��n�]V�	����Z��!�]�Q��K�MЁ`���ݥ��[�d�Xy���k�"���R�b��ׇ����Q����o(&���0��0�U�v�	��F�G���
�}�c}s%,l�|)���+)�5����j����̴���[��R�#gb�S��d*gŞ*�qĈ:���-K%73XùT��:�� �QRj]�J�����1�z%�sSCܖ�4��ڜ�T�JY�@��T9ϚSؕP�^f0F�`�����f���i2�i��✇����au���,%a�^t[zh\�*��Ao���U�:}�ZX ?��~���6q~5��/�cI�'5+sm�#�ؽS���[q�!+��7n�W�U��1\J�}E8f�X;��x��L���i����Y�1C��&���������T����,n�#V���J�e�ȫ���z��Zg�0zy�J����ȧ�8�&\F!(��Rh��sz�vґG�A�.�`�l�Q
Y8�4]jI��)����᫯�la֛#D	pul��0�����З2R��e�"���}g'Y���Dp]	��:�gh�>.'��� @���h���
����F
��buhz$�]qZ3+�|'k�W_}��*��N�@Q2\y^5Q�y�W�	��wP�3�C�r��C�i\���H��`h׬>��X����whGq�qY���-��7_�c��6�<�
�>z�G���m��Z|gxO������������0
~�FƉ���m�w'����ދ�?./��E�Y��%�e���M!��a=���+�l�S�rW�ȇ���2v����vF`�$�
n�����j�
Ƥa����{�g5�4ڿ�B�8tג/�+��Y�)�nR��jT�=����Y��s�������%��e.<�|��|AM��=+}\�R*)�'��6�����u���]s�����Ӆ�@!$;�Ử���Ë��F�V��tL��ҋ��W����|�m�-�C�vOր#�_��:cB���~vuW��C���m��FpS�j���� b��Y0���@u�!����V
L�=��^a5����j�슑�s�A�k��?=�{V/=T@UP6:|#�Ӵ��<�@!\?��.� Ƙ�ۮ=�_��A����#�b�Д�b�Ґz6�2����S�f8h`
]c1Z�2e�ڡ(��y^?��E���\1��,�Ϗ���p��4�Ҝ�^�r_�� ��X\w�vq�\�]�w#���w>{\iz�Al{%}ջ6�q�r�1�E�G�<�q��Me���3W._�X5�s����":ӳ%t�=�dpn�2$�9' _�p�Ɍ`���E/�ڵ�s�~������Q�IMe/!t����ǘ�^��M>=q��qB�$�cV�V�1��)7�������
{�JB�a$fsÙ{ьu��i��P�!���y��TG����W"g�6��n�D(oCW��i�h~/�cS���X���F�ebΧ�]�rg��PeFT�h� �j:"��,�C�	�xL��S���������v#���~_�Ja�j﷿�]on�I��-׮�����5��B`VVR��E�o6x���Q�P��ן��jh�c�G�V3��^Ĉ��<a�/�f&�l]�P7��%��@f��N�b����ל��Z?�@~U���ݏvS�"�a������)f���S��KOh�7��^��2����e��w��fە�tRS����a�p�~��Ejs~6�;��r0i�����ٓ')}�����J&X��u�aՐR��}yws�΅��XY,�i�p�(� %�7��|��& ��M�`�{W��a�^)n�*�����A^M1fU�$k��r����o����͟6?=|��4�Z<7_�3������Ғ��h}̺�!_���<,b{���+<�3�խ�S�gȧ<�����gh��V���������>��������o�T��<On�X�C�!���d�&��^�c,f�S�x~}���X	�ä<=kǔ'��{քҁ�l�@�:G���
.1������3r*�cֿIE29�9r�4(�-��,���JV}%��x}j�J��i����mv6������V�X�"_|���B�S��2��� �X��^+K�(4I�֝kc$����7)^������͏�ؔ����ˬ��?&�O/�:)c�S�(`$��J>hh�����-hU���E�:G:�U�����B�831��&È?�	�:C��3�����I\8��L�?j__��	Iy��k#w�9�Nl�����5�Ȅ��j2��]!�����6�Rqа�IL��i�tT�z3�>fczM,��e��p��
�SM���\g��)m��m��*�0r:���Y>QkՐ��%�0����vm�K��{ç�#B9��ٙg�[ƨL0��:)ag����G� T�`��Ғ�?كw�Iǔ�����g�ZC݅��O?*x�&��R��ʿ����8�I�t"�{�h�:N���ݷ]	&��a�U@�|1�Jn=O��,AW/�Fr�_���|���"��	��	��5���ZC����+a�`3\�K�� 
? ��Õ��:-#�:s��I@w��P����X��	�����T��?ւg�G�a��5��� G��]P��Ԙ��!V������.2MC`����#�T�#�^�!ߡ�ĺ�YK�ʑx����_�)�/�5eM �ɤ�w�6zs|�P���E��]�I�bB�*�i>33*�;��gx�r���S�c�?�t�ꅆ��6>�pPu� �����/����cF�&��� �JE+�"�ݤ�^Q^���䰞8e���sL�I�c�Zluc,nwn��X>$z�|�(x]�J�G�K
�b�����������p��Ø��,�߷x�?=�<J���`�{��٘��&#=|xs��s����͜�������:O�ۊ�zS�����-�[8�{J׬�U�sZ�԰$(�:��#S�Y���|���~~u����]�jNCoY���Z����7G�6fd�l�Ge����Z�E����_����1<h�p����㼫 ,�KiW�����v�@���	Fk�}�����כ���a��)/�^mb �«設m�,��M��?���%t�,wP���EJ���*��
c��6�pJ�̌@ȫ=�2�JJ�ƈ�k�������}j�+��F9HZ��o��������"������ov
5<��	3Ei)~�Z9�t�q�y�c���Ք�Box�Æ����脯N�3�El&4�����7�����q�eZ�ah�u�?嫏)��_o�?|V�6]�;��km�v���ѹ��(ֲV.�)eR�C��a��)��BYȬsY�-m�C�����7����]��)M�`�$���^�C��D��F�j�Ѵ:_��E_�2�Ǒ"f�Va~��O;��X�G��d�kYu�*W��X��Z<�w�E��v0�{�ąm�o)��e�������u/^r�!�{_|1���7��/��o�,ڧ�S���c��G1�s�}�{�rfd�'�]�YP���H&���SD��+A<g�h�N[�(�`����,*���=�R�
��>�	���1����AT  @ IDAT<k�d·mb�X���/-f�C����Iw>�й�p��>TF��!�T��^e \t�{)L=���׵Z�����f��v�N��p�c�,^��f���q��x� �`�4��R���0n�eᆁx����z�7}��+�ީ!��Ͳ"�߽~�yؐó��в��ݼ�פaXWƔ�K1�	]J5�ߐؘ�%� �Z��^��Ow��J���^54=a��|b4�tf��	��[E�b��p��v��X�X1���#>m�p�10�TL����63�\i�mm��0V
���f���3�@�h��
���F��,N���{�� ��`��g��R�N9�SY'Ts�.��u0(?����?~���(`����׿�����fV�=C�W�𬏥T~���YUư���z�?4��fC��ɟ��RE�M�꿺���Z���^��wY�&�� ~)4�Y�{�v.+A������O����?����ZZߏv=+�o���6�m��/fؓ�1�8�	.</ڀ=4�ѪG�!�A\W�1��'͌d���w�G	3S�Q4Υt���_׹����<���2fڻ�"���䥔����(�3ms����t�.�E�?\��P����Ĳ�c�I����?~�����0rV��,|��_�W7��_;��0|<�C���;JP�6��)ozܲt���WH��3\���e��9�L�[	y+�ğ�]��7��u����כ�������nVh�u5c��tXn}�~s��6{)��o���fG?�.�Vlu�^� &���F	c/F̠YmO�)��l,L�ȩŅ笞ܶE��o	��3l�+Es�Ko����G��b�@C��@�� ��I�w:�^�
~b.��Rk�g	�S�#Q�)�e�z�~�6�~҂�ϲ�ܺ�B��(���hw9�,�˂H�z�"��~���,��[m[���R�4�/���h��כ�����yn���(�蟓�aM�Ҳ��͉>�}h�j�_	W�:z)K�|-�������OS����)��Ik̭��N�p|��E;o��\�>��u$<R�0a��;�q����ͭvm���t���+�)t�R��X�ԟ΅�i{]��OXʖ�U�S��ߎ?�g}�C�W�ы������on��ӖOj������pw��o���&�|8y>2�{JN�!a#���Į�zӌ?��^=��KJ�XÈ╸}5Hҝ�NET)u�k����#�O�
X���1��f!����SOqkL`Za�0�\���b��}���(���F�Y�TX��9�I�.Ѵ��g�@S�����E��p�&��SX�kt��@��x]E�~��`ʛ��UC���̈́��qq���[���6G��x�m_��~E��t����6w+z�S���D�|Xl�c����~뙌�)µ��̼���}ڍa0�jo��Mí�����d�	�������lim�[p��zRE��Oco�m��Y����c��X�)*a��:e��0��As~��ת�'�����o.à�o9$$t,��GiI��E]��v��n��������N��M��u��ȑ��Kļx�y�-���[�PǢ�����P�(o6��:�	�h��5X>�|	>�[��a�c}�rs�۟�fx���Z�az��{tP�j�f~���M�xU#��������c1��YL~���u���3�z�2s�b��R�(�K�%��?�C]1Q%Q��: R4)���f�[�F{o ?�����m��3R�X�=Ⱥ`}1t(n&�FX4����Z��̃G�gH�N��Wc���(�9��a�K|�]CS��ۀ4�e��y[�|C)lf�m�tTo���Zk�|e�l��X���3\���������4��Ѣ!�k�^M��ng6o<�b�d�����Nu8ʗJ�-�ǈBt�I���O��h��G�f�.TZ��Q�XPl�^��	n��yR>{:T6p�i֙f�BC��*/BԽN���V���&�+3��)A�}��E�%�z_��@�V��*��~<a���|ލ�W�JE���|B�q���nf��0Ьp�Ef�K�J��@Z������_t�������D	���O�}�`�C���Yg�r�E�6K��x�"��l��o�xɃ�,�� �yf���PsK�����Y�ds6��zL�B/�CZx����f��zY}����*�Om�Z��JX�z�2�|��&-���/g�+Yn�5$�#H���C�W����M���i�7
X �������>�iYlw����8n���p��-T�hD��?�0+�Q6eg�:�Pg,�����\a(h&޼~+�v�r��6 ��1��D����[�����]��#�/gm����0<@��H�nL׎*Чן�����-?�Ri,_�n�+�=�eR�D8&PQ��!�&a/Fluq��=��c���?x��y��7A�>i��^cp�j���SQo���X�y�Qe(��P��������E�U���Gt��ٽ[����=�U���'ֳ���	�e���$Q���=~J��o;����,���rf?�b�Yc̊�;�/�>R�"DV����k�f|b�iS��:�����;�b[�m9P�u�鉤`�>�c&}�K$3�]��e����>ƥ��<�΍[9�$��?��z��C����7{�)��c{��� �tf"aj���{�}��B2�u��Nzя�+�]� �]8��H��� ��Ճ�֖E�>��Bx�������5�^?�G(��jx�3������X7��s=�6ȣ��߽���4�ėa�(1�㔵�/RJ�G��Mf�,�kճ^'�������x��b5(m�#��S����(T�f�2��Ũ��̓���?n���?�Qz5L�8������8�!_�ӳF����d4�҇SD=|"f�7��I��I=�G)�O_6+�Uտ�1�K�:vS��e�p��[^����u��nfKZ�� ���������Y��n�Xc�R
��\Bo�4�	u�%){?�ۥ�����:�B�����IV��y|����x��`���4A ��M��ϥ�m���t�m��c�5/�oZ��2����zux���%��%`/���1�Z6@��x���?tr��胆�^5��Y6Y�f����Oi�¥���г�[�5>�zU��c�O!@ˌ2��E��^ '&3�L�*�iO芋\V\�W��څ=$�~:��P��q4�X�a��VB]gj �m���f�<��Fy�QeS�Q��p�������-ؤk�U�`}W�ݠ�p��y����T�z���U�����S��yKj<�|���,�W����tCw��CK�|����OG{�"���x���x����c� ��꘽i��O����`\j��{Y���Y��D�h�Z���	���o:��$��,x6�&K��~���˜�E�G���Uu婍�3�v�������+>���?l�������_��:��Ҏ�K��,gk�?㉃25
�Il:�]w���A;B�kJωc�J��|f|�J���(.��U=.��Չ��XT+X���#���:�����I3�˾��f�V8�Wi荏��K7j�wǼ;S��#�S�P03���P�f�P������n�BM�H�ba*�ߏ"�]jcM�T{��W�k���WC�3k��[V4~wﴵ��k)
��x�j�O�!?�U�E��L3�#kI�8滅�����_5wn���-�z=ǎ,=�}� �o{�4�q|�v�|~���]����b���"z.�{�wɬ|>=͗)�w!���g'頰p9�������}�?e�b���`x��bކ#�V�-��p�t���Y��,�����`ޖeW�]	�u?�تwF�3�2��ݲ��f�L�[�����������9+KX��M`W����{��:z���N����k�֧��`�v9=v���I9xV/�~N�?�ix�����O0Cy���1���q2��p��$0��O�0+�γѶ��~�FD�@ue�[S騥�5tp|�<��&ң|�^�R�Z�����/�gZa�~ç�I،�!{8)��5�``��_g��TY��q���m�'����`>�<V��m,�V��wZ�L
uU)C���)O0������~���~�,^[��Y
�+4b���Y��|3gM���YX�+����h���ċ�6����\�z|�^�T^m�r67.������K��8��~�5��_%l	�7!�63(S�Y�!��a��ꃈf�TO:	cIq1Z��|(<%���G��6O�/�7�:|���yʔ��f���p�T�x/: ����Qՙ}���,4V�ױ"'�F�r�hج����8�봰����J��E�N�|��E#�51��������wn��gm�Nf�N�9��y�M�ӟ�mQ�+/��B,$�::��&�� W=W�p�:����*�S]�5��*A�V��YOڥx�FNVn�$0yJFD�rT���jG���<�t��b@���"G�g��.d�[��Ŝ��O����3���48��i+)�cݧpt�Q�+�i3�%���&�$�R�S���^�x���Mz@����N[� OAwx�,����~|����?T��+������k`
4�_p��L�~��K��7���7��b�/��7��E3������C`��!�q�ul[smksh�|g���zF<��uů�m`O������y�g:��Uqt�-�����u�M��FC� ����x��_�Ͽ�p|*������v���C�b?���׭��Y��Lj-�`�[XHUB���~����Q�ʳ�YD?��k�I�z,0F�0��X�zOc���@�^>��-)0f��l`(�e	��I`\�|�����l�7�4��?}Sɑ�(�Z�_����9![�F�崯�kl��$ ���g���pR�yP�D����������Xa�z�۷�l�³���bl���Y�}J��O��'@W���6�y�}y޶�U݊3^[�4��Эa��f@�l��aƯH��_�b��Q|j���c�^�T�|V��0eF���� ;8�2%��_z�D��}�5a,�K�ܮf�&��%����l����	f �f�MaT�W1��z�	˽f�+\���	�e������~�=b2�SV�-G@N�~��·rR�,�`/;B���ML���ݳ/��%!? �D����q�3*N2xu�e1�|R�X�ݖ>eY�q���$��Ջa%�k
�U�u�p�,F{{?���A�Y�o�:ţe��Bk>���kY+��h��/���^Š���6kR6/���e5��Fg���g����� ��V�A�-�ɱ� �|?��M���r��Rv�Î����oR���2���h������x~L{?�@-�x6�1R(L����xN�R���u���˕�uW��}�g<6�wz�W���i�$++����a5��ي�����Y��1��T�*t׳�\A�3	��՗Y��E/�+���}�VF���LkyQ�o�m�d�~YGٌ�cCNM,�x!^/^o�U��f~>�|��C�ޱ�ĵ|U�/�<���T����,��Ä�aFB��冇�����Ti�/��������M�Ҏ
�ݫ3�8jŘ�f���K}YJ���/6���򏳨������,Yw�5�J���W�iG�l�������~?�v�I��Ű)9�2���sC�*���\S��>���Sd�,d���k?�?�Fյ�rT�����u�o��o鎜�vKޥ ������\�����[���)��������k��:�i�C���LP�ǖ=H�ئ~&�4����m,�N�x���c/J�a����������f�6C�/�a�e��pOV�i��a�$V�׵�)�/j�,p�	o����:ώ�+��a�_'�+��t��/��|�o���a���|]^+�f#�M��0�a�v����F�|�t�k_.��k�:ǃt0���92SVψ[�ĤS��l�>��h�4�a��p�X��T3�1|�e���R6�`ֆ�tr7K��_|m�w
ع�_��tєC-�0�Y��������"���E�q0]�6�W�Q�z��#��O}�n	��G��v�1O���PȾ-�P����1�
;��a���]��XlaV[��r#�Ӿz��h�כB�!�tn:���4j�iɍ��0�w��k�˺V�V���C����?�Q���uTL���]�u]��ٻ��n��z��+�>�1DНǕF��o��
'��8x����,SҀ?�z?��o(C��w:���s��Q��x�������d F���d�g5��<AS>hc2��=�w^�/�N)eb���<����X�w��v2������s	�s����½����<Y��w����o�I����`𯙙�@'�';5|L�z�Af�<=o==${�.���]&�/L톐�+{
��fq��>����<�f[3/��sEYe-8QṘ	S����N����|1����m�`�򇶳�嚹ܵ|ǔ>�%Z�̪��pұ�!�4�C4>g�3���:����?Z��������tŔ�
3�����~��Κ�qnݯgx9��R�`��x�)Z�����qz��C���/���<��̄ Z�β8,HN8}�VI�>�:�*G-}r#k_����2%�l��~��Rɢ53Q��lC����SXq~Lx��f�r��'�z��+	=F�C��[���T���=�n���=% ���L~�-~H�[Knf�Cⱺ@f������s�s��1�|~g��uqr~���͓h'V�����"kⳬ`,���n���,Z:��.K��E�uPrװ��e��6���$2ҋ���\V���-�r���zy-�m�Lty.�Td�+aJ�X��>����0�߶V�D�������a#+\������	��o~H���đG�->^�z�E틀�h�b�f�����%�Ļp�dYm/T�\d�G5&Xq��;����r��	D�,�Գ��X�)*۬�Q��ID�v�$�����Y�'Ͻ(���{��0�dk�,,B��<ʉ>�&�p����Y��ߘNY�|�@A4V��&����:�g��}���~�Ƈ0���p�r���O���jmx�Jf�ϐm�"31P<Y��ɒ�&._��|y��o�������φ�|h�7���W��Wǁ����Q^/��Z�Dy�Q4�-�p�-Y=C�=�g
\>'������������n=�_2n�͡��V�^��ϩZ��?謰H�_f���3�[]����¥֩���ۿy�����/"0%�*R!�<k�p8���N�S�Q���:�5(`w��H�p~:��{1+5#� �&�U��i��h=���W�C�'P���l�W���i�,��Hq"n�����4�sws�k�\�ح��m���_6��y}|Xx�z�Ґy�tj�12c�|yfy �7���B9��_}����P�<���]*��oWV���^]fI�	1�&�.;,��巋�n�"9�a�b�ۊ�P���ճp����>���,M�Q@'�,������֛��Eʴ�E�uq`Ä�\��{�̰co���k��	m�
ޙi�я*�!e3~�d�H��(�A���RB���r��`+,���Y&����0�K��cci��(�A8tկ��/$4f����),/%=
X���ef)"FKe�ad�Ae��0���a��֐�:�����bf����^n��V���o�vs�L�FZ��N��j/�������^��2���^e��o|ߋ1��d8u��W��kdʒ�蓄���7�?|�}��pAxW&����0�Y�h���W٬	�%C��s-�p=PnרϦDXQ�r���Ļ�V7�ߥ�F���0�nON�bƖ���6�G���X�5�F����3��U��2�=�ʿ({D�8��0
O���'k��'��G�'dI}��ʛ�6V��F�g)�?5$6��<|*aA`�
F����G	;�P��Y�O0�#"k�۽
֥wш���sq�_[��G+�=cmH	:��lt��iGG	�)�_�Q������zs԰b~b�ԜcݡuD�_p#za���b)���!�%,�q�/q�K��vtr)����ϯ��~��:�ў�Y��ǃ��G�@[{߯�,!s�:y>����ϛ�����j�%wh*��^Ёu��4dG���UN8�L�q@�|WYM)y��=���Ҫ\X�� 婊E|Xu0,�r.i�����[��U�X�����-zʱtʯd�3\5tnag�fg��P���;��6�!���������l�\<��n�S��cw��ƒ�$
Ua��E���lx�N�Y���>�����_l�n�B�ʓd ��=|?܃��W�ze�c�Y���Q�NJ�+�N���X�2�7c�������
_����*��]o�=k��K���/��~�U��v��b��t���*l�P�������A�5;[�&®��!>f�ȌTg�R���Xy��@�u���'�M�0I��o_Yk�]j+���.g�P��򵛝�������ْ��S��IBc�	y*q�DL�n)9�
	�r)"
�F3�S-�9?�Fe�W
!J	$���9���Ө��'��c�1D��}��b�?W�5T���4����ې�f�5��w����N1.��p�ey�{��nj��M�4C�LVB3Ѥ�s��z��N� RZ��.��	���O�@�v�\q&޼��.v�[H>]��>mӞ���Mj��O�
���N��m#M���F��s��- >�D�x�c�Ҿ_zi�kp�I�b��d��*㮜�u�;�ա��WH/v��U�B���ߣ��$����Q)�,� ���P%�\�ɣFRoR�������Uf=Y^�#�a僔����>�ˮq�-��)�����7/�9L#'h8z��G�!��:cE�T�ee���,��5H�lu����Ka��嗭�t��r80N����Dﴶdhk�Q* \(�^�O�zR}��
^wۃ��'�"D�yC�6,�I���"~'�E;�r�S�)~x��4V��ӌ����s1��_�~+�M8�r�n��j�>^�p���Qu�1����u�Ѝ!C��B=�����$�D�}W~�h��
����+�oue�,Y��|�ΕA�,�Z����n�8�5�����S� r�[��`�Z�(�������qJ�U�J�S�uH�R���3�6 ھ$�f�����ůC�5Y��HB־��6Sj��a1�m�~	��׃�Ged���G�����`>_�5��b�@*,�t��%��?�zU0�x~��LK���$��PY�g��;}��@��2�� W�~�w���	����)�������me�� .�oc]���ৄ��:,�����+��pЭ�Ԃ�k�L����
�Ǌ�����ژ�����^��f��{闆ʮ���r)���Z[��6��)|������"��Ŏk���W~R�z���a��n��N�N=�DR&�Fǫ�7�Z��V���Z�W�HyZl���t��������Ӓ��"N�%n�7�ï�����.��J��z���ҝ[76��՗��������"�)�%[�ٰ�����'WZ��Z��7[T�V�XG�"�:��q숗R9N��ɺ��aѝ2��D�
K9��� ���ǞɵJ^�1�=�o#��&�8=���u�N�5�1^m�KC����x��A�*�xT��s~3���oR�4AJ'Y�E�a0�Y�z4̳3�0�v*���cW*`�V�P�)t7��zBa���C�6	�����Dc�[��0lh�&3��=�U���q��9aG����)L�ѣ<����4������f#����l���W�
?�C����k �'՚�0P&�ٗ��Ma��m���ű�U��>?��g�Z��u�e�y*̖HHD� �xú]�y�^�>	��~A�^�#�Փ?�yʲ�
~��X��)�N4���E�!��P��pB�I��-4zs(Ji�0Т�u��U�{�l��xb:���,�;̾ag���� (o�%����o��aC�<�,3�603~�ɭ�(^5���h�k��5�Q)����%*FL��'��ԉw5��֒���}]8���/k]��0��B#{�7I#�Q�yk`������=+\��}H�a�Bde�k[8Ð:4��0�~��&10V�Sd˿�"��9��K���F�4�p�&�C�j���VP�0���.�x)P�m�ײ�]��^�Y��M8����uȧ�t���I�e"�e�Z0I͜5��_����/sJ�(!�0��0S�\�3^ºͺk\{�ڀQ�.�$����l�YT=����`�b=W���fKa	�A&LX*�,[��b����r�����}���E3���1��LB���*qBЫ/0j_��p&��S>����$V���I4�#;�S��GAs	����C�!��"=��q1��*.m�:	�F��9<)�����ׅ=�9�R�"��-�+e�6z>E-z��h�5�.���L3rϵOe��o�B����0������Űri':(��V��������V�o6�\$�*^G�1;�/��;E��ګ�`T������Sm�Z[������R�;Y&�vֽ_��7c53X�g�.�Y��n�-�*�SU���}�wu�I8�pa�V�S�W��jѡ�F^F�c�N�+Ԭ�YB��%�"���7�jYJ�t%�YX�|��N]�K�����#~���|�`U�¼�>���C]m���	�q�O2,�B�Ϩq����f��ۿ����|'o��͢M����w�ݬ�ݸu/����F��%�S�f�ӻ�6��}�RV��U`��"��E���F=a��BVu���p������ �i;��F�`�ֵ�-Kc&p����	Xso���ex�A�wJ�p$-p���l�^�BY�Y���h��[�kէ���1�n+��Fh�pJW����)����>�kb:��z���9(���$����L��77B��0O���͊P�V)g�6.����TF�^�2��u���*�i�!��?<�'�M����o�+�6�	�G�X��@B"|�[�s	�A�ѝ�P1��
�=i���;�/@��CYד����PC ��L�M���&�琚�+~����6u�-L}Y��qG	�1��r�>�1OKu��������J@�a�P.i��"M����T�)��)G߼7�-��C��,e<�'l��Ǘ��iR�n��
�.��Aa�u��%yW"ʺz��}���M��wD��,�`��i5Q�C5�-M���0�`?�w���|h�w&���=��4v4kޙࡰP"�7PF#�q�x���@�UZ̲t�A����ù,��W�j�4*�ԕ�buO@cg7B���Ga�7\j/,s~�"�cB��b�3���琞��W�_�f�j�~/G�%$ϵT�A0Q�������Q�H?
�K�(�R�	Jt���|�%X��pѝ%��s�N�(�w�0C$�a�G�s�$���C�@CGʭ`%<B	��UؖQ��W��3S�)��5Zq(;�V쁨�uL�ũV�>���M	��?����Z�]&ꬭ��D��7��ɹج/�A��T>)�#lJh	� ��}+,aA	����h_v�;[e�m�Ug,)�%I}8��m��C�� �)YC�f�4�~������3�NEf��p6%� �2tg���,Ъ�I?�R����?9@�a)\(\�6Zu	�� �=ic�S�cV��%uJ�X�_>�<m��g���yX��߽=��k\*d�1�򜌷Y��(�"��Wg���j��Ҙ���{a��W:��S��Mk�iaV����ee��g��(��\�U���gʠ����@���Kr��a�FaBa�J_%�)˲���u.�	7�]��uo��_|��$Z�il���
Oa���\m�w�k�r�_�V��Gee,yy��-�M�p�/�v�h�Ӕ|��mDO��ru�l��r��&��7|�#G�+�� �q��34��K�nב���g�L#"�B� oK����Mf_J�L��@�w���	��E$���*$>[���"|�\���V�V�ш�\cx�9&��$���h1?C�n��M���Ů�4�;er�`�SYvb6i���w�%�L�&�uDt!l98���1�̜��f+���έ����_�;�nsx�I���bU��zp�nJ*S;��!_EL�o��d�C�`N��8-S�p�9� S�0�B-� �bu`��)���窥��P���a��|��zrLϿx�0ԸkI������E�@�UA~��J)��#�<� p���0po�Sdu'��~Y$��X*{)�EH�$��Uq�qj��^)�a��%�}7a4g�jzq��8d�~��B'u�1��S�H���й��G�1)3h�.$8���K܊���I����7(��4lq6�a��I�|S[h�����
��U >���]�#�FP��|1�`$"����8�2��H+mRWa��t�b�J�/K �7�-g������E���0Z���I��mh�ަ~��w���:� �Ӱ߽����U?U[I-��k0��(%��U����(��.\{�X{&;�+m�$�U�hO|�p�������?�ci��")nغ�y�7OU݋�3�����ԩ��U"j��&�9��������u���(o� `[e�q�Xz�!mbl��4���$s`����^��Ǭ`����v3�7ڼ�d䂗���o�b�k&�q��Njt�;~�ż�Ǒ�g��d���$,y�s�s����}mo�<Č�k����8J���Y}Ħ}'�/��}V�������Y>Uå�6�������3��3hz茧�a�+嵽%��]	a�A�����:���`�YČ�,:c_�u�|�"˷_��R��\;xU�����w�����_|�S������ӕ'/��f?��Yq��=�P#N�k[8gp��y��(�ҿ�^��k��a�g���:ެ�p\������}o�y��X�����w��c[J�>��!S�\��|a�v�mwyi49�G| h)��{ë(.����e�+tn���jѯ���u��?�I�s~������9�۸����Yg����,��Q�2��\���e1}�}�O�[|�
��_Yp�����?iS���[�e��7ob��7�y�Δ^מ�ʕ�Ѭ @����/��8����ܜV���G�8o�!���J�4���J�k��j��y� �8J&>e�(h�BP�@�ՠNFN61e���¡{�m����?�g�f5��|ʯ��(}t�/J'�J�Hp��)SΗ�4|��w������8�}��+�+���G�F�X������{�C��M�|��3?��py'��x�಼��0�F;VM5Q�Fir{e�jX�`p�n4{�X:�Ɯ��~���A���q,�������]�CDy&xY�!(r��1��"�i@�:3���3�����\�y���������c�&�L$6���0^���$�P�2.V�N���C[��lJҴb&���O���\�5,cK�E?m��P�6՟�Zc�T�A�C�۠+8Q�˷6{�ɣtt�#r.���$u�s�c9���:4ӂ��	X+��㍃c����n���	\�P�m��MAՓǇ>��������5�x�v���f���L�i~���toqz|E���æ��`;���'m�B��k�.6t�J�P':���K�&��'��ۋv����Q�v!:��s�ϕ�m�:�_�ˉ���D崅�l��?:9
�1�$�����{ToZa��01/��N�y��W�[�����Om�j�S�j!Jl�-������\E%"]��C&x���1�� �,�Y@N�:Y#���r!�x��|��5�u��8E�`'����H�6Ei�?dr�VF+S�'�9'Q��Oo� �L�MWbg/P��!�^�{�r�_�g�����^_���'��u���D;�U�}�[��x�8�mr����|�\'�cύ��F���U�6�@>Ϧ�'�����C^��9��c�5� ��b--}�_���;��pG��/�)}+G������	xy�
�
�M>{�2��d��Hi�I�I;)�r��Rg�1�ʸ����ż��r���L�mu�p^�#�����.���'7�����ʾ��W�z�e��6�C~�� iۍ2��܄�w��y����_��c~��9�*��Bo�W�*�O��������	ߥ|�}>{�彩G�%^�KAp��hd�t����$�+I?��f���g���l+f\A$���u�G�d�C�.����=V��֥����x
�$��6�7�5���,F���b�]�fc��Ug&�4Щ�!���+KxN����8:�E�8p�޻�����G������Kx<C�����	$�����g�*�G�\tP>{XbVV	��b�!��5=��$wn��xE#���U_�7�z��%�_�������s��?������{T<z�I�/��B��tt���Մ��~f@D-wp�����0r���Ϫu&9�ڀ�_�I�v�`�O�)w�{�HI�с���<�$K�a�nd����Q�t4σ#e&LkN�?�ʁ����+.����� Ce.
��5;��N����H��[ ꨏ�D��r�HA��GtЄ
�2�6�:�f"�������d|$M�Ε*+`!�l�ji.�����]��l.%N�\(쟴����$�,�;�����ӣ ���㧙0)�!�5�`�VsF�L��Kg��+ҕ�MK}9��{���>�r%��i��ŪL� �bc�A:�9Y�K@ e�/Æ��������ᅍ�'�47^,R�+��r����eE�v�&�u�c�ހ����%�$!�>�*�G����F{�ש�f|��b1��{AI7Ў8�N�u��r�Y@5�r�h:���Ύ*j;XW�:�j7��Ki3�S/��+�Z���OR����jc�mmV�P�ʑ0ag*�aO.��nyDTR�L{��9�̠.L�u?���w7�Y��D6G�h��&�	�_:�8�B4}�9��%����Ue��xCo����<b�D�[l� ^�8I�v��Z��RW���CV��O�ʕ	Pm;��*f�~+���W���Gl��������3_HMo&_G0�Jٟ"r�/bS�vV?�zxz���`Q��ɷ=���/����~��:_��kb|'�?���qu��MP�O�&{���>�I�Z�Ț~� Z!�׵��p�Ε���r���A����y2��?����k�+V7�6���_��/��ww}z%��\��;��I��rC�+�W�ydH0����p@���C!�֦�@�_T�?,6(��*���	oF�l���G��3|��:���y�FV{G���.�W��r��h�8Q���g��/�V��'���c9�g�m>4��N
I"�g�A%���7���%��э�������K�)}���[�`.��P�Ci$GFx�2=r�b�竗�'p�w���덣 r9�aT�|[���k?�;>�K2�d���#3�YFU��J��7{��C�� ;�� �P����N�Àa���#�A���JM��!O.��t )&����_2��JS�:�m{��*.w:`��kW�8�7�hP�$��Ƹ�m�� ���ݾaEfİ̀G+��6hemal�cPIi|ʗmP��n?	�BƄ���(��)��
���&��#�rC443IS։HGG]��0��%�L"Z�`���+V5G��
0!s�`�������zǁ�a�k69�"'L�� ��	��y�Z�τC��߅A�U4(]�#����~@.lrĨ9���c��Cyڰ:���F^��W��;�X�e§Qo��KHlA:ڪ(�2Z(pd(˾\�����]�gBں��A�\�XIo��+�쏗��uKF�ޅ� ���z-WFm�0���Ȕ��.Y��\�ȡ,�l�OyT^����E���b�y v�Q�8�N�G|�������x�s�,���'!^�`�A^��ړ����K_I���n��P�Wis�.7�l��5i��Jl�ŅfnH�P1�c׹�?��:7!+<}�7J�8�Ӥ�l��ݕ�ƫ�xq�6qߺҏ�>z�54� \�z��:d��M[n�.����l8�&���t^�*cmݴ�H�Nd��/r�����O  @ IDAT�p�x�'�C�ݲ'��~�g����s��E_�z�/#e�E��>�]R�~�JV[�O˺=AKZ��cu����io�cV�#����>���oL�g?���d��%�����_|O�=���r}��!d�>D��
K�]�_�/�؝~����	�q梍[���D9G�<F��;�c@�q��ܣ��苲��@��ĸ��څ�U� �3���`���mup�9����͖Y��¬L�,��x�8:=�@:G�U�*7��Hӟ���/O����z�7J�U���VZu0�>c�ɪ`��+��c�+6㥺��#v�]�{\N����s9Ox�����y�������/p��q��CA��/�º�n�	�!�1�%���q��������\g"e�`UC��C6"���'l�i_�q�J�N���u�ȑ_��,��|�`{e�s�r�z�T��H�>��Șc&���K�6�<���u�������;8���G���8�Y�3v���c�D�,D4aS t֢��P��|3��"泚7y�B�t�v���X�XѾm�/�*C�	'������J�(NƂ�r�Ib����{)���`�-(v��+J/�����y��"�c����ɍ���BT	�=����J'�9Y�4���:Gm�L��'6�Z\e��&hV�DD*���PQ������*�Hشp�ɾ���b$�E����z���V��h��������1��I����5��N��[Z�i���iu�v1-=�(te�>����"s�bd�<�[�4�v���"m��y�9��R��f���!��[����,�����\���E�?�W�����n�y���9�:����r���[L���[n�x"=�;����+��
��N�"�:�&�Y��=|�\5�e�ON�ù��b�J�^�Ѯ:~?��嗬t��|I�
%����g�U�?�W�� ��ȣAoT�Ǉ!�^�aCG۬��LGv���#�99Z&:��[��&I�K�7�O����>��}���W����ot���΢���cV����>��0��;G ���J�z"�-e�2��`2���?��f�������/���O,}�S�c\���ͩ�����(g'����s���eK��O��|N!�C��>���?�B��پ�3�����G����8^<r�+�z��oQt䌸���.�=^5؊+h�QvO�Y ����7��ҶS�MF��=X���6VZ����ڱ�H}=�����^�3�|�O�����+��\�K�s��!LG^;��2�b܇���b�q�A�\�pl��#�۠?b��/��s>�yޒ����6y1C+;�wK���SDQ�	�O�H����ᤧ̾��!&��aV������=�q��{u|G����3]ϰ�+a~�D��Y�S.�.��\e◧�B��g���Ѣ��xN�0�​2�����?c���8�N����*J.~���jܬvev���<���I�B�"FU�$6���,{�w�Co����N����tp�8�e^D(_�4N_X�lыlV~��T���� �pL����RC/Z?�L�S�����R!}�Ȑ^�� f�����x�(J�3�Vx��T����^�������T��;rV^%s������
?���4+�꿩���J��)�T7�3h�����j��QC�J䵥8慁L�eY�����(�:�r�*&/�<7��������=DW�$ԋ?��R�E/&.�Ȧ|V�	� ���D_�'X^�MMy˖F�p?�T�%b0?�#���f�N��4�V�͒��a�f[��]���t�!��5NOz*m"]-�=i��4�j�]�?v�6�v���&�n5Q��77�̳�Z���z�y������>�4�k���]$��/5<&�&��=�+�w���g�y�G}>u0���Mo���c�زr.�rmվ6b������FK糛�}�h�s�K�u��g17�\�t �Z���1�`���o�d`�.�"�[,�Q>ڧ��9a��Zu�*�P�Ĕ8_����_�:�����ax?g�=_��q���v#?��H�RH_/1sK:��JE�u������U(�l�"�r�0�S�M����yMէ�z�-]TR9�����8ay��+_��"C B��ɧ���c�W^���=ek`s���(Q��)-���	'��Y�«��flC+M/��	KxOp�>�Y�����������I�Cm�32&��3C��� F>����0l|���˗O�+�n�P����,ϧ?��L��9�_�5w~���?�JaO��n	oP�ҡ�!5�QL�lM�Y+e�L�Ty�~:��
����oⱺĲ��)����O�r�?���矝������ς<���׼����/����#�������f ����E���wQ�ځ<��H׻�|w�
��5�]�g��jtB�!�v�ji�Y �ʝs+6o�mL�aܴ�-4�m�݉{J2�aw�~�Cʜ���-$+��=Bg��!s`�C+��-]�إ���>�#Y-Z�R	گ��z��o��ɗ"��?c�@�5���P<r��v�*��b.�SW��
#��h%�Z1JHaC���o��r��5�A"]}D (�v��y�#e��Ʌ
U�F�j�*O)�-��GlE�0Ql�u(|�ʖ��|_1�+)��j�u��y�8�9_�Gi�>�GG!P�/Ћum%,�(�vI�/��h%�f�ʤ��X��X���X@1�ܷ��F� '���|W^�����s�rð��ؼ�.1&�)cNz�>�<�6�47x4j�#we��x�l�J�����x]�(�u
����9�s,��+]a��s6[9����Lۧ��jP�/���E��|�<��3n�q\��=��/.�%<���+j\���}�-��_/�'lF��ض2�#."�m`sV)lw	���*W��k�Ӑ<#���7�>������={V�>�M��鲼*������Cu��÷6�6!�M�ӈ�\���"g�A4��C�}"���%쇬~��2~�>0�>��k�"��:oe���ў�3�D�yK��V�F�p�Pz?� H9�Y��+_I�ʨ/��9�l���n\�X�+F�ȫTi+�����4@	�=2"��^3�j��ý�c^�����;��P�D��H`o|~�3ޏ?��e܏�e�҄.�"Tn�g�"�R��#O�S�D�U�����+>X�;W�X	�+M���WZ������_���������K��н`.����n�!�ΖSe�\�$�0"���h�/��+.�^s���_���şO��o�����<�#6 �b���-�|��~�&��1x�+�c�<��ZF)z�i��lV��0�L��uvN0E��ؖ"���ˎF,�Û2��L*�,VZy��N3�w��2o�=��NO�Y2�u�8���ge�lX1*;��B����	�;n���#W.��u�G�NRh./�L���*�-);A�WO���M��\zA]��\�����.�0iyt��	�pM�$�H�9Ma)U6������)e�4!R��CL�\Cڅr���tn�/8� ���1�<�?R$,�l���Wk/���
�i��HGf�I���g ��2Aw��QohP>X̪�9V"W��[�z�%>�ml�T`�l�dN�k�m`C�i�8>ș�� Q-��ks�7o?��N��/
�j����	�G�9vEE[�o��I�ٙ�:�'�7A�U�8Hض6�	M%�OXW0�� #D��x�aM�⣻�K?��L�nVx?m@��z��t���k,f��_H�?���'�)�v���O��_�W��0����t�"�ݮ!r"����a��2��/!q�.묮=h��ʕs9�{}������ԅ�G:���2k���9ֵ(S���ͩ\s4�ȦB0��P��7�-¥$/�,^8����{��=�%����k���|��c�"=�+]3CI���M+ 
��Y^	���[w�-=L9�R��{�r� c?M�׿�Q4�#G��w0�+�s�a�t(Q0�U��'�Ӑ[��l�!%�a �{u�/٤����cx�2�@���%fz�~'��/7���X�NFq2�+ɋ�õҵYX酒�(���m�w4����+�U���q }[.����_�����������l�g��_C=�hr�� �X��&�E��ɤΔ0�^�|��K���c�;>W󻯾:��8}��/���5����	��|w[<��R��(̤�HU�cG���d�)r�P�4�����E���`[�a�gLq��Y$�鯙��IYi��iA��DM��`a�?ԛ>��Ҫ���� ��Vf�d	�=iy�\�K/X�v��B�Z+�#i��f�Mn;�Ef3��uF���<�E�{�������e�a�bx	�Jf��r�x;	9�ڧ�����CZ��AR� �O�̓g�\WũX �xhI�2i���&Gm9Y�ŉԡ���7�l��K�ȕ|J�SMaI2jU��PJ��N]��RH
��
��mŃ�W�eĥe�X<I��$eړi�8↛�Pg���G\s�t�Oh�O�fN� G�q��X6�����8��2�b1���lЩJ��U�Y�fT�T�m:��.�G}���[~����܇�b��#^����_j�l]�ؠ����?�����t"�/�\'�K���Ψ׹�n`��S��N:x\��8��0�)}�Fye��s����-�cê8�!䐳�u�}-I>�.��>����nEDf�1�]}����Rk"
�_yml���g�Xhe#@���+[X}|��k���w[}�{������B���=��Зi����CW��!Đ�&�%S�W^�̧q�HV�^��i�m�	��(>��̇������M�\������Gyqh��G�]V��$2k�ȩ�?F����}�t�떨G�"y�����C�u���׻�����V�[��S���'�>;eҠ�z��UX� �,*8N1�8`�WéJ�.���4��V�������	�/��+�na�|��\Ȭ|�*R1V���^����Q�~��דe�`?n{�`����~�3�G��',Y�����r�:�$m�H0���=\G0�?;6�����6N����/?��W���W|�n_���o����2��s<�#� �3�Kw��"�ҕoқ�KEfO��e�9��	�O8	�E�;@��e�L�pl7bes�2�L�\(�L�������
���Ea�������ZK�l�[g.l�5x��'�C�ǊR��d3��>�>鷱v�#&>��I�#6P@لq�d&e'���L��-8z�?�u_���k���!��\4�7��� �?5��Es�����RVǣ��X:����=,=�&%k�Y*��F�-Y'��$ILڄ��B�XZ+kO�t�W�LURl�5� ��o(n)�����[�ށ_mkF�8y�&�^\J`�c`kc��0G�Ί@%k? C	�m����
	�R�� �S~V6�>�� h�	��ɩZcI����rk���<������F���pa�����˽�I#Py��)�D�S�	�KJq��S=�z4�xݿ�-���=�ok?�&��d�/�5-j�sBA^�Ͳ�׀[�h�ZypI���M����q��'������ب�cڿY����)UW�I�v�H�w��ȧl@�.�W܌kK_�p�u]th�(��:~u�GS�j����}c�'-����k;�8;�Ď�iUd4%֢D�M���YiS�|��o���4�+:]KF�a��0���<&?�T*��{�$[}[����M�3򩇛�9��m�\�0�~�I˯�]����0�
����.��-��l��,��y�~+Q��f�#VX�E�DK'x�FE�g�:��1�qU��g�1���P��$�G�5��%M*s�@��a�T���f-��0	�m�yΟ5��7�#e&����P�GC�:_"�
�����dH�ps�"�֨���x������ϳ]־�7���Vq�_�������o�yG�K�o9��0�8�� ڙ	K��6�	oufm�$�t0�;�"v��j�#�4v����Dm�B�!�d�L�w�='���+�s�C�P U���l)(�̿�tz�ir�D��z!Ϣ��7F��uJ���M�T8Pm�Ka/��K��G?�>�w�[Φ��ǖ���@3&�@H�]��:#��GS�	��%�u�LU���"���j?5?�2E�"�b!��u�WP%�<�!�3<����S���v�(s��ŋ�"���M�x����cڶ!X+� I����V�G��x8����X�� �U�j:EB@�)%�v�S#>m��<iZ�Y�}�q�C���;�F\���r7?pk�4��>Yp�*f��+�iG=���T�bVW2ns�����>��d��{��3�JCeS�r����Θ��*��i ��]eI[��ہ��k�����.�[�'v��&�z�{�|�H�X�p��3�!�=��]E��e��c��G)��ʬ��~K���#�3�{�n�g�]�'�@��Q-�=�K3�JM ~���r���*�C�~�$N��ƹ�)���ߛ?��M�0��}�͹�jO?؞o���5���,䍓�82VFΎQ�$��Y�A =��W\a��{lv����W��5���~�д8�6����x�,���mWx�|u��]ڥ�W��w�-_0ȵV�v�ssr�d��!y,�!�6����~ k#X�ښ�VS0��{�T��.ʞ	;�v����RF"H6�H��i���V�&��Z�#1�
5j�M��tD�	ӡ��T����WQ��kc�;֙9�*��V��v����b9�L�u����_c��f�<�'��h+�S�\�a�YM���N�@���t\˜Ǚ��i�8^�c+ڭ�8S:Н�x���|�C��mI�P�����4{�%^�[�QQB���A��V��<�|�lݘ�0YIK`N�M���Vj��0'�B$��t��[o�{x�El'�5�YM�,+ג-2X	��9x����c$m'���8TC�S��b)1�G��c����FJ<&���o&��ߔ�[�.8�"�0Q%����u�J$f��X2��@�-k���o��m��OX����h� f��qS����BÊZ��!l�	0���� �"�J�V���bZ�lpȧ[�XOB���uӶ���eR�O�\�9w�0��*c@���He]�ԉ?W��������2��D�����-�M�ǋ4�c�9oB���x'�����]JT#���ٕ�Ę�� pnl��Յ����~�~��'����S�i�n���_�P��q��r�����h�xF��z\o��Q7�~q�"����<�j�1y�l��%��ZP�ro��e�?{uz�':7�q���������x�b��#+Y�z�3�CX����7qƟ�xC���F�&�8E�̢�+s>~\y�G�4dE)�t���'����#U��I��z�{S�J3*���8�5�z�fa�+�MyZ�Ǣ˿�Q*��&L��oG���`X�DCC�{��p��@�_ �r�,���q�˅ӆ���˨�~�F*⌤�sN1d��T�,~���va����pi����w�3h|A&��g�_@:P�$e�y��簷	<�kC(�:���*"��B�����N���~z�#�?��4_��G|������N���<�ƶ�|�v�Ǎ�&�E���@�RA�ڽ�:ˁЙ\��R��\�����Q�i�N�gP/��C��#��ӶO�(g�!�J�,���2�	��R�� +�+������vi��,EJ�sb�:b敽z���sn���e���.{��1-:y�-��8(p� y	'�y��M���*��	qm�HY~5,��a�ߐ�Cyn������=B��(Q�+OV@�����j]Dp��)��K�E���T�8�-NI+պ.�Si�`꣋�(p����2�v�*�Ƅp����BR@ dI��;c�vi_2�amS���)�bW|qj3p�6��	����aX��U^U��V�3�,ٶ��B��,/L$�u��Y��K�#���͉�[��G�M�Z�	���G������q5R��iL&:��3e6>껒�=b\̽��Y^�� ^'V���(o��0i?a��`�~H��ֱ�xK���^��d��_���)_����FqPm)WO�_��c���aV� M�6]�%�x
�>e�8��}�'px�?|ci+�O�����xC�����K<�H^s�}���00�'���1���8�����G���M��/}&������yA{k��i�qd�uƐ�2_h��,� ��/�e�{�z�a�+ӝ���"qQZj�o���i������� �~�Nc�/b}����.���{�`�I�K��C8�*b�X�p�eŬѕ8�O�a�$A�X"e�~�t
�Y�u
)`F�h��Ph9�vR�������x5jZ�H�����L���]#����Ggn�����\8B4�]��	����j���u*�.!�����`x���ד�>=}�����n↥d�r��/� 9_�a�e�g�f`'�����GǖG���f�K�7���@2��H����3 L�<��F,tB�͎���ShPMIHW,9I�rl�]r��QX#�f��(;L(-.�C��:�BnQ+�PY�/�#���>`^����\9hǤ�o���5����L���`SV�\��no8�lr���1B�k�סS\���waRn��q��#�X+ �ڤ/�����G�2��bŔ�/l�V��B���mBG��%���K���س�'t�=��5��¬ �8aSиv.v~��$Bf�rTV@�0��-�U�Ė��ڭeI���~֟��?P�!�^�T��-�
ۨ�S�/���zq'�R�k�|j�B�U��>�)o��XKޓ��EJ[pHg!�����`S�x��a�d�g���'��~�x�2�W��o2/��E�Y�S�����n�Fb$(��3�i��0�g#<H�ڄ�QO�7����e����3�e����`V���I$��/��{�P�.� �0"ٶ���ڞH(�>d�����ig^��x�ёD�+��jy�m��v�_?�+�/��mĲ��c�mH����`�t�݉�IZ��FVEN����袽��|��u�F���!�:2OqV�)k��H�	��B�������kkۂ�\#���QER�#��U��/�E'�YVl�]yD�I� �J��9$)ƈ6��Q]Cp�hpU�8���������S`�Q|�^�Ã�q�xg3�v�@
�*�.E+���G�~��x_>�>����rBC���7t_���v�9����m��X�#�������?��!d���_�C~���r��Y:�W��^�|�=���-t�GW��gƦ��S�"_�Is�1(�g�n#-�����ʿ�Ib�Ħ�QLk��ʓڅk�� %��Ng��-(�=�f�o����9���H29NpX4�$-~�����8���X�**���S,����}���I���&�)�ALV1�j�M�����N�o�z��J4Cgii���D1�֦x�N�j�F��	��0�!e�+cSѿ2�e�E�p.
M��=���R��EUꝜ�'�]�u�Z�
k��/t+H����_��/�X�#y��җ�!�"�Bbc�,ik���6�� ���6�G��D��U喓�1��U�Y1̜�8�|����[��8�!"�8Ҹf� .N���xU�RY$���8ߋ@[�fn{���YM������J$#\2���p��e�W��G
ƌv�:��FGϠ��F����)Y[���#��ί)Iw ���>�ݐҸ��{�y��..Y���v?�w���Y�)�`�qL��k\�7+���E,�'�L�"|�1_���ؖ�፺���d�Dz��u�Ix��.=t(�!�/&�|##y-r������8K��ʧc�e���dB�z���ܸ�/:Ҭ�{�g���eb�+#����N�﫤,t9Ƕ�A�YE�8a0r\���`A{�MI��F�\y*w�&dյU�6����tB^ʋ�*v��<j�@�`�7���]��&�3�}l'���Ȍ��~�O�N���SI1<�tYJ�<���O`x�B6A�D�Vw`ٛ�0�^gV$�Rd���i���x�|��r��e�w.{��N�QeY'�C�k��0��yg,�*����x	�NX��3��A7U��V:��4/ �� 6c	xΝd�iI��o���MN��FI��I�б�L�!��Tӭ��v��'��
��hlp�[��)���L�U����^��Q��&D9���y/*�c�MS;BF6e�K�y	/l*�:�-���g�/K(�V{NYN��V�chYJ
��B`ŕ��H���
�t*����Z�&Y�R`��w�*�8�K���$G�bWz{�)�b�����2u*��0��~�>��\]��0��8clF�#���~�U�=��eY9�]hU��Ҿ`~�It����c������WpCqN��%��6�����F�g�Gr�r�!3aJC�A�yS'L92�f�t�
��ط\��.s0s�+��嗊����sK��Ż)�ȫ�r�xy(�����, )W?���t����P��u���3*��\b��'��r���ǃدh�ۘ�%�����`#�Hm�8��K,���_�ꔸ0(}	)��N�E����� I�~��(�s�T�a](י��`�"[c��s�Rze�b�ѧז��-�I�~����! ^�Y�cm�,�lmy�OrE��$�
���)^,fbaZ��� �F�Q�կ�&��Y�͵0.��N $i���&�(K��9`{QS��/�/�q9#�΅/�se떲��a\����f}���+sǃ��U���_AL��[���Z&F�+b����lhȥ�:"vT���\n�᭳?�WS��^�!�QX6��yp�]fc��4�����G����8�#��C�u��`{?���gy�}���e�x�#�	nq�⌁�{�0��#2��FH8�S��q"-^��<�[+��R���6�����02�'���0�e2*9�)u�����Y�����1���I�U!ek����+|�aC&!��@a�N�#r0 ��q��d���g=��8�!4��`l֠��-"e2��@���F� ��VQ�%��L�drs��Y'�%�8����WJ�;u���:���$-���V���S8K�+�^���¢��Y�a���S:�k�j�K`�'�Vy0Rف��8���C#7Z�k�M�0�t���4#i�� I�a�1_������+�w��o['Iy�e:�%�(��1ds�#_�-�ĕ�B	��<�I*��#|1-V���#	j�P�s������ǒ\�!�
��ٸ�)]�H��1�I׶2����4!e���ӫR��c��6�MVy4�qI��a_q^u����V�(!}ȄAG���w��
�A�]�:u��^���e���B*t�5rV���:)U/_��/�����b��=<K��yU����`�+_�;��K%�-4���SV�%���{��&˙ǔ�y�J O~U�����ol��s�|�Y�4���f���c�$:���Ȳ�TC�uOPdz��� �@�W��;{h��a�P���'��C.ܑJ�"u歡Ja8T�]����<�|���l�T�
?xS�Rb���>��3_#�Z|�l�@Sno��PB�<'���d5�F�0!A0o(j���^P��+G�A�r���;���y�/'�Q0�8��c�=�)�	t���L���6���t���q�d�c�)�A�2+�wO����ݴ�.���M�B���ҕM�������d�¦�X�۹6޲��*{-\�'q�끹�|�dj���*s��@!�ӆ��k�v*��]������i���ShHG9� ӌ������F���� 3��L�RD_���FBq���]�O�V)C✂���`�W�R�S˒.�4�舗`�]zȻ��-�@�x�D�F�i��P�{^���Hk�ܴX"H�$W@������z#���v��Y�RS�#R0#���n�&��`���b:�ԉ���Sfb�)��n�aU%���ΒE��%�X��T4R�x/�Z$�p(ʴKs���(ٽ�Z�R���S���Lj�_QV�A}�wiE�:H$-_#�4�9�pl�n�Q�$��(X�a���0�Tu�f>�dQl�N/��N���N��
����ɴ��L:>��B��8v�-��p��%n^�
���J�*�#o���:#%b0�Ϋ�t�'u��B�>�.ļx�'�Y�;~0������?z�E�7YQ�	T& ��qH&Zɂj�Px�CkWe�n@�<ؑG��n�|}4�D�K��K�}�J��F��ӱ��N�ѕ~���Җ��۶�=��w%��U+�z��/�U��稬��,UA3��ϸ& W��5�AĆ���
��ԣ*ъ-�gE��l��_��AP󮄱9�z�】�b��AV���sV�Q�҈��`�Pƽ�PVu�lv�:4��m�X3O���*7}��RUj]~�	n�bB���6>�@3FWpv�3��Z�M�2�@�x�@^q"̊YyR�-��SvL
�X�M�aO�!��;�8�c����q��2�h�)�TV��n�!��l�I��|�g+a��56P�PY��#,�i�g{Er���H#eH���o�)P�%�~p��Sk�e�(��RNb�ih-�!\�{n�1��[aFF�nZY1� &��5\�'Tsͦl2��
�x�N��=��Zm���f�pL����0��?r-�R�r b�����v7�&��d�S�sQ6ͯ{�����M�J�<�W�,��z���E���%fV!�DD#���m6Pae:�,�Ԗ����Yn�˘�(��Y=�ˮ��We=�Vy��2t�(��,�u�I	c�K���L��6�i_5U��1$:?L��D��&&	U�pm�r)����'5���A(Gi4L���F -��w�9�y=��:c�k:'�f��\g�=q���gO����Q��/&ܾ�|�ggU>����@��oY�PpHnT�<�FA,���Z�"34�����{��kXD�sʕ�]%���
�0�� lgv��F8�����;65V����n���b�.L'�/! @忎��359����"�����Ag�����/D�IH�&�9���5��2
9�b�-��@s�O�W���ء����D�qg�o{I�ʍ���LC����Gxgv��� �f-�,h-!���0W�N�r��$���f���1���5�Yq͇Xt�@�	���7LZ�cX2Ď3���`��x�bJ �UXm�Z��2[N0N��I�B�!R��C}���Mq���Bb���L��@^$��m�i$���2leK���S��4��{��W(��i�iVh�M0rO�xS����ت�_� ��6�Ej�w�٧/�%S:�0�C�xqI��Km�/�^䏔ϫ��!���Z��8g��/�i��b�5i|!S�d����M��N�6.��Aӄ�b�l��'K~���Ʈ���޴y!���sS�QuIG.��K�!�`N\o�/��r�d�M�|Jq�������G�Ny�²������֚�ta7����Zq�g��5�-�����F�>����ߌ��ȳd�t�قKSإ�'�d�7G[���`�4ȍ떲��н�`k����_T���s>����S?T~�V����=�yvz���q�x��rPf�6�P3�����`4n��*{c)���/6�	EA�c�_�{]�<iW� ৫�{�>�W>s�&+L��n�Y����S���7�QzdzE�lD�!�jmq�I�����t˽�2�.�FT�x�Z���E-DdP�R;�[��pK��:i�qV��Ug���靼4t���c�}���^�,jq�Fg�Cuc�Ѓ���9�=ҕ�h�5g�`�D9<�/`�a���+�od���R���ITV ��ף<�O�!�hP��I]P�yg�V��%�v���Y�Z/�*�(����\��\z��6��m)Ru_�0�Y^�������v�/٦b�4Z�&�`�ca�6���
D�D��F�\Tc�e�2tZ0�G�M���G|���*�������$�;��L��6x�[&U���Mȟ *��;�}4��[gz`&>�aT�J�>����+&Xv0�&+[%-+]�y`P�B�ca$:�>:Ya�xqdaz��-���R��k�@�=|h� `�Z�8'2�[<2�N���o�SqO\�N��k�7u��؄��xK|;�-B��
��c��l��G��B��R-��0
Z�!ⵕ
�e/Z+��Vd�l�\�� 
#�T�Դ��TP)�-C���/Dj"�'ߙ���7��c�����������)_�q��5�O/�f�?`�W��������H0b���W��q�R@�bɖ��R�rme���4�,
�T�8=�������V�J}`�/��B�{����c$G���&Z�ڐ%����'J����s��uEk��P!m61)sбq�]3�Ҝi�Ͳ����j�!\S�q�c�������(�q&%�Ik��n�\��]�z�:R��������p��|�xߘ�N:(�@�6Jc�b̑���RQ9�d��:|i,͡m4���MV������ԉ"@��n%�=��%F�m���m�lx�[R�2�"������n4&q��O���>qUh��ӎg8d��6ٵ�����J~�Y�oGi?q�3؇8�>m�Ʊ85�6��Z2m����ƣ�u-YT5��.�]�N�2��7��v��j��L���Yf�9��g����,92O�e~�J<}fhLl����Q�~ܖ��~�^A�󶒠��B�=7�r�A��}I�AW��a�����0[:�M���j�zrD̸^*���cxO��tb�)��;__�e��t��v������l���6h�D�R�M��o��Δ��#�Вu�+Mf
J����\GR�	�BZ���_�8�)^r֣�9�k��鮲��5Tۺu�X ,t�����2�!��xs����}����O�4���ĩ�c�g����ї��1��)4QI{�wNn��6K���JêY�rK�okp�E�g� ���)^�Qaq�q��B��`������x:�����@�"Hf�P0#���8+�ƫ.Jz;B�e4�so0f�aئ�8 ��z�:8.Q���<�H*���I��0m��'�-XZ��2�#a���/״�#�������?s�`�ԟf勸�xKq뤕lq�����g�Qި���%D�Bu;J��=�m�����=��F�����ơ#�BN4e�@qV�X���GT�	Xk��*v�M�P\��\����:�042H�O��G�.ف��X��.�C�c�$�c�z��H)�:"3�;�0Ғt�GleY��rЃ(�t��2��u��.0b1�JL���IO|�$G�c��/NY`?� `#�D��#ސXMt?�;J��Q>A/��3�3�� ��,���X�c�c��޹2}��f#�_�Ba#y���#�IO�y��C��{�������my�ns䱗��_���:������S`���������M�/%�<J��K����2�?.�cU����%y2�3/�׊�v����pi���!H����H%�\�5��^C鏾�e�H�
���+�7�p��<��˾0�˿}w���oy�'y��J�<�{�÷�|uz�7��RP�]QB�<�#+��&�P�G���Z��ʌ:�<��_�}��@_<[{����s�+�u聪M�y���>��5��#�U���CVd�e�H֤�NR�p
CU�H��x��f�XX%�Y=I��p��$_�bQ�J`Hc�v;h�Pк�Jg�%<d&(���v���@�B��e��M�����o���Η�ݾd�2��8����g����O�?���yyŧ��ݾJ�����4���/��J��C��z8��V����kSn,���_'5%��q�(MX|C? �vж�p��x�4��5�9/���@"I��	=�K�~j}�cKs���> vr(��{��r�����P�?ۿ6��I��0��dH�{,��%�X�$��w��݅�.�<� ]îk�'<�&�v�� �!%�NhYF�=�������X�e�  @ IDAT(�qdT����و�U�t?����<�;���?|�{�X�#�U?�&;��oʏ��N�m�/_Bh�-zK���Q.�̧l�<��ŉ<�[?8�e�>h��d�����f��R`��8����LjH%��u���`]�bc�69����G�st���H�RԩSde��pTC<��)�>�q%9J8��f�hYp�ڲmS&غv���ʥl�F��(<K��Z:���Ʈ�y	��w���O�L�ĈG�����/__��+��~�����;}���N^�&_r�*��|�tyS�+6������\�޳ų�]mi���Y	f��Uvev&Ε�Cq]ɺÑ����(C��]ĕ���[��B��׼��߅v�F�8r�oНoa���8b:a�+G�,#i 8oaIi��+�_���Q�u�"U5T)�Q�(��n�Ǽ��y-�oY�s��eXŋ�^��Q�ⴹ�񁛆-g�vlu4��j�)��B�Y�������'?W����oO���8��aYT�h����_A�B>�����f`�2a9|�L��uT�Q�0��w� �7�Wʑ[ٽ��Nqt�R����[��4K���t*��6{��H��6�����ᑘ��_bN�����྿�˙��g�7Z�b.���,��m���s��6�����.N�b'�c����͛m�p�ZmR��=�u��1�p{��P�Nد����R�#[ ���J���):XޢJ��qL]�k������o�;]�(}�őH��C~�AV��:�?a����� ��oQ�:�iiOV:��eT��?��S$i�h栖P5�Y����`�x�Cp�\�ߙ�o��N�Lت�2�^ ,���A�8z�U�#3�K�pl��A{M\jf��)n�B�	{�H�.�p�t3w0�U��ɁM!Nq�x��5�7���ʜC��_�B��V�*&�<]=�.��ɛ���.�:a<�c��+���X�z͵�U"����O������_��u}�����7�����7��__ް/�k�Û'�;���xX�AO�c�_m�X��f)� [�#sV�X�z�cFc^�����[�v�x=�u���T>%�����-�����7,4���$���O��C�0�q�X�j��R��	Z��8a3���4�v�:a����T|����tw��C�^���T����Wt�T��#\�I��mB�e�>�;<���\r�b(
A�	��X4:墀�8_>�u�S�����;I~ǳ�?����?������;=�����x�f	��Qܡ�߲�ӝ�'FyK���'{������v�ԥ9�F~T$U�v��/0�C��'�;`*GPd�j��3[.!�ٌ'����V��ua�����
�e���s��'Ζe<��~�MeQw��5y+������7-v@6B�U�W�Om�i�S�. Ǯ��LnG="0�%"Y�΁kE�Ji����W�1��(VÖ�ȏ��AJ|(_��ŷ����{o�4�%�3����I����\H��:0�g��3���HGrCcb�&ؚ�^�e�Әi��&���%����6> r${�q��8��-�GZoUN���-���Q�����>z�g��w�M{r^<έr�`၍��wv� ��2oU���5qz�Ħt�$5��l$�@!tp���hX���1��4�!���y�^��EN��s}�&����*:a�h9��a�J�7ߟ�����o\c?�����݀��)�]��	��0�p��ӹ�Z�Wbb+y,ybs�۽QZ��� 2O� �S0�_@�Ֆ�|A�=�*�'M������\)��=nW��^���ن%�W8a>1���͛�H�V���Z�0@�p����d����ڌL��th�[�Ch��8�G *�ڀ����}�o~E�2}Ń�
.{��z-������lR���L�N̦���D�k��G~6�s>�������~����߰�͂�����������G߄��i��e��"���`�"�LHBI-ఓb�d[0�-�:'j: ���_�h������[V�_�$�R] ��&/x[0)J�$����v�N2�e/lw�O�:��K���`�K^���G��K�RfE�V(��jTo��U�'���a�D6�e(^y8�w�7:��%2#�eʲ��r��	��/,��_LP�,��?A�ަ��I���8o��["��m�}�S�s/�*<�ߡl�1e#��Ǻ�}Yw��;uq�+���#����䅹ܛy�9�eGڗu����^��v�����>�M���0��G�[��^X���j��oa�m� �H��#���m��@�~Sl��,ի^j{(�]_/ˆ�^)s{�p���"!8ɓ�k��Ԅ���ܕ�M��*Ѿ��G����o�>=}��7��>~r��g<]�Q��ʅM�>n��1���oNO�؜�j�~|z���|d�mA^�	�t��\y�\�s��%�{��y�.���
�;������XRZ�J-��3����/<���1�+����.DA�
�_ᑏ$�i8t���Sۃ��WdŶ#��a���Udk,M�tf�KO/��kV����J��ŋ5�G��9��p�!�c�|��#�w�+��r (%8:������47`�p��E���Ek.5�SS�A�3\��~������ߝ~��?��������eϫ���?�G� �U�v�[��^젷��m,e����T{�S�XZƊk7O�
>�`9Z�Y�N�)�48��m�X "l�����Kj�9����������[��8�=��,Z��I�m=.;J*}xWə(m�h38�:m�@,�b��%}<�L����nL'��-���䱸%�>v1��d�<е�@{ $~(�Y^�{B)�{��SE�u&e�%��o�L;�?�Sj,����z�S���K�Z�X
�j���9���&�x�h�J^ʣ�����IO<��Ҷ3)����CJe�.<lp�5����,����VC��2#{Id�������}��e���G�	D��M�O�!���
�]�1�Qӱ���NGJd�ټ�rw	�H�Sw���	/*/�nm��E���_����V������L�+8����
������0+��ќ?$ˏ�^�p�S���ԧP��}��������W/��>��%�(�ľ��J���6������y���N�>�r48�n�ޤ�~��o�޿d��%N��B>��mA:d��1oo���s���2��~!������K���O􀅨�k|��|��]ˊ����%���Q4\��
��H�������{;��V�	�pj��'HY~�	 ����t
I�[��Q�e|\��'x�,�ad1�3%��?��O��R#�,!Vvxied��F�h��~�)�?5�����2������������/_~�Q��{�C�>��eX�>�,�
�-+_��K����!5 ^�Mg7��˦�,\k�d��kf_��rA,�V����3M������T���'F�s��-��L,S�|}�2v�i����*�
Z}�W��c2�*�v�ŏ�΄���`g�8ȼ���y)<8cK���z�<q)�`� ��Y��DkG���|�ٲ��ԅށ�.�2Ӌ��_i렸<��4L'������_������ļAR�#ȅ��J8�{��ty�|UoQ�OzN?1�K�� ��S^�Q�.:�7?�}��-��a�1��?����Paٔ�����{m�0��]{�!���f;�����'#M�9ɷrSzO��c�ipJ[gي����'�x��e|D�t��(ee������Hm����>�E��U6�l��P^ɤ��
�<Is���L��8���˴������� �kex�˂��Z���C���_`]\�n�Sg�Mw>�"�E��o�w���|�5����x����>=����>�5�v0"W����C6��}�5>�׺f�a>H���3������ώ}��?���)]�F.4����a��c��/��z�|��w廾��n�2/.��C[�c�*ƛO_�!�N��+v��׼�Ǔ�;�����#���- ��~��/W��C?�����_���K�=��eUGI�"!
m�#]&��"�/6޹��/!n�Ru�nX��y�1�~׳������y䌌8E~$1#�:�5�2���[�����tO��Wu�W�<z����t���_�����s~u�X��C�lV�x��'�8�������6�as�R��Ѧ���5�v�	D؄ؚ���1H[0m�[�7�ڎd��*�\��m�a��īB��@6+�^/�)V�B�%���X�)3� �d��+y�T�m��vx�h!�ӡN[���	4�v��: ꢷ,�7/ e�`��~�ޫڭ���֎+,���Ű��|���=d���"�j�%2A�"e�Z�������>Ń?�@V����V憟�	-n䘚��#m�
��	��r��76Ծ�^�z�M_ZGz�/�/䇈�m����uP-��->���S�Z��#�t�ָx��K ip�Αòv����
�s��S��(�t
��,;˟H'LG��~:*\�Sѫ_d�`լ�Ŭ^�Tlj��sp�ӆ9@�L�$��ٲa���V��iV�(��{B��c3�:?��"S�c懶��ڃ��[w�ٺ�(1���J��7����Ͼ8=���?���k��"�"ߒ m���P�5�5���ts����u�F�|T��n:]R�~�=�uq�Y%Ιp*�ў���,n1�b����#|i�����n�B5�w��ϰ�㓽+�G�����
����x��䀸��E^q��g��<�}{�G)_�����>�t_��W�*f�˔�&�@�6���`w8O�Y���8N����~xz���q�tĖ�ZE�	�y�*�+�+��{���;H��o����}χo�}�3� z���Q�����ߜ~����|�����}q�Y��8`l ��ro����;֊~�9�<4;�9m��&�]��	�JNZ�|�-�0v⤧���X�/�&�j*�&�r;�H�VҚ�R��*��i�t�� �Ge�x�_G�D����t�/1@��ұ�P��mz���Sl#��ot��/Y),|k�t����~��e�t-Q�Y"�&eT�^!�PD�T;� �ѷ�$���+�������c�e��(�5��I�h����X��J����R�����~*����$6˟��y�_@�r)���X��z��sʷΛʝ��wh�of+&]{��C@�#�)?������+s�2�������\�	Ȕ��m�&�����i���`H�@tPC����3�!�-I;3kbs�,y� 6��0k>�
$N���W<eȕ-�7���s�yN�+Fzj\��\���KV�|���4}�~�����W��Y�x���\s}䇿�/��隧a7<s�K���d�;�B�`eXb.�<@SP�(�E�h����ǵ�+	�_��yE	�t�,S9ü�@	(�:�)^�[�*�Û�~�#�W,P�y�
�X^� ��㡕z�6��L6�A�-��4��^���6,N��1�S�h�*]ޖl��"�_��0�<
�
Gǈ$�b~�ɏt>˦�7��灎��nm��e@_o����<~C�l�����W����ק_��������_���J���;�=`H_�������Vw�|��w[i5V%j�1��`����4����K�5��R'Co�ۧгS-0�;�de� �T��(�Y,A�����ȉKFz���KGڑg�\
W�.Fؠ9r�ݖ�%QE71�|Z(�To������cq���{z�7��Z���0��
Ȯ��jX̛P���:U���W�9�XU�P����l۬ܽ�*�з�e��@$ZĖ���T��Ps.j���&�m�����8ھ ��@E�A4����}���5q�䘖O��|d��Ė�{�
X�I�k��VI�ԍ�i��ky���u�;8+֞������n���[�d*BO�G���5�h������y`G�������<�3N��w$5�Qv��̫�J)�d���塼M�5E�SeH'Q����t��,}c�E���F=$<��Wqې�RWiM��R��:��Ѧ^z � ��<�����~��|�莺+���a��ő/�~z�������>���M�ON��S0V\ta���
��
��!��h��|e�9i���c��Ca-���8Ҫ�wi����\��K�5>��$I]��cN�ڕ��o�
M��p¢�P�Q6:���{��%��*�{����}�+��AB9�e��G�>e��)�)+N0�//��Y��T00(R*K�4kJ,��x�����3 o�k �Ig~�ͳ���}�_��Y�^�wA_��U��H:����+�^ ��i��ἸU�|����_|}�����8��o~�+��K�H}����}$d��w�������>~��M,_��������-DL�4�7�$�X��6�zL��`��<z��٩�׊v�I�v���a���G��s��e��L�t��"_:낊�2�v���aA(Q���ȳ�J2{?�ij�Q��Ioho��"���J�đ�ЎVp����JiQ�W���9!��)�]p�u�`Rng��䱘�N����� �3B��,2��ch��yD�# �0�� L�Չ���^���Ğ�T�R�"�w{����Sc8�6����\y'?qJGq�V���,X�^�XY��W���=U�+B�&��ꛪ�M?k�~�ʡ_JKU�=cQ������r�2�t�#�R�۪��{��R"�*#��Aώ)�W�U�ɤP�^�*�iƢxbS�ꚫ����f�\-���%]��ՑRvx�� ��p�8T�B�����\�����˱�k��cl墳�E?�{���ɢr�N2ׄ����a��/|��z�!m��F���&�ag�%�H^^MW��>z��)cb���@���۳�t�"����E�����[��7/x�����ߜ���7���_������~��G�'����G����y��՝���=�t�m��8<qL��ڋ4���f����U��5�����&�4���X�u�\�2<T'|W�ڻ?���՝Fq2�x��6߮�C��g������3c��ￋ#uC���H6��8��x{�%9�$=3�L�P����#��������ث%G���u�1����7u���DU�CZ����Y���5�=<\��{̓�:��uyp�j��cV�p�S�l� ���U	tθ�@�d�|�)@�{u�ߌ"��ŏc�k��~l�0�H~}��Kh�,�݀��|݄����s�=�d����7��������n�_n;����@�̷0>��W�g/���#��K�1V�\2���6;��㜰�q���9�Rjv��	R��<(��R�%hR�_�'���H�8��Fe�>	�R$�9�h�:������N�.�K�eG�N��ݲ����w�u���3�^��F����jQV����.g�ت^)�F���WiR�6v���*����X��P[��#�|�)�)��s��:�#HT��# �C���C��k8����6�����E��8���f`k�'`EJ�C��0݉���arC@;��X���_ͺ�q���]�ud/��A��őW{�����J���t��/}v�/[F��s��H:�;��^�������XXvA��̪�~����УUsaV^CN�vx���x�o��^摝P���i[�c�
>���"��A|4�ʶ�/G�^����0�v�E��4�&n&`A���Z��T��=u�h���o@�GR���zN�õ�oC~�n�w�{>�B���^��O?ݼy��2rK��}d���߱��?��6���� M�L���9.6E!�I2�(d��9�G��\�3i"&�	X?8˃���_ �1y��/���Zݽ`���K �"�w��|����۟��,�<�O?��	�go��,����~�x��$�>@���H����߼ň8a�黿z�1W4-��-9��2�1,�M��1����g�wk6i"E�����j�z �n��d���{��0�$�&k@t�� �����������x��n~�����C������7���3`/_����� Y?�y�{BL��ڵ�	���!�j���Շ�vF�-�����(㛀8�Wz�F	k׈[q��۰�-A1��T���$P���"n�h�e�Kx�F �b�~B��!zbwص��7��?�������^����M]*(̎Y7�s�t��7�B�+���n�-	�ڃ��rr��x�V'r�^��6�a�>�pb2�_�g�Iw�x/��Ӿ]v��J<�f�1�����o��h��fl��1��v�cr��[�A��q�e=�[3d9������2��1uA/`�����EI���N=��)�]�:��D���O�#o���×��t�����Ə����c����蛺:��ľ�9��Vu�e���9'|�Ó��b:�H�S�3+�$h^s\'�]k�9��{A���s�]w���|D�d�+r>�[�w^�J�����w"�x���g^��F����7����_yG�_������_���_�ɢ����7��B	X�}3qb��ռ,
��k��'Jk���>���}�hd����S��j�05����τn�9���Q��t1)&\.Je��8T�߄|�B��$`��?������7wo~�����=+`>���K�Q��W/n^�zE��n�X�������2�L 0�1*�Z���9Q�l����Ӹ�L���� 3X��	J`�'�ЃHP ���[�ˋS���Od��]_�=+_>|�m�|����-0��z��7�����@���2&��l_Gb��~M�v�[Z���K��v��.>���ц�ʯ���O��=�,E�4*wP�!'�]W��6��t����G�c5ek�A�l�Ҭ��������%~d����/��=�s9>{/��Y�7y��9Q��ս�x4O��Q^���nυ��ñFR8���.���z�rq��+�:�H����{H#N�v�c��Ks���}��7s�1�]����x���1�]Ni'V���g��<^3�>��3'|�i�Y!?yF��c���ߴ��c��@ʵ��+2i>���}z��;v��w��c{ʂ��5�e}���Bo��]�X��yc�K��l�X�����꣇Fd��X`p��#��U\�9�m������#�%�6#��_��M7���Y!ew�w�!�^��5�\S�)�6���>P�?ik]��bA�3?�����>d��cC�Cd;�X���Ǣ����[�Z�x���$a_�f�(T�Κ>���E�b��f���&{�2�<?�����q��/�����vc^ ��P�n���cK�\@C�s�JW����?\�����s8,��������`~��/n�2x�n~�۟n~�+�����&\�_���������o���;�,�6�a2G�.����@:�����$�"�VF����$�BB�d��m��Eq�XW��;�f�o��N6�o��J�;l��I�����������?�����y]�Wo7���7/���k'��H�oX��g�|W�A{��t�Rqw����)7˂���6[Z��?�Ʀȡ����+8�,���p2�.��hX�_}�XbNbZ�'h���h'c�O�X�H�X��5|h>vΑ忮�gS갱	�'NK�t�~t�\�W%�(�gXk=E@��r���ӖD7��ԿC��XraPLK�"r�����1��tH�0�3�?"O���o�򞴗��h��}�=N����ζ>���9��_��������A���Ѣ�QZ43N�rw�
��k{f�R�c߱��

J�0.�;�feH��XN�I��Sm\��xw颁(��j!L�����j��|��=� B�t[����`mS���"�yS��{L����:�����6�v���m3#׾v?ii�l:�:%��>ʮ\!\��ܩ�/H�[V����a��(�z�z��^ϟ������0V�>s�E�<������ݼx�5��Ǜ���s�?�������v��뻛��5I�a�����_q[�oF�������%w��J
(��,�6�+T���A�$�c�;zX��|�%�_�w�Ý�5Ѳ6��cw����'�|yg�����C���$�o�G*A��U�������y������Mn'z����H��W����sb� �@�%�w_̧k��ֵwdcp�q�-Z��,%�"Ac�攣�N(q�ۡ����L�:w��I�U�-T�X��=�����n�����g���o;������?߼�%^Y��_&[����

�/e�|�^��o1P��O[u0�ԧ���{��V��,�*��D5Cq�jȊVO�Rj��^[Q�*6�<!9�-�e��w����r`*�nx*��X�$p����m	]��]�:G>�kGvK�IkL@�nJ��G��"w슘S��R��ܘ�v�P䛄~�q��1611>u��tSq�L�����hG��>Z��u|z��e�>~�=�iÍ�ѳ�;�Z�u�Z�5om|܆�����(v�;�3�96������<�7LFYWs~�h���L��q����S�4O���1�-�P-�m�c�(	�ǆ�?�ж%�����҆�B�X��A�c�����U�g7�S�½v����a�˼H��J�m�2��5��C�rǇ�}��b���r-�Hb��2�8�����h��$Q�mOg`�-�5�j�%�q����Iw�
�_��u�śܦ�5��e�_��_7oH��)����� ��᧟o���/7���'���[M�^r���_��x��4��cR&G+�U.�-i��U0�D������[dhwb�sBV���;�77ٓD���y�	���F���\?�����W>ׅ�;_Fjt�j�_����/$c�6�����/:{��*1����('��0j�G���|��B�U�3[/H~��<�\ B���<�vGp}�Da��Q�@'�sߌ���eeJG�2���7��_o���?��I��D��	�}c�G�_s��._9��M����u���z���{���mKo;�����?x�O��9_�
h}��(-'�Oۃ�r�V��2�
��5U@�s<��|qNnme�E��1z*���˃
��/F�ి~��G�-븲�=POE'�^Ћ�Ԛ����a�_�˿�\���)�2�׸w,KQ�g������ݯm��=�?%�̈Pʈa6β�@��9s�$��Zg��)���$���Șzp_)mN�_"z7z�~�,���tT���fy��3rl�6��G����Ɓ]����14�sji���9�Co�������4�����z�?�7x�ݚ�3zw:���i_�N?�����b�e2�e��d^S'q���yf�h�z�y-9y8v��Mlx��Ŗ<���#����:��� ��IТ���#��B�r� ]�������K:��%�yK�<3A�5��o��k��xߺ�­����v)r�wy�����e�r�g�9��X��_y��]�z.	�|���R�FY#��8�J��y��$PM�����ަtL:.�ʟ_T�	����X��[L�̩�cil�5*�qc,�Y��!w��c!$�2��w�~�u����2Q�җ���@%3��u���b�m�kXjL2G�QQc}΁#�:���/^����Ky��9_p�6�:��_H������o����*�W��|ǫ$n}����mG��ŷɼ��SC~�o��'��a~�B���yFVm��	��G{��֔O\rb�Ta=�8�8r�$2J4��v�+`� �Wڴ��SC���j5�W��V����Y�e��{�7𙨫/�muNd�"�P{��^u�~P�{ڤ�lc�t�� =݈��od�'�U\��*�^`X@1�y����Wl�>�m���T��6��I �O�J����`c̸�y�]�#���1uĭ�>]��h�	=;I*�l���Wş��pY~�~I�L��a�������Sv�z��!ե=�f.��9��ϸO=4{-n�>�]���=+��Kg(��� 6��`#'\�����\�ʽuA� J�;�ϖ��v{�C\�Z���t.��<vFg�Ȳ���!
\�4�S;~���ۯ3�๛��r�*Rٳ���\{�}+���ZԬT� B#@D�!2湤+6|�}D}^������q=�|��]y��{~e����M5�[�\�v��7�V��l2��Vϟ��֥d��$��Z���	� ��WF�^w�,�[��k�ga�R�ç�4+h$`򘀙|e��g�_�����r�x�����q���g,���W&5<3v�?�x��x��޽��>�o�4���3��m���ֱn��6�U��ױ.����xχKv���%��\y!��m������Ш��*�p���$���3^���=mz�� 0�<�Ƥ��4d��:��� ��!��S�1���w f�m�8���;�	xn!�z��8)C�`�=8�Y�9h`lk�����D�{�| ��G�)���pm]�m;X�I���T[��jeKa�����H�j{h�n�IwҔV������|%Y�����e��ꏭ��!�!�C{ m�ࡕ����(C`G8o��Iq!w:�7�9��-7�;ng,G�^�����E��:�UC�<?Kܶ������`��
>�
z�fB�N�'�1%C�D����M��ݨ/�1��C7���L���ǋ{Z��}����������g�ط=��~���7qn3o"(h�N�9���S>�9k�m�2�.�wm'F��;�ʾ.�?u�avw��]��,�*�y�3�`�x�$z��-�D��j��OY ���e$I@iILL�R���e8��5��W�'S��lȖ�>��9����)'Ux'.�\�5qܒV.�>y<ً���5}�[y���ڨ�V��_�7����Ѽ����r��"��g��6
;���ݰ�xU{�[jz�Zv�5c���+%.{�1���S���#t�{��3xѬ�*3��`���e���m�6���}�;p3Q������Oe���X5�p��W/��e����+��X4��$:&]�1mj��>�Ձ�R"6�0�pnu<	�K�oYi��8k-�2���q�m;��� � @�W��3��H���/�����fP\���/��z�
��?��=&�"p���`�+KΙ-f��S9�`[�٬��f6����;�y�ˉ��@C�B
�
'1���2��`�b�c��|O&�/v(�1T��*��~�@��K�ե5�wu?-J��ZB{��]�:�����B�6���~�MC66�?:�je�U-�V1C�Q�n>ܧ�E��:l�]	O��>��|�:�8o�Qp�_�}�[��v�"��_���FB?v�a��F�sҦuv��1}��´/����m,ړoyyű�8H=��q(Fc%:�ݍ��?.��J��y��m�S��mS�2��n`Sﴵ�j>,�v�]94©�<q,�.wcK�z��s�:ؔ��s�f�����b~m~<����c��a��kZ��:b��ɉ����pR�}V��N���nYT�5549�͵�$�*�9&3w�#��|��viy7i�8$VC:hp^ǥIn��DX;�F��rK`^�P�9���,6���+mr��8�SL��D��ק<�S��q���p|��l&��Þƞ����ay�p�4�^���WZ}T�:U��E�g_����v�;_F~�ìp���-�w<�n�m;�X��y�h��7}��+t&_ނ�"c@����5	(p1�M��9�	&�D����ӑkB���-���e��>��_&`������H��=���۔w�K}c�-~�7��/�=ɥ����^}w�ҟ�ʟ�<�����Cy��`��>,�F���
�X�@�m�	ȪC������Տ>õ�A�J���9��VG\S�o+S��nW	2ر�y;NX>ɟ*�N�c} OQ>:��ʉMS�7��e��?$`��k	g?!X����X�!	��R��'I�� �;�JcŒ�);�&��w{o���q�B���c�/�.�Z���x���Wz��.3��a������S?&�ڮ�y�׼��u�zw�k�/�w}O�R�c�ߢQ��N=���čS��Oå8����:Bu=���2"�z/����y�贆&�\	7���ڗw����]���D�����l�mӿfN�,+C|���K�/���*��wy�Bq.r�I�R���<�G*<)^���=(�1��K˯�$�L}�)F:G�����E�|SP�-纯ͤS~��kW�x�������@)����+(L���[�*a���^��5�Ď��JQޜ@|��������o�݉$�ލ��i�A5��u]����u>���蓏@}��u�$`1�=I�{�c{��$[�X*zGM��	�[V����M�u�� w��X��Ή��,�N(ؤ1��Ǵ`"��j$Q���T9�GqV��D��$MJ�<�G?M��P�W�35_5������{p��L���O��2�Ws����G0�Mm�1w9[���713!bF9�s���ӭ�M��c�~g�j̕��c���Dw:���$1�V����/&�1�E�X�\5.ג�t�'�i���;۫H�[b㴩�E��+w%4�����+F6�Q7��@	��,����V�Χ!��Fï��Ü<������Z�T����~�~��^ �)��yH
i̯�:zǭ�iЗ��w ��=b�j|��W���~��ZЗ�B6�&^�<���_'�1��`�mxJvǩu�@�x��� ����T�DO��	)���#l��ue<�ڑ�(�m�A嫤C��n�M�c0c+�Tù{�b���m#���+���`�b�P�F��}8\�p���.�/�f��hĜ�v�L��&o7A^6��ʒ�1Ҧ�� e�b�,��4_0���.�p��ɤƟ,z�Ő\�Y�Ɋ�(h�E�GQr=�pd+����M���ڬ̹M�����_�Եd�J<�$'�pE�WZ�b�z��IH�#�z�#^<�u��K|�oJ��������oɰ�x{�>��=_���jR^���$f�����=��xW��!o�8�'�=�2���
m�dZ��Ϭ�#��-�g�5��!<���dp�^{܎$ �}����ک��o{x��7�j�3+7�f�mn9r��@�#����X��Hb6p�F�+qNTlD%���p2�q�'����E�!�!�(�{0 ?���%+��a>L�;�vh��D�vh��ׇ~'1��+΄rz���9�qw���nh�ʉ30�g�_��dv�РG�	��yS�����Y�q,�~D��.n���O����2�+���~�FY�ݔ�V����v;��Lߦ�S�����qj�q���H���KN�;���#���w�[K�	�`�h�S��%�@M�U{�2�Z��d'�ǱyO��O=4����eM�O=6�1�ݝ�V?��1�/��4[�%.Ud,����O�Ѫ�Ʀ�3���XVƪ��Z�׀�<I7��F����m���������d�=�������nt^ văFdMp`# Uj3�MXrĹ\�놫+�A@|~�{�F����nކ��B��%�s{��5�~�6Z�}
T��<`�}���qMZ>.Np^��9�!<^�+�g�� j��3�ܩ��5�����/������u��k{�1ZM�ё.���� �`;��8� $�|�	�ڮ-�?�m�O��E-Y� �0F��o�-�%	�`r���	��w�^�α��8�i�oR��WV�\�2	��t~��{�(B�=�0�N��p�#W���b�>x��-�.Y%;Ѓb�Ë�m�n� h>'��70I6Dy��_I�^k&C����q�HV��u�ަ$��G�7�u�}��G���Y��!�|�o!�O�Ua`�<k��D#����霓�˔�X_C�!!R�%Ìn�lJ��S��[ҹ��+l~+�̺IXf�[�e�+w��U��O/`�Ol@��.Q4G������0.ntG��!֠�^����f�< uV���ix �X����dQX���A�0-	5aD\�V��h�%Хw\��q����^�p���/y�C���C�QfE�D  @ IDAT��T)���b=�i�1��t6i��U?*������P��~9�1~�c�ԥS�F&*`����tdd���~jyF���۪��16_�jp����׿���v���F+�������C�?�;������+;v�*_Ƒg{|�⊿5��Lka�ڻ��y�R�Ѕv1Mԍzq[�4�O-�sKƗ��_Wǟ��=�Gv���f�$���3�Z��ے��G�\E�$�����-�,V�3��Z��2�=���gQ�:^��ˑ�hpdb�|^Q��YMcj��J�ḵC9�<Bd$7�Q$o��:�/,������=�,dp]���V;cD�ד���B�11��c>&�l!�,溃H�M��y��/-x�;l�y}59��Ѧ<p��7:���}H�u�>��U�9�B~��_�vi��|p��~}P����N?�w�N�ߊ\_���e�Ё4�:�n닃Ёn��7�
�n��	W�r��Q.[�ì<�`����Y$��L��>���./M�E��2u^)A&�����k���EH�����N�8�1�S:�����h����f���s�xP�o��/�s�=;���DN��C�1�Z�eW�} p��D�M3�sr��:m���g뮎.�4mJٱS�1��q)N>�Z_�&�SD�i���ei�WĨ2������Gm�C=�%ch{�ڝ�E�$�O���3%t�;Icx��n�k�*��Zl�6ᕪ�񷪆ZD��XtT�R�2�3^O�>����:�7�)ʟ� ���UP���u��؞�@���n��1~L]+FQ�9��]��q����k�U�I��u\ƿ]����m���Ў܁[����O}���k G�xۏ��c�C.�Y�B�=�ʔ⌧�w9�����?���Qa��;q=6O=��;������i�?N����
��%�P����\C<\F�z�-/?�{��e�\C<K<�N�y^��Ÿ6���y��-_��B�=���v��՝'I6�T��c�o3Z��!S��V:Y]�a���(���G4����t5G_�M�>��y�ce�|m֧O�����p5�~���u`�pmЦ�L�[r `���ج � �-Z�Ng�'r�F
lx�mR�'����W���K���[W�E�]�C�	��Г�������g���sF��T${[Y�_��i�Z;�Mcc�JQa�X�h�J��$�����<��u���	�$�i
�\Y��w�$��y��d������d��2dK�ZU�Z���b�O|��+-�Цv�B�nʪ#���˵�z�`!9"	25�4�;~���.�M�
�y�*}mV.~+~���y�T��F)p �-�2�~�� E_�d<%W�Y���	�lÖ���C'�����!/mm��BJC+b*�8-�_~����_p�i5VFgAٍ7�Ľm�Y�� �E�h���r�ʊ��Qi���j��!X3M=�mRO,���D��$����1Oj��ًo,9�э�@e�\1}���i���C3���!�R��nXA�1)9,x�q�(p��^e�Z��lUٛyj��G���Io\�I��E7�Ӟ�R�C>a'T��-&@'b�}�9q�dx�}���Z+�m��,���>�R[�hl+�"�%�O�����]	<��?�o	[��B�EWs+��U��D[cY�tC[/���Q�����鵣g�_m{��[�~��o?޿�ݙ�o��+7��ᖋ̫ׯo�����Ϟ��>�E5�}p�TH�c�e'�R��f����4S����g�8\�߾��s�vV� �o��:���8z9��$}���I� �d�9	� ��E�&a�&p�M}��J��ҏ'��u��2y]�R�<�h�J���f�b�BF��Z�X�-w�&_��"!o�Ũ��s͌��9ω���o���D��`��[���]��r��(���qH�	7�,S�N� 5��&�r�o��t���(�!�I]�cD��Z�~{�����d�
#��4��F��; ���h���R�kG�Ýpm�?vi�Dꁓ��~}o�U���k��:����?������1���w�����ߔ"����]On�2/�������5����6ir�]��v�[?�HʕOiF�2�E9�����%
�#i�+k��G��R�+>sMq�7Q�#'v;��6(�Òm���t��������_ɗFĎ�16.��˅F�rF0�گ�p"[�zK�&z2%�"]Yÿvة$�u�Aⱐ:U���"�+6ۢ�-��L���2rC�×X%��*y��}�vn}!����-�e?�y=�<���6V�W���Pׯ�h<%Y�V������9���R��p/��o�s�.��5Ih_�i�j�R�fȨs\2����D^h�a�����Ƭ�W�l�V���^%��J}�;_�`9�h�0�3��u����*DBb��=2+X2�T�A,��9��>"�����0��z,���|u�Ǫ	U�G����^� y.Y�Z9 �eu�;�/8G�0c��=/%��o����o���Y����O7_?�?o����p[��;s���[�y�a9mh��sN9���A�G�+�^���6�k]��^���m�E���3#�sJO|�O|������Sg<vL@glb�<+t:)ҵn[�!��L�.J�k��)��pr�u�L�L�nY9���\���k�<&�lW�|[�_HJ�몥y	���4�k��y�����AV�n�[�+_���|�Yy��uLY+0$ ���=8��goY��Gc��^`�:|z��E�%�5�tԀ�l�$��u&a�k@�=>�G�(��&a�U6jVj�z��nOw�ʌ���@R�x���	]XPϳ��~2;���o�a�����O7o��͏��{ws������o������{י]c�b�ȡΏ�ה�B˲����7v��޹��&��lh��'|�R���L]�����މ٘?F��`��M�6"�i_՝� �PN��C��+AG�m�:�5| ��m^#�:'�̋PV@�K'��YZ��d��>;�r5bJ::0��/�8���ʛ���)��F(��a=a'g��.#�X�A����8�Gc)}�
�O��u�?�<���\�_Ҟ8N�m]���yL���	�����'e}�\����0��yl4=省�"N���]�ԫ�<��¯j|��>�cC����0F����t�]��]1Z>JV����f�k��<-���䌼�>����
��F�sE�G�C�@�?�-�&<��`�O^r|�7��Yy��o�C����~�V�˛Oo�u��'�f����|1zW��s=�<�_�����ߣ�}���e��P�:MX�X�k �jg!��Ny��;u��CB�����J��͹���F�4���FiFoe����f�:���E���k+��k&��Mf�&O!�l�� �t�5�D�r��$&	�_���{���G��%�j�N����ݺ����fu��T���\�u/P��ؒ$\���d� ܝ{�����%qB"4�.%��JQs�V'�V3��X��hO@��&'�gc���E����ɦ~Pk�5��Ձ�}->�u˯��Z�oo����n��?��@�J�/���q��_���7�@r����0?�i�"��������V�����R�"\&S�ׄ��.���wƎ������w�����d�ԫ��t�[�˿�HU��t �QD_�����i��!�A(�|ِ>z�Mj�1K��n��/Hv�����G����W>�v��/4{e�_���l��6��P~�K�&w�`�X}8M�#Ov�K�ˏIZ?��ZՐ&�����)�,�]�7���\��X-�mڜ��Q���4��2���^C�`E�c[ɉ��t��OL�ch#ܘhsc��96N�G���%���`G=�Y�8f�Ί#FyaV��U�%�귎�Ӷo�V3v_���W!����]�˴�<�o=�	�,��P�o�c�VT<����|ͷ��ɞ���9wP~���o_�����ׯy������-/Y�/���ɷЖ;Xs9s!_Ch{��6��m�o�Q�X�I�z4R���9�i:�KY*���6�wW��i����,>�I�F.4�#_a����dс�Uyə�3V?s-��;�w���|� ����s�4yo�
p�v�˥Inf#�F�oyX-�]]��
S3���?jA�b��Q��ek�b-���Mwb��	�b��\&}l�OquO[��S��I]IʐRv=;�FwI�5r�:P.X�a��[hI�g�����6�4̊_po�_q�����O����<��`s_?���>T��;3k�T�ð�ׄU���֠���k`'}�>y��'F{N��[�;������N
�BU���P?��H��XI!�}�n~��2�22T1�*���1ȷj��xe���O������n�&��Uz��.��@�b�0�.M$�=���.ťH�����I�sͳ��.\ k-�f-[R0�V���/�	-�RO{q�X�N����!�ktD��9HcF�ŕnN�x��ë�eӡb��;��gp'_�2�-��Ŕ9䟼;��G��nȃ���������;$tl�اX-�hO�L�9>�ơ%b�ң���)!Ep�W^E8& 騻1ΫZ�S��{y�^�ҫ�G���hWX0��=*����7�������;�tL�|��?-h���y�'�I�g��績��w���5�C6xt������{�� �6�T�BR�#]mY�(]0�O���:���L΅5e�	�����,��C�0��V���oq��o]�"�qf���/�?���w/��'�n>,�,����&����j"4o��`ȅ�l8�fc��4�\E�b_�:�<���§
72T
�2t�W�R�ؗ�ɶ6�5 z�{���[¯�C��Vm��U��F|[�(�+(~k$���`}�r��_�V~��υ�ۈ�yP��o��y��O7�9�~��w7��_�����Y6���[�����r�-���	�����%.��l�*d�{p�Ӷ:����o��2w���sR�6���_�5���E��w2H"	�c.�B���w�=�'d��t>E��,��9��|��~�)��J��'�Je�ƎT��BGJ�iG?5	���=���3NE�>�� RT�	n�(l�t���@��ӊ�ܶX�CQ
a[U�Cx䏒5I����R�⢜�����$I�;�2K[J��v����a>��s�;thjHǳ�Gګ}���9��zK]������%d8����[g�îx^Iϖ��@V�����!"�Z�&an�	I4�*�j���*Ǯ�F�H��z�Թ����ܴ�9�_��ЕL����5�c��0�6.�UWƼpM�n�o��r��k6�V��u���!�k�I��x{iJ|B��q�݅���֏�_������/B:�=���`����4��74�u�Zm����b'2K.�=0�#ϊ?ڑ��y��`3�]�^|3�9����!t�J����C)UYh���U��ZI��Ļ�x��{^�OM�f)�����  4�r@�ի��
A���72���d�d�Ĵ:p�մp![�*y����36ȝ6<��r�#�������^�<	�I$\��.����g,���[���۽�C�a��t�?ː|��8y�-.�B�f�$���_W�Ͳ���GL��~�,K���$������d�0;�N�`;��CE�VXzɽ�>�$
�C��TK�+~ ��$V�'��s���{���!0$�`����ǰ�
p�!(if<䰸?lIg���'�"<|�t��}-X:��_�-)�8�ퟸb)�*'�
4�k�l��ݒ�~卯���X��4��E�/�����H��4�B�`Y6�>�����.�#3����N��o��^	{y�y!g$2�d<*��ڮ���*��6V��R��q�Z��z4����IH|�8ˉ�`�T�� m����m<Tw)u��> W����+]�Y�ߣ��hS異ӎ��6ܹ(��ײ��x��{����W��3��{�d���˯ӓx��|>J_rs-���]�e\Po��o��gsF�Un�[�Y���:;��@J�1!	�;㑾s	��݂3��|���)Әz�Ԁ�����"$�9>@Hpo���k�s���۸�Bh0$��D�[�J6�>���5�P���3�9^;a�	H���_m��GK	%��i-�t�T��񁫧�G�,5�*e5�җ��1�:x�H^�K^`3�����C��؆R�]YD�����FG@Q�j�	�[����9�m�O���	f��b<~|����-N�Gɏ?����'~���~M���zo{�e�2��һ%N��-��76��B�\1�ኒ:rA�N�A�tNZʳ����v�����P}���{�9&�r}8�J��f�צ_��?|
3�2{��ϹM[љeh\����HR��+�z���^��Kvv��� 0�)K�e�z�w��trFsw��Y�Ц�zy�/Hʣ�R|QIʉ��Ն��>�
��N��ث��_�
o0+�I��/�S�̩��P����m����R�2.���Ա���/��D_��rƇ����_.�_3-��B����a����XR�0\���!ҹ�D8�����mIr�uз1t�Z���1x�[@��Wt<����8>3�h~ c�z<�f����F��w]z����\C���˯��y����O���#�l�J�=����3�H3����69S��mǫ�y,�,��2�_��m��6���P���:�=�%�s]k`�d�\4���xa9�D�<!%���l� ����>
cl��6x}��/�Q��S�$:WV#���#�5B/�T��E?�_����tq8�*C{:<�r� �?��nY� ��X������f,���Q�99ѓѿ ���6�H`V�$OYT赥(}<Ћ&�����B<M٧���EW1N\�s�p�#��ׇ%_�t�н�����|byO�e��w<��R<<��zii�,�',cvq�9��7��]�m�\j;	���_����+�1?
�x=4��J��=*�v_ȥ]�2dAщ�r�4c�;��v����THv 2�B1���U���ܞ }�f� oȵ��b�HhbU�����Z]�pnRl��U�)�W���&fh����,��F�������R�+�����K�џ��TZ�O��:�׻�# �>eIw��e�䩶bB�nt��i�&����yO����S�hѾǠ�N��Sh��C��Y�؂.y�6q��!���ꑺ[����'��q��G�vc���sY���׋�zܦ�j?�I�\��r���e�+/ Ѻ{�����oo^"�#���Y�[^�<߾�g���k	�R�;
��7Fڛ3�:�ie�R}�I��X�	��{.TF �.�d��Ҟ��#�n6m�&BJ�@�tc�b_���DPxM���)y,:8�C��&�Ҵ�w?|[C�hKU�ӆ//� �&��[��.2����M�nn?�(,���b٭�R�%po��ݖ�r;ӄa�_�d�g�T�&AQ֒�t�&�,-.�3��;�T���@��P0�%�!$4z�j��ʖ+��pGO���>��j/�Aׯ,k3+(�G����������9��6�t���������|���ӌ���H��G�;:�Pb�����ډgSc|쒗mo�5� گ\�"����Nb�ӣ;eTΣ��KCo�K��GROZ ՒA�V}����0�����	 
n5Н�_�J_��<�Bz0���%Pxڵcl,xⷓ3{��#����7(�x�ByF�X�{�؀�x��Gn�Y��>w�O-~�R�[�4�|������o�K��T��<b��-���m�$�t���:�*O\�ieM��_==ϕ�}���0Cdl^2V�J��P:i�E��m��h-��V܁G���!��s�D�]1�䈜����T���Nd���8�y����5�b�w���5-��{�_>õ>UG�����eڽ"����_O�� �)�����4߳�n^��_n��x����8&`^K>z-��}V���rN��jG=6�w�b��@]���#�ϼ��L��ִ<᫕���h�NtV~�Rڇ�;�k���}�%-ϸ�/`7~p	ps�C�>���%}*H���&�1��Pߦ�<�KͨU2�͏]s�1/\%������%W�e+���& f񱖺������P'(�`�P"�`n�a��]֥[hS�HV��ͬ;����������c�N!B�Vn�>��X�kr�Ƿܣ�� |��K����O-_��~�������8?r�(���܆��u�eu��-�t�,s��84�(�1:A��ˋ���'c�V����ǀ�3�7�c�D�?�ӆ�#w��Os��s1!��x'��
����S��;f�  �~�Ϙ�L��#;����J���G��[�K@�ݨ�IIyGqL24�O��,�P7%��a(z:���{�-��DL��C��\����UwEվ.;*7��Sj��e�W[�d��.��vm7���t�_~F~m�9((n��x�T�jS�j(����eq��B��@���l���ј�W�A���|n��f��eC���n���y��@(r�4-U��<�
qqQ�@ [Ү�`0,"�|�O�ڿ�6~��-E�~�tt��#z����S�-�?��� �M-��Es��)�<f���p��g^��ùo�w��;'�<���00�3`\Kh�!�C>��Z�Q�����w�-ĩ��u�Ѯ/�c����]�i�O܂,�]�h�F%RR�Lmgڍ����2ܯ��6y�5j��7��4�k� m9W#�]oI
9�l�Y]
X� ��k( �Lΐ�a&I��r�;�Y��˔������e�GIS���u��6M��U�=�ҤLz��SW�UC�@�4xq^�ĺ��<f�(j�����n=��kVňI�����A��]�ӍG��ཀ~0���/4��ۯ��Qo7z ���- �ɠ�s�&<6�r�Q�o|�3:d9�J�c���/Q��z��/b�Y�B�V������W�#�2̏�7�țzC͌Wl�dT����2�sR��W� ���6��v��/�Evѭp�0?�8>yCs�O�C,�������QǧI�X�K�юNd&n�%F���O���}#O��cR@E-dI��1�!�����~�V��'�/�c�(�7v�;u�ʉ_���"��_�$�x +~�:v��}(���Ѹ:� ��=���A�G�����2 �p�C  ��ι���9K�C�ܔ��m|�����"�A!�j�l/z��u���,�a�_v#��@��	?N�V�J�x�o����y�K�i�)[��p-���6���[Q��W�v(C�����<d�S��m��O��p���wP�(z=f��=�˳�^<E�?�G�����z}��_�a��|^;g#���x۱O����&03�풁��g{�O^�(�M+�F$��D����z���U�� �Ms�np�a�r�-p����(��m��I�]�K��z�_E$��1W �f ��*��<��M�1��	���WYy�����u�Ր�v�a���d���Q%���%��I�aO]�5�EV��*]�I�«\-Q��^�Y��,��O�罨G�>�W;
_�4��-���O-�^*l�QXb_0&|�n���m�P�6�#�����7���E> y�Z�H:z��fK�e�1 i�5>��Z�P^�8:����̗��{�7i�v�n �CL �$�fl�D.�s��C��>�z%/�)�"NJ3s� �6������	�eW´���b�Ъ!���=�r�q��מ�s��GG�`�8����o���@43����DyEEi�����. tb�@�T#��Q����U�yDE�d4̡]h+l��qk���iYy��j+wm���6��!tft(�]ʴ1�cS�ذ������6�.�*�/��Vsfd�#����.u+\"=��y �٩&���Tޘ���ꩆ82~��lǄe�B<��T��[��w�Ey��۸B�&慝Ȉh���<{�a��[ʷ��e� 7�[�z�qCC�@��U����[�����Z\��������|dr%��}��u�k��s&�5[Щ����)mז�C�*�e~���C��\΀�VM���<���˳���Q��,��ӫ<����>��\P =&"'�v_���S{L(c�]>��.'d����K`�$`�֟����o(���$�ַ|�M
6�;_�$Q�׿�e�l�s����+��\�[C��EV�P��ڊ��0�J�_uā�{�"��:(�5��:�Bs蕸p������]x�ז�Ԃ���R��Y�͍��em@�� ���3����率�3nP"����Zu���E�:!��˝���G�q����_�c{���E�89Ú���l�V,6�Gu��'��";�;�p8���MK^�ĺϾ���:�EW��결�E�l�à8F�˱bc��߿hN;F����=K?��G�";W���q)�LI��^E��c]t�gwEWCjmefE+� +�B����#��$v�kbdS���9|�z�
]�B������a�����n��(��Kwlz<���J,wlO�:�H����9\�"|�0I"/t�[���d�\�g΍��ً��]'���ۊ��ˉy�9������XH\CLǵ�b��?������-5����xZ���������M���[��wS�̅]�2Jxl�f�v�e���h����=//yN��wi���A¥;V?���!t����M�r�b5,��RFC%�A9 |l�X�����Leԑ�,����Wꒃ�ȜZ|�(K�\�<U"{έ������ΝԂ�qF������Y��!~�dZJ"�;Ċ����3.F��s���]_Z��G��D^�QN�뀙-� �X�"%��_q�,Wj�d�[cCz�"bY���/ �����`Ac�&he��ړe&F�*�r��T��&�z�EVV�¦���r�X��r��mLW�k����tŦ]��*J��M\!rlz1�#�I�	��=y�
�׆
T�>L��
】��
vKС��LL,��(��Q=�1ֻ��o�����ʚ��N���_�Ǿ���
.��8~p=�H�j�\��~p�䕤2ʗ}�,x�ʪ<etsn- �����8V�� )��<�.�ұ�0zѦ۝��2�ֲ�@�QI��"�4�a�E�8�mq�W:ن���JOo�a��Pe����E�ɀz(N"ˌ�J���[q����~xĴc'����Y���\�x���>J�>4�ZڛpW@t�Y)O���Ws>�:���cst/[�e�q� ������[�M\�}�ܲ����9�u*s�c'�1,e�:��#1���Z`�R��i���x�9���<���� �Ҷ��0r�k?Ub#���yw������&Mɍ����iK�q�n�U�ۀ>�Rޑ{�AN{] ��/_��*O���!X�[�%�X���]�v�'b�*@yn�(֤����wFd����!���O��;�9�,T�7�ڏn嚄�P�w
�>���o�*s����\�}��OI�\���"Wd"���s+c�x�n�a��Pq�oUڏu��^ݜ,�O1^l,:�����R�mR� �	{k�va�3i0�'����R �������(�.�{e����>*0NJ0t���f�������g���z���g��3`�����3W�|(��O��:wL�f��H-�8�lb�l�A$�HH���:YG���|�~��h���Ȋȇ�M�����BN�;�' ��;3�Z��"�Ǵ�=ji�
��SE���]�h��p���o��S�QE4�W[9����'q<ǘ=9h�4�R�E�Zz>����R[R/V���'�Y�y�,��s��*�G�:&�/�|�{�H�e���]x��y/+�OB6�SDE�G�SШ�uby��Z3��P��`\T�)��g����JA�NDte7e5�v/�����Ľ;$�����9��Ωs��Ո>�+��:�#���!O��?>���͎����6�a�t9��H"Pʒ��6�浪�����ǼX�:��wi����s�kæDgzp�6ʖ�Ϯd;�Hq�L�|?g/E�Y0���L=��*瞎8�+�x�Kl���3��+=�Q�JNW���Ԧ���5d(�b\B�vT�g�&"׆����Ⅹ�z����c�zu�h3x��k��Ԟ�{~�4+8�R;�;2�����g�X7J<8�����V��sW�a���2l��z�䎞�b�1yd2���bm�εcwLGئ8���A��/���K�`�!0�Q��� �XȒ�2+�}��В���K`k�G�#�*�@v�"���E��^2��<��Rٖ(�Y��S�}V�b�S8��r�7���Ռ�@��;��-��ZT�.1�.�Z���Z}��Eǉ+��9&��~�!��;����z�
�E���5����W�bK�GnE�-n���>t����S1-q�%&r��'>(�ǌȷ���hZ��m�_�"2��jøK?�B�Ieq�����-]Yu�"�����o�]��^�K�0�R���|ZXS
�y-��x-�1Wb����[BLm��0��/�L7~��W��,t|e���-�u����5t����Y������F�R0-b��C^��X�ȓ���e�V5�N��R�q�1�d�樂f�/�4�����z%��$2��]~�=2
Ou���H�`��N�|.l�V�ȡw�v)l�����b�ah�K� o}Y���b��F��t0��F���4oi���.бkt/)ĸ8s	��&a	��@��hn7&���u<��|�Z~��E�������Q������B7��DpX/	����a�����w�غK_3w��"�T��U�dG�fL�!ֶ���Rg�sN����+&�m�ܘۤ��� �ؐ��|q
�9� �0�Y2�~"���O&���p��\���tS���!��hu�"RZ�!��W7�d�&�+?.�&� �,;�h[j��tL@��7;�B�
�<��tL�Y�=���������ޱ����<��F@aʴTF���Hzm6�E��q�cgn5��)�>}$��!WzN�p����[G���Q![;$�:^؝,�z�ꈐ� @������Q�>H �Bc;%ʖ΁]�
�Q@�8�.�BX�^*�尖����fc"��7iT'Kآ"���(Ɣ�[��f���l���/�c��/MļYub�
�c凉%�=6���eB"wtD�=p �[�Q˛�g�T%_�O#!�;�x��F�'^�����1c���fL�qu�ze�z� #�ȴ��N�l�&�xHkrB���0�cf�F���{0��?Ys�I]�	��{���ӺI���{��FE�.���'�ɘ�l���$�*�C{rYG�V��î�b�P,"!���`������K�� ,Q��jOlnQ����l,^r��:Q@���]�޵�yw��J��PV3�����
�,8��s�[h*��bg��i���w�5��	
D�P������Z*����(j��`�-�5F6ѐ�B?�
�]e��]h���g��� ����1�MI�2oSQi�.���	Q�}���M����=����%�p���:s	�Lal�Wb�mr�/4�࠿�UX��u
�	�A�2u������b7��M	�vU���Y*A��8�H�z���]|I��羹 H����I�������)*�Oy#�F����(A��~'�G� �:l��D�k_y�����,�ٍ\�m+�@HL��ht@�;9)p�������i��@�y5a��'�=a�2˖��X���`�Z{�	�*��[|&
ԑ(��O�ʖ��t�b�{�ڦ�#+$(�f��@�'[����J4n���f�%��aL��%��E���I�!Y4=8� �����t�豳�K��1^�un�,�ĕս��Ki�����[ 6��Y������s�[����$���q���fE$&n���	(��C�MF7�	a�:cU"s�]�����c5C�[H�jFe�~��	��iO<�, ��V}�=��aMW���^ɐ\>,qr�T6�!R~���cm�^P�I�E/jr�ò�`)�i2������C�<#,
�9i��B���ǿ�� K����|����n��9��k"��%���8U�rkǪb��� �����0�C�^A�O�μX�S��I>6D���:F��p'n�Kie8��~�\O�ܹ��1$ˤwݎkg�@k��Z׷˱lhe�ŇV��KM>�OQƺ���)��v�f�gB�4��Y��)t�W��*gO�ǌo�Ր�/��G�`w���k��.�h�O�'�������{�&_���qV)���Wq�����y)��A��6jC�٢�!;�J�xuꙷ,a"����<�<�6��ߏ�~�y��g���[�\�{<�v�������!��IȞ�:
�y���{p�q?Y�/��tgh�D��P���ǯU&|h�`�ҪE�\������Gl��AG�>�Η�;���A�^?��ܔ�Q�i��m��"v�i��	r�w�F]�OK[���rۥ��aYt����T�,g<sg��~�t�e�9ρ91��E���R{t�~�l4M��F@&�![VJ.���.���]��Y����Q��G�_j���klt��*�e�2�JӸ5�.^/E���>�fJ��W�}E+�<�����1�Α$�9F�/3Ig
G��p\c��&�E�v߳:j�3v�C�˿ew����4�V�����v`ֳ�O�D�c)"��ѕY
�gZJ�?�w�H��H�B&��y̲��y�ӟD�A��r���<�`̡��Պ�g�]F�<=���/q�>���g��T�;�F-��(�-���AV^W{��7��EV�,qD/��;�J�Ly�����~�n�6�r��l���EFϱ�{�Y��'s�0�v��]ٍ���h�:�˿Ԣ��96�\�i#H���ǘ;��L��s��Ǐ�}:+=��,%*cdWO�l��r��}�����Q�_�16�O�o�g���K��U��^�}P����qz�I��#G�]O{R��
QN�z~)�{�fXVm��yt��֒}������\˵M�h�X�濘��1�C�?�&]�[=�:Go�����Ӯ�V!姭Ψ�}��{��	�w�ADiCJ��w���mf�����0�6�ӫ;~��o�PW�6l�'oz�{>�z��
����<�L�J@��h^�Y3L������Ƿ7��	�������x�<G����D!����d�*��/�z)1�psR��|6c�'|��p��� ��zB�2�Y��6Ґ*�[��x�I���	��PBڮ$92y�F��\'F��Ȇx�{Y��4�VWD_��ZpíOS�n�(E,��Mߍ1��k|�r�m�6���!c�r�q8�U��C'�>��_�D6�>J7��Dӹ��)ó��qX���ԡ�&��F�!ι9c-6��==��(��OT�����$_������àz��޶sQq�u�@�s� �/`i�G�˱��k��Z�شZtT%H�ֻ�H�-n�'a�$%�ա���<n�9��v�Aڇ��Q�,`�w���'R��#]�;ϥ�hl���M9d"���R\,��ƽq��R?��tr$:�? �&�u�PYK�XȤ���V��8��숽���&�ig��.�������Ԟư��$q��S�^F��j��SВ���Q���JC�s��C��Mpb���ڸ"�G@�Z��EIP�K�DZ%���U��,���	n�Ӧ���D��e�yѥ����~Ss�b-�=	laO�kad8>�@�g�w�T1b3� 
ӷ����И�C<���o$�O�l��-r��]C���ݰd��3�`\>�OΡ&GYp�\,s�� έ&3 �O�ј[ b�-	ܭ���#��EO��.��2g���'�snpnj��5��׬�Y��P�uޥ��t��?�t���3�#ex>�y���ޱ����[�/�	]	�������wd��a���~���[Qo����dq��߁��o9�?�ѡ�<����޳:����j�&����vl>���M�D{;���9C�����%�z`�o�  @ IDAT��)��=W~RS������� ��Y��׃XU�����Cl'�c_�� �n�AH��n�g��^��KQJ�"��#Qq�����!�r��3Xi/�k�4^�� ��R�2F ք�h�h�/��C�>������zdN�a}ɧQQ~AؓAA������L��R�}p@�h�R9��7�܆c�6H������(������5i�J>�@�o���c��GV��2]x�]�;o���e����;����44���п�\���K�����O��	p���cG����s~#Z��4�dŊ�<�-�0D�\��~�f��kY���|�x�%�R߱��0�*H>,)�2�!\�=�)���s����r�L��?+5��_���÷������󭱜c"��Ġ6�:(mK��նڿ�Z��7�Vጝ�f��wF��I�a5n����/&�� )��*:� ���9fV����E;�Kr%UWj��wJi�*ͼ� |٤��:mB�c)�fT�mVָ�8%�*w�*���(+����*^��g�PhPۮ�l���8G	:/�n<�M}��ĸ�Os�FF���,�>z��M�p,�.(���y�}��՗^��m+�R6��w�K���F���ZK��c���46gi	��-@P�S�IW�>s�t|����t�
XWȼ�u��폎� ��O'"2��D�g�o�~��&_.2��8���c����	K�2bz�Ķ���~{w�/ٸ(�gf��W7���*yρ���L�}������L��$�$� !������_>�|x��{ŭ�[�@^w�쎗�)Փ�_��ǁ�8�)�ߣr�p˷�L�H�|�,6£�ޚ�ȓj�6 �|{ Y	�$`X�{3Y�|S���-�~8�k'��di�%;�Djڵ�}�)siv�V��-��o=��hd,J$�'��<��:2۶�
�6�KO�hX����ףCH�۾	���)��%�	ߘ*S�I���}��*?'�ŵ�U���kcb[�B-����vw!E��֡j0�jN�'��,�p�~x�����C�+��=�8z���� �2�b%�?�k���ǂ�����Pe�~���]_C���������/�p�E�M|�C��+]�U�a��Cqu[7M�r�s�Gq��N�ؖ�!��bw؜"Ha�?mg�I���`��ɛ�������ؕ ���/�X ;�=WOw,�IR��{d���Yi���wss3sss�#<Zx.��èR�)8�2u��TX/ա�GJ�üS6BEE�hg���3y��%F̊�t:Sq<�&\'��R���ę:<ɟ4U.^�SF����D\�
�Gn��G�I]oWa
gOgP��݋����5q��<��1�<1r�,����8a�á3�l����Gx-Z*���2���"E�x6��`-|<���[:&ə��Ɖ/�Q~�77Sם`ܛQꊱ˻E[�OUe#\�렡a|��t�&�u�#��##��8�s�{҃[�r���1v�.[�׉��ȧ��5�f�A�'���7��F�\4�k��	��ɮGc|b@�ƣ�,*3H9�<��02ӈ��:���dF��M_�3��"�a|�~���ƽ�g�g���ݜ�D�t���ɺڝ�@`�q�����y�^�-�����6��M��o�'�,�^��Xص�a$���%Ӗz���:c����˼dt���E�����e�lc�7�c��哞d�"�N銝�Is$��g��Ae/+�A.;st:�56�a�D�v|fD��z�d�4�i�<��'7��+
(k�	so�C��	��VJ�Ц&	���S����G.2�
�E�H����ki^���D�2zm�E\v�����@�t�@Yq�a"��S>����(8��k
Y�Z��L���c���uJ���uG�����=u6~�Od	&6�JY�E������V�ڡ�����t��5���Lʺ�*�
#!���(>|��8`�YV�� �a�:c ��i�dԏu�����t
츨Cw:"V,�3�WƢd��_��qM���4Q��U&$L�q�w�l�K��61P�V�� �\���pF%�A�D�ʈ��j|ʉg�J��]%Ϧ�AAc�+a:��G�6a0�^��U��h��_)4-���(��W:f�g�P��gg'���7F3���X��hY��,�#�\�
��7%�M�<��&�.y���٫x��s$��_<�~��<ư�8�����ʔǔ�ɍ̵��KF�Ki��c�{=,��,"My�rAy�	i�L��	���|��h*Wa�%��[��[�(�_􂴕?�H,�Ŭ
KP���Oі�/�\��!�!U����;�yH]��<��g�i���uD ��Ǳ5�Oݏ�<vP�n�q�P�������:
q&�����N��a�6KQT��Y�B@z�*٧���C�!ʌ���z�L��Ӵ�O�s�.g���Θ��2[���r*�KM"��t��������U5Z����_<�/�Q��Hyp'빶�A�N�sM���.��ܸ��u�����·Ŝ4.��b-�|��=�)��8��+��e�=S�[4|M}wg���T�j%���FȊc��� ��]�k�a&!�O�hu�������R�J��go0l�z�G �y��	�)+)l�[�ˆ��WB}-t�[���,`@�W�YNVU}���G �}R uW��R�I!x�w�Jo��|��CXAj���m{�@V���)����I�:���:Y��|4�������t=���%9?�����"w�&3��Ɵ5���nr��������V�|�݆�̬���ŋ)(�#��r�[��MN%�#��2�����p�`G_p��|-��e���zx�&�58�Y����EH��݂K��/����C�'䅢W�#�G�k#`�a��()�z��I=�ef�♯`��<�E�o�����Vp�N\�6�P#�p�jO��8m�uP���/�L�:�����ND���q�����G}r��<\�@�p���5�8z�C:�����yH����jX?����rJ\�g�Gp���[��8��O�^�ֿ��g��"�e`Sm:}��"�A*��=|6{K�4bB$�7�xmh�G˚���(E�Mӳt�!�I� W�U�4��Q����铷�｣��{����C��C�;f�
L(����t�����+	��+��i�G��7E0�*\
�z��`�\�ϳ�T��Y�ɑd�8������\�W9B��r`�s1]�h�b�qC�u�2c ��,��c�׆�m�ڥ�崤Z�g�OBWp�Zjjpɯ�Q��m�#m�%�jNٚ��ԥs�UXt0NW���1É�R�S�0u�5'�{�0�8ɬ��~�j�5c��1�����غ��w�+��ԋ���ag�La��⊩I`�Vq��BIA���t�W��8_����	�I4{�� +ͅ�*�0��u$+8�[Q����Pp�6�05��T�Zo��i#��uw�#��3�[�*�W��4!��Z�%�(GWF����&�E�*f~��C\	4�� ��	�",���T�;�4>a��$oPV!�2�.aӄ�ɘ��*a���N��RJZ����H�ȦaA�v����IQ	�t=�>�*D�;�T���1��F	��x�͓�U�hH+<�i:�vT,*w>�M���]�_�b�3����FA#`�x{s[���&=�P�z�t,p�a{s�[2��;�p���"]�6#A�/������hIU����b@u�U,�FUZ�W���Y��A���p�8,�A��k2/J�p�s��>"YKG?��N����r.���0�S������(��=X�W
»ś�y6��]�Y�e,�J#x�o�f��w��Ƚβ2�a�������(9�ɴ�0L��������2/�'ER������vc3�K�J�Ht%zBXV���Z����/�Q�^�\�v��
����Z}��V�V�iFt��f�,�uV:.��9��h��% dJ~q�Y��u�!I�cBm���G^I��U�d��I�������!�b��v}�k��b������:�l��@F����:�(ϑ��3?^s� ��`L��a���9G���kF����J����z�r��L�Ϭ�C�\��ׅC�y�m\�����ӏ��:b+��m����nǞ�ġ�*�t���V�#H@�hq>r�U'�>�N�^�\����들����͂ܑ��Gm���/����I-*�ķ�ѝ3��ҭ-�2\<3��xq]���2GI�EO���i��o(\Л�1<x�0�O$e�o5PflO:^"a��i^y��LQ��XT�,������W�/J����j�X�<S��6�����-����Ϙp��\�o���|�|꨹(����6M��� ��>�9�E��9x�Iɚ&��m��O"�5�c�$=m~p-��L	H4r]�j!K��ypD�Q�!��x/�1ʈvo�"�/���X�cz1=Bߘ�/ݬYh _DU��X�SY���[��hY�:^����+�l�^E旣fT "��-*�C�%
u���B�ŽjܘՏ�,	v�~�g�H4\`��;�ZH&zx�+���������˅�[���L�Y���p��@�]0uo���T�3���Ac��<��3����ˋ�������Z]ZbG���	�V�W��R<Ri^��C>��	�e���hpk��S�z'�8e�|�QTx�B��2�8zo�ڡ�o�'��ް�2��u�GQ�t$3�H�R{�8{Ze蟲�>�
'�`�#��^�����&)�?��ro�T�\�������U35C�a+�0�5�
���7���a�Wu:�"<|I��笼�u���!�*�-��)Np�		.�9a��^e�������s�������H�E%S����j]��G�e�yhb�_��O�E�1��KOc:q=||x��$#��ׇp�Y��Y�J[�C�se"*��K���!8�u��
��Y������W9�yU:��/p?�/#��N�cu�(cwY�÷�-6i����)Gg�̆���x3,�����C-����*=Eͣg���Q�r�O�Ti��цz�>6�i�0���!4�//:��` ��ڗk�����-m>|��2��{��Z<�M6[����`�rC��k=PV���\�#D���*P���t�P�5�
��F�ק�␑x=K �2����bJ���g�Ly�SX�k@�ұ�x��W7,��po6�bb��ap�f4y���4M?��JN>�6���iL�<-�RԮlByT\��0W��qUar+��JqTT'"x����ʉ�ܛg�oR���FT��'μ�+�F��#<&�LZ��A&��[����G��S��Z���;�4�߇�!��_�(��S�ቮ��ou�0;��0��/qN�+����Y]\��^x;��p��K�5��TM�A2=g�,��3��9u�=��]��g���p,����-���a���p�������a��!�
<�;o!F��;~%-�s�G�K^���׏.G�(�z6�p�q���������������<���l�W�>um��!���7��{��ڼ��g�+-XH��D�1Xu�N�d��t��NK�9%(�ـ�74�Q5i�v�����r9lo/���]�f���F�7����}�Ӑ�u��G\׬����6M֚#9�e�"�:l�ϾܠA�BN�p�E�W�.�q�����О?ҁIi��U�����q���:`W������� �㒌L��zCg��q$�9�пjVK������'4t:��6������q�M��{�����x����2L=Qw9jj��8H���:a;�,�͵qN��9u���k�x���22b3#�c�NZTx3�	�orL��̒g�)����ðI<�%In�a�P��4��f�ZZ�r����91̜%�b�Cˣ�]z.���k��$�m{!W���-`�9���I���抮�63o���iI�n�l�YW�o���ݧSz��͹3�9=<���X"�=� ����oڪMH���1oۢW]�:m�^I����%���ҕc��	�/��ɦ���=/c�|��<�U>��''��G:�T IlCTb{C4��� ��9S$��b;�k*�)�)o�룟���LI��D]�:��Jm,������W���p	��K�-�N9^1O�A0؅��1�u%��:����½�������ZR��r�xy�qùA�N������
Տ��u*H�#i������봑u$Z�(��ѫ�ȌR����9�X�LgB�5^�.E�@�h������m��c/������Ȯ���}��S�]W�|�P��F�C�D��t�m�j��
c&�0GS]�U�魰��P�}��4D����l������e3⋬�L����Qtdn��\1"{A�{N�i�]�����pyz>�t�H�c����lxr�;�z�|x��o���C7���z�J�� &���B�Ce��1ޫ7`A��,S�L��av�
G�V�����ߑ����19��y�S�Tk�
ne'>A�\r$_�n5Z�c�l������^��"i��N���'�i42|��[�)2,���Xp�C��vy��X�6����]���M:��C��׌V^�Ϗ�:���c�h����E�W�:#�8r�<6ӗ�p��(�g�s��W�§\�9S���':c���s���QV� ��Do�p��vnW�E��Axט�_�-v��.#b0���q�L'h��*OրZFb�~k��i�ā$���]]��9bA+q�m��:d�e	O�����Gy�!N�p�]�]wu��6F��Ĕc���⤑�iuqD�"�x.�㓙q�Xa�pD��!��;@U�7����aH�+T: &|�|*˖ʇ��3|6�f;[\78bE5�8��q	aJK[;1�h7�R�����=�ɯ~�� �H�t�I��p�#[��aH���K�2�ԣ�s�K��&v`�̀3 :]{8]����;����ptx0��逹I��eP�@&Œ��aZ'lZ��b�[Js�h4��n�Z��[<P�ҹ��������~�A:�]^^>~������&��0�AٯP���B��
�z�䰇ǹEo�ڞ�3y��a��N�R"��շe�"_�鰿�#y��
EV�Uf�>��ZK�y��)������k{�\r=��~z�	�)�^\�p0��b�K�cy��&N�����hÈ�ԝ�^v9b:aR�W�lT����:�<�,� L��T��Lml�M^�#\�Kd;M�W�͹�W㳾G�u��>=�ďʗ�i�u� CkO�߇�������"|pH������cɠ�����M� r��������Q.G�l0����踮���:e9����Ek#�	���%��b�6�l�ً���q����F����8CTJ�;f�����O�_��2���S������م9���;��'�Û�����c: ��kR���/�a�P�b����u]�w9���K��I%.�.1.����9k?���������#����ϑ�2��qݛ�c��K����Jcd�2��MQrk)B�������n�\!��GF���Őw8��f�����0?����`g�Z��<�џ��G�ĵ~Iy�~E>��F.���#L����H،Q|��7 ۤ/�Jfr)<�!�/���Ӻ�fs/�45��r��˧�����6T�O��nrn�Î�ꀩKWvb�c�Q.��^��6@���Ɯ_\�޳)�'�3�+��[�Ѝ>Ful��S~Ҫ2]�j$��T6�H�b��8k'��N��~�o�`2k[io���c����B�eK�X�ƩK�_���?�N�{Y��?y���1��1�L�#w�{t��6�Оz���}�� *����>��	�,�$�|�#��TE%(9�\9�Z
>2��2�Y��_��K;uȵ^�8��7��3�lF���-Ge�<��.��Ϟ�_>���������m��r:��X,2��+uƼW��l�����z�SZ,�����&���F��� ����\3�n�i�H��c�t�}�ԹK�l� |xΈ.��/cQC�1noP���u����a�,v`�9��=z>����Y��-�LaHfr����AIũ������j����`�q:,��jqy�BR�LgNcqE�����/�O�:c8_'g��������	�.}�BsŨֆ
�(�@��~�Xh[���U�:��2*ؘ&�TW���b!v�+�E���*e��
� �\3-i�dPU@#��_�+��"��DV�	��%���`oڑ䍛��	� ���pH�ϡg�m�{��244�c�T�P5_eՕ�M��f�#:_^���_��l��N5�iI;�$�ET�7*�������1J��`T��%Nْ7V|1���N	ݒ_w�6�ӹ��o�χ�S��\Ov��|��.������{�G㹿�9��\�fPki�������rȍ?u��I�bH��!;8��?2󏃇�6��p�p?2pV�0�#�W��8�h��<Ia6�H%uK����6uթ����ã +�{i�*Ov�|v�/:��L��o�ƪ���(b��Ù#yp�c�B)�(���.�d�DƵ�af�S$������+���Uc���e�C^�y0�W��?kQH���i:|��r�]S6w��u�Ĝ���{4Z� l2��h�ۜ��mP'�,L�#W����St{�Qۻ'tl���.n�qr��Z��UYJ6�2��ڜ/��^�!�`�7��[��̆��B��fX?���\�:jjShL�UP����d�@�%V~�ixx���'l�/���\�Q�zgϣ��M�I�	����s]��Ƨ�z_��-U���u}�>@���+���s� �V:����'��0��0���`��=S�m���d��.ڢ�����Ö�/�O�|�}�b����c}��Se�;H���[wU��j��]�q��A�a],��Ö-�^d�ֿt�ïKG�œa툸 ˑ\Nש��0bw8��B'CA���4#z� )#�ˊ�3Y.������o��ްf�9?HIيkrO��:�b`HaJ1���m
I��x��#d"�m"�4��b�����p���)�%�:bV�k��5~�����������?��~8�<'�Q��e�۾cZՆ�7�\g�d�pu�:/P��^��GFS�Ѭ p���$�`�9���|̦�*2S�F��c��p�^ǣp�hJ��N<�>�o$�K����+{9%a�A_�7��ô�ٯ%��=��B+Dm�F�H �C@���]�a�JI嶜. �^f3�moj�i=߸�a���G�t��6�׹�'���d�[�0����q�v����]z;4$8`+�/�3zic��g�����p���܏��BKN�`/�WԱ��9kQ?15yZ�S~�a��%��p�i�éL��v}���1:���¨�G�JR�� M�	S��]�Z�QZ2ſM]]"����&��⅐\̈́�H�0�6D�щ0��U����3tK��`4��=�K'�:���#hnj$�t�-�O�#��l��:M�'�k���g��#�,j�E$�t
gPu4�-�G��s�(W�)�WH�O(���	,x���(��
G��Xj�H,��'������_/��cԀ�:[L�l9�����0IȮ� |�t��͋"(����7L1�sH�%0mv�|2�*o���(#7��#cG���)�[�񓧙�<g]��f���������G0/�ر��l:���>�PXa<O�D�N��|"j���1����5GJ+e8��zTzgL�_��<��|�8���5� �W�\����ga�?�_2�'a�V� �P����V����6�	:໹�:5��Y5RG�w��[֎�l9�����s֓�M�63o�����ۗ���O���=�5�`��⺾��>���5���.k�Sٰ*	�,pH4�5��X�9����8�*�:{�Ħ���M~U� r�Ǣ��Ӗo0��A�Z.���O�_͒d�㔩��::�r�/�E��-v��S;:z6s����$�T�76	q�d�LkzA���f	5�C$VgO朊T8VJB;�Ԃ7�a���cfevM����C���W��SI`��)�����	sŇ{���p�~��#bg�9��N���vF-�Ȑ��<��mԦ-6�:W�"���>&�Ftq\)�o+W��w� 
�#%�?C�A;G�rs���a��c҉��L��'�j�O�`�q\�3A-0w�#�ǘ�gX�c\_`^{��k���2}e5�Ȑ�xX�s+��/P��U0L.��O�WϏ��^=����[1�v�ˊ�}KO[�m�^�m�P7#�� �^�@1��Kp��p�&r�o7��g�)?��� Mj�Q��?�w��k���9� ��?tΨ�~�K��֋0�n��' #ڵ��ҭ�&̪�Un�L����miŚ���� ��� S�w�͒"l���YII�뜪�S�=�W��:a�m�1B���JD���C��B���a���o�Q�|f4��HY_�8'{n����^I�qj�p|GG;4�\x�t�M�=�%j�CF5�!S����N+yb��7bu��sZ��`�s��t�|xK�_���4���IW8$L���,Rv�G	�6�#3
W^�}��9����t�n�B����h�^kW�a��8l�]q��R�,�	y���p@���s� ��M{@�c��?�|��[ ��	F���N�؉?�8�~1<{�rXи�1��O�9��������i��1Vn�i���xԤ�2�UM��FQ�GiS+�1ԛ�EX�i�Є�%J�.�_�x������"��� 	h����K�ò� 3���Y�QI�d�x��$���&�Â3:�ΐ�Ⳃ�-`��e5����{����e�~�������xgtvW���.�}�z�����W�_O��I��HM�2��vZ/Ӎ�VE"M�7�L9%n��Z��tX��ٍ��L�2��q����Af�� l��˘\	K�&^�|�s?Cd�y]�����W��gð��?l9�{�Ȗ;�oѻ�|
ȩ����������=z���.ƛ��2a@I��IgUh� �烒�� �*��e�����@�|]R�Ti� 8C�z�����r�(H�րq=;?M[�(S#@FT�#[��W���}�v��?ҳ���������6�ao��Q�;6�]�#�/w6����#�W�A�UB	�r�4 ��\e轏Uy��I�b�Ucc2��HB0��(=���o$���*ȹͽ�u/���L,�b8�����3��E{�u/nQ�cz��1�+�H�|�`��֨��z�'�U��9��4c(��ct�`a��l|\���~������f��/�oXW��Z���>���7�N?���>a��E���5�"PP����������wi��� �*�|��2���|���85EÒ����4z.���ܮEg��2��0���0լ����ص̼�D�uaP�2U�G�H<Gi�Wr���������\��z��t��3:�0��f��W3Tb���B��-���/���f��z�5�D�Q���M�h����4�yt6�+��k���+��/�<�S����Ʌ��"p��Jr�	��$eC�ɿ�)��q�HqH�t���}��1	�rN��ab�[�>��D4F�Xp(��j?�+S���5*�nhV�����t�<i{-�8��#]:[�4��ٛ�dԉ>���p|�|��?B8n�o�u#e�[�W�8W�R~-��`��aޣq���j-�~�ɻ��aVY�I�-_h�#d��F��CƋߒA�#8�%�}����O�+��PyJ^��$�kݯ�$�yN�_A�n���������ѯ��P����?䛴�!�nA�ɟ isc	u���z�V�3"M������:UTZS�i�չ���퉰�Y�Pg�b�_O��i�;�-�龈l����3�c���W_��ś�뷯�1FX���\ /c��Z���s��=s��y�����et�u�3� ��v�5��_q��9�)E�|Ie��0}�Q+KyfD,i�Md�Igf�R� j*�l)�M���N���34�����aΛ��o-J��_��m?�X����������_3�rL /�R����:�~�jS!U:�*�+�=�Â��F�8�EK岀�Wcd���0
N� 8�F�ȥ4*Z����U1x߉|�2����a�}ggxBE?�u����p@/p�ъ�x����ƹo�O#H��R�rL�&��;*h'�;ZҞF
�	��)Vfu�w���)�,�4���OU<�`U6�%�����`L9�K��%��5H�,b�R��We�zZ��h��Ea�DU�X�
�2{�+�n����d��|�'��Ux˳�V�%�qV���'+��ќFy���Ѱ��A:;�e]�b��z�Ou#�m��`j���^}�.X겙D����Г/�Ew���N�P�3�$뺬�y��������:��F�\�m!�	,1ʩ5��˳	8��Ø�ت�����t�u�#�[/��{�Sp��t�`�*�kt�E��h�ī����.TQ�)?hțS�m2љqJ�Ƽ78����"�&���+D�G.�h;�i��D��ǖTT8��!(�������\�z�9���b�_;��95Q�˿U�d B��#N'W"$�G︝�wFՐ��bb����xt���2�Rթ]ܴa�&�����A�(27?�����\dL�0,�l�����,�w�',����L�C��5ڢ�x����Q
��0���ν��"lo�糖��¼�A�8$�l-5˥4�+I���I�[�����ନG|O[���AF��y�PԓޏniC?}D��l��(;��Jo4����^Va9EXQ<T��ǏZT�Fuz�&� +�~�3(Kց�9r� P�|L$���xo���ˉ^�f�5��n��Fb{���gÿ�����o^O���fꜵ�N7^_Q����Ӟ5��Zq��e�����dԠ��L��I����z3^P�SA�xv�#�bή�.UR�5��9�vY!8�Ui5�6:�]�>��>��J� ��N�E|��Y���!^hJ;������WT0zFG����8岿�ҡi)��e�7�,�x�!@��N @��)\��B/�!�8G�$�ڙ[��@�@����ao�r�PY��r�`��ҩ"μ�d>���ŭ���&���y�G,��~BIò�b�_����|�K������?�������#�kE�z����35Ox�LK��Nw��0���)	���<$>q&����7�Ҧ_5�񠱕?$,����<�	��f��Y�����|�u])'��4&�w?AȽe�ռ���>���������~���>4)����}�$��C�
�T��1V�̃?eb~N9R�1�T��H��.z���]�K�H�6ӊ�������t�������}]�.�p�B�u���<��%�+�S{-�:_���]L�H���.��n�4E�<)�aRZ(�ɶ���y���B��?�+����A^x��X���CH��G�u.��/�GFp�p_��р�'N��_�R�m �.�r��9G��	��Η1��4��ru���-�	��&�ts/m��@�f�3i��13�b5�*�\�_10q	��`��9a�ߧ��[��}Ȍ�䃼�喺��*���r3��A^e�]�Z�{��O�`�bz��|,������鼁TyX��ꬂ�����
3i� F�K�Γ:�EY;��ϊrpz==w;ŌBܰ�?k��=u��/u�)��X�̧숏�K�d���aϻ��f��U�r*pN/�Cr��'9?�0�B�F8e-��W����e������:ڶ�=I� N��Q$6:�P,��s5L~���9�#8�a�F�)'ʰ�>"8� Y�'²���g
�е_��-a�M��#�L��Ί'<����״�~V�7����C}�a�>/������믇߰����}P�\�x]��8:�Ҥ;t͙:���70;;�Kvi8��v3����u�V��7���Xkx�[ Ai|e�����;Y�w蓿�/<o�9���ce�Ea�5��q2�:t^�9�d4��/��?�ﴀ���'��rx��C�J����%�f�.�֍������C�k8��B9��F
�a4�8
dU��7�<2��9�}N'c���2�D�4��RXЬ�q4�ŀnh�(�kn�ҹE����.�e6d� 4g��1���OÇ3F�xS�qH
��ǥ�n��"'�O�Ґ�KoO�JcD�J>�t�Q��2`%&d`� �(�#�ex�SN{�0Co�qfu���D*�x��x��T.r6�0=^M����[��������O�;�Д=�	��^Dx�~�ZoU�!Y*��3Ϣ����&�z�Z�Ę��z�+�J��ܠa���*�5Zy��^�AX�^:m<V��W|��tb�?a�S�xY;���pA������e$Z�  ��)ZF=?��=B�??,u)*Z*^�z����s
W�R1H�pG��T�4���W>e�r�s�+��m�7?%�Ga�GEN�������	<���q$g���'�$�/"3/����#/�I?�љ�n� w�;{P�7�8Qŗԍ�&0G�Bg��w�/yd��ў8�[9���vCõ��>��:25�rC��)�L���7���L�/�(�;o���<�O�S����@���Xyk3y�;�k�wp eĢ�t
C30� XC�zj�)31���ts�%��΄��r�H>]�{�G�O�D^��|�e�u���m�tX5��SR���"1��ţpL�E܎��T����u���D��\Tn�q��
��� թ�u��(�*cd��z�c�)��96��t��n�FT�jx��e83s6�P7o;�kf_���~���[v[8�!gM�itl墚��z�#/|X/���ml��I���GlQ��̞u�kg���O�,)9?��;�Z���Ɔ�� őTN�t�/O���O���0�'��!K�z�����;��-��0|�%3hsF����v��i܁��}�;������e��<M�`���x��8"`o�9Vf11��F�U�>�� X�9�,�[`Ąpj,��I�M���T��p���`=5h��bM(�\���޴S�¹AC`�P/WWx��F$��!I򅗗lp�_���{>�-�.	;GYnp��0.>�d7�����3��m�>����r)E��P��(l=�d��hhJ?����t:�eʬjV%N
mC"���NpI.r쟤b�T�83�|�
!r��[��V\"��|M�Ļ�Г���A?�����Ch�_�&��lDj-a�����JE�zdxyV_w�XIo���R��֊|)ǰ8yg��5����'�q(G;�O�'�%�ʶ��is��'���B��p��Ѳ�5�a0�d5���] w�G=D��A���Q"�n���?G��Ao�����qrWk;Hzw__P��u���G�2�`�I�|�Ӹ��q�0�v�5���ާ�+����;�~�c�|��a~�7[�`����c�H�Ӿ:g� ���V�7ВO�1�'�z�J�:���H�U�����d@�:�%o���ӡ�^q���jڵV�);u�p�>�|���.��y�TJ9��8tT��ﱄ���;�8�l���Ζh��<�:H����V�_#��\!�����]�
0����B:��H��4.�[b(G'�� ��V�������ΪW��=�$M>�uE/9���e��xKy�.��4�)*�t爍��i��T׺���w%��o����i���%��/�4ʿ��t��Y��)o��ZY�	�SR�z@�����	�~�"���#;�)p+� �t�%	�R��A�]�&��d6@�iG��$�K�Ns���b5�xv<�򻯇_��Û7O�=N�(iGl��[�V�|O�ͪs�F��%6�0ۗ��/Э���LwV��C�\��\���l&}�/�w�/��:��W���1B�T�y\:�Lg����1 uP~��~���*h�;G��_��
C��>��1:��u������[z�fV�*:85nT
N*#Cvmآ�¼  @ IDATq��V���e�"��*�^�XwQ�0�� �!p�ܰ^�SJ�zh��`�ס;��捝}o:|'��00>�wb�U.�(,��<n�Gp�=�b�l��Z�a��7�W�^���Iv���O0��Q;̉�p<\Y�Ș^94�bN���5�\�_�{i�}%)N#�<T�8B(��I�#�=�WryᙴV�4��^�<l��h��-J���~�C�v򓴅���"hR=4:�'�׷*�(+�&����S0%� �4�a��@v�����\7���Ȝ�LNqVm�K��SN;:�Q�6���(u�ڍ@B#V�9���6�Ŕ�<�[ ,��������Qyu\���Y/4�'{���Ax	M�3���Ņ.i�T>Z 7+v�g��;��E8�e��ӆ3�4�C�bК��td�X�C(�%��!�M�������2� /�m2�u�Ǝ,��G�1�5b��	�Ҕ�v�mس���z�4��rm����[V�kS�!�>
=o6�T[���&ɓ�o�1������v���M֯й��<��$`����8�%mK:�8vW|�7q���Ơ������C:Rt��e��u��s��R�>m~:#)[P�_�E��{��6`�;�,�NmZ^��"������x�OJ[q��O��]�<9��UǺ^�u�� [����x�^ݯ;:�����[���(�K���pb7�����d�����`�!��5��ږ�v�tv$��ږ �i�<�̶I�T���k�A�p�L?F�F��x�TƏ<�sA�����/g�r�n�~�y���8_������:4�I���up�ѡ�ԁ�2�����ëWoغ�	� Sx�VM{;c���e3T		m�,6�N�%N��u$/ZEX����͎ ga�|�B,�?�0�h�Z/�oy��.K+�u;Z�8]��O�#f��H�Kc�'4n�Ѓ
Z؃��%�!;�朧����X���"8����$N.��ق2���c�v�G�Ʃ���Q0	��}��	��p��c	a�+�H�����@@���9�>}~���U�j�j!5�d�s��cpb<^�(�����<l�W����?��� ;��\0�礑f�������Sv�,��M4D!>"!>�Bݏ���;5��:���4\�����U{�h����,:��N��|��	ݠ������!I��f<��������UxB璵	{���5Ð�a��z����C�P�|��Sh*Fp��� 9-��B�X���Pפ�Q)y���ccS  [cI�BcnB����Y�>��+�'����C"�c��9|�P/��F���WH�9L��`�'#V�ԫ�p��� ;�S/7/qLp���#��EYS�t�{�8�`�F�H��);;_��:<��Ο��.;���L	�&�C ���5�.�(gK��':5�|S�䧨cۨ{�6,����V�F{bc���/���|��յb�m��G��+��E�=�$_�G9�!�:,�!���-+��A�6��X�م�ph�Y��0�>�7��E���Cx�.��؃�&��T�u�r�&:��֪��ٙ�N#�|ltU�3�%�/kì�����EfQآy8���f�)�JZթL�S|)c��:(�:�e%a���ᥢ��r&�A��go����4=���u
S��w
+�i�Ӹ~����Ac�)��r��V��N�
��Tl�n씣V�'�̡9!Zl�����΍i
/�V{h�R�Ȓ���Uo����d�x���@[�T��w���)cѽ�^����g����7߂�u]?d E|��E�oH�5�83/���>{>���&����^�IN��*�T��wCp�f�� y��#^�z�w�
��/�����L����L�2R=�� ��)�H2�W�{�ZG�v񫎟�}{���,贇^Ǵf��(?�� ���%c�$��TŠ9d��x�[`K�G�z�w<;�dE��xù3�p"��j����"#_�'�����v����)Bz6<C�������(�H:͓C��0O��#g�0��P1�Lu�U��d5&?����-<l���L^�N1�l7[�Q9XG"L+k���BC�OA�V�3|�j�ˍ��d�M��A{C!���lq:���B�	��ƅ$Q.�* ����g���0����L��D�a8̏EC�FVc����v>*Q��ݘM��x��"�h�����,��s)��1��ƛ��?�^��ȁ��Tl~�����DX5fⳌ04�w��fer��-��*�PX��HnHm�O�ʸ� Uއ.�L���9Hg�<�"���������řmN�.��D��5�%_�3N����O-]1��6h�E��o/�/ԟ�c�{�\g�Y�^M?,�~�Q�[*�;�iy��k7��hg��F�ih"�l�dFr�l��,A���̺���~ZJ�����FL^�n���P��8�)���cY@_�z.������ �c}�R-և��d�F�<G�ÉZS�hz�nu�m��Yyu=��Ty�M�p���x�]Ǵt���*��h�P~q���t�\ܼ�î��넺�%��I����^�i�t8m ���c~�DTݲ�ԭ�@J�Nah��$+�鯄�[i%�����FƿpX_��azy�Ob���t���2���S廆��}�(�r��(�m�f���OhV�|� �� ~֝0�v�G�r���1�
����´O�7\<�v�l_к�+�����hD���Fw����V��'�w?�O�@�{�~�Nic�����'��ׯ�'�k���y����(�!$�O$�):H�Ć��̤�0
wŴ�>�9�o|q�
�MS��+O��l���$�䃮�	�Z�tJ�<:z���v-s�	�$�$�lGM�/f�I���ò�� ��vV�8`�x�����Y�3�(�N�3@V�v�*����"�̙f/)�n�W��z�Ǉ!~�+����7�pcv� ��<��H<�7�w�w}�������{^�H���טڣ�-�-��}�~�.�����|?��F����V$ӑ:2n�9����(
]�+�B�tE�U�P։W1L�u�`�q�8��84Fpġcf9�pR�(�cC��x���ada �C)R�(���	C��('���G������JT7Iߢ������g$a�~z����0���Ԁ�'��4,�>Wy�9��c�~DХ��� ��4us2�̆�F�7k��Ȩ��;��j5B��*e��U�呷�kB�ej���y'�_-3+}���]�k���/qc9T���Z&����I�2�w���<�Q�4V�JɅ::٨���Ya�+uR�D�mY������P�� �[�-���]W�>-����y�T�5�_wd�Bm�������J)�E���BD�b����5�ө��'�iS���KH���O<�6��1��O,����2QO22@Z��m�����ٌ�5:��
�.S���i�./yI�̩PG�j}nf#`��s�D?ec㦽yYe1�e�GY� 80���oYX �����ûN������M:Nٜ�-]�]TR�)��vz�p�m؜:��G;=�ٵ�L���G�nˉRC���	�ʺ�,��T�@E��'j��\p���r��l���YtX���&x:��S��Ї� ���t��S>|���9��P��[����q�ґJ�X�FG�%��?`2K���{qiG*	o�Ws�_��j���`�k�,���o}�q>��_���;�4���k9�c��T�s���u�;9Й���-uG�R�%}XĥL;�^`�%��)�휙-�3m+��p;"�x\}9�)��O^��r6{1%� �-ZXҵˈ�k�t��Y�Mፎ"_[%��ɚHDH�"�Cg~�{����ӱaJ@o�Þ�=�*������"��-9_�W�|~��d���u��9;��vf�8l�� R�9�ȯY��1'���H�o�6�
'��R�Ξ"�8O+���c��
���Gw�=������&���lM��$�V$��C���ǻݹ���=�WU<%Z�ӱ��@�d%�4��i�0m���n얷��%,h����t0��!9,a�͎�#+BU�d��s��0��a6t9i5ڊ�s��ƙ_�ϕgAKWL��6�K�0�r:�v���:w=]x�X�A���w-.
�{Dz51��OX`ė���/��_		@`l|t~=�0f�s��`��4�KK	UZ�MYy�meU�'LJ��Ս>ҰK~u����_[ܿ�DgOޑ�IX���dН��w��V+�H9"s���hu R�#�W��K�a8�����	5��1�1�����hY���cF.��Q%���4�0�f�V�ɶ�J��8#<:*.]�}���b���#�)_�1�Fa��	x%l�%�G�� 4��1�^�t ���jo�踺0�^g7Oe�ۄ�������_@;���a�~qu)El��ķ��i8�fo�u]�F�p��R<�8͟3wԭ�7����lm�_ӊY�s�֩e��׼���u3��W?�~J�:5�)My	^~��~��ƣt�K�i��S(��z/�c["��u���Mj� Z�p�kzt�a����=�����i���㨫r�4�3��uR�S�[��ڨ/?�%�'�� �3��ަ����G��:I}�9�S���+O�,��-z�*�zb@g�FՉO��2(���{G����*߲��_��}��N�M��/����5��Z�I"`<�m�/!D�**�����WG/n�qGn�&<ɐ�Pv`ε#t��-�ת簎��:⹲]F�n�.���=7(���F�/;hbG���5t��Q�ĸvX����3Y�$�!$������s��,���e� ��(�o$Wg�o
�5fG��XOp�G�q�������f$��p4�4B2�� �����nG�4<(!ڢ�]��7���)á�8�Xh��M"�3�V]�՛�|C�t���_x����q,�쉋������u
F���\R�gA�P�J���2��L��pK�ӎ���6{P�:���.yK��rګu���[WFn�ܑ���\r(Oe`|S���J�/�	������s��1���l��1�����1tDX!ݐď!H��ha���+P^r
�]��TJ~LTG���$_-B�M�ޥ?��:N�v"�J@�,�ú�����+Il�}����VV�,�.�PJ���yq�����t�b�l�z�a
t�w1Ʊ�(W�a��y��f� ����V����p��F�VA�-S�{�S�"ɟ���H��U���A'͑��N�.(�����8��NӾXrA^V,N��p�]��W�b�1����&���V��m8�	n���Y���f��<~����qZ i�+��|\��LሦΗ�ԕ6��l٭˭���ʎ�=r޼x�QEa2"K��m�jT�}���0�D{p_��4:}a 7��Ω�*Yl;�ˋW~4���N)�S�Ꞥ���V���/Q��/v]����ͻ0z��ty{�Jw�v�^��0Lz�!mu"�+gI�����<Ɛ�Iݛ��ƈ�#m=���:����eD!�kZ���H����	��AA����)et��&2�P����[�N'׈�/�s ��|˓Pf�:-�b~�_isͱ�%�����	@M�*�s:1G�g�:�Nݣl��5�3M��ҁ`9�N��񲍎�ŋv��z���_y�� �mjuҚ�#i[�>$�S����m�����&���:����*C�8�#�#�"�A�.8��~dZ�r�(�%_pD�E^郤=��UWv9x�i�ړ�V�lH���H�2�zx{���#���g��)!���� o�']X���+�,Xc{�qYj[���
3�hM�&�łt����1"Ʃ|��Z��DȂ�Ez��Ӏn9��<��M;7��9��)��FO��Xۈ{C�U��2M�?���A�����~�P���/!�^��{�m�y��^����
���!�+�s�x�L��7i���i�7R��*8=|6��ʻ 	��J5�_��nW~��_��f��4���%0��&3�y��W�- ��ńkdZ���\R�Ī�.H��o�,1p:WgJ^���E��ݰ���\q$l�l'qj�P����Os՛te<�a2��a�W�&������:���x�)'��q��BB0�	]���Z�-�`�%oFb4u����e
}�T�r���[<���ɲ��MǛn 	3N�>C�.����Z"� '��3�cOX?��O=ݘ?&W	K��֊�d��͋,�T+�g�7��#�>�~:8�-��(_ud�S(��i�y*!쑬�	�>�qg��E�N��S'Q�&�\=�G9av`=���Ё(yױ�\t첮NY
>)_���g'�C4��M@���?�<;����~�tk��6��+�������O4��<�ڑۼ�nۇQ�CU�'��)޽O�K](��OB��OP�nM�M��;L�^3��I�\ś��*��o��m�M�DG��lM�C��m��k)�C3��c��/�؞l���щ�h�[�~e`��m	=�j�Hg;B���4�E�PX�Rtʗw�&X
!#`
F�S�rL�Y?��8��R~T���A�OO�40ڄ���3�B�T�K�ܾ�QV����H+�6�qO:�)��W��WYO�<9��T)6���ܱ��oRҁ0����I���X�r��}#}`W'1ӎ|�Ag���<U��8�5yvjiG2�dv-��Sit{iG%3B�֞`������޷���8� ӑh7���0c���-�V���L=��{d{	��M֋���pdD#`n��2�rj푰	đ�
�漍o.�Ӌ����0`X�mx�r�l%}��0�r��I։��ی�)��5),.�J^��ԗ�&?Qlt�n�$�
��7K�y#�^��ۡ�0�uÞ(~�=B[A��7�W/x{��ܛMz��he�������|6/e�}��~����yh1A��^:3���Հ�¸)k$u'܄�Jg�GcՑ��6�=��N�9=׏��t��6Z"s�1!���8�a��0b�ƙ��: d$3"�ਟ��K��h��4�;O��NK�)�q�T?�b��� n��UO*��5y4��:QI/OA����'0�������n��M��68n	��-������!3�ۚS��&�m��	���P?��S�@����W�q�t���Խ�F{�,�C��1F]!���KF�C�=s*`��'��nws�6��c
n�����nh�cTʐj���@�����gy�L-S�����l�����iyGR
R2�݀Na�j1jO�F��:Jg6�i$Zy�#�v
E9�3��O��ݓd�3MK�zM0�%/�̆ذ��=o��7��<���>ca�����n;�#�}�G���~^����?��,��-:	`�2��0Nu���Q�uV(�D�c�������D�=��-�c������a�\>�@��y|8��8���]X���r�����w���u�>���:>�������Μ#����'����2�`g���tHRO�4C�-=�y6�h����D�$�+/�9H��a�/�<d$�o>n;B���پ-]em��CȠ��[���e]�,�A�jʼ��bk{�@vZ&*P�����5�@đt�r��:�����d:�|˩T���� 3_X\0ڵ��>/�I?H��r�ȗ��t�hH���k�(�H��{Q�O`��j�[�'
Ǡ����Yl�^��1���
��	�b�xa���Y<]<Q����a]TY�c�>!�ߩ@W�����%Ͼ��N���q]�aO2�;��;�� '��s޼x���Hޒ`��ޅә��]��M��V�=k�c� E��?`���������\�4��N��8����}<�^�&(f�M@�]�o��|����l]:E��s	6Z��!�>���md���P�}�
Q�e��06�*����.�I��-]���s�6���!��$M����WT�i��4e��L������
b�k��k�N��,�k�\nz�^�d�ϖ��R��k"��A�]n	&�p�,Q��!eD�ђ8'&&��x�#<HQ�T��7Hl�-��{陎��eUr���)���N�F���F���Hr}Z1B�BNל�.[`х�e����}ס�a��^e'=����r:j����9�[:v��'�l��+�E��� d�2+�p�5�Si���ٙ��7��l��F�OT�42�^�͏����+��o�t�SgC�	D^�z�ӹ�Ѵ.�.ld���#�	�Y@O�Z��o�2y_;�w�	���.H.����ϔHh�w�$��:xv/we}9	�
����|��t)O�R��,��+�,���-����_������5c�ПO� s7�Ζ�P{����s��"��Czڵ �/���,��R4~zzc
�@㑴a��ۣz��\4vZ��=�����u�?�Y�y�ΌQ��*/y�Rw8u�8�wO�t����9�ɹ�sW�?9-�WlR_�R���^�i/�N3�c�{��_ց9 .mX����X&�|��ԕqg1�N<��g�L'l�=�3C|_���.	���Q��<��3ټ�t�ܶ��`�]�=�<�����E��a 6G%��p)j�,/�\�CQhJw�;�G�!�=Dk�n�v�0����(A=�'�� ��-y�s�y5�^��/��2�f\�eģӤg;����!�tdǡ:+�C�NQ�s���#/�/��Upz�LI�'�k��1��N��
e\?��������F��B��#g���'�3b�v��RG��vࢁ�^�����d�����-so2j�u��/M�g��Hk+!�|��P=�`���k�یPi��/>���w���v��ßxM�t�3����+˯����Hs�|���Ȳs ڑ�k�f�؈�GYJU$���sJ�Mb�JX{n	��э֣�C"�8{�40�������-�SӴ��QY�\k�� ��9(W���k\�)�3�XFeI�.���(�O��KGD��{썘\@Ҏ·��`��!3��4�"���jx�|���!��}�{u�2*bS���x{s��}�N׈QՀЗU�Gݏ�DC]|M�Io�������=�z�H���k6$���E���Iri�Ӏxqny�qE��{�������;�4Y�I�?'\U�9���2���̷�ً瀺���,������L�"!�����_ud<��%4����z�nx�##L��S&�6A'��NuڐTX�W��Y��@�V񡗟2c�΢�>�iW`M�q$Ƚ�g}{W�Z�8�4^��ī#�;	�*'�K�,�V�؋R���0��)eQG�� N�g�#x�6��Ǔ��Y�����|�܆ܼ�n��c=u
��hS�esQ 6��7ZS'�0��Yt��fc{Z���B�3�+�) ��l[f	��'����\ƀ�e���w�N��x?���e-鸷�O�@T�DV�	�p�ǭ`�ݼ>"�]�g|_q��|sڼ=^2�4=���}���E��a�bT��4��W;d�G��kQ:@Y{��rc=��^�%�W|u�6�oN�ڱ �N��[|��7��lE>7���5G#���"�-7�v����m�Q��`�� ��Fft]��f��0�>�ַ�O��\{c'�?�[:��AԾg�9AT�P�P4z�9'dhGr(@�4+�1�~���0�		�a�H#YY7����d�TXT���p)�0�vpĦj0�9^Ƒ�l�*Uɴr��'�D�22=�� w��3��$�$-�,T��3xܙ2u!/F��*�lx�&��^��6��z��Ҹ:UiN�5nG��T�1 -r�d��(wQ���6î:bg,\=eS�?�4\��kz�n��d����1=�樝�t�eH i���1������Ǿ�(X�l�S� ni��t�66k�i|���Z��+\�P�ǰNO{��vL0O������Jٳ�0��׈��#:";���GeW����
�(��5�c#>M��d -}�`|�i8�h��
^�Fں,���'�3�L��Ux�-��`�>|���#pΆ\]iɚH���N��@G�VG
�-�I��vx��_�����_�0�C�y��i�׈��B�����^8=+F�.�f� �C�p�#�>�2�V2���\������9�-��jx��7��_|;��lo�zkw8w��	�3��K�_��`,~�a��~x��?�?�ȧKX�B.KE#_�ۆ�6:�m�{�<�X4���<T��y&��=�CG����-�� �z5t�����aa�>A��Br���Zn�uq^}c�F����:��zƈʅ{%Q�v���c���q5�w4̵���������V��d\!��]���@�𕛤l,\y����l�Ti:��6�Dy?@�4ܣ(HyU@#����ʻ"��GsK3�H��U�y��J`@G���76����L�M{�#��Y�]q+�[:4���Whc�&8y����R��.ys�^�ɐ���0�Mhɵ�dD=��!QI���7��������v�NH�;tl�љq��uj���+Ԕ�uG�ֹ�U{����z�y�y�6����DWO�z������Z!䋫#_�@xh�7�"u�����:'�G���y^�T)j�Y/��,𑰖�!��W�=Öe������6T�AVA�A&�_��5B���C	ɴr~<�(6�+��)L	�x�>Cw���2������3c��������N��Xd�"�:��s�􅊁p!A�AΉ&U��_˷R�����k��Ju���������K�SO��O$᜽|�4�(��BV�C�ɑ��wn1Vh�4R�5Q�|��YJR��,>�5iy���ʰ�X�"�W#��2y6H�$)DQH�D���[t5!X �qMbp"��܋�iD�h�:����~��������j�o��b~�B���00s�қe*?ejZ�X�D��e�S���-�i��7l�L7�u�����г�s�-y	Ў���Gh��O`
a"{2����L�nzNj��6(��C#���b*���.#_o�����a����hy����E�+ivT�^�&�� ���o6n�	:�����[�Y68���<�f[8NLWޱ}���v�q~�+�l���׿�~����%�p��E!���?����R)�ff�(����a��6cT�c�3%9!!��=d��S�)?i0 �F3R*y�K�t�G�%*ݙ�)�{���?�E�SN/���R�w��5��}6e�H!��b�Eg�L�mtϴ��<~���wt���b�oz9���Cl�z���=O9(��*�)g-��mfx�a�P�(sȄN�<w����k"�U�O�1�:#؈ߘ���u��l� ����e�o��`J���&�^�W�#]���Z\�)w;6��Y��ٔ�v�r��bg��x�)o:��~��[<��δA�g�y���BkT�r��k�A����;G�e �zd�k?�e+M���E|�����t�(��)�g�-�=�,��!���I7���G�H��
Q��n�ݩ�[W���䛛����[��軸< ��F;P9���E+�gd���{��@���W8�{�)��ً� ���K?���]#@�AiˍK	ě-a�6�g����IDJ�i<�2�@� /��`d"Q0�K�OC�)� [���x6`J/�
/��޺1�S�+n��6=Ɖ,���2(*���'��g�9�]�f���+f$��+�t��
tu�|��+_�x��5�`;���/��0���3�g56d-���CʧG�l�<�����=�JO��4���*�w���K�ٷ䑵Ƭ^�ǹ`Tfc�i+kbĄ���'����}�����(��Siԃjă$�����b���0A�`��0d�F#u9�1�RC#�4�� 3��ܘ�Ѭ�/�'8@O��f8x�:��&�<v���K��v�zꛉ��޲���96��n8�Z�O.2ft������Şm��b�|����ā�c*D��%K�#;�5šM����&u����O~��E�'�j��������z':��g����,�-'GD�T>U`9�#3���Ο� (yp�:_E��e�M�,��3�kF�L2��$UI�g��9��L��_��gZjM�KU�sc��eD��/�~#$KR#¯���� �Å�'��Oʋ{x���܂�t����O1���o���1؛��u�OOe�Yϙ�}!�)���wf��{�u�-�����yk^�/X\�˝<����d��؋4��1�t�C2ty橴�C�t�����uf�)�|�-��ޤ�G~�� ���-^f+w���O���0\s^V-j?g;Ѷ�4���u�N�l�G�E����ç�`�D�)��W���9�aߋ��6�������w��N�dVi�U9�x���F����2���(Q���M@3
?�Ѩ�7�ӆ	B�7{H�\�\� ցK���
�f&a�c���5�'�y7#�+� {8�����,פ�Ȁ
cǳH���L��#%1���*:��<�Ⱪ�!�����	s6����J"��0�T.v�93��%�fS\��� `/f�l�����]��M��K�7���5��m��o��܈�Q�����Ï���GI�y;`Y*��\�1�"��LA4�JA~��^~]��G'�4Ͷ[i644@���a�i������'n�jx^�L���
 xl���x~�.g<�nP6]�N4�x*�<�G�.LpX�%ґ�R�����l�Fj&#�i ��ځ�F��ɦ�m�d��,��������t�[n64/3�oq+*�~�Hfؼ���A8S��B��| q���7)<:��Iݷ9�����K����͌�ˎ;4٤������ �EB���F�Ŀ�`�v�)���?�|�/�7������Ǘ�3��@�ǟ~������|�_������X��(���դȿ�Q��[�ز���ѹ�A�UwxK�sx<d?�w�?�|�O�ss��{t[a��Rg�#]��P�.#�yO�lt|����:��6�1K���p{_���d``��"kG+l:D0�[��T7���g|��3^/^b����cdG�8S�c8���]:y_�r�öU��g0�I��Q>K]<�|^L��)�L:�f݄��x>���1��"��Ձ>��z7�3�̯�
�������)��p�����'��җR^����$�;�9@� @￸1���E���Ic[c֞��)��L�8�SV�!.���9��X��˳0	r��z~G��& ��蕜�w��Z;��̵ˍ��6fߛb�
13����5.eh�,ic�����Ww��Y��v_��B�=8(��C��� &u���\29/�dL���>�ϻ|L�&�4h���	�IE6 �:ʀP�Y10d���TT�ք�a�5S���z�]~&�V�t��'�+73���&�k�7f�T���0����1�W�E�qXΏ��H��i����p�Z��3�Qγ�����,y����=oa�i�F�}���e�C޼8�Wx;jig5�)�*7q�#�Д�(���@�o��xf����%eC&f#�׿f�^�_��M\{*Y���>�S���\҆���U��#�`��{�t�S�����j;�5��#�u _�o��D�w��B*S<���	��J����-4�1g�d�{��o�4�񋿿It��g2=���#�����^%��h[���z�Ob,�����љv���
˿�Of���ɬ�9��@�W����3"G,1����x#��.��=6�����|�w�y����܃6=K��ys�<���kE���'?дSr�������Iz�����dzÖ�z04Bp�����D�"(�֟zތ�F2%��.���]����ɕ æ���r�<4k�O�t�BcR�%�p��Ry��w����Y?��O��������s�zL��Y��ȣ��D��Y�
�������0d� fq�Q߶��dHa���"a�S��fM��5���H���;q�����
���	�N��{��O�	
�x�~�}x��ŷ�2[LYP̧��D�-�`�Rx����}��I��|�,>v6�����m�}�I�D33VA��bȂ�l�MF�S��!y��2 c���J��Ӧ�k�7���w�/�'�"/���\�w�eq���c���Lʃ�!�{��g �/��c��w� ��@���X]�$��␧|΀]��y;l۟���B��Aq���Ss� ���,� cf�ƜS�i�e��IW�U��Oc'_�>��?_��'a-TF����0���X��+�穤ͯ*5���~C�$q�2[❿d�?�B:�;�#+���2��ˏ?�"���z����ɰy�.�����WnH�[���^lAgX���h�$�� {�^a�0���>o?�ĕ� ��y����g�oF7�-��	iP�
L�K0����`�x�T)��&,�ش��m���ۦ:�m�(x&��ϛeY^$����wa���S0^y�6����u��ܧ�^`�xc�"���y/>4��@Yo�ӷJ�ؑ����ߖ��da��*a��S�:��e�K��:��)a��q��S��V�"���p�uW��B�dϘz�vu��Ǜ?�_�m���3��0cf�|�Gp1Ύ��	�e���r�����2��fZJ�v��v�v�K�u����y����~�aJh�7c/�uf�E/n]��B����!����AH�j�4��[�|2F��%�|�xyI{��o��]}�l~O��Հ���]�+��c%�0*�N���"�6��,D_�w��%.�e9��/�}��K��S�*��Ue�����ɍz�!^]�*��U�2kԔ��F��z����z"�kabܔa��H�>_E1�Gz����"��-g+�+ld��1ģ�4�r1Ķ��4RVʞ�̷8Q~���}����+Xh��7��Ʊ��N�fI�9z��Jc�������M�f�?�H���N�N�g��6%'��d��u�₃���4l�,�{���vq'c�Kbԙ`��R>�~CM;��}+h�k�t-O�����)� ��S3��G2��n�ⶈ^	�����qW�f�f���X�n�F�6�d.��@5�$s�?��/\Jt�6�I/ĶD��w�e���
�����2��X����QPFv�t���:�^��N��c�B���n�k^	I�m���Z��l�y壞�!�s����mM���]6�T����!���d$�$�k��B�^�	���?���4n�h.���,Q[4ְ�[��7B'��x���ӭ�I�-#{&p(���	x2��!q�M�	�5Yz�%a07���0�5�e���՞��+܆��VHg~��2C;3`��6"^x��H{֩dy�\�R�Zv��P�����s��**Q[_U6\�dmcG���s@�Q� ���/?챬��v��}3K)E5�ٖ,� �E�l�� 3��v�I����uH�x�A�a���7�0�0("����� ��c
[�)ȏ�o�
I���d�qw��7�?ޜ<}�y���0�]�X+����́�W]xA���i	S�I�X�Z^Sfޅ�S�)=�Mi=4<�F.�9y�Ω{�>��+eE)nΙ}�`�6J�1��_~`O,���lG��2m��o�=N���5��D��V���4���24I��f�k^E6��]�1��|^��_�@����3�'�>K�D˟�ɂyz��|���7�fz����V��l���2fߣ�F��[alO��{.�#�y:�!e�>��9���=娗���6�(R��P姜��bV]��r[�4Ml ڧ�㘽i�M}�I��L�94�֥,�'�0R�C2>�G7�81�r��SJ�N:i��W!
mxur�D���*�<_I(b\~�D���M�g�ґd�Lb+���L�����i,�\(e?���f���e��N�U�Ϙ�,~g���f���4�S!��2/KE��A���ي(e*�%�Y%�!�A��z-z�ZYX�P���e;��'���3H�;��T�oN��'t�y�=oH��R��g�L��:�&u�V�ȓ�V��4Iu� L�*��~F��V�R����C���wv�7y3���8h7W�,>����=L�Ae�c���8��Qw��|�v�,pClI�~g��  @ IDAT-�i��q�8�|��x�t��R� ���8���n��d�%�=��������;hB,�S��`�+O;�1�2g�ȟ�WX2P�m�.o��q�7�Y��Qg�/�3�"vD��F9QJ!���ӑqd�R3X�-��ig���4�o�u���l$�,�Aڢ�^P'�+e`��-s�N2���d:�[.�{�8��ȷ)��m�
0�2q.~�"�U߬�ݭ!�k��3x����ٙ;yK ��`��[�U�oF�(�-G!cX�$y���~�N�s��U�9��R���o=�w�{y�d>�����'໙ەO߷�r�Z��s�쳿�v��'|f:���H��dJ�_���Ыq�[ç����I?鏠��J�'�[��A�[ �u9�p)Ô��Ż"
*��c��_�P=�n��<:*ͅ��cʕ��`|���ʇ�i;��b�\M	?�M�H/l��c����S�`ڙ�Vg������u5�w�
���0}��`S���i�n��"=�~�<�� H���b��KR�@��z���!�n'���	���?���~<%<��4�xj����`F�W��D���QZf e@D�ۤ��Ӹt��L<���ss��P����8�>e}�?����ng���s��ӥ��ř��\�b=ʀ
�N�� �F��RfB�ԙq�ِ�#tfh�\x�Ԡ�(D8�ŎXb���#��뙴$����G��iYA�����~*��p��_[����y���0�F�>����
k��,L���5_���_q	�4E�4U������''���8ct���]�(��U���e����22,�r+��4Bl�pؗ;�Y���LG���p�!x�a峔%!�Ff�m���{hmGI�Us:�L����5�d��57{��uY*�t���eu5��2�J����*�)kO�?`�.Ǯh��r�@2h#��]^�>��wdQ�Rb�Q(us�+�Bo~Cѥ7������x���gͷx�	�k�=O�w�V#�J�:��i��I�ޖ�aSv�B�&l�'ަ�!q�j�7O�/�zʊ<yn >������.���<}�o`.��I:sbY��/�8�j�5��������7Y^����+��)�+Y]y^l3�m�m����^��ȓc�q3�6�.��u�ż���+G�v�#3�ޯa��F0Q�Sk�y��QR�ٷE_@�@������{Ό�w�[z���6K��W���0v(9�{��7����d�u�l�t�@�x��o�|×]0�33����{��㟼�n�۪9N%jݮ �bu�v4�/�-�uU'��!0�
#0:���4.�|��f�0�����,jP�M�A(-��}�m?�K��؎�N2��ϫ��V
�c2��f��&�[��ܸ��%�)��^iǷ>N�J��' 7��3�!�����ʅ3M��5����h*�wt
'�Ϩ5��	�ɳ?=V- �n%��ڊ:R���;��37�y�W*m��3ry_ٔH�L]�l�� Gu�AN�
�6~+|�NZV��'<�_�|6.��I���@�7I� ����Ӈ�8�I����qk�-��ԙ�(�T0��s2����"y�L��/K"��i�=�|�!0�U�t��Ci�rاLe��i��w�ق�#&#و�>kYy�U^�~]���:��R�t��bǯ�~���$��f�͆n�+��)q���}`����	��"̍�X��4��fi��#��q�[ڍ���pd�l�~�������@�Κz��7�������й�r�'��-{"P����
w?m��7"{���!�~�X���"S�A^>����r��{�>���9��.FD�	����B�S�xS"�Y�b�!{��6?te�Qm���v6�Q}�'�5�	�,��3�#�(e��l��"��D�8��L�����dv�rsv�%Eg�x�'_ڸ{O��d��oc{p���;f��7#;���=f��N�ӫ����"��װJ�g<^�C7d{��ڈ9��$q~�,v�x�������'1�����zlXUD��Q�}&b$Mx�nƵ�O
3��r�2�i	�?߰���)�3f)�`N�Y���M�a�3h���lC%ϔ��#-7�yv��2���X��-��q�zT��^�~���D����vh�hl�=7���c>Qv/sfL1W=���>n�u>��:���3
-<�0����N�����n�>%=�x��{oF���}u���')����M�3U�o����j@u:�l�z伥|0׎�@�g0eǂ��od��1���E�2�W�G��W'��}��Y�ifȚ�>�_~)��ӎNT�.���|(�>������8�G%	N�Jgׄ��i��c'ʔʅV��(��I�$<���������#]F/�" .-�DDI���+���2��B���(��Gq f�B5>7�LE�D%���u7}�3Ґ>>����5���7�2���j�S*�l:ƀ.�RM`=mG�%,R��S���l|�gysד�I#�x��\|�M��c̍�Oc^ڦր�r�	�D�����N�?q���B�~��Zxi��UY��?��wd���M�`�&�3���韲�Y"��p�9SϿ��#%�e���s�1�Ԑ���v�(��-fpvYv�C�
����H%2��t��SZ����
O��a���o2��ì�#�΂�<�-
Yy�d�������]��b�yj����$�ׯ+_������m���%�����af���ᐙ,ar�����7�ǅͷ��;t��8K̬�^�v�6drYh�M�ߏs��kۄ�J�?W�2�m�M�z'�D�U�LX��&�18a`tl��oҁ/���?����0��kő\�R@�6O��_��}3�9��ܤQ�_J78��t��C��F󖣑�����j}���ey�}�}����]x��Xp�C�7I���6�^2�������9�o�E4�*w�ʼ9>c��'���ᮞ�X�#�Sy����FX��O~���;��7����µM� ����o�z���aO�n�0'��þ��L�{.5��mE�Eo��-�C�#X�p(����?3�GN"� ��ԊT�f�ꚉ`(R�����	aV뼯I��'��v�M3S�_S�t�C�
��W�/0a>rt�����޼�{g|���]+�g��ӄWE%��I��PV��"����LL�1G>���l����;~SA�`R!9c #p�$)͙�6�&:���")p+>y&*�<�k�a�� �W�hC)�N7��v�U�$ע��<��*daB#�T޽Pɰ��92r�C#�Go�0#�T�=��zz�$��/e0��oAfm8D5z�9��h�4�9r���z���1�SU�L�/�y
��Բiy4`;J��d	~띳u9I�ve#/{�\��MN�W��W��o�2��JE�=���;�Q�P��g��S��S��6�
~@۽�L���m�|���������7���m~�ӟ2v�Ѥl�����ߑ��IΤ��o�	c��O���ᴜv�t�C�5��-O���D��1g"}��W���~���
ACׁ�I�C�M��ƥ��,ze�^6��n��_�� 3�������3��3A
�03��; �Xs�����
�+��<9���9se'������9	L�ҥK�� �s�yx�7P)�m�������t��UW�<@v��+���z��_|��ߙC̀Mغ#�� ���l�f�:/n�^�\E"��.��濲&>�b,>�{���U,ao!%�����Y�ª</������3ܼ/���yp��{��,C���l�6i��Y>�x��i�8#���o�e�\�
m&"EO�~�%_ 1��ǫ8���jg�"k�O���!�+�Sfj�t�y�4�/�ah��'���W��ոޚY� g�N�|��b��Ox����s�����Ձ���|�{�g�x3O�rS&f��-c�iX��9-CK%�a@��;�����{N7�X��٦��mv���>�j�fp�&6�Na��L-_�[�YFAY���G>��c^���l�.�W���iQq�?"}1���2"ld �v7��xg��ss�iE�k�c���^��H)����GX׍��)mȄ/�!>��RI�4a����1�&�
[:��!a76n��M�F������qz��I j��"����64@<i��z�$�Cd5�L��A���~�i��u�ƗF��`.��O�Gf�#/��*) �u��e�R�)u�ƋSܶ������#��4� �_w��<��+�Ż�	�K���8���5B�ȼ�˥*�lg��{ڌ9��`�Ջg�O�߼~�ls�U�:K�7_h�9�b��A��v�g�r���o�M�n�e}�l)���T߽}��OY�d/F�r��;��9W��Y�X��`D�C�3y�g�͠�P�~�X>���L;d��<�Їb x����r�z�@�!�^@eT���ʞ8axّP��)�Hc6���%E9X�*�l7ͻ�4\����0y�x_x��q3A��O��m��)�H�"r	m&�~������*[�W�ѳ|
��]��u��o;��g�j����S榩�,���pw���"3S�����l[�A Ղ4�j��`��ޫ	LT��N~"j SD�Ŧ�p�Q�덟��q쪮:�ڭ[~U��%�v��C�k�U�Җ2����q��O���C�Ϲ�dD&�NƠ�ON�1���ޠ��m�p�,�3ej~��P]e�M�M.H/g�������6���z�����@��½S2��;�Һ�Ȁ�� l�NQ�;�}���`��J&�y�*��4����V�Op�P+Fץ�����&�}������g�3	nt�n��UܷcZ�`3�ɡ^.x�����6�Rt3�_��ezp3b��H,,����w =��e3Î{�����s�qt#]R�,��N^d��TUIY��{<˳���ۆb�'-+�wqy_�,��?��M�sR�3X,ȵߦ��ґ��ޫ��a����9����#u;]��K�%���%�PYgyR\�Q7^UD����'�ؿ�{�g%�}��#�M������z��'�FE=���@;	�s��<�[\�Bt?�X�i�HY����OyG�x�Th�	�ٯ�\=��٪���u�җo��I�`���̘�������>�n��a �ɷ�m~`��+f��+��	{���>3�-�7�C+A�� XO������_k�=�����ϛ��Y�̄e����m8gѬP�����T0���h6��@ʟg];R�CϊФ�X?�˻������'.P3��qV����K]2�����6qh�	��z)���~���'��]�n���C�c=x�&KN��f�!�ȷ!��F�g�ɛ�.��d��H
{�1����6"dI�;sJG1;�^�Ɣ��٘��w�9��L9��!֟�����Y.���0'0��)㔑�3�q�J%B1s����¾�7O����why	�p?�&N�]�&����ٱD���s�i�Y�NÓi�e䀆�8z�����|!����2�����V_~{�98f@%1��ǟ̚�\.94�:���g�nv�+M�p��m��i�8Åd2'Du�L������3�k�L8mCN��W�G�[�)˙��;?��tM)r�	�p�ɨ���1��`�7(Y��j��	��ĵ��B�[289[��f<� �]O~��,���*�@TF_l���u̍�6v+�;��'_�^��R���ۖ�O߀R�{��5�?�?ޭq��x�I�<������MAax]^h`f��FF��aa�>0�ѤOŊ����4b������'����N��<���A��0�	��T�7zI7n6F�
S��ʐ<l��yF��B�R�/ B|�N��8���qw��ZO'q�g���ɭ2M�;��"JEt�ְ΄a�@Ŀ�Q�qe������v�u1$.����4T�k�A7�"_^ʑ{?A��)U�t�����A�檃:�,�X5{��:�t�d�B�����2su��>���8//ȸL̒.��H΁W�=�}�q��t8���f��>�|�����:��q���q����t�G$��V\J'�z&�>�i���j�ȍ`;���#KAo��R�R��H���4�f}ՠq0�t�,Z6�y�o���Bu ��fW����e�����2�mUqf�$��x�8e�V�Bm	�^s��$��_*f��p\+��W�+⁋��7`"+�3�T��4�	�b ��%x�g���[�_C��7�W���|�.��@L����Ac�(+���{����}����0�N{��W�j���q������E����%=h�z��V]��<K����'l�y����ε|p�����>5<8�u�ځ��C7�+�5 o)��K��\��%�����+�yT�c �R ל<r�!m�e�.�B���p�au�J0�D.�� s[m�[dI�z��r�،.�[鷼��*��eCtD˞�	�,�hX+֨<T߀ru�}!�X�{^4b;4g�Lu��0�?q���fp�mņ_6�^b|��X��2�F�
�i��l���9�A{���m;{$0�4�\�t#��3S��d^Fj�4.����X�����'Q[X��D�����D�����枵*�LA�9U;p�����[��f��PkM�<�R�a�8��=>�5�I�����nm�¶��	�-�מ�[>LU��A ��{F���)Y�U*'Ӆ.p�E�3e�ed���.;��ś�RQ*nԾ`�����0g|��f���l���K2چ�۸̨�0�� H��FZ��}�&U�IF%�"�g`��?��Un�vV���-�;�MT�d�%訹��(E��uкg�}���e�m���liGَ@���p9x�m�6������E��#�U�<��^�����E����{K6hKk(��qyԈ��9���拿��͗_�6o�9#�6Kz�I[��6�0�~�����>A�/T�>�Y@e�'p0��'����2�,#��΀Y*�@C�3mq�N��x�h(A&�����S��PWg]7�F�3���:Sy����������9:U7s��;��=1�����s2���`1���	��M�<�N�Y6#ל9���1�B�Ǒ���%�L���9/>ۋ�Ylh�@��h�V~�Y]p����1�e���G�ݔ� �@��٢��²�	�w�Oݴ�n�om��o�����G�1i�b8��2�#*�[��/dXKʆ����O��ND�-�y������P���i�p�2�K�g�o���ͬ�g�|���7]Ϣ_mD�gKUgA-5� �-8���������U@HUgl!�x�τ��+3���B[ �q�Au�=b;�>^�3 �<u����ː���P�W�58U�C���m��M�����,���^Jif4*R���+k��Ё�� ��鈃��QAf��F��6�(���_h��-�S�[y�����r+? �OɀkǷ���?r��g(�9�t�T/�l���^�}�4�{"v�L~���_Tl:;+{;ȡX#Q�,'��~�`�W�-��PHo�4:J^��ӯ1��£�:K���ٴ��v�>hn�o\���I�i1��'�o���d��wN�7f��ҙui�Y���f����1tƘnP�i,�u��/���]��r�,r��n�׈�I�:Z����2;�y<p�����C�4�Ҩ�����R���V����:{1�2R�m�6��5�WE+���)ڦ�<,��+�>�۱mT����ɺ��l	�ަ~~`���S�	������fc��ͼPg�����H�B�|0���Ӡ�Uh�*��!+��������� Pc:a�_�<��3N�w�˷)����%�r���K��0ͥ�l��ػ�<��p�F(��HפE>pI��̛��s�#�_p�o<O��.��5���d�I�,�s#z���(�e!;a�M�R>�}!�M�,�Q~���ut�|���P]Y�gn\3[������E�翗y�yKM',A#�8��W��}��B�y�튭!W�)�cxVG8��	�Cx���6�2ܐ�o���J���V�^�R���&� П�����n��<������G�(<f J�8\��� в�Қ��vʛx�'�C��F���9��##��]]�r�_�Oѿ�z�y�,ؓ�/����/��h��Y%>u
zy��n�߿�G ��;�g�*Zk��N�a�<�%�ɴ��)\�}�� �c�9q�KA(���k�s�f<�l�i9N��wVE��!e��}&Nԕ��0�td]Q���=���s�mFdJ��s��,p��8aF�-��њd�b����*�y-r�A*{^��`���03fW�,�D���;�.���Ե�ś�-#p��2���d_�y~�#��G������6�����	Jkשuf�8�q'3`�`�~���b�<��QYG������
��rlL+v2�xb)<aD't���F���7���?�r!���b)wC��/e�F�L��}q��<�'��Y��[���ķ��
/��On!=�VR�H���r�mCi�����0��递�2����t�X.�I�Y��n�t�x���6�-�rD��и�!B���(� 0i�f��5�Y���AK��#gv!g�@'6{h�1v&�<̢�E�l�r�[���O~�x,u��<L�,O��R@;L��Й�O��Tf�Q��Cģ�8\��v懫5��0|���@�,�;��Y�����X�+Nf����O��^�rF���|�[x"�Z���&
�!��>� {���,C� #�I�kɛ�7���z\���8oj�&�Y$���#q;7'neKO��²�a��5qo��\�r�'��z/��L����..�@�+��C�1k�L��J;BWG�_�s��Y7�˪ ��{�KW��)?���7'��C�^��5:X(�~U`�#��4����U����k���	%P�Kxq+k�Ǹ�K�W�����|l��AHg:����bn�/E݄Oq�o�)�8���;8"��,�����|�.�ɿ�����8aV8	zI�Ȃ���y��*��>ې	���Q1Ը',��'�
ý�Ϻ ��(����>T��$�i ��,.�j�p�l4���1|8�	��/�n�׿~E?���o?��e����57�g�Ƿ�:FG�u�7,o��+�����i�<�wW�(!�	 �&<휾�9g�����W�aY���7�{���ց���:`�O֩]��X`��Rh����m�sɞU�C��A�(F��]�%Hr2d(���ܻ����$� �g��Z�"C4ғ�7��2��9E4�����1�'dXg��;�S��[w9	#�O��?*R�(��ddR0�h���
���#�>O�_1:gyĥ��O�O%|����w?�ظ��eǝ�.����9�;lķ����pnWP�w}W�vH�&�e}&��ϙ,qH���.V����JhB_ᡁ����c:�p�w����#TZD,��>h��P�5v*���y~�SwF|���ydMKxdCl �	�"��@�T����*`�Ye��ȎO�F�7rt�$�i�=:K�=v*�9��jʃ Q�,����ۆ����v�h�ט�iALXER�KX>��Y�&�t	��_C*�<oy�����qx*�"'ՂӲ� g��?rV��q�lT�r�K�'j��U��2^�}-���ʮ�	Igj<��}o�ն�6^��VE���H1m���7�\������:3d~ҶH����w�N�M˥����S�I�H�5�alR�D�K8B'b�3D���6`��<	8��H�c;e ��w-#ÓC�-\�s����):���5����=w���8�z��
�.v�)F����P7/@梨�,F�7;!l-���1���S��-���yˊgb���9 0a�51)J+��X	�	r�B`�}�<T&�WO�8��*_�G"8�����+��iq�È^V������E��:x�!���S�F\�+�̀�I�R�ֿ�W*�i�R��ɋ]&/>`T��,�9������7?<c���<|p�1+`�@�P�4��ax9��O{��ՙ�����K���,����|F��wt��_�B=�Q�`�V!ܕ1��i�+O������sfz�͖P��v005�&��Ϡ�*���ڙ��,�}GY"�@�c�:S;�S B��`���^`I��f���#�����w�#�6�!q;2�W�"@�?�'���\�ãw�{���h����4�L�D����,>/e�h(���J���/�p�����,�^`|�����
�ʉ�_|*��'?n������-^m��ɼ|����pRc�sj��h�A��(_�#/N���)fĸ+ac��E�3~���#D���#A �Q��t#v�i��h�Y�љD^�MƯ2_8N��	�&}���5ݔϼG�3���G�&���O�Fը�����,5"�~�o[�����tZ�$��fR4<ӹS��>ڀm����Md�������y��dF<���
Ѵ���9K��m�
d��0��c7I+�d|�����|
4~�?�GzEۀ�*�<K9~�>MK[3��+�UT�P,�92���D��m���.oArr�mR���L�~ YJp��=�J�� ��XN��.H�k��zg}=�����1BZ�Gۢ{b�s���8J���g���?7���=��G�my�0H�D�i�5X-ƴmh�������w�$�;�PO�)��QWŁ[��/��&�ᶼ�l�����:�,6e�t��\�x��,YN\dFY��h��$L�3܎�0;���oz��Ϗ߾ڼ~�l���+Խ3�=�퐃���ep졮F�i��ݼ�5�wz��G���1�F��Y��<��^q�(��������
�EQm%aSB)�Ȼrm#����7h⛉*n�z׭��YB�-	G�LD8�H{��;��2�!|\��>�~F^�D��>�!�FQ�>*��^P6j���$��~��5�3����'�4�I��j7ʜ��=�lٱ>ʜ����cfV����x��p&��Gw�Kܻ�U6�9K~���T�/��qvɳ9ݓ}���C���ș/�Xƭc�������3g�N���=^��-��/�C8y%(3���:�Nf��rg��I��_Z�/��^Ύٺė�ȣ���+�	����~K{���'c2CZt��Ty<w����O�3e%�(����5�`�@
c!j�e���ϧ�D=(�C3�����Ng�T)*%������0�~�^������,�1KO�ң���Fx��l�'d�-�|�y���ޑV�3q̀�l��"O�f��Z��{�c���<A�w\��0����CW��c���/��[��Jc��fmp�@�
8BS��L��r[�L�W���ж�Jiƅ?qA+i�=I�nb�a�����&_����Q1�GŽ��tA,�q��\�+�"�+� H����ȁ	�Q����6:���a��0y����K:(��}9n$�LA�#+�v^nBv���]��[oB�?���#]yhd��F��,�E�$RvqKZ�Ǖ|��.e�`�=�2e��oÉ/�g1!Y�)�7�@I���@ҳ�c+����:ك���O�2;�M[.o�=�wG�^n>��_{抬�#g耧ϟn��{�����w����]�H}�h�G��-ƛysO^�Z�7�D�t��d��dO+w�5����MN Wo�SRh�<(��p��[���LyV.m�[�B��&�@dQC�;UG�Q�zL�L>�-Hgv\�rF�u��s���e�����gC�} 麗R�Ӗ�� �@o� K.���34�	P��l4$"��N7�yt�K9���]��f]#�.�i�2S��/���#;�$I�Xr4�� u�Tl-��2����|�iB�����ꩉ˻J~�e�K��V̟M>�G� ��T�F�!ݟ	Us\G���i� a�@#>\���#���ԣKW�l���,���1+N�S������-����<'�e�]f��`�X���if��E� ��^�eq�Ѽa=f�ΰO���>�Ç�B�`�g̊{�ӆ�f����1�ONM�����="�6���x�N@��/m1��r����%3ɗ<��-������x��!�� I�QfH�K�#xG�5�<v�gg�I8E�ʩ" Mt��%�I��"N����C�Bf ũԯ��Q��Pvw7�P���zqX"J��d�\�FOPf2[�v�*���Tx�2I�� ����&^o������Wߢ�}�;��^4� QJ��s�#��7�������BQt�PF�9��5&���\�\��J�&��t�߬$�̒w�D���OEU�4mq�z���P�O��Md�P�rQ�hiQb<�ۆ�����M��6���J؄��<R4�lN�q��s��,\�Nؔ��V�#]C�����Q�<��Bv��uǽ���������<G�n���ԙ���"�:�O��+�Z�S^y[���^���$dc*u�T:���(p�tK����V�Sj�(�kR~պK�$C6�"ct���!�
�s�l�紹;k�!�_�N���N99z�x>�zq���c��x������_=�ts��|PZ.\"{����)'�w�.��>���ͧ�����>�aʯ#�W�����s^��na�%���#�۔%
�oXZn{~ ��7��R��.���<�'�|[*�4垔�C�	k� �.F�BLY(7�Q!�,u� �e>m�p�'�*!�69	�|��LK'�.4o~��2q m��ssߢ����Հwo^�)1�@���1tH�{_:@P���̾�/�x`��T���c?z %#{�i����ò>�tf5`�{v��͓���!b#]�����[I$>���Aʩ�@�Pʐ��,f�Sv-�ϺI'⟩��ɒ�$l�R�,��5)��7����EFx�v�_	"L�^�5�	on����0�=%I)�?�?D��q��������Q��dd������ 0���i��	B��>ߊ�������6G���D���{�&��iO���!�\��̠����ca�ܖ�~�8�??fYѷ�;Io����?����W#���߽[�W�>H���^Ń6͓��c�Y�݋4��$�1 @��4�K�L8�@s�����<��E��\�e����C��i�7��˞6�&���~��X�<�n�5G>Vd���K�Ƙ�
�uVY�G�s���oq6x��\���>&	�ț�f.�x�LS�o�DL�7�m�ЭrD���р�@�
>�b�jUw��%������7���Ϳ~�ˏ.=:��E����_���X�?���k��������xb�NH밮Jv�K�Z��0�d���0��0��a\�f��+)"gC� ��ؖQ�.�#n�����G�9˹������\MXqN|�BM��Z�B�����#pb�N�?��-�_GH�Uҋr2�L�G%"\l�68��K[4ԼnO�VcNE����J� mF����.� 5��@3ے����lE1�l�_�YXl­<��8	5���~��y0@��	��f˳��g�tH�g�6x�v%h��/��tN�?bs����6o�<e�7Kd�P�Ψ�b�}�G��&�G�����'�1���1[>|���9x�0���^��/�́����#>����M��Ә����e�|t{��Of�0������c�Q�@Y.������q�#l`�or-�nͧO3T�q܅H'���˫�����9.�'�`�^L�����U���c�?v,�9�vN]�W\2y�4;l����w�pVӃ;@������Qw��D���#��6/W�=$^�L�»w�5�/�q�y�l�3f���o֛���Y�J���L޻u5��Mz�4~�_�j	�a 05a�I����������g@�����o��g��q	O� +3Ҳ���7�J}>�)�<�A	7�֬ЃFS�W�� �/�?�7e,|�F�M��n�x9!��u��ȁ�@�W�ް���:��Y�����l޿�y�`���k�xF�������p/��;��i��e��
<�&��oR[�Y>O]G�g��:�A��0����-Һ�f~�k;4w��4��+������K|���&}g��(�Z���}�Y�d��o�8J���+� E� 5#u�e����@�c�0�(e��]�!V%᠌��<hQ��0-�|���rF�6���Z���B�Տ�7�8�1�;Q|��&��C�`�.vփ̣`��g����V�)pP�~ʞ�'�^n��?��;�(x3�)x�}�a��M���,�kξ�y�a���wD��2@B
|:��I$���d��lKn��
�,��{�D:.�i����6�V�M�%l�/� �Ԡ� alй-���g:
z;���� /���R?	7���j�U.����6����(�_���$�Ә��V&�v*�i��>�ߙǫP�NY׏FC���5�(�N�I�']f��7b�'�W����yu��-\��J�«u��ޢ �p��������5G:���ޅ��5��7;;"c��{9���5!m��֙f;�Ca��.�us vd|����o����K
/�Eng8Gs�dxL�~�������o���K���!8����%����6�����!�_>�hs�3���:���^�z�yʉ��q����0�������H=������_���K��[x�	����W돇�zY�2���⡙�Ԋ��T�����啴�с(�����2ek[SV��/�W4�4�f@����C��zs��.��vD��z�8�0r3��P���^�=d�+���c>ςδ�8g��T�|kZϼ�$|d�}��DA�}r�Ðã��Y���Vg>��*�ٶ�~0���x������������=�Ə��r��k	mb�k(o���~BdbW�_���X���<�d���#o���1pM�w���T�S.�i~�"4��g����G�O���#�r+�&�ȝL�^�ߕ��"}�	��Ѩ�?�߆.7��9��l��=�ȘG���|���3^���}S�8F��mE�� ��>Q�m'y+�z���v��߿DQ���oN��N��<v�����y����pf�\�@�H��eyhv����򩇎}�����'u���gO6w��s�#��b���D]�#�'.�茋�#Q���WF\rĿ����d�!T��e2���r�af,o��N=�Ҿ���Sf�P��};v��q����ė�D��?���Lg�,�b���%�t�㏯7_}�d�g��~�HV.v�4�Ƙ��>P��PB�X����1�kV��d�p���O�6��>0�A25�ŭ�uҚ��!�b�I�Jl�%���gރiF.�t�3hhԄNԂ��7x����1�'�'�k7����}�6�r�� `����i������ze��S��o�x���Y���䄺Ƴ��n�ܡ�< ģI\r�3#�U^�*<��1��rYMq�	/8J|1�g�5&�0�{h<�˾��)��WB���k� o�����?xO�&Td� ��L�J0�&,
�v�&X��3�����̻��|����w�������"
_�џ���sX����6����nn����$��;>c��v��GO,��,�v���'��<�K���p�����?�1�t�9ia�R.��z/@��?9ρ�*���B��Y���<����ʸ�.�x�n��I���8�"�%=?��O���/�; 1�R�Z9"|��.�p���X��Z
�tK@�c��:7t�m^�p�A�wt�^�ڼ{�n��v&����,���63a\P���{���I�6_�^������[oQr�XF^lL)���y��Q�pʇ�ƒw�"�[Yo�M�M�~�>7zrj��_^�I�����x,g����5xF���&1��У#�~����*)� (�KtP$������Z��&?���P&:��%} ��Us�Z2���<OS[�D�gy�>�z����d�;f�hz���/}�gF��=V��O��ۋ�d]�]/#�q� }��S���y5M%����W�ʷ��mX˾e�f^��W��B�5��\C�A���@���  @ IDAT��3�=t[�۪�_�|�+��p}�M��n�� S���� �-z.�y5�e4����U2�4K1�V��P��%�pȳ�����hs�P��UN���tF˷�T�)Pa�@%MZ�<�y�M�
T�ѺgԼz�)�/6�˷�o��C��ˎn��G�u=����#N���톺3jL�Č��	�da���5��� Z�+;P��e��V ql��A�\�~��
1�(�@)�@VoБ)cfT2�� ����)\҈��	0���gv��P~�o��D�o�x���I�5���/�Z�
v��{�3���w8I��CҶ�.p���''2�r��´z߄Im���`�RraOE���4�P��5�dm��g(<!>�"���l�9�� �r�>	|�$�4|�+�v���T��z` �(x�֠r������AW?D��5�X�C�����10������e::������l����o����P�;f1���V�oE�|@�X`2�;{����>#�=g��e�@Bg�s��#f�<K��ǟl�9d�]�K�|}��Y�<�H˦[򗼃b1�@�n���ua^ ��:n�<ÛT-�y�4���O�쒣2eșlX���#8�����ٱ�Jݱ� �Y =�Y����x�YN�G6�1G��{���e'�u�O� x�FaV��zɛ��'RM;x���YJ�þ\X���W����I�A�{���V��4	�nq#l�h��e����*/�����:�\5J,��hLI�n��!�3z�Jd�˫ifK�.�.����X��O�C"�ű�e��V5F����v�j�G��w��H���P&�Ȩ�8	`:asO����h�.��]�n>�G��6О�E�' έ
���s�j���׼�#�`7��x��{�v�Չ��Q��0�jwX�;��>H�
��v&wd
i�u�s"g�@,���эƥ����2!��^���ұ��	/��z������N�ϫ�?��v6���GG�b��2��M�+�#���k���Ja\C�%.�MXo��Y��L��iLQ�*o�J�[��sڨs`#�)
2��%be���*>�����	ni82֠���S�a�������|��|����
�b�Y/��9,�����{���Q2��L�o�����֧ �F��͠��+�"п>��<V��f@�#�)��j�����r�	��M\�Q+خF�G@aC������m�֍-�Q7Z�>����^�]p��3�J~���BC5����nL�Gҹ@��s6 �9�&<,�Ԫޭ_ԽFp}&���&_�'!o���L�t����f8=?��h���v�A4d |ݔ]��@�(@�����5������|�@�Q���s�C>2+f�F�o�yb:׎zF׸�'``�Mh�#6x�:�-m�Ӵo���[g�sz~�h~� ������E^-7�Fq'��)3� C��]���Q�g�����0�|�Zc�>K�9�*�L+�A^�ǂ�@����	!�\�ZC��#FTss��oR}���9M9@��,��G�'��<����c�ɫ�uL�β�a���� �X����bsj�RQcL�s��\�����ׯx���;��;Y�Uv�g�
t�]v�Y�/�yS�;]!����\�(���r1�+<y�r܄��$������a`����Bƨ�]0�9�o��?�g�M0p���V,�i�Ev�M����"�[��[���Z_Z������#�D��{�/����^�!�h�_�Ľ&]}k`�4DDa�n�������3XzO���f���.��qrƗh�t�gs�Gh9������L:��7�6���硧�&���g��*� �O&��+d���g�l��x
kZu��@��/�Qn�q��ζ����3���%��cl�!1P�2�Lhh��%DЃ��%�b��(`S#�=
��}�m��_��)/���QZ(�$�}$��H ��NU^�	Tp�s�g���BC婀<�C:�����y�o9���'/���%���a��*>p���v������0����X^k�����l��°�@8NY�rK��I�D^a�`����:���L���a" a��3r����G��$~�Y��9��⹖ddeb�},-C�����߁`��ּ,�?�8���(�L��vTϒ!D��:� Ľv�T�o:�!
�D��G~�8���y�у�#*K3����y�9�-��m�h��3��3�򹖃�l��^FX�wJ�lpK�B؊�M�_�J;N��WK]0����ʡq<',��Ф��R��$'�Q~Ҥ�d���/�?�\|�#"� � �hR^��h,
�%93h���D�r�N"J���˒����<����A�BE�8�%����Wxߤ:Dg�px���M����r�Hϝ�!Mz(��o�^�}��i��`v�y�����\FQ�y̎�8�D�W%j�c���W)-r-P��a�)�<[����#��O�� �L<�V��B�?�˃YUƤsP���wV<�g6���H:�P����l~�^|`��Y6�5������;�Es�����u_��\�h�i��3&�y�%��>.�3|`�\i�����pg��a$^ Ir�L����+1����Yg�����P�cD��V��5�~�~!ƌ&��Vy����|��x\A����`Mh��nT��\6D3�Ĩ��e������`�z�8s�����m�gܕ�I�߼�4�7Ǽ@��I�g���d����x�f�{wx	�-T�E����Ŷ��I���Cbs0��^,�g�5��=t��m+�CԷ�)cm�`$�;0���:)�^߰�L��V���㋴Sb۠w�"�	K���M\��������.v4�@@sL�MeSY�*�!h�-Ô�4����idE���e�xvNE����"NB�g�8�ra)��)E$q2�܃Xɩ��(H�R3�~Ź_Ϙ���'���d����Z�%�c|9�����;�|���94|V�n����|J6�	/7$�,9�.���6n܊c<Ѵ�SB8<�[1��;���1�O S)M@��1�������|Z���=y�N'iWD�Y�$�=<	�[�I?A$�r1�q?�d"����`kh���F�}0
3�D3��1
���~��F�>�C�;�cFg�;|k�Y�t}Q<�S:�!��y���:�ڢ�W��M��$N�L�����r$>��N�vۤ胛���	�D�Oy��@�?K���T�
,��N_�޼��6���<`pst�^۵�X�N���,�UA�`���"fAR�Z_Ut�ȸ���t|C��J��l����F	
��2r }��r�� L�L�?ڷ��h����^�������yq��z�c�y�%%uG#�oV*�Ag��U�c\RO~��/�h?aE^#����8�@��0E5�ɜN|ҕ/�e̡�J1�HSTB���^�ѡ�2���K}	�>8���G��s���|'����KA2�����e]im;����/��\&C� r;�rS�f~�	� &�>��\�4�� �ǣ�uvٸ:e��g@�'��@@����3|ݏfY)(#�ff��CK���>� �,�2#�^	Z��Xi �20	�4�(o.u[�j2]��O�:��z�z=C5@��Nf�Hv]��'���y��9�Y������g��v����6�$�g��"!�uǺ�"�a��瀺}�2r��[<���p2�!S�4~�笱�G�ܖd��'���%}�L>����]n�,_�Y��.=2+lC���7�9S�����BOq���͘Q-L�	S6r��U�6���C�k�*�ʚ��8��%��cJ;���l͓��HV�� sWq҈����3��y�����c^c��{�^�`��5���l޼�3',Cbe_p�o��q��%{�.�r��1�vX~��0C�ó�9���+ڷ2yo*�����Y��[�F6��5~����o��!���Z���4<�X�0��"A4�$�fN�O��݊��26�a�������w���4
0w�!��5�[���k.���a|	�̢����	��U��!6&*���dm�.�uy��B?f����=F�v��^���z;��p�A��i�N�"���c5P���@n��+l�aV�SJ�;�	�?��K���ϣ!āOd���-7�-���$�����A��M+dD�y���9T� Ck��ێ��g;�IZ���/����[��}���ѣ�BE �.�dF�r(*�0�d'�MM٠��	`�yb�����)3ma�=�����Ͽ�b0Ҷ�-�ܓy�Z�*(u�ᐂŴ��]�M���4o"T������6���g�I���E;q7���j�]	�ܡ)]᥇��i�a�|:&.L�����-��ų{�ԝ�^k����8W.�?��϶��94�7���^���p�s�7ӭ�.����T�<���k����3Ӿ��s>n�8ˏ�;#v`;�<�F�kȝ0v ��� e$�̈́����m���z��$�Z�K���*�A�Du�ݒ]x�|��Ad�-tFR![y����UbfL��'�	�?ւ�)݀DL0�Ig�+��:`8�A��1���KA���&&פ���#����p�9y��D"~koL�xlf�/{��=�X>�;u�}זE��=ܝoBZ�.����퓙
��|�-��9�g��"��P��ݩ�5��A��M�Z�0y0�������q�����H3�nڛ�U�9�&<��Ӧy��t b��!���H+�i�}����5I�c��To�I��܀)��,V 
E�2���tb.��ld�%��3`vD%�[�6B�C�F5�ăSX91�F��װ��#���#Ø̪'�3v9��e	?O�Q���Lg|��{�^d���֪S�l�¶�.6�;v��i��:��G��臶�o`����[R�a��+p �Kc":]��z�ܟ$���6
�{��,I�� f����S.�M��/�-�����D�<q-
<��,���d�ְ�n�#,�1��$�b���F<�S@~&�'����`��"�BJP���Ɍ�H�C�&�r��E�*#d���̮^�ʾKg��0�j� <�௑e;�|���0UN�㦠�ζ�@H��<�w�.�S�	_��eAXd>��N�8���B�\%Ap�#8F"��rXf�TԦ��c����������_0�X���$:�8�:KӜ�HJ~��K�����G	C�7�~����3���ޮ�O�r�bo����$�B�<Ю�\�Q.��3<ؗ��N9bxEgq�؛o��<��?2����˪T�0�d� -sg%���&��)��*7|�a���;it�?�R��2'��!yқ��J��)u5X��1�Ɏ�g�h�)�ěd���[�N�:�C����q>�?:��܏q���.��jR�� �\9�<�KA����+O���,e��o}�+̬oɦݏ ɲ?��6Q��|�k��޸��0ϫ,�7q%��t�E��g��|i���G�	1��o���22�(
P�L��>�G��J�-��ߊW���l��M4�Va���T���,FK�x/��`_���k�|ڴ�K2����I��o��3�CW�����&pF�I���.��+w� �%>�	�\�Ja�5�>ǘ�[��(p�S.��ن��ٴ/�m���hj��E}�E�����F!��[,]ݹd��ps��������]��05���Kصz���gv+��F�3�&�(D7�j�Ȟ
#6$�Td��_�l�3�t֯�YC^0����������P�Ga��X�2>;gs߹Ɣ�Θ1*�(M�{ʮ%G>�D����GN�A��O�˂�!	_V��e�3��$�u
��ĸa���o^�k���C��|���q�U�"�<R�`%DŢޤ��Z�Yi��P�g��6�%���5�E���i�u�F�`�)n�����x��薴wKK5'�����΢�	q�~���;A���c�w���t�P�=����=����ٕ{�Q���Rp��S�c�AX�G��b���N#%3�U��uyF#n�p�o:�B��	Cd�R�Wf�ҳ���&kZ[�mm�KChe�7�G��i���v.�7�������?8m����?p��o~����Վ˅�����p�գ<X�����M�:�Q���ޏFsF�Kf�^|���=�6yUos�@�����_l��	��M}��̈:CDB���#�W�ֲ�w1n�3�.���_�?��y��ā�?d�.�]ԟ:f�2���4����F�	A��������@�,9���S�y�֝��i�څ���c��M��zk����*A|NΧM�c����k�d��9F�[V��{�\v��O�/?��JA��vR�o>,;pJ׺�>Eu�Y��s��La��]���L�j�%jq�*C�3.e����#ƭd�|s%��k����
ob�ǫ��Yv�b�������O�W�Oa�=uV��"�X�(�o���G�-�MD�7q�g�K�AW�ҧg�%�2\�h��d�t��FC̃3R���
��d��P�"�	{�/�-)�|r��RGINL��0���<�k]���~�9H�|~���i��5a�C��>��F�_^ �hO�S̨cs J�P*��֣�Ǽgy���s�����Ӈ�S����kަ�����W�6o��s���8-�(��P+Q3b�ԕ���g񚉬��W����!�@:qڑ�.U�t�͸����	^���b̑ޅc���ۨ�� ��$�X�\�d���e!�֧�̄�;#���U÷̹J;��hŝ�֊>q)�g@2��BǛ|%����4�7���Q6�
�4`���G�LT�Wej@p�(i��Jw�%�
�V��l���zO���G\n�!Ϊ�-R��<4|2A��3���jyNh���,�CJY(]�݁������l�M-M���|ڇuT������/�.�k����<ɯ5^�xyY�!ގ�M��������0��d6pН��a�w�
'3<�ʺ���o�O�x2-Χ�O���+;��Fr,=S��5���fj��3���/���sڞ�ruugVfe�6J$��y_�T���)���� \ �gG�E���Bw��p�8a��ȆvL�8D��>�̴>��.�ₗ�YH��8fI��%[v�m��:q�7D�R�����ͯ�X��i��C�wO�Q�gK��S����<6Je�v�D."�0�7�g��N����O��z��Y���?/>���b�[�g�Lg�ox�U�igd��i�Փ�XF�tnZ��d'��3�Z0���Yǧ����
�7�J�c�z짒��ڟ�e� �C�$3�S�� ��إ1��p%�{{��~�ҝ��ئ�y�F���v&P����b¯���M�r.�˗p���ﰥPE}��!�SJKK���Ux$�gmG8� �X����/PbG\�#u<v�܊���)4-�b2�}VPaG0:��+x�	 ��)W`gd�S��1���7�8b<���,�qG���IR��y��T��HB��=)�� �%�;Q��<z�ƹx���|����ʍne-H!�3u���C	6ϙA�'�)�Gid�N�I�	��UCN�x����W|���L�ޛ�/ڙ��{��)��fh�nhѠ!ub��z��fI�7�f���>%t0&�'���}�J�Eℬ��n�8�����C�DD!��B?'/�� �N%���#; ���K���sec3��g�9,CX� �h����*G�U��D)V|�v^�L�p���9ӓe{	Zg.i��N�w��F�.���l�9�y1�3]�:J��/�� J6�&���f���7`�����	Y(���k��-5��Z�����@՗+�Y��){�\Z�14��XB+7����&1���y�L�s�p��"{i��}0n恞�L���LL�9�3K�@]s���0�	mh��k~��[�ߐ�/<ץyp=���چ%�=y�D���������<+�6Ɍ���5<�	�ʡz)~m9`��8f=j�΀�15��Gu_�y�)��Q�؆�*�A�q�0��+��#a���z�yJș����yL�U~.vW�4,y��yC0��){��sxxɌ�3W���.~���k�fѿ��?.^~��4��-�����>f�z�32���5�@�������/Ρ��Popʘ���?����7|W�ǐG����m>mTˏ����i���#���8�o�q�7�7�������ݰ�6��ZV��O��EF�;:?����ʢ�2X���/�<�b�v@�@5�-2��B���y���-�zUTy4C�/��5r��x�U�6�]�s^��n�<��Z&8E 3����7J�A8���+���}��/�;�-=�Y�qJ����\�M&�����/��&�[�.�&��{n%��G�k��c��[��$3���=r����ԟ6�}!ጊeN���u�����g�2�kE�t~r� 4���2�Kt�O�0fdLz��e��(������ĉ���hgq�ц��;�c�83��"&��ۈ����n(p�^��bHz�"ԎS���1�-�P"m̲�Bx����h�(uҵW�Č�1�bIY�tk(߈�F�k Gl��Ҁ����.�rN���6~�!u��;����>ZL��ꭇ����7d�ǔ�hZ�Y����0�6�5 ~�D:�!ױ�p��8k��ѧi+".��c���M�.�ۉ�Q�)��'̕��@��%ڣ�-��T*��5�u|"��Iv3���$��/��� �!�,Fc���!�3�b,��V �
�z�7m v:�8Z�Gt�̗������t�q���!A��B�I�-����."�,ab��zE�|Wy��(?��7��N�*5�
]*��:;�4��id�0F���bJSJ�z���3��ӹh�!}�ͳ�B��,�őbfc�ȡP\ΣhA'M��H�{_�Q��Dl��@h��a崓��s�L-�߃NLP��9�}A��\܌E�[A�|�2��Yi���&M��F��1�獂���6 ,O���&]�)�Kf�jA&\���L%��N�gIw��gi�1%�+C���� {�и	ҫ,�(���{�JJ{�RL;G~/qX�����z9�^�Ns�7��{�z��Z2��<Ko�������Ѱ߆�g��G���'�!�~qN��ۆ�����C������V!��G�oV̊��W�݊"/N�����Ku䑚b�e�Z�����ǿ���'n���E�y��d�l}�Y�t<:����q,"�lWq��v��@��Ѣۆ}E�^8ٶY�]�M��T�O�)_V�``ж
�f��#��,V���I��t��Ga�2-�xmU�ղ����>����;�},n]8G�^������Y<���Ƽ�%�9���:V~��G�-@��<���6@Q��]�u���C�z��D��A�&�����LN0"���$�K)�ۨ�n�??8c���Cx#���HVH����&@��l� �8�h��枏T3W������}B�'8����/�Q_�۟�+}��L��k�f� �yLK:�����}���rK�#� `��.^���������13]�~���u
�a�(�]����x3�%o�1�r�gF����l�˚�f��ZA�� ^�͟��j���E}(K��Q��,K@lT,��8�����%��_���F���49`_�- Dy-�ډрM-oy�3#ў�����8L��ʕ�KlB
��
�+(�#F���Rlb�����Y>d��4�����ř���f!�e���T�bj���/��<"95wM ��T��C�Z(|0J��`��t��I�*iK�^5�KhҘ�����>(��+���ct!zM:�m��?�&�������<��y�	ݳ�5��qmLG��&)�p?�LE��0_a˫yt��������(�WJ8�XQ�T�b���	uԕ�����ݒO��O}�X�F��rK���?��٘�VȣK�i��Νz��9�"ξ�<�I?�G��k`�W������A��	�7��9K��2��m�h8��쌷l5p{�����u��_����p~�%q�6Y|�����ᗟ�lipΎ�>��E�=��Ɍ�W_���?��ٖW���֒����{�}�6�C_��#����]A��o���������b��AKp�^�H��7��~���K�N8�3F80����v`J���o?��O���������I��������m8��;۶���#�3�;�5"\S����:�/����Xߪ}!��iñQ�&g�V�A��y�(�Z������:���?ؖ��'0ĖN�͵�vN{��r<C�&hZlՎy费Q�U�A�V��k���6�)�݈-�O�<���\��KWس3 �����.��d�,p#g��M`�:��ڠ���g .��ͯ�㨘����y����^��)yo[3�ףe�Ųț���3<�9|x�}��(�0��2o�R����o˷�y��c��S�����^���q�/�A�v�?9b��}�c3�c?�5�`���U��g�^�N;i�)�8��)h�ʁC�k�R�٦pA(-��O��Dtn_�ma�N*PG0H�:��93+NYlq�T˷٫Ce�z����(?e�&>�����A%Sq��q�� _V��;֓�M��EyAK��o8@_:3N�Y3u�#�b���ct(�у�s>�tdf��#j�`ǒi?�O�3I����3ם�1�?�F	\D�����4��`���U6����	S0�MZ?|xXN�����fh�����p�8e�d,��W�&��̻d7�F�{�4��`�zb���a[�׸�U�4T�}�����u�����A"�6�0���Q8����/a�6�Ƚz5>�Ly��s?�pdJ��I���g�C������F����+>u`���ýQ:6�O;
>�O��P�+�9��Զ�,�Z8�Z26�ď�E}edc#0	!��>
r�#���Y�v�M}�:��%�8d(�fɲū��X�9�h}����D6 o�rM�D��������q�%3=�>d7rE��:D�7|ؘ��8{��
��ǡ�ݰ�%���V4FG�V��q�������/��g-&�<a���͇Œ�[��my����Y�u��uB�{���#8�C���Sd��1���_7~e��=��7�G�ǞO�|R�G��/�\��L���J��0��woxT�I����m(�U���Ro#'u)��9�Ge�`�J��l���n���Kx����)��ߨ=D��i��xp|L�ߍ�	mM�I`0�#4�:�}�y�gU���&��۶��Ƚ�eF�v��`�%P��B>G\�"�y�`l~�,�&�ϔ�S�S�%�,i׵�� ��lDZ��_�v�rr�r�{&x��A^��>�8΃_�իrOP��{L�En�OFЉQ� ��Y�G�	d� ��ܧq[�懂��,r�`�Pc���^{�#^��2 i�l�c��f�cN��Z��b�0{L�zá�]g&���L�N�vH��h���R�G�Y�4JG��Vɺj8�)�r�qΑ�(��-6�ݪ�8>}�j��#b"N
!0eZ�e��޼J���q�]D%�n}�fD��\p�42�_с��sf��v$�C� ���q���UEޟl]嘌��la0��Di|����-Rr�KK�&�z��a�8c�[L�L�x�l���CA�=��&˰� o4ri����ę�Nk6z��C�i�8_�k�#�(ؘ�M���a,d半�.����0���1���̐�c���)�xa��3�,`��a���
d#�D5��M8�>N.޵�h��H�󅬴��2C��^�#t�J=�6'���y7Cc���L�\���9����AJ_�&㔁�<�/��h�/���9�6�
�!������\ȷd}{�G~'t��`� ��	�0UpH���G\�B[�0N<P�
��{l�����Ip�g{�Q�]�`�ԍ��̺��|�ݷt��APX��y��������*X�rY*W#�qjg�:�ڒ�h� G8�:��0�$�T��l�l�a�s�bn�R<C�f�8uj�3��+�{����'��ݷ�oyx���N�z�3f̖̤�X��a���%� �ݵl��,&�v�y��-+68{�]�3/o`J�5o��Q�rq�L�W8{~j�/g,����Φī_A��el�2�~�lÌ:):�@c:]B�S������[㾈��x�eJ+�G���`��u��afd�6���1��Aa�}OPr����V��J{YEk�I�e�`�����1�gF8;��ɸ�DL��:m�ًl���_\Jwfd�S��]u�욵����u��U9okW�#;;_��<�J ���W�)� c��
��E.�Fh=W^՛4z7��n��|�>�L
���k\�B��u|�T\�_!$Gˊ��o�va�k#5`vhc�ƻ�1� �s����K���N��	_�P_�l$�ǯ]�in�*i����23&ƒ�K�T��4����ö�3m!��@BK��c���G�ԑ`�G
�
���6:�y�Zo��-��;:	VJ">K&R$Ȕ7G���u�+���+���=q��м��G����U��݆ź tM���V���m#6{0�dq��F��(��rq���b��mc"ma��<�L����٫��k`>�jI?��+:� � ~���"ou�,ſ�XD��N:�^�̷�t�ҁ�z�rZ@�;	���kA�p� smTr��
U&~&�����,���k^��5�le�\\Wt���i�|BG?Z4�"r�K���ِ��GB.N�����o�=��@oS+��8+�A�g(��Ƈ���:���3��C��/eK�ģ�d�;_�GL:�����SMŦ�Xޑ��c�m�뺓�zX9G.�g�\zz��Zx������B�mn68�9�V0���5���($�ؤqo��:����3�s�q�q�"$�V@�/�`3��??ѣ(D ��3q�Q�&�
�sA��-�<���I��6=���$�li��H���/������%1�l�$K���v,X�ể:�8^�A��5��6���O: ~oҷ�q�������ʂ�^l)�f�t�С��� ]��k��.ܳ���yu��w�7,�y�oI�Z���?����! }���m��Tn��cqLy:^�m��'��m�OF��#+��:<���̈���*'�$�Ag^�E�$���NT�HA�)�v���2��g�!��~�S���%yT=hh�"uF��Je�C�S���K;�2ipV����I�E ������?e;��7h-]j�s��En{eIC�2��0r��O�@�|�%�pO�җ~�����)6М�?�%����gI-�2��1�Ǳ�3��`�v.��|��3��8Z�pp��K�M:s�oS�/n8yB��6b (i�m�xm��o�k{$ťi�7�5'S֞DT�s§��GjY�r턈�D$^*C�xX�{��k�!.�	�:b�	 ��G������0��ŮA�v�aY!����-���R5IQ^L
]U���%����@A�+����������#)�� R�΍�DcdPEٹx�Y4 '�Ȣ�QI�o�cd���2FR����#I���)�Lc��4?;|$�}:Tx�&�S'ˢ���r��I���9T��)TA�Fg����}�1�`
C
���>'z0G
�]�r�: ך��on��I됹���oQ�y��bXc�X�����|Ls ^���F�,�����{Rƅ�9�yzi�=� 	���;+���X`u�z���c�?��7�����J�einZl�ї̎M�)1ؙ�Av��(+�=*��ړ&][Q�s�h����1o?������Fup�g݋q�ґYv�C~l$��bff�yz�f��(�C'),g>�� -���3�;K5�P�O%?�.h#ʃ�'�8�d��������~Y�:f�H�n��G7�C�	Y3S�����<��pF�8'p�����ݬ3��"�������w�cg� �:������L#�N9q�.�$��8?�qǢ}i;��8���t������j����V�n�b@G�^�@�+gW}=>ߠ�ޙ�Ά9��g�\��K
æM�F!0�9�R��� >����L�z#ho�j�#[Y��]pf��2�L%#�8����y-�sf��s���6��Ƭ)���rM$,q�;m�Y�E^?Ɲ��hw��5�:aa,K��Q�pX�������Y�l.Ni�Iɇ�#��#���)��}"���dʙ��?���!���u:SHd��s��"��'N�	�b�gLΦB{,3����Z>\�fe�qt�Bpĺf?��'}>���{ٿ���5�qvv�x������X�z��u}|�Xߎ��\<"&rѝv�^()�P:>u��(��V�K�tƧ���K'xZG&o��VF� ���z��sw��t��F� �)a�ɽEE�\�\�F(~��=^�O��R���"��4�G��L/4�D��7����?�3�,R������Wôs�������.���yў�I	 ��#K
�`a1r~3Q�b��y�7D�1�1��gύR�TD�(B1�7���J��ZY�c�I�8j"d$m:`�MN���y�)u��U�)q)\P%B3X���H�W�����p�}B��{�0>��g.��,��^	� �@���<rt��-_���_/oiԁ=Ca/�=��#�1�|�f��錗�;fT��;+y�j=�-�#u�9��JS��I%O�F�>�Ce�����!ס�����8a��,ׄ=0[,Q��ĩ�4��� �>�<�N3�=W�6&�|\kW���ށ���v$=��q��9��bv�\�90#�iE팅K	�)-TL-?��a��e�|��A�d ?���L����C���M�'sJ��P�"��i�#@i��｝x
�t$����g��4��\7$BX8[�MO1L�ou��{v��)k�R?KOlּd�#ppѱ���_�&T/~��G�N����ܩ���Գ�m��|l�Ù�u3�<�������Ĺ�B��sv!�E�=�fq� �bM֨:�E\�A�M�	��-g�7��`p�x�|��*g���8cf;��0��6���{Q�wF�r�jm�hW'��|x �Rf:E 2�6��MqA�����a��g��p�^y��1���=�YG tP�)d�y��+n��Z�Neu�e � �m������4�N,�#���MQ�����DM3��i+�ýrɅI	ZA�Q���-,a�I���	K���<nMNv �6���@Kv� S����%�Pe�%u�k��z}A������g�3�O8�;�~mz��-\�m�[��-[�>�����i0�,_��u�f"qI��W�#'PrC0�f��0@�k�YL��)kȏ�d��Y:�E[ӯ�e�:�H�o��+q���k�hJ:����8�����;fA��G�И~<Ԭ<b?�9�+}���^�-���p��sԓ�.(�q��4�FC����Q�� �%��2*�@ �#0��5���Sj�U&X���-l�H�iB��`DNx�V�pb��c��ͯ3����n<�Rq�$%N�i����x "0� ��QY)��R�{-?f���r�댵%�����ϋ���r?P��������6!��c���Q�-������DQm�K� ��]G@`S��x#��w�<40h�~������5��:c{�mS���z^aB��$���@Sn���a�lb,�-)�ɷ�p�8Z��9r-��*<�eRq6��śEN秃cKw����V6�#��g���ƌ=�xv^����Sq������J>�r���q��_��j��LF#m~�y��������y��U�̐�)�)�$(��Am�c�����4RҮ3�Aے�a�,��YWM�� ~ivv&�B��_�R��>e�s(�Ӱ�T�Y��^�� f/�L�eJ�2WN>K� ��ƴSʍ�A�c|�̊��5��A��t*j+�$�sf-���E�j�.���9�w���b���gCG�~X kڠ  *LIDAT�šÕ7(���탼Bm�]��e_n��_n��8q��|L�_����t�*_X�v�;C�c�@{r��ܫx]���ȃ���������m��R]�F�fO|�r�,��n8����E�<�T��Y�N�����>9�eZg�����o�\����[�U�'y�gy�5��/ι}�0ѧi���vI��Y?-G4jJ��?QФx)
���`�g�8k�)`.��#ho�Ѥ%Ñ��4d�-]�`�<� r��WxBfh8+��T���Ж}C��=-_�M�������{�1�-|��A�oJ����o�r}A}���]1 �I��:�\Ә�3/�%
xe�`8��"���;2�8wdA���|d$f�)W#-����?%@b�|s�zg��'<TH����=Y�I�l�&g	^�zax�Dnȝ<�~H�0����U�=m�;�ѾNh��=�����޼�#p�y�5P��Wa���5b�j�R�x-ى̵y�!ȼB�?g�#��`�V�� ��)�r$ �
_�r�i�(����16E͜��C� )���RR��D�O�rcNe2��Eh�5��BSg�\,�Ǎ�~]��]\yOG�f�o�������|����}^��\}G�z��DǽD�΢�\t���lBe`e�*��/�FH���+�x?d#H�y�Q�ʾ�l�If��ר�����M�u���ׇ����IcM�������`h�j�g�-2u:8�G��p\�H|L�GB��C:Uv���������*؋����l����O�:i�u��,EQ봸/ԓ3,Yl�5�1��Tp�T���<zɬ��R"��,���_��2�0�=��3mjXl�z��������a�k�"���I�ٺ�kd�}��kZ��6!�*{��H����V���8��@���7�9?yq�w���A"	�J��}b��N`=���z�.<�ulJ�7NWL<��K:!�M~`�/}	��3o��ɃT�<�Q�����y�H�I:��E;&)�Z,c������r�R��A��R��X��ppptT���Y9��S:m����t�����	ʧ^8�u��}��L��H���I^��N����_\��s�SҜi@���\��ϰ�: S��Dy7�A��*Y�@h�?�JS�uUI�Y�C`�grYg|a�q�K���2��x�N���@�Y�� �sP���m��?"��C����K+1�Mg�������b��bC�K�����x:�qdփ��M9�?�q%Z����	���33MȜ��E'`f�>:p���C����q���-�s�א��)"�;�&�~�l˲*e�T/�{ʋ�{Ԏh+h��b"��*���r��=v�Z1Q����\��)����5[�/]-*0�J��œ�7#Q�iD��]��zVike90N,A
��0�D8ШF���I+�a�=�W��A�eW�j#��kLkY)��B4�b�o~�K���4s$�ye�К���D�&��V(�� ���U�pGr6�+d��Z�+��OQ�ߟ��+u�xԵ%�Foɣ.���KF;g:`���FKeR1��4(���|{&���I��	MT�yo�k�gБoDpJIS�.��LJ�ا����ɮ�!��B�i��U>e��tu���A¦�o>m�$%g�\d8P�K��8S>&V�KXm?�>e��0�{�)A/�����t��e�:�3'��d�J�5����Y�����0�G�I�6���ˏ�����YN�e�4�q�hg���quN}�0k �Vf℗tbF����`��U��j�	�"W@8=��F�t��D���>m��M�Ȕ?��mV3�o�BFYn�;�����5'T�S�[?]�0m���3Cv\�x�3te�$K�C�틺�i�5�~;���9���2��ʠ��Oڥ�#yeM��5�Sv�#^�s�6��!���v�8;圗��� ��k��܉�8q��<��u���"��h�]��.�Θ����g�P�e����3�Fp�Xc�Bv�TZ��\({�c�����E'9m m��4-u'��i�J��M;�H;6���#��y�d�3���Sd��%n�I�ϙ�Z�vVC��m���U|��%�$@s�rc�Z�d��-s�;�7ȁ��׌�i��q���b{�#�v��\I߂D應���lǂ |�������.e���3d��p�(�M����<[?|7US��A����%D�Jƺ�}d���y��[��l��8y_��8M8��>�Kd�F�R��]�S�7���e�F��<�w���>hY�a�	9�P^��p��9Ƞ�vw�Ӻg�%'�~�X�3|�x���oZ�b�C&S���G-����(���u�u��~�.��%�(2�&�Dɤa��VI�z`zr@��&��\� ��X(�(��5��_���J�l��E!�:��4Mk����#�y,�+cs�u�9��D�3��o��t�'��r�^'�/���z��K�n^�c�ҡ�;o���o���X�x�
C\f�t�:B��M�ya���H�4z�SϥZ)y4���O�܀U�#�����<{���'>��%�4���mJKM��w�����kMMVg��py��Ǝ
�cTV~
�&��ʽ[��=���|{�����k`o��# d�@aA�X>�Il�n�#iӮQ����R�9�"��&s�^`��?�*x�!���k�3��'|d4̛+�Y��?����}�c�
�L}��5P��Bn���.��,����><����Kʤw`�,S�u�R r5�x��{��#օ�b!m<�H{A~�@�vC��s�y�y�,?D$D�f�B 	^�G;�dl-��s��6L��2At�䯞��zb�@��ë��b������BW�Sgi{)�@���ZZZm����2c�C�}���q&��G��|������ɟu���HG"�c@�K�/�),�6$Y���kC]��t��f���'B[Ҿ�NMy�]�����/�)Z2�@�@�M�&�%�<eN�3���r��}�t����Y
�@ ]���G2��S�������An�jɮn%pO2����ٵ����B��7�B�
^�<��v�d��}�%�Yv�V��tˁ�Cֈ��#�W<MY�-�����;	�̾z��l�W�K�&�4��2�R84˜�������3���̫!�~ ��2,����K)-"�tDrhˊl:o��ľ'UfS��^{�Q�svf� Bp�t(O����!�h��-OG2*�&a�m?�q��b���׷o^.�����fo��y#i��G4:[���G��oZ��>)1p����J�q�X�C����A�ЉN�3� �_m�i���V�BP�R��?�%kI5
?��يeIf��&���II�����%s�����~��8��y�'.�F���]���t����o��J���k�ƣ������X���Q!�����o˔Ύd�^�@�dY�9��
1��6p��֫v3�L���Ů�o5�R�a��.ex-���z8�#�'WVLi���>��Q��cc�c�����6��U2��t��_=����`����O?-~����O ��x���5x��� C	�[����c��S����wK�S�6γ���egcl��3��p�������0�ؔ��AXDq|b�_��|{��y�������8G8a���� ��1ΨtL�B:(���K$y���툵�:�Ú"q�K�$�iʫ8��NǬ�2�+�k�H�n��N=6���{���"��=�~X�N �-X�B����>)�gʳɑy˓~���Y�-0�`S��Fr�!�6`���ն���]ֱ)lH��P�R��8.+fQ}�*�O���ZzC<gu�����I�Bi�)����1Ηߵ���5m���؇�O3ays���h�1dy8}|���� �;���q���{���`q���|��G�w:dOl��M�~��ku�2 �Q:'�
f�nyM��f=s�����8��M�^������Z8b�|�C����2AQ}ki��)���;��78u�` g��۠;�5t@���nH'��'��<�7S�����Ƒ�cu��7�-y���
�y�AB8�>~|��|�~�fq����G��-a�p��P��؇�-P�]�6�EۚԦ��pR��'R�``5m�H���J-�i&R��6(���W��;$ތFZD������60�	���سr#�6��Ĭd�uh�A��zm�u�`i7���9��.���L��⎙�OT�P�����]�~\���4��ϱ-?|��0�r-�$1tvɕO8�P4HgXP
%Q��t�є�����A�"��5TKx/��_��li�F�L��⦁����t��N&nK�EMDK\<x�U�b�@%�a���U;y�&�?����-�<<�?�k��gY= ޸�`&��X����O<�:BY��M�M:�j?t|���D~$�W���{GC���d$|�1�>�6ʌ�?t��-�-����!tr��w���� ��yS�	ܫQ����z-���%��8��8mB38!b�׺epi����]čI�Q"k`�y�r�go�;Õ0;K�������??��o�/~���|��)�,Ч���NAˡ@ʉ]Zշ�L������1����2��`�د*��h@��Y���I;S�<�����֟ʭz�~#A��_��u�MGŊT��A9sD܂+dl��*fi��c��	��8J`6�3N��Ә�l�W����_��"��,�;c�F���%��ї��YL�YM���ǂ�]�^$цS6�}X;s�DG�C&�^��]��!YލX���J+gaC�"ˋ�<�9I���,ИY����G�h3s,�`] N9s�u^0����!�{�v�/�? س�Z;�a�qV>�KE�r�R8@ɬ�8�S��f-��O���A�ْ�x���C�J>��6#�,)oڡ��I�n����IG�����->~b^:2g�u�\G�G��X���l�W���yf@� �cf�t���at�4 ]�'��E]~t�8dzN��9�|�y:�q4J���6V#њ��d(�n�-�Z�t�2b6^Z�zD~�e;vd���KO�OA��C�;@G�%b[��iC�8��h�����Q<�?o��w�e:�s:�+:}�â�W�\���f�5}H߈�>|pd;���#��ip��q�]�jݲv�K,@�p�"N��6>lQ��d�:����|E��DZW��"q\#E`�Cґ���mS�O�������WG���#���dv�8e�m����휎�x�!mq�ɫNƑ
��w���ڥD����^��d �5_�~���o�^���Uަ��|�E=������B�r���ޝ��y�!���Û)<�+,�Ά#��
����o ���h�@��@��s��A�`\j���#i�����8����)�K9�\,/>��J/N��y��yxmh��{�f�d*v�.��5�-���}b���^���j{����,FD+*���˼A��6]Z�Q�X���y:����7�%�HA'IR��)��8��K�p�U��� QoO��#r$��?�9��,H��g^���,Sx��̈́��4�|��/z���?�b�T08M�
��@�=>�-�٘��,w��`���K�{F��a�/6e��l����t�x���o2� v�}�F����9wР��F��������9��F��1�_����kfXP����.j���)�hG�FYeSvF�C~�5u������C#�qNM�QS����w�3VY(S?�<�ڐic�C��93Oq��IÌuwzXz�(�}��j�3���U��6l�U���!��AŞ܊Ŏh�_;S�К��Fgo�c6:�r%�pN�ڂ�Ȇ��D��n�#�H05��"���%�Q�[�H��_v���D^���#�v�ά�fl�)WU�U��Jy��ox���9me3$ox���ݵB�C;�N��;o��=�S�0�ہٞk�:ʚ�m_v�3�����TҔ�) J�䵎<�6e�<un���4e�����\����ҋ�ϔȹ����gəez}�-^|C���p�6�g~�Y{S�ܴc�^<�Ð��fK��2����"�-W<iv�9��ٯ�\����.x�~P7v��O�
�]��+jB8�G1��?\��#�pvՎ�����R^���m�?���M���v��9+�7G��v|�l䧏}S���5�7�8�����Ҷ���g���6|w��x���>3�L�@���P>
��!�YO�$t@"�����5PT�d�AD���݌ۭ�3G��M6�2��X۟�{�ZG5�2��.ɹ�i�mJCA��C�m/��s[��x@7>W��n'��*_��kMAJ���S���C�,O֯�10ڂ����p^u����1�CΎ�p4�y����_�������8`���}�ݷ�Љ�a��c�z�|�'���6��Kc�3��Q`V��Ĥ��Hk��Q��D��(1���z�A�?�"�#A4�J6�R�_�y�B�5q�f-D�j����\��W#dd��T��v�GZʁJ�0^[��8���+�B7eZB1�F����a�+�q6��菆�]�Y�w�t�������ѓUD���%��ۯl�M�s���̢a�iXP��49;S�9q_��[�S^%Tnc��s<����`t��)�8e����K�N����!�8���X�]��7���ī�ᅿ4�T����F~7u�ଛ#�3�T(����f6�-�l]SQhx�QDR����8`��vΎ]�%��O4Z���)���H������]֩	�A�?��~@���.bԡ\�(�/i��>�� �g}��}��8���]^��.~�c՟��#G���3�0l_9Iw�{������F�"^�$�[|����s�d�1�*4�M�8��
��*Ӏ��$;���=�%��!+�w����'h�PVt%��H�	���a�)~p;��G���#����t�_�0����߆��]��~����KZ�8�ҁk��83��#�L��;�ヺ�ɝA�־{Ny�M��c�i�����T�K���7��z�tG�i���I�:)�e��d�-ĀTmm~n��5n�������83��r�.W	[�r�'Q;5�dfx\�O	��H���Q�
k��*���Ǌ��2�M�9"R��#S�"���N�Yi�>
��i?�o�8��ԡG�mg%u���
�����V̳��Ou鬄pjϴt|�7i�c��;�ș�m�v{� oV8���E�~zFGCGByE�r�eZ��|$�Z�k��~j�58�b��j�E	��>}۵6�n��GZ��c[�u�>�#����POEt�|��]L�T敻�|�-|�U[��٤��f)u@�bv�����I�N O�u�: =+^�Yv&T;qЩ�5�\A�pq$�ML}�#y�j� F��Jmٖ�\���˳�����A�|�O�}�K)�^�Q���Pf� Z6�>G����������D����R����gnO� �C���o�ÿ,���Z�x��|�'��_�˾ߕ=���!�^��>J87�����
���:x}y$��0L��Ӑq%0Q�,~�UvG8
O�5(�8�!-���
i4\�G�Aۘ��O�t���\�1()&?i���>��vh�m�T�ę'Ό��$l��ʋ�MErsHs�s�gC�T���g��O���hd���oq���b�$�-4:*�8_�}|���#`�a�3���� l���6��UC{�9tDү{�G���~�������i(��bC��r�F(��\�8:PXT
�K[F~\+˰av}�8*�Q��ͨ��a�y���!/m����=�(�-qH��{����p�x����-��B�Y8��A�a��8��8�7��}��I��Gw�ݤ�١�ʧ!S��**�O�훝8��V׊�c����eq����`������-�����\�N(��u�6}�!��x�C�Ҳې׹��*oEW3Mg��E��e+�ryd�'��.ξz�ˆ�7��v=�h;�h�:��E~�;[$L;���"ę 1�FS's���}eǽ����]��W!�En�؀�޴ÉO���x�nlh�{�k�>fs���������
�:��؀r��6lљ��y�'�vV%k�,k���Q�kμ�pVP>�ڤu�`7���9p���[���,E��De9�� O���b������as~���!4d�P��϶Ⱥ��6��9�,��r;��#{��ޯ��b���P��I^<�I�w `�v�BOf��Q(��$�ʑ�^u��{�(��忇ylw�l�3�
}�i�c&�R�(J�E����<}%=�g�;�����"/�8�,�ڕ4qJ�I�%��t�g˫�UV�L�l����dҨ�'?u��;zx��:�.�[�%��K۪-ESb��Y����G�v�y����o f���Gm�K��(�S���5����: ������N�
�v��'m�ɿ�2�OW���5�u�z�M�*II����K���<-ײ&]�Jq�z&M���>*;���a�Q�^\�#m�Wo�,���]��S�{���|����{���5/&�@hpl@�xXF�Yy\�i'��f���(���)տ�T*�7(4�ʂ��˼�F@[!K�Tf�KG���ťbUZx���ct �oi"?!N�ʶ �9�S���v�TpN;E�M��-��C<��)N�wƮO���Ye(������o����x�\�"�NUk�i*��Ɵ֟2lA����Q�AjE��+$���QǨ��^�v@Vi6��V�C_� (/a�T�;T���b�he�F#k9Vh��a3Hm�X+־\�7=mD����^҂��	�]�G�y���8`q���*-;��������0��FV��Υ#Uq�����]����^G�~T��aE��u�00P��Z+;hb�����}�@��v�,�_�9�1xx�C{�>�Ϛ�n?�c��t�i����Ӊ�#Ϩ{�_�:J��Hg�|�N�`��u���v�Lc�*8�2õ·M��.A0�����:@�s���u)�7Ζ8�-=�]j���|�K�E��aQ·�9�M:���`��V���E�����A^1��!��,d+�p.�8b����dv��	�p7qy�S
�uW�:=�eHl�2��~8�:��B�����I����R�tD�[r��:�!P#f�5�5dlG.T�wC�7y�>V�����Qӳt�e�a��&��K��cyҞ�V���[2�u��_��88_�}b�GNೝ Aω-��SS^�K�bNdQ�_k���J�N��XՁ6sB���%�I�����/�N���!^�ڷ�i_R�&m�w�Nj�LȔvK>�Gt*�@W�� m�^�D��M�T>����t2d\h���y4V�X'��=�9��x�|�_��A���`RQ�%�L��}I�C�C��:�FO��6�<�>�x�w�-^y���-xl�#���խ�Y_m�cg���^����A�~lGt|�8m/u�`Q_Ca�ׇ0q��Kʙ��
Xl�P2���<�t�G^����I�	��p�'�Jm#��6�E^�����1�����%�]:_�Ϲ�� C�N^�����y��[�M^����.���`$@�C�w��Ӓ�!4
�w�ʢq�Ph4�dR���@���Zy6��gp�UO#L	�ā��U�p�@�Q�Fn���X{B�K�2*�
�`K�H�xk���c�LzKW��b�-y��
���ؤ�x�'pQ$r�Z��P��r�l�LE�#��`X��<�v��F�-iCfCXK^K��_R�u�CZRI�t����7�=t���üY�,#va�K߆�H����j�6�s���~.�I�,�xq��yx�ڴi{nz�(Qّ��$+�VFe�;�V� %^=9��[���P.Έ�L�|�t�:;���U�8:iL�!�:Z�mx</�>>s��������ۯ�_���u��ǃ�+/˦� �	NHt�����A�,J�:��X�m��)�?����%rUf�Uf6��۴����UG��Ѧ��ȩN�K��HÉ�
g�į}+���KLU��334!]8�;��g̵�ktrǚ�#��2�6�5&�̐�wN�Ǩ�jݠ��;l��t��dk��x�Dm��t!����xK\�h��c�)�� o���xYA��Mj����hf�iۦv���K�Nz���g�u�q*�<r��5T�-(4m�?)�f�ʗ�߲�,���m<�Q��":xR�`���iێ]R�z;�-D�%��a�w��A�V�ڕrf�-�b#�{���.̗!���v�^'&q���ɯ�U�����7�q�n����P���"O�d�eV�v�7�3h<�}q�.���-X��+2D΂e&,�����C�S�L:q��c�̄h����#�I���98����o�S�qd2S먌�L�Wa�% ����*�5��{��~EH��T&>��c=R���J��� ��g��A
v��Ôwi8�Cڴ��������Vڸ�oȗ����_�l�k�+.A�Ҕ~�6%�!{e$_���/C���I���f��M�+�����:l��	��S��?�	i
�$    IEND�B`�PK   (}OXإl˨6 �= /   images/734bc482-36f4-48b6-9076-7f88fee16b3e.png�z�W[M�u�B�"Ŋ�ŭX��Sܭ+��x�R��k�"!@p�w$wwr�{�����dB�ZÜ����w���I��ٳgx�
2�Ϟ��"_�Xϑ�|�yk��m$U%�=�M��3�@���E����3���J�s�%�KzY}i7+s[g':m[G�g���	q��������ҸT}���QQFR�'k��e"�+� �����ӳ��,F꬚�,��Ʌ�#�hIି}��b�z�EK
�DP������b�A�P��n�����m���:eW�ν �>j�Y�>����F����"���0�Bh��'��KL��w����ۅ�7@" �]�����d�dr�!Q�/�Zp�;+��6�͐���ú�t#�ENR��90f'Xo�H:N(d"?�φXs�u���y� RB��.��i^�&�/*:�g` ��@�7����q��X>��i$��4�~��VH1���J6L[<�w��bH|l�����W>��#������:;>"g��_�%��wq�s�7�"6��&<�����w.I���"}���M�׶vΨ ��Mx1�F���lEf�h�59\Α-c�_x}�����A��$5�5��w?�oj��"6N��_�@�o��5�o��/(���`�Qo\m�:]��{�|I�(��M�r�s{��;O������
�	��&�'6�-�}�.(t(7R'-��F\T!�8�62<	���}]I	KW=�c�WM��pE�7��߽:��H.�k�;�u ������6Pn�3
�~x��� �S�Ťvl�)睝A,�ԟs�$l�ӔJ���#�����^�߸����Ň_&n�ܰ�g���e.S�3����)��w� �އ���Z�˃E�y�r��C��c��a�C��Hޡ�,#��m����DY��bdbSN�h�����`��{G�@v J}���5������^Y�f!͔�����M;T�,C��itu�<~�҃���8��;sp�y6jӖ=�'�͋������E�"�ע��/�~�t԰����K�}U�a�x��'ǲ�.��+v�=
K�{�wTA���y	���"ȧ�'�(�}F2��i(Ac�V7��Ѩ��ӗQg�*���+ZlF�'�m6�g5�����±#J9L�����,�!���#���ߎ�V�߯�u���#E�O8n� N�	4�_"��z0w��,�E���^{�C���K�SJ�þ�[�hTN֮�O	�������D�1�i8� _�j��}�ˑ�]�٪�8�۶�LR�{�<��x�����Q6;=�G�/��t�u)O��|�]�uK��9~�ps6��]*�" %���������`IYF�Ed��:"2���e�ܳ�}��x�{bJ�3��~�|.
V��6E	��A��F��x#�^" Λ�0�򸨃��5�&�z�LGz�:�הi}��P���Kj��*ٴ0Ǳ߲Jd���{w�K'J�/��0�
�8��d�F<�xX�%�&�:��i��_09�C�����H����
x���>|�sj��(�pN��V��T��BQ5�}��{{���_w��'Q9��:iu8�m����H�
�_�泐!��wj� ��?>"����&�k?�^�{�q�ήQ�k��ؗ��q��>5A0�p=����d��`ݔ�Maۚ��c��)���xҫ��T�6��V�]v����v9*�¢�B�h�S�U�I(7E��a��	�i�v�$�hp�Ĳx����z�|\��q�D`��p��:����c\�Ө7�%ٹ�b(����|8gFh-��W�����dA�^�D�O�ФS3#5l�p�y% ��>Y�N�\n'v]L:�zo0F��F��a�MFƑ3��<�_X|Ll~e+�:}m���t��Rc�����DP�� ���0?���'���'�����J]�셿iU��1�j���^�w�I�?�ޞ��k�̥�\>�N&�ʚY�Zqsz��
^�a۸uM��	^y�}�����K�:�4�Z�J����x#�a�{@�wV����U�1��P����T{����n:�2�׺oU�]G�pf�]be��6��Fʾœ�;�����L�����	�������Z]���J?iڻVˁ,+
�)�"\��/���xŨ�l�aע>	fZsr�
r��B/z ����k����MQ�s&%,6 �;�
*�F�lǷŞ����C*�pr�2�z��i���z�����ƈ0��|�7��Z�6���j"��:�v�1!���멚��	
`�_��i���y�@
m8>�M��d��`M��uL��̨+���$(dq�Q�|���J^���(7x�����3OϮ�{khK6D5d��̱�zU�Q<�<h���)����k�"���V¼d���jh��I�k��o�65�Ww��tť�Y�^�9K,���Χ=��J���AL������50m�~�����l����� Hm1j�S/�[(��S�?1��#��5��gr��ۋZ�}kA���՞ 3ׯ�����@f�I��E�����&����[�VB�(��A��qR�[��L<�Å��	�NNy�|�p�GJ.����D]��Z��U����#�ǪfᎺ���9�yV�cg�'�@�M���֖՗�Pc��.���Neޔ��sl_���$(���݅��bs���W�M_�S� w��:3�\�f̽���0�Sj���ME�J��|
��a�r�㱹�UNbgO}�()9���翠��d�QJW�"�5�2��,Xl2P�'1-��d5�&T$OXQtT�w[�d�T3�{���� uTֆ-_�	ؠ�'��4/ֆ���u�o��h8ؖ��yQ�x���L��!բ��j�4�9�V���m����c�6����7�ዔ��zGyɯ����He�"��v�f�y���r/��V�}��l�r�n��ͭ=��H�0@�j��*E�A�Z�k���-�s�6��"̓d�8<f"�����W� 2�T5�Es!e\PW�+8�"�w�;U�Q��oqyC�#����Z��D��Ѱ*ܫ~gmə���!V�g),��DN�F�/m98aǅ�np~s;��h���/B�.��'&��cT�C@�=~gR�D���1�90��^�T��gɚ*˼<��=�ё���B3h|�$�7�0Ba?�h�� p>(w�;�嘃�uRS�}[
o'ܼɐE�MF2�1�'�����2�Bo��/�?ֈ8����e� ��Z�}��B;U����\�4����R�JV��:�3���4������+�| ;�)�Lƕ���٭����`�n�DTj��i���]퀅��*�P�$"b�W�[k�2>��6�b���u���f�I%�.�Ȫ�5�p����=dQ+���7��Ww#�ijdd4�2�𻁰& x)6b�bG;d�-[L��MI�X�������o/�Enk�:�����Y���?���$�	��X<^��'TX��]��.T�[΁���zA�C%#�*ĺd=�{x$~D ���ҟ��Dܮ��c������;�"#������{hm�4���]��1�)8@�x���V���6e�V�KmDӌ`|<���>��2��Xzw� �K-��5���#-s��\�(����F������F�Ƭ������.G�֋��?QF1�Zi0i;v��|�|�
���tN2=P[L�ݿ�#/�3��5�/�iJt����G3�Ԉ/h�ݯ�W3j�����=k�v!gq��!R����V�#���	c����E��J��Z��l7�f7H�I��� ���� �x��\���~�>#Nv�pi���aS��/hA{�l\aW�#������������� p�\�V]J�Q���� ��F;G|��H$Ha�e�t�#H�Jj���6��җ9j�}�8aʭx����cp����lT#�Y�_R�_
���8~Q͒�6�/�H������h8~�*�k��WH)&��\�[-Q��5��=29��l�%����m҉�6w�-p|��]R98�nR�x��6Us��й$�Z��Z�(:m�ʙ�����Tg&����G�ru�%�L�;;�5#�ݎǉ�Д����ۥ�&���6�d��>x�����I���y�3o<��4{_p�]���<
V��u�B����L#�\ĕԐ�g��\C-_��P���u\�S�)�JR��D�Oλ�`C;�}w���D/���&
-�@d<$� Z�;4bY�®��y������.Z����$]Ԩ���{>>K��Y�Mƹ}�?ޝ�"�u�81�_j�*^�}k�O����\ؼ1��tŝ�|s���G7�K�w�|�=�4i��+���ʾ�ޖ<R��E�gG�x{}���\����X�N��W��A�U�!T��gu䲢l��`Z�"I�q�|l��iU��b){�QxH�s��Ԋݦ���U��_���Ey��Eo�~��b�Y�y;2d��G�,FFtb��Ӟm�/��yImEh�Kp8IXa�*��Jz�W��e�{�޶'����8b�4����J2��O"�GX)�B>"��J����8��_�(�S��ң��y�\�Oq�˥)�3��P��3fd�X�
�MιTl�K��T�;s7���I*��g���[!OV>	�����X2��x�o��>�K+M޲��R�C�����W��]�I�XA��J�;BCH���-_��dѓЫ0��x�Q�F��O�F&G��	��k���8�Ϲ�|E�\�[������`��9��f����a�Ͽ �1R�; ,:���B��Ff����rOՅ��"Y�rv�F�3`�g��ӎ�o�{��� �T��*���H;P�~��w�Y@.eKj����IͲ4X5��$X��ݴ*90��x�,�,�]��]9ѹaj��1I�<� ~��z8��:���q��f*�j�$Xy�uV���m!�iH|)�#��hIY�Q��'��ɘ�N��XL��X�c��8���o{��Z���}���;�}�Dn6~u
�W3Gq+�I��|8����$�l�����-�tx}+�t:m�R����)	�����)�>��/2�<�����b�OKw@�#rH�r �� ~�erA:����vڷ���b���b�k��W��o�������\q�*o�����'?�3��*&�0�����wq\�\񇌐h����yzb�m�gn�Xn�/,�xt��sdyM�6����ʃk/�;\a�$M�#�ϫ{?#S�?�ܪV�JX�6��{c�_��1�3U�m��/3����"��F3��t����P�i�c��錫�ϱm�Y奍��#�
��&�(L�eS8��ؘ������4,�Q$�w��O|%�t���a�Zz�B���)�_�3�M�K>_Ҷ�����[ÿ̣O�����:�e��HK�N���H��Y�[ɸ���.)\X���RX���|�0̠dZy�N��]nlq�(�hD��o/��j�e���~%�g΃�����]����=���FĶ���p����r����|�gL '5v/�gc�����b��|܅ qȬO�;�Jؒ�L:�8ҹ͌��y�ث�����e��+�"bmO��^E��}t�Zp��4O�3��SR<�^��lo-���/�7K�,�Qd;2r�a0�Z��x?�.h��3༮����o�p�27k����:���q��F4N��������2����d@���I�d����@��VU�)ϬF�������"Ȩp�9.��t3DI��)��We���l�r���U����P�w�/�廚�ØgH�DN-n�W�:e2�w^+4Ȓ����l4�&��A0ͣ��#TE�j���y��?8ep�w�|��@pu\^����s�z8#�շ��{wc��TzO����ޜ9�����r¯	�S�b�j=]�ֆ��l�q��Q	�������̬B^�������C�)��Pe�Q�&�©�*Iw�нS��y,���<���k�0D*�YvK�+і�H�$�1��
,T�\L��p'A~��`���q{�ned���5. ��A��0kZ.S���0k$�w[��n�k����H�phuc\��N�U޼�Mb�%d�w&�x�I4k�t�ԙ���kK8m�7�F`��uJ)B�N.��"��7���`ӄ��-5�jy��h��ч�S ��������,�Zg_'S����^?�z]Ž�D��j�>�fx<��lS8���k����O�g��� *��kq=h��.��|�#"�S|(�~������!��Z���U�m}�B�&|ܭG��;�g��F>8�;x@�tb��'{�'���Hz��ݟ72��\b�čE@����Rj���R�1�`qαm#^�QG�N�����32�b�"C�(�`S8$ ;��W�v%�F�u'�jj�����L�Z��\FKf��n3�6��ɴ+r�X��z�g�!bٖĥ*�#�{��8=i�W�}W5���>�Q`:�Û�U!�}�$G�޸r���R���w��f�V��A>1��!�v����b�Ы_z~eP}���d����㻯�WO�Ln �(Ҿ�p����(D�v\BE������}n������q��Z�0,_jc�l/�e�w�
���ڟw�}�*S����b�u���|���./FE���� �!����{B��5��C�;�R~X�]��ɖ'6��#)m��5��FfSǾ�-qI�����X(޲���6:�7pmCA�W�+A�WV�������.������1Caȧ�?�lX?�i�<7%�Da|�+�`�⾲R$�lʝ�._���o$�4jl��	d�6d�+�$Le��4N9F�D�: ��,65f�'�h����4���l�[>��3!�>�y$8=��Ǆ �C�k+p[���Uk�Hb�U/W�G�5�������1bBY���/���T��p#��x~n����h��ݚ���K�e=����צ���N�@B.G��m <�?�3ÌY.[���أ���".f�vrp���nr���5

[0=N�D�,I�}��F��12�0ӻ��6'�,�����?3���=�#˴�\���c`Z��_���L���Ɩq�m�"�JRD��h��ˢ�*�Ǧ���3��m!ԗ���˓]C_�����#�~(7v"���+۶U2��qMK&����k����@������c�p0N�;V u*����8ק�������]��49g5�#h��K	3��$�R�� VpfQߩ�ӟ�p�+�5������^�3o��|��;ݖ�ݧG�\�F�C�܅;��ʄb}f�����f-eǂ�Ҩ�@�Gͦ�V+�K~3��XQ��L�͕pk�(CN'��k�<���SJC<6��g�ϣ�Hlo�l��A��)��]�P'�	��~]L��޽$m�ۃ��[�4�# ����o.�)<OG��Sv�et\-�㶩c���Ϻb:��!����)� �Ś�Xj�+c�ыL�1��������܀��9h��*-�N��&sj��Q���O{jG���1~fv7tR1Ur�5����O~;\�ADC��=��At���n�2�H�K�-H�c�~�E�k�+��	�_ �Ok(t{��M�U+�9��� k��'�[>U�>l=RG"ϪM�W!�G�[�{���u9��b��5���iQ ���?�c==PmJz��1:++���1~�ŘA͑r2�	}<�D�>-�n�<A\��&�*�wՔ$ �B��ӡP+ab��`.�g#S3����7��9��F�k�7���il)�`���9�s�8�qr2�NuM�5��0Ŏ�O���Z6J[o���r���DB�X��E����9������zh��jG���ZGQ���'s�>��&�r{
b�w��;���R��$3l��;U����a�I-Q���#��.��C�q���Zk?/�)�%5�9A���ڟ������a�T|-�l���}�
$W�Z��s�w#L { ��)ᚇ#�����
@�LW0�$����	���-L��N����m����t�J(�gm��_�bT�eH�U51�\!���)2���c��M�B�q���ۡ�,�.hݷ�C�[���0�e�l�/���(X!5������2��ᐄS=.7��d��>�9�#J��f���z��#�K1ȅ��ǣW�������MZ	F� G���-�We��f��D�9>�����O����z)�����}+}��~��`v�*��})�ϿJ+K�L�*�\�n��^S��M�+��\�1g���}�!.x��"�Ь��u�u���5����wud|�ah��;�?�gЫ���5��F�βF�rK+K���t2&����z��lԻ�����G����Js�'o����f��������8Ώ��iA\�H�]Z���1��Ȝ�m���>Ϻ��F=���[ק�BV�q�h���*#De\W���]��C�Y�����py���6#����R�@��\�P�2�)<�Mg����G%���Ge������CEyK�|�����GN�8��+Sk�?u,��԰���@]�<l�hM���g�F�,��1S�ld�&_����'��oh-�1��`ib�F
��p��\�p�ߔi��oj��SZՆ�a00Kg���+�?R<e~�(#����Cd`�m�"5�e��)� ���az%S�հF�%~؄�����!~�

���5YV�̺�Iv�׍�5t���]��"-��O��6��^�T�#J���L�V偲!MlQK�p���H��uc#|�A�d@���?��l�q�o>VR�N�D+��Ʒ6��fY�ɲ惘��nś/�5�������Ċ����8�Z�߸�l{Z��Z��O0�FOcw�U)�1+��B?U˲}�>˼�+���g��VBI��8��ӗ.p�?�:�5[]БilQP�q>�����t���^S�����aD���wn��裇��9�@X���f��p��2 �<�ͳ�Q*��?�����7�5_��GUH��;[IQS���T��U#ʴ����~�2��L��!���&���܉�D�%܇�)T��!R�����<):eT}��N��o����A7�io�][.�����lׅ�޴��R���Ph2jM���˱@'���yk5�9�bƄmG�����Loxc�K��N��A�%�&��F���f�!���$Z���� �z�KM�y^�����a��/[�;��������Ƹ	S3쒒7c��>9���v�M]wۋ�����w����m�,H���]O~�՚��JTcu[�Tm�y���2�?��|�������"���b���O���=�畬ũ%߉�C^�������:Z�@'����!�ow:$$�`y��v���t:���ր���y�g�b�F��{=6�J�뜍%0��c?�ܝLSTV���
�ɽ�Ǚ5s_�dG ��A5��9uT#���H�CZ�K��gK�Ɇ��65"�ubݚh�YڹK��:���D�k3�Ҧp�(d�s�hM�2(��� �4(^�7w�2���_�H���4��{����H�|��~��I��b��և�+��X�]�0�qV�l��(ټ�?�?u+-1Ͽ��&��]�� ��1��n��	l�F�a�\��kYZz���������{w<��R1�cΜ�8�'�WV�8�j�T��oԘ�)k���фK��L���̎k~V�#xjT�Js��0da6߉�u�T��bPcɚbb*b�̐���**�俸���{&��� �{�=䯓���(�|r�����];R�F�h��.�^h1��c]��U1_��tn��[��H�TjD���+�w��
�����$7g�l�5G�����%&�RI�w�Cc0񕎰�!O[@K�`��Z/F�+��	�R�r+=ѵ�OA%�tKb�/���0Hm{l��9�zh��(dB ��(�hZ:q�|D�B��=��)�u=k@:�c�J1{:�Ԯ��f�N�a]�#�ߨ��hd.JYP�������_�8n��ǂ�T�Nfҟf��5-6���[�?����������«ȓw�wC��/�;�J�y���|̓���I��)�/Ze@�K�fv\��ghs&�t��$��I_��(�F'�	�CO�����q`��C13���
��-����C1p�m1m�TKM���c�~�U@$�'5��b�;�'��K��aC5�P����L*2bB���׳��?<��|��Ķ���-).y��Ȕ�;�S��e���KC��iё3�}�1?n���﻿��+�Q������8�J����8V��C����JbJX:�(l��$���7	L�C���A�i�	��)����j���02GS�p]�ÀU�{�K��Oυ���L*��bާ��ݘM�5B[��剈��9UE
15T����ew�Zl��@	��:9Γ��O���R�#��e�Ҫ�x�B�+`�s��2����*�Ȯ,,�
�o-���-�������1@U㳯nhh,�,�;�5�f}��{?�v����X6F�!7m캗:�d{��%�U> �AẦ{P��p[3����V��_)�tP��G������щ�R�k��,�n�Dֆ�k`�5EBꃞk�pM��Gy+]T5��I@ֹ��G_X<�d>�t���q��v~�bw�"d�o��݋<�!�߾[{j¶��{ʲÜ��.w�����>$������h�I;D\t�
	=�4S���!��j�7��O�5y�5�TX�ӥ�Hd�w`�f�TbnS\ ��\ƾo1N3�YԾ�x�#m$��x�3sv���]�����S�^�^F�A�2K�����S$U����͉��8|z1~QI��k�b�,Yl-f�w[~�e�aŘ��l$���^Ĵ�r��n��[�\����}��}��O[ݚR����}Ն -��w��t�m,z�����`�a����o��~%��_���譙ϛ���A=k�{�^��m}���1�\�pj��C3)&Y��5�����s�Fl��[�>�#$�Ӎ0bk{P���W;$n�\(���=�-�nz���$ݺx+7��;�=��g�5?�Qy��-�_x�#ٰD�2g���a����^.;V>A�ק�IF�	�������m��z[P
�c�<�Q��+�f��AY}�.��D��Z�x>ԎՆU�'���mv'!�G�C�#&�w���;.�(�
���ântQ�G������U�ϟ���v!ta�4����8A�O���Ҥ�ZPW7���Q91�(�[�o_�l��j/ΜȪ��LN���.�][�A��A>/JH6P��8����Ǡ���2���{�B=�遦.��)�e�( �X��~��&���Eg3i�zj�_�>�5k>]��?@6���H�G�����̓S�U>{�s�����~�n�j�/5���X�R@�!�.��1ү���,��G�+/]�ۯ���(��Ú�{p,S?mc�" K^�������3sv�^~��˻��qH�Q���uql�N�C{cu��^WO��c���2Ũt#�m8�*K����%h�RƟΨ���@×4P���}@NCv*e�~.������������p���5�ͩ���#�]�T4��8�i����e&��1c���S��{3ã�GG�I�"�hvE���SxAX��&Q��.������!F�G*^��q�L�-���:U!����]b��c{Y�)~���9#����
@i�e�^��`ixp���"��>|Aj��F?�Gţ��aЫ�.��ƁM����ʆ��j��.5_��ޗ�W��dy-��R;�Z\�-���L�h%_�l���h��]KU-��R����gz�M�G���D��M^a(�_��?�!��
O�~_l�e��K�畞|_pıN�Qq�3���1���Ѓ	�W+������'��N��ߴ�K��-)��@I��)���b��l�k��|�����wv����m�r -��S8||
Vk����Q^�����tȤ��T�ۼ���(\�s����.�%��~�"���3U����u<�{����rv�;��Xh`�=�K�� a�r���2��Ti��j�K޸��jkٴ3�11\B[��"��`��iL�D�{<��*��*���t��.%��<9!��VJ���Or���2"�o����$к%d���Ӹt�Uݴ��:&��9��<Β������ �)�3���k��/3?)��L�~!���Ϝ�ޟ=�m����\���]�?;w�y�a4���x���D]�/�����jBؑo�䟱D���&�^�n�����D�[����&�E��j[3n��lh��׫zmV3�F��O�����T;�`$�=����c���^H�!4t2�ϔf��#b�F<����`a��[�Ջp¹bC�`�3'{�� ��E�����,`�#���=��6|X���8_��w�3Ɨ`O��9x+��1��J��$�ch��u�#b�Lؾv�K3~Μ�����:�\�0q��?pŬ���=�9c<kA��R��P���v`0��l�{s���n}(�7�Ǳm���rJ^SRBXC��6������Ȍ��d�-G��y_�zN-��?2���"�/h�m���r�դ��~��M�@�G�*P�"ʠJ�����pz�}���-`}CR��>�6��O��:Ψ�"$��G�Q����.HI	E6������O�N�}�YOBM;�c�E���l�/o�������H\����:ǿ6x�򩽔����1=*���=�w�ƞ�Gt�,s�y`��vqv��~���>�gKXy^U���\���P��/���Y+���rǌ�<��<>����%���$���00;9�<�{�.�Ԛq�k$~F����KM�dv��-{bA��RuK��� aouF�Zr޹��MT�A��B��(��H��%66�����n�D��GKd�W�?]V���o��>�Q����M�6���՚*⠌�S�>S!�ur��1�~��\9نxN��v�Ȧ5'�'b�����@%�qs~���3����T�g�)�g��j�~c�]��G&�Z��:͖r���$_Ѭ^��Hl��Gg���&d�/�SF<^���j��l�T��k=�c���������x^��`[���N��T);}lf�w�����֨"��qV�8�q�ڧG�wP!'�m�����^�f4=� &Սª��}8�J,��+̈ѳ���C	���WoZc>�@6 ��<���k	P���(P\%lܕ%�1�Bo�_0�����oܾd������ˎג�/���z.��=:љj]M���A��F�h�����^�^����h1>���S��3����q���<�0�+{�'�z�~a� Ud��`�d%g���w�#���C]����ѕ
��sj�"o$����i-"�����H�殪�2�L���-vѳ���V�G���	P�2�;U��PJS�
�4?�������r�u{є�1��ΞoX���������v�-=�&�=�6OY���P-(b*��V���Y�䅁okDf�L}�,��������R�B�3*�����5���1F�S���X�M'��M����Zh�q�[.�A��h���ٺ�k_�J�q�0�;;�~fܯ��3'Z�z�#�q�H���5�f��.�Xl|`�F@.�Q?�i�y�8����N��t������+�v�ӣ���|�Gqr.�'F;��.d$<`��8$�s`/2�����"X�a�N�R4���a��q��i�
�@�W�\�6:�w~g�kֱ�����v��h�gZ��y�昫�����e>M�S E��c�ִ!\k���s]+
���i�6������[�������O(:]�g�l��u/5_t�d��	���y��"g�hӂ�#�����|��/�u$[.�0��=��ܛ�i�v�_�L�ї���z�� ��?�h��b;�>����>E����N����������]�gi����?z5�7��,����c�����ܱFh2���O�V*���L�� h)C��B�k�y�G����/ܧ^*�,�szSdZ^�{=�_��/�]�l�?��o��+�������֨�b�;R9-��8��0/q��};3k���Z�fC�ޢ��}��;�_�~+�[���ȎJ��6�����R�|0Ɔ���+�2m���{2�ټ?���X���! ��v���Gf�F<���o�=#�6[xjbBۺ> rZ���(\�9�~���D��f��j�[�� Ŀ�j���&mb܅$����H�oJ�U�0:�F 8���3.�,Ch1��E
�o��e��c&�t�t�pT��b��B�HL��^yl?�h���;��t�-�$�~���o��U;�� <Ӄ�I�����	��f��m~>	ٹa�+�#�+xp�11� w�������7��$�.&��>v�5��$6��~�V|�Hƪ'��f��{��bS�����n���`��S;O[P��2��G����jN�Ŋk0�X��۽�7�(��y��`�r���%�m��2"����`S�V'�%
�3��Z��:2kx�#e����eV�/�@�3E{^�R�;�Fz���`)��� �^3D��8|��!~VX�=.ߒ��w���,�q"p��f���S�K�c/�O�tM�ô��ǜ�����s��`���J��}�n$��>)8�bl9��5��~�͈��p���-E�}�;�`1��q��^�o�%�WP��.F �۲��>�j}�	��<B�$�RdD��@l̗�����n�pʿ[;����A�"&���XN]oKzӅ�*SG�G��UN����H�hTM ��еWY���T�w�V!��7UJ����+������ZN��[/ ����;�K�*r9�]и�v8o0�uNS�Ź��������g�l�q~Yz253�$$�l���[O��������tO؏�ʿo�Sc�_S���K����
���i\B�z���A$��Ҧbi?ay�9^;;�Xs����>öU��<� [%�}t��gTW0�i�A���'�}��w^�v��/�"��pc^�X=�f�z\݅׿��<oʠiǉ��z������$S:�I`�c�7_��P����cbK��A�u�B=���^z�|6���iO�����Z��Z���T��e���Gzf@"�+�B�KC+��=a�܇�����\8����8|.ZK���u>�0�=��ڠYr@��G��^����%�v�а<_��P���*�_�^�R��@!�gp�#��}qS��hǽ�s[,�����/��<.N�K�1f�;е�q!>kN��P��a1�,�Jm�V��
۳�'���@�.�n�?.A�>+=�����W�z�X���z��f'�z{�G���?.���4�l�ثz�Ks� ��cp��TB�aȀ}0��nwd=/ZaM���������龜�lsX��?�.�V_��<F#w~, o`���X
���9�³X��n[㝷>dT�P���'���m��b�M�Mq�uo��7�ʠ흇*,�t1o�Tik���틦��k�[���=�W��5�ŪaRA�lz<"��.���q��3x>��f_�*sR�k?�yՔ��lC��=}1��at+�w
`>yK����%��(�9ϛ�,to������?����R�3"��&�ɠX�9J�,2���򻅈���G)��]b��b�M�SU�pe�j��q�6�r�Ç�|��r�T�j@�oK��i9}����T�8N�/��`��~��iG/�K~ț��	����iS��S���|��"�`�x*��.��U&$��&Ĵrٴ2|�	8
"2�^���|ب�
���E����8+��[��<&,7�$��A�e�����QE�=ZCCKŌ#5S��
,����d�V��aDi}9���6�B^D�E_�E-����/�N̂V3So���rH�V-��{�g��~�^ʹE�i����կ{�p4GG��jYhf�cdwk�0��pJ�O�z)��4�S�6�'}��Jx��0Z�c�j��݊$�j��z�X|�v+��lm3�q�����)�E����2!^LV\�{�.Fi�kt&:(JJ��%�+���K��p6�S%ߋ1�M��XQ*�	�cJ9�kVJ�Q<nv�L��vկg�qw���6/�3r�vA&à-�GO-�G����֍������s �Y߇g;!��Z�����,�h�S��=�EyI������gWTPg/|ڞG]����$�tR��[���<��rJ���a'dє���z�fx׹}I�{�FDj�WU�U�z6*���e�i�wf�{ �����B�$"jR�U0rlg
Ď��hf�<5���f�U�x�jp���aH�
�(�H/O�
���qa��]�����^�Q�����V_N�O�"��@SK.�o����|�6]��4��g�<akH��=���ۛ�=Bl��-��9�{�Ϣ���6�F{���l7wr1��\�R$�ɼǄUs�U�>������.�l���L�^3W��,�������X�j��M�0&[9�Z·��6��Of���,Æt^4��q;.S�RBbh�iV�!�@�0�W%U�������6�K��Ҳ�2V�\6Nnu�:Y˶m-��m�ԉ������~~�u_����d%�R<c\�`1�9D�j5a�����YH��#:�,��G�}��,n��!y��y�9�WF²�H�j���r�]Ɍ7Ha�[�T2~�5�VU¹F�h��7ֿ\�6�/ضed9�5 �x������C5ڵl�]�T�;�U�-m�bAO�i� Z�E���e/�9Rnu��{*�ۦ'8*�"�k�I�E�(S���ش�!��;������u�����+�g���"�{[䄃��9��Iy2?��x)���1��t!U��0(IsCiEC4!0Ecm�q3X�B��.�v8����[B�ie`������n|���Yg�K9�@nC�ZP�z�+YXc�_�����䕠��e�~f���:����JuA���Y{	�V�j��ǘ_�C	gbӠ���U-��.{�4��=�`\>.r�w�Ȕ�ru�� �,k�Qc���޶�t����V�1�fp�Z=��e[�����:�?��.Wd]{f{'L�G�|S}�DnA>w��i�m��ro����p�,��p�f�9�ţ�!AG��m#���(_�((��I�C]�p텬{�jt"�`��n��'��^s]/�sW���	1��|��.d&�侑�|����5eA��]A{I���3D�L���k�x.�Fz�b
¡�	G�x���!�c��(�[L��g�g��J�&��2��,ג����2e��8�3×��΋ͨ��+�\�������L�8
-���/!Vu��23~��X�#�x���@0v��wt�E���WsȤ���1B��j_M�MՑ ��[����!�NW8�ˈű�7�$[6='`�w�Ξ)�8�M�͈e�
RR��J��p2?�~�DU�@�HִNI�|��Y������5����v]O!���<`�|�C.����e��p�_��r��H����H��lW֬,�_&���766ĚO����u�.��n�VæQH�����#ҥ3̐�D���USms��k��pި�e�8P�w�``1)���!L���	Q�teU��E
9��yI�s\+�J�ԉ��J伎-'ck��=#�{�BRJnxЄ�?J�^Vz�� C�괉R]h8����M�T��]p�\��V�+��u���Ԝ��s���å	��W({��tl[^~��U�J�miN��ϲX+V�+�C\E�8��U�;�Y�3�ߟ3Vɀl;��T$�CI!;��:���<;�Os�Y���f�:��<���J3��Y,��oOD����7�|��Y۰Xbd�,>�Zښ�G�U�����܈z���(�hp�ew��bWG�%W`U���|X��u+�lk��S�k)ˈ��:�x�>�^���mϺ�����d��˄�ocFլ���B�l�+��J�tY׊��쇇�׳�����¼v�5��f|�(�`�zξ�i���i;ޙ�m��ɿ��bk'��Q+������P*S���߼�P
7�D��pZ��a�uVN�L�b�)�z�(n����V#��F�����O8����YO�}�#������G�[�i �C��.��}o*�HeN����4/���'�� k���NDUM��&�ќ�X����).d�4�Ĭk�YJ9
��ݼ�&�YR�X�A���_��L����_Wj�˛�L�W�d+�z��	 ����0���-��(�	�
�<�%Xw��ʰ1f��ܔ� ⅾQt�AB�U�	mgNN*��������+h��n��k����|ު�w�oMDY����ܥ�T�jE+z58d��@�L��Ӏ��P�͓�\DՅ��J�.?.;^���5M������ʍ׽|��B��Ar�ќ�@^��Ɋ?�B�
MZv�Dj�&�T
�l,���GErr���W�4�)�p�3`E�,]��["{\��ّ����X^�8�>��ý�3�T�7r���q��â�I��`��r,f��b2H$�!�� �o�HQ>�{��<CCV����7ʇ�8�hV+G�Hw�������r����a%�u�Ll���{�X!�e��L����Y��O�H���KI<:k��E4�T�F� ����?yC	F'�˻��1;����`
�<�����p��=��]�	���A�<��+;�n�����̊i%qw5�w[�6OE�b%-H�2C�z"�{\�:p�Ҟ�fL���_aב�*�T�ّ�DN=\���S�U�l�xۣ߿��s��-4�;��!�S֗��c���d������df]�*�ٔ+�Ԧ��C�-?W#��:ᒖ6��_�\濃d��[���{S�	p��\N���0|�E���6����"f(����|��eы�k�0o�@���D姹<|�e-t��)P]>������\�B'���4�"ޢ���$���&���OI���Jk�!�����N�ǌ3��	c��_�:��T��mRY�8�F5M��m�p��k���VcX|x ^`�]��z[���P
�y��сz����F��B?qq��pC������cf����`�ݒ�h1�C\,�}uO�&��'�P��^1	E��/���hY���j�)p1����yO�$X�}�T��3����I�Z�.���Q�s2@���Ġ��e�&Ơo��$�c�|������v�@�,$����#�;�s�������q���q���[rb��a@�<���O8�C�$c�Dc̱�Z2��tZO3=S��f�7|y <m=~ڊT�fC���^��0xf�򺦑�r�j\3V(o�&������+�l��f�Dޫ\@�@�Iib��X~�w`���@e$UE>�'R��I\�<��dyXVu�z]]�nR؎~�}��օeֺ���Z�������fj-�8�;�Z�=��}d*�
|����O��s��b>��1��������#��}+>'�}l(�>���d�w	����@��g����^Ӹy�v���en�t"E��}��k�cI����
�3�?~jao���F�H6�j����!�Ю���8��^w0��;8�¡��J }�(C�
l�m�;Q#��k�� �Y���&Z�ѻ9nS��l��^�S�V���٠��b��Lt�Ht;? A����A���C���#kV�,p���q��_v�\JwZ�Yt!J� �/����{3�,��Jo�[���Y�:h�(��u�a�&(����3���R-���n�'�^�N�y�rr�6cNz�kxT���6g���wG���=�1���e�1��&���5_w���P��A�� �{)����t��D7���:���fA�CJu$��L)�$&���
�~9��Ex�5�O7�85�;X������f#׭R�����9��v�772�]�O,��HH�3:��l4Ř�c%�>qՐ[���������XAp ��r�]^�fz�;C�ρ ����b��s����C��-��T�u�w�Dew���O:!�^�$T6�}�*M�����S�P���>��Ui�$�?��m�n ��KG�
=W�ko~���@��xğA/�[�P?�ѭ*�@�L�Q���# �US�Ui#Qj�Bcy��fDx�i}�]<�x��7c�逎� ����c�-��u�)2@��h��ɉ\qhu�i	e���|{ig^+B���O1��9ԃ��_{(	8	�~��1�8��|>4�F���װF�ݍ�Ǥ�\ױ<Z���7��@��@�3rs���5��)��/C�K��B>�n��yv���P}�a�b������q�𛖺'����zn-^&+�w	���p��z��Gw�b�vԕ� ���i���t�pӈ Hĺ�0IϩC�2�{uZ���61�S�^{��t�h��@��ų���Yg��;
�/#�qS�e�ş�{E�\&C22��a�\a��1�w�0D#@)��8�DJԙ(&��^w,��:V�Q�ج������ނHOj�S������O�ܹTyO�	^���{�IĘ".�$ԃ�04�� b��P��T�B�H��+�
?�*;+y�Z�>rK�k�~��88&3���'u=3������||O_����뉷��'k.k��
Y��3eSW�[�t����J㻙�`R�%I:-��Ֆ9�l8���&�����LDU��[wmæ5��$��|������G�֒��l雷��虮��H�P^FR��{>��Oc�'�q�N�=+7��=�4eSG�$Q�V�*���Fq��$�R{Ԗ݊�̾tx��7E+��o�Ӗ?h�v��l���1�Ԓ����Ӿa� �����츙z���!.T�%��gƫ�˴n�D:C�{`g��d�Z�����|q��-kI�y]�
�_l�J-�w4���Y�gu��X�w�7�q&�l�)��q�����R�8���dS#��/�P�>[կ��To�����9��҅�鄴bk�v�OEA��d�3�~���U��W)����?M<,]�l��5�^<W�.m���hr}t����v-rܝ〄���m���PQ���;ރE}6�teYUZ�s��u��b���ā� �����&l+?�~��1+I�R+����f��e��5ʹ��@��D����b����9M��3\��Bce�z�T͗*1_÷�?� :"G��Yx}d��H�[���$�Z�B>k��0|D`�|;iKf$Ap�򼎙1K�Ig�8kIa�v�uЩ�oW'2�瑂f'ރ<Ls^�E�ҍ5�K��0G�"�\�R��x�!����(��m��s,�~��gN��1��8�5Ս5������-�XEY����vW�pӎv����Uw`d^߾�#�^w��i��Y6����S�O�~���ԾT�vƂ�n�s�^�@�<2gLli�g����ƺA��*�oC��V����B��s���D��E�=b�g�ԟ"}�q�G4�LDJ�-MI�T�M���d8�����X[�l�?F?YV ��~`��uZ����|}d�O�����|]�x_�;u �c�ж���ee=����E��!d/���m��Нl^J d|(����4�ܾ3����t �*i��8�P�MI�+0��e�/�Y����v�K9s� P�lG�I
á�G�LT[��k691A�/��-:d_�Ę��`ךbͨ�h��l�C�)PFr��AB��]���y_�m�>����b�>�.�g�j͹=Y��g�d�*fH&����ro,�,�p��XE�T�jj���#��y?$`Te��(�9tcqy,2�O�C/!�v �6��$#��bQv��ȫ�\���-N���DEVux�Q�sSN썫t�~�3ފY�T�0TT�Nq�*��FD�F���̟�.���%�1p'���'|�D���Gċ��\ج;�I\n�D݉�\>��m�^��roQ�W��O
�yҊg�����	�M5X�9�CxZ_��*�u:Er��
$Yd0�sx��DQ�
��)�cN�l����+��U��Kl!\(���$v�1�3�D�p-l�N:]�xl���p�w��:�`pD.]��a/"�'	|7t���
t���{
��,��Ql'�.�������j�$���chb�Yv��}Ў�Ģ�`�I�W��Z�X\yr'�<˹���J�T_��ر��Ȓ"���f6&k���tKj���I�uՍ�,��}!��;�$���H�{o9�7i���,[�Z��fU)+��� |�M�JT�=�1,"�͆�=���H�� Ǜ��|�4E$�h����������Ħ-���X!y�����G1���DË~6�P_>�aV���?����h�5��֏0-7��X��������xzldZ�\���%PB�3�Q��m�f�����ٛiQ���@�B��Oq�U���+��!uO����xT����z;������?�ʖ�~��P	�G:�P�S�������ٵ�D��	QI�t?��F>��V��vM��,�mdܫ.��{pE��]�3�G���ѐ�.hxH�Y0s�}?c+L����2$2LsIp�6��H��fR�<~A�cZ`*_*ɯ��!�0Z�U-a��t|a�8Zs�j���1���`�ȷ�[sՋ���]�SFRk��/�4���EX�����E3�//7۫<WRl=��F�� �?��v&�k�(���x.9��T�-��y�G$=���05�<i���L�X�?*iĜ3�z��; ��X�W�bt�2q�� K��/bao�	�fHn�0�1�[?��i���9���[��������>��DM����w�[����(���5}�;�F�8�ӧ$��OO��g��/:�����o�.��p�N�olٽÊg�ܘ��d�s��,ϙ �Q��If�t	�ؕ�u\��8�ޑUds?9���l>�w�k'��Ӱ�I��+�&j�y���.Td+"ߥw:�.��l�T���2V5�x�\�n��A�����x������s�c����N�C�'�}�X^/?���Q�����T"lN��Ig�]U�(�sOR(�G`��o���������T>ɤʈ��"���<��\m�� ��WG�ǿ�=�|�\��c?xE�.o�R䳔s̽W�K�o�����P=׃*q!J����;b�H�'�Y�v�+6�I�Ӊ�[�u��f����->ȫP$m*��{{>�iά���ðb����<Yڍf�۵���A֮\���mI���+IEl��G+�V;���4=^ɀ��hI;��!51�a���E
E}��~H�������I8�.;�uF�UFy���a���&>����LRJI���[:��Æ�(n�%/؟��g��J�<��V'�'��{���.Iօ�KB�my�IQǙ�gu��NDu5g���͇�M8��t��/��B�3]5�9ښ��ѿ7�������,�wTMx��9���?��bg�銐�Ct�7�q���v���,h��H���p�4�3YW5�|�1�K�#��,r=l����-.U���@�<=Rsi��d�IНV;�u�%�(��-��C���iH;6�Ti*9�!���mc+t��M��G�bST�Mb�3"�H�	i@��L�fY��,�8�O�<�]��6��	2�/�l��sh-��� �����J��}���Ѯ�LWk�$�YI-z#g#6����"S%�����P���v���^X��%x�ъ��|��2��wG��#$zf�4���d7�� 
��V�W&C5
!�3>V������ ���	��/"��)��v�Kj¬��N]�~5�a�G�zt��;}o�����N����v��2�fN�wdb��鯼�<��IN� me;�yH~c���H����h|�V+���_�G�E�º�v2� ��إ�@�fӾ�V)_�zB����`��2�����WL19Jj_�����D�{瑳d��o�)쐁�����uo���Z}P�:~�q
c�����PIkX�0�$ �1�]��s���)�j�_������[.W��T�7�D�^�xɩ@O��������юQ� 7���,4�+��a!>�n�)7~j���y���g�K˜��� ���N+��W胕z>�1��XpC�C����[:XF��U��D#F������Yg���8���U|ޣ;]5N�kd�Ue%���K�^��ԍ�)�S0	�C"�qpd�߰��#aN)�8l,�S�ϥ�9Q���2{&�i����E��C��\�ͥS ���xH�����?	�M��������a�a�9����91��L�(�����-S�8�#[ߡ�k^Sբ���B/��{���n���z?�r��ũ�n������*w�g}��`pڌ���e��D�D\K��
��jB%)�)鿂ǯ���E�����^T���ꕐV���t��������v_×}��U-������xBoH�_�=����^�z��f|j�+�L��i�/rv�V�&`5S7�7�hă���+�?�h�&l�c��`��:g�;X�3��ν?F�i0����b�Ym��F��-s��*�`Ї�_�ټ#c�	3���Py��3�8ۄ@T֫����è`����	:���n�-��qӅ����߸≺���e瞇Ԇ��L��s�\fv&.�/�[����,%���^r��J���uIu��Wh�G����@^N�I�����K���SU��ߣ�X[�L#B�_Z�ҽ��f\��_�c��%3b�h��Q{yM��V�ߙ0��ug���ӗ=��!��]D���ܾBd6�k|@QV�뮌A�����nP&�f���nǍ�"w�>W�{���_�Mx|����K÷p�{��cI�1�<�;���,N"�)I��i?4�j%�-��_�\"՗ud��b{gQ��C ��I;�wy�S�z�!�{Q��[�2�U���Vp�}��)q���������a4%S�V�W��gͅ��4�N� �)�e9`���6�8ɽ�G���{dW��{V#�q�Ļz斾"F��F�b\���!�!��sS��2v���y�mj'93 ���):}>�
d� ɔO�C�Q�Ğ��)ɣ�~Td�ޠ7�=ddb�Dr�����w��QŇ�[��m�8z�9 ]�Ule��Y�sk:-�78Zs��l*����,qݵ]��X�;ۀ퉉��%z��:��I����#Ⱥ�76	aBe^�{m×X�g�M��z��С����fG�z��ls�Wg���[����.�gN��#�l��f�=,��@ܽ�� �J���-�6ꇃM�Z;���9Ӫۯp�����d'��x#�R=g"��[�1�}�:=�@6I�n���j	����D�NW)�k�՛�&��(G%	VS�[p�q�	m�V�}t��J�gy����滂��r9�tYF��g1M"���	�9�I��r-�%��O�Np��e��w���ܙ��z���mc^ڽ5�{�)��/�ӱ�v�y��bwMNf���H+��Ӧ\`��H�����5��h�y����Q��Dj�s���������k�n��a9v�x�_����dB�N���[��C�<-���#��d��G�� k���G�Fq��f���ب�Hubr��˴r�q�6H]WL�"��c=5pz
�Y9`��o�K�^r�ݧ��{��[:Բԇy�1��cwQakP��B,ke���i| ����\��/[%o��&i��5b��}(sV�i�;��;� �o��zڪ<ԣ� k�A��?�.uz$N�0	~u�`�)ϻ�<�V_�b|�y͉�"J�8�ԟ-����1�t� *���?��X��4�(�M�~�ǒ���z@3�&�a��p)�`2�~��?�p��pJ@`/��-���!|�K�M��GSM���7ߤ<�=�b�6����D��吵���8[#N�0�{��\6�bo-�X�G&���<���=��bV4��(��Ҿ���縥}����J`O�V��ב�y���_Р�DUM�C�|R�������4D!���Ë�����3�4Ԡ��i������!^��D��hI��@F.�4{'β��5;mE����AY�泿L�Ф�Kx�ǯIxE�����V��4�@!��曈:�'�7��"R2=��<
C��u�TBBRh�H��+4b�	e�A��Y�U�7Խ7ߣ��m��M��	I��e莉=�ܯ�;�Q����`��a��yO�k(�%�oyE�@Q����*��e�Rݶ��͂�ݬ��~��_�4^�@�.������|V�>�D�}�[8z�ҭ�o9*_����1�23��(�������O2C` V��������jġ;��A���I�3�}w�,	2/J�O�6������ߝ6�X�DC2NWB�D1>�	xɱ��`hHóa�J�������܉����^��r���}Ӹ�L7�Po,Yݲ�ŋ<�%:xrU;�?E��Q�Co����<�%
��[�;x��P��n~)F���x6S���{��j���z�'�bA����0��B�P~J7�/��7 ����{�hW��8�fr �i'�H��6޻ўg�������[��
��ϧ���a�|���I�H���v�g�"����&`-j�҈�+������4��Kq��e�����dԧ�k֮�"[Irhb��CB%�@j3�<5��Sq�^c�N%eӴZ.�HO:�Sv+����qq��(���4Q���v��C��%��\ʽ�7/$E�F��#%�?��ck�V��i�e��D�u!��ܟ5'&��R	ȣ�8��8̽n�����)�������y�w��6�Qp�c���^hC���K�2}t	�_9p�32��-�5��Q�e�f�t�H��6t�^���sT�]���2�7�'κ�b!�b�Zq�,�����2�j�'�C}�Hb�[��E�����2�]�TT��Q�y�
Fm'o}��S	����������D��w��3]�u����C$`�B����:;�A�C�yr%}9[ ���G%7� �k�kL{�T�D�ݾ\=}Sɢh�0
P�K?�Lcm-Ӓr��y@��2����9�Ŋ'N�8g����qƪ�E�(]���Td��:��_v���"d���SL�Ś� T`~w#	����o�r��P�����75��1�p|C�b���z�� -�qN��c¾���^���jb���t�j���dU��b��SG%��E[H�36�������X3w]�C���K�������Է2g;�̱�ZhjƲ�_����'�Ý�c`�2g�y�=���?�t��hWu^�	_|�s��R�G���?
*/�-�:(�NS������\�Y@+��ȯ�}�R?G�xz�"Ug.��*��~E��歲�*�f�N�_�8�uڨإ��j<�O�@k��X�����-{����.0'��k މ\�>L�|�;,�[S��;��߭�U�p1$�^}*Ӱ�BS�f��/�PK6o�����|�jh]�ƻ�6	3|�lw�ﾯ4J��՟{ NSn�����a�M>($iU�~,股��ݘ�"L>���}�c�~%����W���/g3��{�U�e�̋��|��&��|�/��gSc�}�3������^�	�ݣ���s�{&��3���r X�����
.y�'��͕P�єp�+:6�]{D�;��a�����1��%f�A�wP�����H����|~!����"����+a���m �+:.����
q66�W�htО��F\�>#���z�ݿb���ԣ��)�Gi�����PuŴ]2�Ϙ<����XF�^A>�E���t%��n*�*�_��ӱ�l��`�}4��X�������^l�)�?�D��a�nb���7�۸��K��C�00�"�a�{�Z�|��Э3`�����޲%�� ��ix�H�,*��qJ�D �7.�%W�9��Ѽa�`{F��+�ú�I����i�(1��
�뫈z��{�1��iy�6���wj�ZD�X/Y�Ɵ�\�_TyX%a�H�J�1�#-m��Ch�o�l����ݻQ�����WI�5|-�L��Y�@�z�h�B��1��e-ś�]d��J��w��<p����T�2<2�\Xp���0N2�'�SK��+45?�����[���R��XL"��?�@�<j�X FC�A�G���NZ��D��Nh߇ZJ��$�L�?p�L5�5tZȹ�I�����ʢ�u�]�&��^�Mg�̖ӌ�p��	�j��O.v�7Ɠ/��0��
��
m���퓵�I�i��s� �L~��MB+��_R����� /E�J���k2���� A�Ew�F���)5�E�жK�<�1"�:>X�2�c�*�:d�@��tԬ�v�1�5�ҕ�'g�����F�:��Iҁ-[c��[��L|a�fC��/�y�0Y�S�v	S�OP5K�a���ak�Q*�f�N�S���z��ˬ�t�����|��1��
t1�R�j�jk�S��� �2H@���|���8i�,�*�4̱� @�;���^��Yo�Q�B�����> �E�Ϙm�h���bL��$ЅAg���x��0=d]��^�=X���>���K��o�Y� h��7Q8��X��n-3>�����/R���Q��/�����^�`�!p���{�ѯ?C,\O2���X{�?r6O��@r&� ���(������%�Q���m��q��x{��Gןa�^����xne��s��v�<������;}��	����tA���x��,a8#��Y5�?��0H�-I����6ݦ�_��O�Q�蘅;�%�cD.�5%���O�,�I��%�hިF�ՈJ[��d�� ���5�Y���SP	�q�q��nm�5�^х�Xp��s���
S�pZ�:ڼ�'b��A!Gw#G�nOY��H�9��I��z�H�/y$���0��J&����/雦��FgFz�W=~�����G�����qdEdd�������njJ�[u��&����Pw^1�7���rd���$��P������y3`��y1������؂|��3�knQ^�W-.Yd�ص�'c"�9��Ut6θ�˭&�h�{\���P4���$�zZ�L��O���-���?���7S��u�Q �������iĭ�����8EZ6xؿ����א~������e~�\���|��@k[�� �K��Ƭ�u{�r6g.n�� !��e�Td;�b�#��'t�	�͸Q-�)�?h����T�����c����آ�΅tb7��rU���Ͽ
(j6s���=Y-�5��^�;�AN����Ntu&t�"�<�i	ہ�'��]��,��אV`j���o���?J�v�_�5$�s�W��f�9���^-��a>��Ά���z �d U �ܮ`�1^����"c��]�yh�\��<բR�,�y�k��#��_���I*k���>�ן@n��%�k��>��ai<��Ժ�7Ψ|�Ez�R�QOqd���0:��$��Ik�u��y�ty��e0NimKS�[~R]�Z��^fj��Ɵ_�)
D�t��s���D�H�|�ξ�
�$s5�^���b�X+�r��ҔƬ��U5q�6���pgd�$�q����t+��%��{��we]od������h��e�@4�X��R��OfԆVp��k����o�=�Y�L0V���H�hM�('�"h@�6Z�V�NC�=����W�C��D�7%|�.>R�ךϻ��/ɷ���m_�Uڕ�r?�=`l�l�˻���%�9�7�<������32���J��'�	�y�=��p��2���ec��(�C�;)U���Y>��[p"�7Mh�pl@���TշG\��T�v��9y;����ˏ�q*����<�QC�f@c�y�~��$�>P�$���i=�������?+w�=Iiiѳl�_2�a~՞���U:���RF̩�����2�p��A��;�nλ�l_�QYU=]�M��@P�)6�=��a�ʑbbCX�a֘e��B˅V���@���%Y�qzwSLRǝnG+s�ªi���NN�As�&\̃N�-�e�oJ�a����ÊW�V�D�n���������O3l�����g� ۄ={KwC�]�8��X�0� U��Oؚ�?����n<;#�=P?�������$}��<�3a�5f� ���4zqY���a��HMp����w�ΛW���ie#P��������+��2��P:�>����Y鍭��Zֹ���,k�ER���wX؛D5�(��U�V��N���0�Oq�	�&��OFC���_�G�cT8��+���9Յ�F���ȳ՛�(�f��l��'B��
�~���D��w�z�7�^x`I7~�'��ڹ珇2�1Y�1
�8�Yveu!���}��נ>�],��'#=������m��p�)��hY���)�tcExw!���v��sp�6������%߃�Y,���jPaC������fo ���q����{ni���m�B:ꥍ�Y66�x�C��-�&�6t��5χ���dxN: �0H�~Tڮ�-�U=��$�˥7'h]�s����	� �KԅE;�c=��SS῝��AG��v÷��n.%l�B7i��D�Q�|T��A�qL�PY��s�%���hZ��B�䂗���`�.�c��35�E$�����N8:Z���DPe�v���hC��L9au��#ߵ �Z�ߡ�}MQˌ������������'�-���U�{�����I(lY��J5(RB9�Ϙۢ�g�K�d�b�/*�Uø�j0\�uwm���AE=[���x<�ض�{��5��uvw�O�\��^���_-[W1ӏE���E��/�ѧC��]|�΅�\UYO���2BW�Hf���W�v����^-�ԁ��&/N&Ѡr1�$���R]b��B}�1E�����7mx_���U4�˯����71$PR�^�����0��5�J��F�n10�q���Ϣ�e@�����Wj�����4΅�p|��ʑ4�L�)E�|����ˉK%�����9����$^>���Vc(�A��J|�����G���
��0�,'֑=p�����0tR���Ol��d��7F
�Ln��dX�z���]�QD�Fn���ijJ�o!�m���**0U���	��7�T��,��l-�]�&�V2���/�f�$���z�cc�K��L	d!�V<h̓Ȱ��vw��v)��z�
Ӛ�i�n�A�M��V��<�ϝH)��v����^��U���xfoM{(�<���[�Q�ί�����F��Y���k@eģ@F��ܡ�h��"��F�:@{5Ze5C�]���N@�f�����?*u��/�Tf-U�ıHͻа���_�T�M�Q��;F\�<9�ָ�#	\��Y�O.�v1� 1ݩA�v�oY���&�J�)�c-�a����M�_545-�-pg�����LRլ�Ą��`�]��rvH���W�32�LQ�F��M�P�}K{ {p�;���&Ԙ�o���>�!RN��7�C'���tl�@�bk}h��飈�9.iv�}X�ڲ��M���j,�(��dK�_y�Jv��0:��@Ŕ��Ѻ�-Yb�tJ)Y1�I�G�n	����4z��'�l<�y�؜�&^G$�!v�!��[��@��pC���#��g 7�{@d2Y�\��R��+����HU��@Z��|���`�f�"�Laϼ B�W(cō�m�S�s���݌��Ǧ/Dj���S�%�m�WH&C6EGuR�Ή�������sR:�1���cJ�%���f��O%�P��䈮	��Y��x�Q� ��M��'�����ϕ��b���	;��� �2#��z�@���)\zlul�_�T�-2n�c�zm�b����������^���I�+�Ljk��4	5Zb�~kJ��h�܎�Lo�z�����h�����ȩ9��(>8aP��8P�y%p8f��j'���$l�x���*��q����
��V/l��j�E�,�M/�0n���$�	���o%��d	��(�1=�65+�H�u�����d�w�)-;���@Z�ݿ�[�&�RB(`��h��#<]a�,;���o�7p%�E� ���1���@Сl�7@={xU@����i��Mzx�J��o�_��s�a�i�c:�.���%�����ja��V�*��Ѿ`0%���[ٵt��?�w^�r8�a��?�2-�6U>$�X3�Ӫ0�uB�efʣ���9h+B�Q]"�����9�z�d�=����x��+AyȭO���yj�kٯ����/�U�XS�Ƚ�<�[��I1e�-7�f��;J"\[��y�^(gA��rXSH���?��.����E"�5�֦��j�Z����8��~*��3�b&���%iv�YLt+o��^�V� ���z|	��Ep���k��se](8ŉ�4�3���WF�b�M׶�C!�5���?�N������
�0�9������p�9/���.�:lɢ�5�+�N�ڜKX������o*���5�8.�,-S@ãG�P�Ԥ�����@�{�N4�]����}V|�R\W��;�<M ��_�&�jr`m��#3�dX���(�jh:u{*\9�&���Vb�7��4���ҤK�
�2N�P��Z��t����-�h�x���S���}ә.��(M^�\�} �.@��3��4^`�,��b���I	���VHy��2���[yF�%G�����g�/��W�7G����Q�����K��Cl�"�$����T!*�vّ��S�/�N�cn�2n2�����e�����-z��;�l�ֻ�{;<}\�&J��#-�F���]pm:�|:��{]��aq��yp�{4M��2[��o���&����=�yU��	9���2<>��]��xR[n\E��@G�g8���)�-�Q@��@��y�ؒ��µlؾKb�i�Qm��.����֯av=�����>�>�J�5U��A�u��=�Я�cڱ�&�b�qcQ�$����Z�F/����$N���9.]r����\���zL{A��2�x���}q��7�{�]������9j'x!�i���[�2�17D�vd��s�^{��|ڥs$�3�a!>8N��g�4c�2�t9GT�\XBY%z�٦��,��rs��V��C{�\���#��Z���;�r4#nb�#F�p�!;c�Qm�-b��]]�}�mU��	ݵ�X�Tf�ϛ��9��GY�0E�X�P��6���BF�������w<�"��/�S�����N�bQ#�M�R��\udI�|a��O4�&d�s[��V5�U��'w=�'_��D��㵣�}J�4+���=�����&�F�;Xs�%���[����tj�}j����3]�]�st1+�G#%���~�:�f6F��o<3��
���'A��H��HH�A�a��\�hӈ�-�U_#���h|w�p�������懘ݫL��]�j�"�^��^����o��.O��`���Ɣ-և�z(��Y �u��KB��e�8�[	���+t-��A������=��t-�;���c�}�������Y��0L�ᐭSO4�4&�d�w�p�I�o�ב��&��v�̀�����'�j�s��mOt��aal�UME�~94;)��"vS0�%R��[�	c+I�)YWB.��NE�����I�
��?�0�+Y$�O��cw����G1|O����W ˀ�x��t�vL�긹�J�[���Ｕz_��xKS�*�}�����e�m6X�7YQ������m�s{N�A{�n��@tر��h4��d���(H!MpI�������T1�9޶W��_6p��?��Ŝ���	�������y�/���U������wXt�Y&�7�z�nMX�o����힭=�u$��?'��K,H�|�����?'+2�	:��'���Hil� )�BjѪM�dpm����&L�k	UZ��]:%)���g~�����wf�?W�w��H�/�����?��&��0�y��$r�tm�iI���r�ZR�*��r��z�h.�C�F�*��HM�����N����GI��G\���&F��KA��j�����z)*He[�D0�ȍ���]��B)����笓.�u�KO�n1�����ז>d�M�_~��ɢ�uz�3�P����L^r�ֆ������>�p�Y�o�_¯����8F�t��h����K���UC{a�ӫU�j&\V����Q4����/��������mn{(S�ڳ[�mT���vL�j#L�fM�����/�Ä������蔈W���t^뵡B4`�h]�I�pI���8i"pK"��[2�3�.]|;^~���>:���~�Q'_�Ֆ����\߮�!ᓔ4ox9�\�k	����=�#��|���<G��a�̿���܃i�,[��VqB]x��A�3�����uH��ky�(ZFc�ǟ6q�����u�����/��#L���Xs��q�a{�L!WM8���|Dq7�M(�C\���8���#Qi�S��3o����Q��e����X��Qs&|��Ħc&�]���t `�����Hu]�@�"������!{n�}孿��v�8_|��B|�-��֛���&k-6Y��ŕ�H��G�`i~�#<#2�%:�ҷ<�뷠q1%�A��*}_vg8�[[��Ca����. Lk%�����gz"4�iA����pYm����>��qk�螗/n�ύGQ�j1��9	y�W��#:V�G�C���֫�[��S�{7�3�Z�������C�\��e�QH�Y����И��ugYe�����=�������������`����S�D�ۋ�Jq/Y����oas{6�,5���#]\|��$.~�b����>�+��#�������i� @EF��1��xZ"Osxv�v��hW��s�����zy����ۡa�ɫc�m6�gf!�E����U�o(�2�] ¡y��f���x��Xt!��ξ�.�~>�����O�	W��ڭ�Igi����ra䢓���&��H�,�j�B)iN�w�%7Yo��������'�>���x��<tX�f�w]�P���me��xs��2�	�Lu�$UF8�0�zo�Y�$��B��W��oA��!��j%�8c,4"�熭
��t���Ѓ-u݂V^�e��42FQ�mn�+��^���b^躜�x���m�Mv����`NA��DS�WI���	o�b�q�%����wpRU�����)[ �WAAA��`��-�7T����j��ލ�b�FM�1jb�b����]�m������sg����,�3��7�4d�}����<��G���#W�����dd%΀I��Z����<��rҥc�g�a6bQ���y>�|�w�/�����ś�~��3�G�=-�h=:��u�u�L�GǹE��ap?�k\vӣU�i�� ���vĎ�T B�YP�l��`��3dH%VI��X�"�kp�YW����������o��?�1�LRn?��Ygp�TB��M0A��>� =��j1m�X��ז�,�͂����7��gTK��2D�~�t�j�w'2��ܺ�K�xm� ��	z%=����ۖ[<����'K���.�B��"�&�k_w��{�+�ݢ�ȅ7�ddV���p?H�\$1J^+
92Hu��_����r��������.[O��[O�A��Ϊ��6��%La�Bn�%_~;�w��d��Z\�Acÿ3*�i�t��I�;ߓ��V�{�bb�[]�������[��r6����в � ¤Y�t��Xc�0:s�Cq��2���7ZR���"<�����Ҋ�ё�5��TP)�a�L���_�g��ˍ˿�_�0��+1��i�D�_��m��Iv2���8�!^O��L�@�*���(\v�#PP�oXuD�Տj�(5dm�iV;���}��Y���<af7�?��\y���j������Ǘ���썡�5�z�4��9,(/�[��J2Ê���Z��@+v��T��W�{��>v{t�,����1��7�H�\�L"����Np�VI����|�Ɏ�}8����_u�~�<�zn{
���8("����k��<t�m�mL5Ds.�"!쪈�#B��j@ѝ�_
�rj���b?�������#qsG�1�W�|VX�?j��8�D!�"�Y~1G��[U����_:��(�&���_OO�~wF¿N����Sԙx���#�YW��i/�`+@��D�4,*gp
D0��q���O���5�<�b�
�n�0낃��D,��@�����σ���>��ւ��lL��އ�ï�~���������~;��m6�(ų����f���z���lH�4�sv��.<�}��W�߁)�)G�(S������Y�ѹ?s$���0��u���}��ã�-���c�{�fX�(p�{�Z	/�pFz� "����-@��f�)��eg���FَpyF��)�G�܊�����''q�e���,�,�3h��;7w��뉬�,߫Q�r����_��B{�s��JP�1PD��c�^�M�d����'qج	CF/4:�T��$P� ��dun!��d`:�R=�/�*��o�R>�1���k�]x0��V 	�ZM�Y���u����.J՚@VH��$3�a!�""��L��`ctF��_�r,&�Ub^�-ׅ%���IU���;Md����--Bҡ���-�%.��B��Fl9e5Ќ����"�
��)�G�5�A��R�Y�} �N��DyMmX��2��}p���M��}��x�_w��i-n��D��KUEhZ���Z��c�s7׈�R�����g_yT������y'�=&���C3{�d�)ٲ/�(yR���x���m������__���n\��}���[v.�#/@Ns9�O$<�cp�?�=!�i;t���B��.[��[���r�^���G���;sWP���U�B�!��9����3�X�-"{��Y�5RM҆uW_y�ݷ�4�����G'����)PD�gâ]p�l:f�,JF��0���sd_2��i��c��HMN���g�^�d��8���P�`��Z+���4�a� �� N���hi�B�f ��72��8�$ئ��S�#p�P���Me���A�6Q�ñd�lg�,�=�^��o�/"K���D<�xMp� �h���-J�*�0��1�hV]�~��q�O�Q��B4֚0�߂\!D��S���Y;mhy����w�S۲pσ_�Ix'�w���ϡ�N1e�5���ʂLq��h=�Z׍m��\B���7j�Pg�0�_3ܬ���fx�=!����Y���p"�Q){���G���o�'�O�KoxN���q����EL$n�����-�5aA�} L=��7
DԷ�6���t�Y.�{w��h�t��?�SԅB�!�3��)�)�Ӭ�?�E3�����ր�}��m��5��^x�f��W=(�("�3�f�E��v�]���Bs����Q��X��%-VN�U$������e4W<'�N�҉��	�"&v*���
N8��#x|��v��D:@��L�a�ёw�D�C�?��d��D̊����o�k����a�(�Ȱ^�p"|�/�j��)�j��p�ע�j�s�e������hh�a�!ێ����m!��(�鳘�2�:"��`�H>�or�BoȠ
1�w�.>��ȸ��Ug�+[ �HD.��1E�n�E%ɠe�_$:͹>}�«��;�D�B���x��`���	�ZECjaX�I�E�"y�Y�0���+����p�OnS�DA�w����9=��֕�c&U#�XB�	�G���ef��{���-�$�|?��q��{`Ġ��a�H4v�6gc�x�B�A7�睴3�=�N��֙G�uΜ9��ОPD,8ˍ�̈́u_l�p�~o���&m���nO��8]]��^�s_z8dWL
Z&�:gF��	ׇ)�;���Kt��"�=&���c�۾17`u���?�&+,mQ�bqXU�>�2K�d+2[�	������9N<�~I�~�n��6� k����5��N�GFMYBX4�)4z-S��68�C�X�h`�^��,�{�⪛�0�O�=Q��;������Ͽ+?�oL3Ӧ��1#��Ѧ��C���3�TA�G�?C��D��Efd L��j�g;3q��Gc��/Ti�u�j�b�+!���
LC��&K6�'N��
�^�Z�s/�=Y������|:��k&�i\�n��5c[�P:�
�nB456ɌUU+��7�z�jB���#��F.(�3��)�h/֚��[a8E��Q���g
��ys�������ј�J��v���p85�;'�r����6@���'��Γ��5�>~'T �
���e���W`�E���Ѝ�2�A�<wB_�Mű�8f��|���Ч�CEƗ{("���|�y����e�}׍��cBU�t#8zZ��˖$�
�7[и��㥚I�O����wޟ������]oNH���ۭ�i���$n���q5�ĆFG�6��Z�	]O��:�$DȘO��x��ω|?��*Dw������������3��DL��2�Z	�O"Ka��(<h)q���
���V A��`f6�ȧ�G+n��0�v�e���%�<s_h�{�3��7��e�-SlA���W)���Ǒ�]��o	<Ϗ8�&�p�Ah�^�Չv�&	�9��p"Z\�<�:�p�P�o��p��#I}�4F>���p,�d-��z6��t^'�sk�>A�>�م��S��VPtق����Dd������E�sN�ǝ�Y$=�T��������쀕��kxD*�����h;����f��0�����"Nz��j�ڻl���w��2��s;���j���<p��u��r�6vb���R+�{�!�d p�pVxՈ�~���'��p5��N;N>��Q�ݑ�'�®D��R�a dd�Bz�M���ψp��9𸹽��>[;o⍷��܉�[��L�����cچ��ݖk�o�E�U�wB�8g6ʊ�T09�8h�y[�5��7��p�?��^UM{W�TES45�̄TgA6�&�O ���i�rhظ��'d�8�>Q��{���ġAkF�S���n���umjE��X�����z����9ؖFgCr�&א�ZHy��J!�Zt]�[DY����j�_^/)���/�'�Ĵ�GU���:Y[�ιR�D�0�B�52�'6��e�w�̣���a��}��1��N�mH�u(td�?�O�U��IS������m��]���W�O���@a��"�=��1q�Ň�"�E�.�f�
�w'��X�Z��n�[I�d/Є�n��ᝏ�"~'ꑏ����*�pȾ�G��S�*�&b"dۖ�|Q�Hw�q����hk_�|A�jZz݀J���]t7����e�����'#���o���S1y������C7�E)*�~sb�*Q+��Fli�л`���w�qgކD��:��sN�I��s��2��x��rs1�(�5��Ͽ�����4�{:R����&��
F*��3��!]�.	gТ���$��c������g��zE�����hjnD��M*�sKI���yJsE+�YjO��~�]�x�_}�_��j��Pt�g�5¤�EC�%!���AQH���6�E�?ң��>�N��w8�������Ŀ��t���K�qHi��LW��'hG��Q�B��0t�y���q�U�kOУ�����,�w�q{�g�m��I�^�r�V��݊V2,+'�_m���Xt��D��/[p�Yw�mޏ��:hk٪�����-0�<m,.|�ȶ@�9)̦�t`�	R#���O>�6.�����r�W��(���Q\u��p�5VHDW��&dA���\ht�eYz��z9������{m�Knx����p�8���t�L����o��%^F+ �,\��?��Z[�����W�v R���S���J��ri��l����zä��t��P��p,�梍(���!�ץRE�*��T��^th��3/�5�~�8t����He{Nv�Y���
: e�NS�0i�����k������'�A+4�`�U������5��xd_������ǉ�X�F��s멗�6#�΢*Ai9�"�=���;v㕇�kiI�hV$�ĀC�0�(tLN�K�W�/SPS6�us�p���-c�ᜓ��wނGVV�;i�|��
)G����A���b��1Q���W�����r1v����xN<d+�7q4�V�+��6l�{�gt=�V!��B�(�l>y5��އ��o�@�����!�lV\J�E�õ�n�4u��o���r�������Qk��2�z�C���`�����$��6fq�H�6v�-�﹮��묄Ǟ~
�N��i����}�����3��E�xou��ډ���2L̞�F͵�cg�CO���m�9Vһ*`ƚ$2M�Z�1/�v%�cڿ��hEO�Qg܊KO���4@�=)P��}й�+=*��|����˹����?��ZM����}�!}�6�Mj���4陲ߞS�7�h@���O��aY�Jp��t"j�h�٠`1��J8���:ҳ���c��d%��N�P�CG��kĈ2�x���p
&*!�Y3��T��X��-��g]�'�2�K��T$�B�]�ȥ8��0n�n7	���u����ǁ{m��^��ڔBl�Bþ{LE��(�F�qV|�Y�̬:��$�E���t\}���Ep����?���8����"{>��@���Y��4��b�.[b��Jذ���k�i��|���z*����FTJeX��x���IöqٍAVC$�|I�>�w�|���Gd��2�~ �4����֊%{F���8�;�S=�[����S��`�= ���?�� f��8�1��2t���p�@X�w�>;���s3��=��S�PD|���t͹m
-�陛E:,�n�3�02�Ļ�8�`iLz��mȸ���5:4m_nee�ڈ����a?��Cu�N�4F[n��P���08*FЌ��u������e�(9���!�<��ou��/`A��C�oA�瑱#�+H4�c!�h�	2.�hz��k_���3/��9#jK��whNQ�in���y�4��(��8"�ل��o��˅>j_�+�7��꣊H�Hּ
���39�6���D,�*&��)V
{b­�_�+m���mhB�	���i������;�=�NM��N�~af����e"u5�l����@B����AP�i6b��Fp���{��V��q�Y�cP�QVDfq7��R�|�Tq�n�E�%���Ҩ�kil�
)ʙZHz/b�_��uс�p�5�t������_�Al}�u��ŵ�`~��[��&�)�{���Q˩KFJc*ǑME]�h/WU�5a b"��1��|��>^П��}���W(��iȨ ������66A[�j�M���Kz̈=�� ]ǡ3�#�H�j���~P�V-��g6=O�暱��&l��h<8�M(�F[Q�k�Y�MV��d�p6x�d�\����ǳ/��Z�K����c6��_-;d����R�z/?�!c�> /��	�ƍ�{d�%d���������,g�V�����S/�������Ŗ�W�k��<4�V�lt�Иز�8='�ާ���{v�gI�g^���ٟ���L���5�~ko��9hn"#�
��D�
�J�?h���W�4���?��J�[N���������l2y�Ɔ�Ju���C�U[�dI*��*��5H/-�R!��r��H���fp{���6��422|���CN�Uz�MZ�VmB�H��Y(�����Y�1��V�l"�Z/�z�y=���w���Gs�߰��'�t5D�b�Z�x�Pp9�ށHJ�;��f���BD�']��7���[�f��A2�}zn�`��j�!\;�J�*4����Zǽ�����]���b: ���!�t��V����x�a�֔u�fe��>�2R,vԴ��y�3�:���Il���5�Yb23 �Ϥ�<�>&I$?�x�5p��BO����pf]�/���~6�R��ȯ�d�D�}N�ÅB�!�#�QA+Zဩ�����_��G_���>�����/�h����O��PK�F^d�3K��R]�J���*��.���e�|�V����܆2��|>�RXF{{�C�W$���;o��m�ܶ��##�-�pm8�R[lۅa�(!v=��D���g0n� �^�/t+FK�B46�F�V�!�X�c9�z;D�Kp����d\���A�v��a���`dD�S�(�MXг�WAs�	�s��ĳoԅ#�{����\��R�Z:��Lb��I��K����4vJ=�~��!��@m`e�N���#���壺8U9`���0�� ��H��T���A��h9�<o0���j�+�~G��M� &��@Xsi�h�
�v/taӢ��pm��Y?�~��^ނjK�6(|�PD|��E���9i��\��$pu��?گb:�8]}[�8ew3�~���[�O���mD4>232,yxF������I8c��q:(�B�iT�Ô�b�~+����.�Pz���ٯ�'��|�~�ݸ�W���egX:ʥ6RaLċ^�}��Gr��m7[��W���ј3e��7Y��[Ű�G��,X���F�8�'�/����>�#W�H9N��wB:�����!o���������H���z���4�׆�/���!���p.��8������R==3R��-�1��3#Ljc'᫘~ĵ��� �"\��8P�3�u�.tT���,N,ǈW�p�;}�-LƟTR�wEė?p�e�:��h�����+�B���$�F�������:�$S&W�Q>(�P���&2=��J�G_E�!�r�m��m
�M��PN�\.� �!X9���t�T\g�O���QϘ�sN�"dd;�TdӲi��D�]Q�M�i�ဝ����>��M��ws��_��R���'����+��RMܴL<��[��H̦k�k�u��,GI��>ڑ~̯�LC4�.��k���ۧ(U�-���1Ms�Æ	9O��5����b������~��7�{:9-�M�����`�6 �8�t�4L|�ʰ5��3����h�lkj�9�vT��T�6x�v��^�i��~���9�iʤ�+��ܛ_���{P�N����^}
ڔ����YX,ܮ��1R�D�PD5�+H8�("��H$�(C�M�s�p^d`��Y�~�ѿ��VZ�V�C2�z۪*&��A�!D�2Jc���S;�����񿽃�	� r!�J�!m���4Y_	����눈+Wsm��
M2��ԫ���̠y���'�k�
�4>��~��>�k|��K���O?fr��~���}�������FY���DG�ɖ��S��G�-Z��n̗O>?��F
a��x�y�Y�tN�r�p��-\���^MD�k��7�?{57^z "�\�Rgd7�-�Z��r��)AR|�a;mz��W~���.��-��wEė/p������4�,OJ��p��E�;L��	Ҙ��$F���O�q�V�=]B��\����pdC{��/Z�[m-Kpm���ց�!���[C8U�׌�)O�$BDs���ܨ]�_��z��ZT�H��nҐh���$�h,Z�:�4ۘ��0<��GP���F2��P��hqah6��v�/�4�=��97�?zu:���j>��4��Fgē�x�CF@io�1T�������*+��� �R7�4P)�����'�IP��Q B�V��R)�q,y�dNmaeD�i�|T[D��%~{~n��GD
/@����h�堼�w]B�xC[�nM�����8�ZVP��]�;�"���N��v��[r�$��B�d;��2\�lA�����7+�����\��`��b�0�4ړD� �'9�����c"C�!']�j|����J�W��
��	1�MH��)��k��,�k.N��z��$��=�#�O���F`�N��$��5�R����6�;qU<��E�k ���(�E�v��x��J	znVh曲n$<|�i�n9��A����[����H�
{5a�h_�h�D�#�?Zj`̐q���C%^@+�恥��,J�]��}V�O��z!��a;��"r�2�C<�t=�G��c��#�4�ɗQ�`�갟�g�)͉���uS�!�E�jFV�Ⱦ%��Q࠰d���A7�t/���4��R������iӱ_���k��Gܺ@��� ��/`N�4�~��;o���E���ʬ�
]��Q(�7>c�L�3!��r�}������$ .��>�_�z[.M��$S�g��kD�4�b�B�4�(�e4�G/�:�����:�s*]?�fU��%��1QT*%��1nU��2����B�c�$�L���8���P�jm8W�v�at����&�@njl�B}�X�WKv:�;5�����c��zC{�R]/��C�8�U�Bv��ID���1�Z�<��.��n�����Fd��V��� 
K<��Ǌ;��������?m��^s���X�1_>Pԁ5N=q�]o���np+�����وS�ޡ+�`7r�1�� 4e�Ό�dGh,6�Ti�O���?=�'_��oږ�_wY�'&L�a��,�-��8D��Ѻ(�a�8�?�V�c��#�b�MVE�O�T�dg�fiRl'�y�sl��*x�o�lVg[OF�^L"������k}�:���g��^����Br�K'E�����D�{5+"^/�m�� P"e��Z�W�4��^.ן����j��a~gb��|uI�5��z���sp���n�oTu��.�r�$�a�y:GU ��a[f4��#w���c�
ͼg�V(,S("�݃�n���z[�Y0�����A�YyN?gϩ��ᥰD�Tt��s*�.���L֪���J{�%0���q��/B��A�~+:U/~� M����5����)'/��j=���;gc�MW2&�ȏit�`�hǲ�
�.��k��A�z2ry��fB�Π��`!�fQ���R�F�)����d�O&㝮
&`)�Z���B}��X2�Xv:���7~xa�E;������l�NȵC{I>�p��cP�~Xo��%�aE��7�$@�W�%�=o�AhqX.4�����2e��w<>��|�Ga�A�����8����MYc�ޮ��|��YH$�S����uR<(3dk�8"n�a@c�G��f�����
�zH�����!}ah1a��lX�lP��0������]����:ZJ�64!����0�1`��ӆM�Ё�P��v�	N��~3d$�kߑ�ຼ�|�ٿ���S\�. �B��ϿI8��[0�e-�Y4_����tZ�:�j/��0��Ä�V�W^��-3�2���6�Zfjy�v7�p̴^��^�|!��	��eEĿ[غ�u�8`�M�.l�5S��l���j��j��e0y����4�\ђu㩦ñ��ǟ��N�:��o6AFuCpc`�6���LY'��&�(�D��7>F��[��r�8r�vRxH��f)38m��)�,M�]�æЃ�{!��}5�s�X^ܶK�?��9�l�U�A�e������6��{��Vv�?�L��,=�����4ё1��LU�5y�0t:7��~�������{p�)�`ؠ<����G����X�`qMߏ5�
W=l��p���̥�����_��wEĿC��O�o��l���A�YF�a��Ry!rM���dT\a���]��qd�(�`�����8�;	�/1�"vhfV�p��6n�ʖo�Fx��uU�^\�{�=��O�I16[�d��;ddx�;,l���뭊��x
=m�e"⮼�R��-���3�4����둼��j�rkHmm-P�p���;��;��4:�X7 M�s��mU�C���2�F�����У���z�Ǟ~�8k?�m2e�fAf�*t���O��R{��I?�g��/��!&ⳡ�L���w�V8q܀���|�I���I�-f�\�6�eAX��@W�e�4��̽�ٯaY9,�_��� ���栞�D�ۈh�dV�R5\�m2�b$�.��ޜ�z׼&Iǵ�g&�-$	�LO7i~�e��\cU<LD�>���ֶ2��-�X2��U�m����b�%ۮ?"��&�~��B��T���}�[�v�ֶ��r�HG3�"�S��8ix^��z��rr�d�?;��?5I�Xk���>;�:�z�:� �ir��Ь��#��6��ŕ���6�p�����އϼ4�]�x.�L��"����Z��}���:wXd�/,����ɏ��!�*����H����l̈́��(�!ι�v"��Z����hj�M��@�
�ˤ��kF5ݐ���L�M_}瓨d�[0J��s$��Q"�
uX2�ѡ��kh�u��p|��<�6.�h<6^8�W�l] N2��eHB���ￂ�8�a�D��!�U4.����|�
�����`t��L7�āE"&��DA�bxj�W��`���,X����]	��.�·��11h�p/m� �Y�Cg�i�މӎ��\
�K��B�)9�;f�Ï9�4���KHRڳ�U����+C��{�g�t��D?@�\�,�� ��/{��Đ#�|����f��D���D�:0� y2�c�Ob+�e�=��?i�)a
��T/&&Z*׏�g��/���W�����ZtO�Gχ1EC�;�b�k�L�(�h�.SmG�4�����u��B��l���"_B$����P�|�ѧ�r/�aTU��8g�y�v�Z������l�>�{W[���LE�d��X���4�T�����,�`�l�g����q�߇i����@K�t��BKe�u����P�]�R�����q�ܘCgl�ť��3��q?_%�эPD|٣y�5o��zc7K��K�&C�B7"�`�y��Bh�<���q�~A�
�&XeĊ��{���F!ÓϾ�&���eH65�г����]����f��p֝0�(,�n]�Ùs768���kq�X�i��=�y�/�W�x��/鶯[���,ݐU�I�����E=a��p�Bߧ��:��T��	��4Sֈ�zY��������/~��ǌ=օ�^�p�� t�D�y��»
�+K�R� J�X&����t��S_|��7�x���/ �.("�l�)���s���~��n�IPb�	�(��9<��k��/�B�a��oFģ:tK�7g�L�C���BAE�{<�zH�C#�MƟ����v�i���鬐q8e�<�܇5O�9Yf�5G�,���鬓Щ /�ƹ�g��ԗ�T=c��Vp�lGʇT«�i�72{؎�Q����9��-���Qhk-�W��Em�0s�^�1�h�����G�t,��ַh5�x�%���֛����MFoLuӑmC�+��q
������uZ��_�M�>}��x��^���UEŻ	j/;�)4��6ޣ_�=:"+�la
�
�n��с��x��\y�P�f���}�����bC��� �1 ��2U�K���� �0�<�t?�V1�J��a1HݲF>�r�F%"���ǌX�dΈ;�r�)ɒ�	�[U7�z���0Mq�&����̚b'g�葎uƏ�{ͯ��*>OG��ɡ���"Jq�0d��F\6�e�0�A����W��$���#z��Z`�M�\K��@�n��PXr��.�&�Y�|�8�H��տ�3�=6���[�×�T����/;Xux��6�`�z\���%�/g�ǹIP�>�������
����?�#�T���8�a��:z�76����悅��DXH�Zf'K&��%LC�j����)��5F[L�������`�ň��n`�vD�`�,j��UgLUgDHgm�B8�]������ Z,Ϡ��W>q�p��1XB��y�d6�2��4DF����'P��?p�yw������~͈C�3aY����M�l�-4â�9���#��L�L�4S����v��S���_�`!��|��Eė8Ck���l5�k]0B#r#�h�}�-�;��8脫����-߾	��CQ�����3��{:�>����e�	��-��F2���nˊ��L�W\��JW����G-����d�!�M�T�p1:����'㎉�C��������y��2��DcG�N�)c��L	��α+�mj=3pʤ�pAH$<����UC�b:Jh-	B����/B�� �ŏz3���Pm��P*�'�.U���)ȶLg�As4��ې$�k�t�A{l��ѧ��!��y�:
K��/<`�7ѿaR�n!�<$���6ɔS������ھT���Q�ͣ:%��7Z��96����m7��D�h$�9A�fR��4Y���>X�,�֛����G�2��l����i��br%S�|ei&�Փ$�ߞ}
���}F�O�g�&:2%L�d�'	qQ�&��v��T\���r��k�k���F8�:�@�Li�P�*g�z��O���`�Kn�y3���ڐɬ���5Dq
K�f6V��Lˑ�p�\�~~��~���y�������6�*�~�уI��hҤְ���2,� M���jΒ��ktC��A2 S#B��p�w��9_Aa�P��+�mC��yp�#��j��a����/o_�.b"�����k�Jt���L�i����Dl 5c�'��0B�M�K��lAO���=Hd�1[r)���jT��,������
���?k'��@O*�XJ�1G��08��k�V�cݵ�׿5�N�	κk#�ӆ�[�0�Й�mUS�LL��'�G����v
��~�g_y7�9t��G��N�`E����W���f�N���4�j��o0E*�6Cՙ*R�eJ�-���+��������/Ѭd5�K��w/��v��춽��cu�t2�L�^�,k�:T���tt���a¤��Jz#~ߓx��Y^R�I���2����X�5�lOԙ�Z_4�x��N�	�L�R���^Ͻ�1�?\f1ED"�aI�����FQ"ۘ٦��w��ڃ���O�E[7CI��Ɛ�w&8�iH�V�gV��+�I*���h}J���^��Q&�l5ϵ�|v0	7���� }W�M'��_�x��������L#ؖ#5%p>Mj!�K��&rd<zeT��t���/��βHpw[��]w	����N����n_�{�}���>�=U]uf֯���4����gق��^�`O�����4seE��"��,�0�Ǝ���tr�x�3�ѧ�d���9�r[gY���o}3��p�J�e�t�<��M?����/{����vQ���C&�ǚq���!�)��������m$��&��O;���'��\�DՒ�yR���Yx�M�`}�A�3*�$�M*�r���g<��Ʉ���f�����3�st���ӫ��ѳ
e76�V[H�l�p'qN���0d<���W��m�ՠ-z�֮Tu+�A/D[��x�~�-
6~�gs�+Q4�{�}r�Kw��U�hb[���O�w��l_�a���E�2�
AE����Ca 3�#	Á����
,��s��'`�� ����;���^4�YRG�R]��P�ހMMO�װG$�-��
�m�͵EX%�����d3܁���e���˳������$)��y��.�v��xߏq=��h6j�:�T>g~�wc\�%�� +Uu1��|��Ͳ�Ԕa3L�`LC�r`�(|��_2r1aFb���K�K��zPSP���C���T�B^�I4�f%���%aIr�3χ�a�� j�G�G�n�s�sP�;@XO�_GPT�\���3��?�hb��:��9�n/!��f+�Y�f\�y��T��M�D��9��
-��ʨ�.�F'.k7:"G،�l����ó3gau7�ℤ��&�Һ\2�L��� �"��"�:��6�sxO�<ޕ�K*S']�$�������T.Gz��0��s*s��gm��]���t�sߜ��R9����d�J���Y_�F���9	����^���J\�,��=o�D�$�������Uf�!O� �b�Sղ� 0Ǘ]�h+!������B?�4� w�;�S�g�V�5玎$�nBcw�$y/��l��M�>��N��ȍ����5����l}=��'0�'��f~<3�>�K��V����{��c�c|����1���#���`j���MLy������i�}p��7�&\~;�T�_�~Z|&�M�������#�.�E��r�%���	9�[4l��&������%���,�����`]���KP,k���-p�%��q������ �����:�����0�I��kj��1�h�))�g�K����#�'�c�2�`�ࡉ!���	��@O;T9Y���se��W������;Mk*��c�)���8R����c����3��o�ȠH+	|s��UF�ϻ]K��Ȭˬ�+�R��� ��4�{��v>��i�_�[��;!���9q�&�"%:��mJBۤ�:;�l�<���)	��c���ڔ��CY��b�i��i4E�[N�O�i�]$�Dy�T���n2r�\��S2� C?�Ʌ�/0��o7sX�
P}���:�������-�
�#���<F%��鳴�yy��4G�ݑ�5&n�6��cG�yz��mwz?>jG�X���EBq�U����~KJ��cM6��65��mF�N��#��--�r\�N�d ���ߊ�c�|d����]V��� D6�8a�����5Z
�l���"�IP�<���\��y��%/����'t�ʃ�%V`��7�-��*v�K���3�|��Dp24��a>�ε>�ُp�o��-�P���GN�_�i���&���-�cw)g/{��[���B�u���f�b��A��֔����Ũ[��O��?~�Ù9o`�}+]��k4J��jݜ��9Ӷ����#,E�5D:K���A�⿯���ݩ�����u`��<7��P�D�$j�(;HR��Uś�]��#�QЅ.p�'����.\E��_��O���p7Z��̎�L�m1��"���4�����%��I8wSAR�P��}��t~��(��?1��o��e��EVT����O�}����=n��<���%G�=\���/c��;�[��)h9��:��W�Ъ2톄����qt��6T9��|�J~���L���Yr�##��-0+b�ܑ���y��7���|V���z`��Fk�Jo/Ȧ����%q������<�k�'koBء�+,�OR�ٗ�7K�h����]�[��I��_$�e�z�$ӈt0e�\�od�@�p'�| ��^w˖���86�d�ȋ3��,&����fk|�+,�6q��M�p�(�Vtb�^�c����mF��8�(��4�C��4τ��0#�)�d�D�͆�/�6����?O���:���_ �Idp�D�%�h�x� ��U��i���2���;��;�4)�de|<l'Nj�JeHg���0�A̢���塺SQz��|���PFX����px20�#�Q�܌�.�>5���.g�ۛG9TW��զ��_`�=��oP�A�?�F�Eѵ�(��=us�s=��^��L�*?1L�D�S+����-d��b,�A�t��5�gY 9�Q�U�@P���!*!�C��Z�+J_���^)f���iN�� �@�~\ֹ_��a�@�^&�ؕ�e��a�r�T4j%*i��[:A��Z�'����6��kI~�	�Y�����dY�P%�w�:�T�t��?�bs8㽇���P,n������[k�?o���iZ�m�'��U��t��&��e��>���ӡ�Q��윁��9��1A��k�ȅ�"���{N�F2�xr޹$I���E-��e��9zg&
r���,��wr�Q�=�˅m�P�f�2��r���~.9��Պ�����ު'����`Ǣ�pMR#�B�!�DTa��H�'qa<Ì�	Q!!�����̫;�8����^�}�\R�[z��-�K飇bV��U�O���Y��.��|�����IV���}(1��̭�����m}=����^�X�m^������V|��
b��l�v�(_�'�� �����D�Qiv>�TRh�A_�_����E'�/#ߝ��~X2��/V�d��~yBS<��$< z���/uS(L!C�������IԎ��8���(,%߈�2���~�n�����)׫�(G�ʉ���!^Pb�IÏ����P�x�ιA6�6û
C8�V���>�w ��^0;�&�](��8�|�:\����C�����}�"���8Y�����y.�,JL��4i�49�:����Ռ�I&ti���}�s�i��b��9S3��qlsD�U7!N��!x�:�:�����1v�KĊM���DH��dn��ú�:M� �77#���ŋK�Q"�G��\������3Ug��t��.��\�%�՝�.athx�?7��?�\&�n��Xz����]8O �i����vCq��F�M������":㚿cj@��8���#��Ox�Q���E�~�5�� 7T	f���j��o��5K=ځ���cn*�1�?������z��G��]��j�e�R��bw��kEHY.��J(P�Q s��q��x���5;�������ߐ�ϸh}�qfK�H�DӯJ h0���i����Z(i��.6�_]7���r����9��J�"DNJR*J�X�	�_;S]��˰�$��������?'J�T>�:f�o<D5��A�G���~U���Q�J6�xާ8 �=�@��Dyȿh;��m�qJ����������v�I$`��*�d��5�/�/S�~��G���л�&5h$�e�nJ���	[K�Q�5�.�����3&�9 ���vD�*�`6;����r����D:ۢ0)E�B����N���j��x	�槐Ϊ_.�]]�:��K�G��R��ј�r=�.��K�6U����b�������޼?�T��|]�b��r��,sr}��nh@���ȗ����s�G�1!P%*		N��l%sm�6�؎�!�o�{K�ty�GȂ��KN�e�`T3{�����~Z� �v�ys6�l�E}M�pζ��L���#�3����UqlnG�o��s�Q����͉zź�r��!�e^� Y�{�;p��a�#*���D:�W�������-����5`�Q}Jl<�r"����xLVX;�nD�D��q�3ޟyVpߙ,�ݘ[/�w'Rt��(�u2�ue�3e5��5���� Fc�G<�[C�R��u�o3���>rb����E�%.i椊z]\�k�b��S��&M&x���x�|�}|����vr�c\����H�hRm7��S�H�(��K���w�"�1�%���E�y�x�*��GU��ő<|�_y>A�"��FJ�u$�%�'��F�]1<`��1���mBÿ���iK����y��&�j"w�Q}�]\�X�/iH�+��|Or��bpٸ�rk���7�'�����R��4:m����䤌݋�����]�ǖ|���p��b�GR\����ye��o7�V�1�9餔�z�s k�)�i�L�����M��_�!��&6a�8B��%S����}"m0U��o�M���[�@W��f�wD�ǂM���T˭囇���&<�le�?Q���}n��I�Րq0��ž˟����m+�՛<���v��3��f�n� G����c �Q�݀���BP�}��)�21��O?�R�D"Ol~��ͬ����d��:*�P�$P.b�p�q&(Imv�N����>[��۩���|x���K�yB�5n�Ǥ�{Ӵ0
�%�̗�J��i�A°K�)�(*�c�j��W������;]��EiQ��SH\���Ij�#����~�!��>����"�}/E�G4��<�F�J�I~���ڊ�T�1������)��,>�٣�"h�*�L֎R���X����ӗ#7�KI?�Y��5`��(e�g�f�������7\��@��,���"�eNB�R�Q �PUY}�O�γ��4�&Q%3ǭp�#2�2�R��!�u��?+:��:�-E$��wAC����p���jx0(���?vy0i�8 (��gg֬���h�j�a�:�X����on,ڵO7mD͆?��]ݶ�liX�ZHW4������2c�R#�hy,�3kHE~�n?�PH�u���me�fI֊JDD�����ǒ [C�J���m��?%l��F(�%�� �sAZ&υ��#�;K����t��Ʌx=D��ʪ �~/]�BQ� <�i�q��ӅR�5�9��g�7��ڙ���.�Z��2D  |��P�INL��zq�d��u��� �kA��[�G�i��2W\�oT��ьJ�F�n�qįty���D�=��ṔOt��K,°��&�`A�7�.�f�}�'t����͒�����7�%���[�.�?���l?���S	̰�uXc��ff�2����`$a�J*QEi}*��yv��3�̷��l�2�1�.��ey��7)2u!<���O+��,)�l�wM����*�o���z��7���8�C�G,�/K���J�^%�����/,�CO��je�Nf��׬K��>�������j9F��W�C��XO�at������>��O�2���9���w)�o�5��%9�Z��k�D�
��Ѭ>�qH��Erb����͉�����#R~=w&^7�$DY�=ĸ#9N痼�'�MPZd]BPo�r�6�PY2�R7���z�i-�(��4�$M�E�0�yn��4o,{��ʿ���x�`��B��?<�gt��VT��&.� /��N���hւuƦ���6�h����ȟ�8�n�$��s�[?c}��ߋ]��<�G�4x��c���%��j�R��Y<W�"�U�?�}��V���c�xbV$M�п���-�Ԥ��=.>t�h=��..w��8���(Sb�$��QUn�DN@R)(R�c��ؐr��#��>'3��O*�l�e��(��CB��u��~���5IdqjF�A��0��W���QMwq2<;�@\�d�1x%���T�?)!��vW��1&hd���v}E��w�F,�B<�i9���alɔT�!��h����i �PYi�FV1_���>�W��1��Z�ȇ�v�m/GvƮo.F�B,句���#��n�|SQ-C�Io(I��H��l��&��k���< M�#���8�@�>����!y�F�0�q���tz@0W�0	���<�F��ҫ�R�(�D�Fn!c5������O>�/}�Q����w*�c8	�-���&hB��f !�DpF*4˼�R���>�"G��(,������ϛB������ϳ3uj�ي���3q\���z�Hc<�&k*����$�,>��XlA�f�Z��e��i��1��|��`ہl�[P��d�+������d�Q8���}AD(J�c9��kVMO���p�P��~N @'�Dne�^�҇M�w"�1�*�>Z�Qwr���z�GX5M?N���.]h�!���F�$X�T�12v���cD��`!ƫ)i�C�������55���|>׻�w��f (c��cxԃ�G"��G�[#(�h�'A�~��h� l� �].iU����5]��l�O�����GH�n�βդ͜1���ꙺ�rdr��<�W�8m$�uZ��b��J�/��o���b� ����(P��\ �\�
���(�moR�#h��~��D��t�����^6d�-�OW�a����j�8"Y��+�6e��u��z�ƽ�}Ή}j�ԉ�Cs}Vya���=��>�������J�8����6�X�d�1�n�"���c��mt!Xxֳ�	C�`4�,)K��Zq��|�*�^�]��Z�WcA�0���}�<��XA�%hb4k��}�xֿF���*&q:��h<��Bd`�?ɀ���lc�#��H�I�e�
Y��L}1�f�Z�9\J�-U�/�������P=�Yn\�:����������*���M1c�y����Dޘ�������.!3��sz�<�?�˰y��ɲ�#��Hc�xU_! ��x�O�aX��M0�5�g4��3%���y'���EIa_ew����n2~T�d��,s��3Ж<���9u��3�K�Ғ��S,�F���
Yf�,��U]jwl=T�'�c2�IF �Ϯ$�>t`\-�A�IX��̢�aE*�X������ ww���g�:Y�N�� oH�*��$�Xm
��o(�k\M�H�i$\�"}Y�<�v�y���Zh���`:��X���sJ]�`�v�����B���������_[hB����^@."C��@�^�~S����upIT��)2�{2NNƯ���P��)D�5�PE��La7-�=`���+�7>�T�r�郱���'��al㑤#��!�[N�zނ2^>l���"�����n+��`�R.[5Q�)��#����H�Vs�BE�/�&e-��y�})jTq#�e@11{���g��R;bb{��^�sm~��*Y�|0�
L�0o�̉E��@hA��Ry�ڜQތW�`G�y�a�V��^����G�Nυ9OO{�
1.��L���[�(@��;C�Զ 2��nKKl2���5��T��1�ڒ����l�ǧ��WUH�h�u��{7�e��4;ޔ��j�z�=I�8;~�}���Rʯ�I7�$�3�{�0f]N{o��^&���r�0OlI�8�#v^�A��[y�����8O"���[T��o<u�P?�*	G-�g5-��՝�1�֦B����U�BE�n��91�� ��:�FFM�p���:W��<$M'��]"�F:�ЌJ���JFǕk�&��?��|��R��+Hy�~oGUOSQ�����o�H̃-i�Y�/�k�gx�?��M�k�"9���#�'{e�^��kvvR���gc
ݮ"��&n�)��
GU$�=h��]�9�EZ��ۓLA�fJ]HM�Er����B�/"pO
��B]�ֱMd�H�m�I&�^\l�-=ao��(���!��q���e���(<��l�B���
'�ٯ�[��H�E騷� �Mr�"�G9�!�s;lP�Ր9��,<E��_u�5��w����n�A�a�E��5�n�I�%pW�YA��KQ�۷�Ob��g|ʽ��:܈�)�\O��� ����P� �Q�R���s�x�+�*����
R�&���S������QH�XD(���]Mc��]����Ms)��_�f�������DH� �J�w{�x�7���fq�}vm�咱5n]�e�2�_���U�%�N�B",�7��|F;5��<��l^�M@.��n��ߜӃ,�ůFU���9ܞ�罯"C�7C5D�x[x�I���>tdd8H�_�m*M0�5F�k	�����!�Pt���m�A�4���IV[�O�W5�h��|{^���W,�#�l�'0>�A+��Q�)\���X��k/}+6[�w� ���xYMw��v��#*|��t��?���8SH�߽��L2ՠ����"O�L��G2&����c�Y�ܒ�dU`�؝�9ǵR�>y���a�ſ���␤��\�~� D8w�!��+�p��E9ߏ�FdGH �$�� ^s�'Q�yi{E�]6XT�EKD����b>�q%!-�8��=���Q6=���������S�xu8�x��c8>��r}��4s)������@*��͹��A����c�����ES5��16�5�pY.y?����V�\��4T�ӻ���`e\��o�� >�T#���O^��^�0�W�w߻���~��yq��9�����\8}|9�蛁���P�D2i�dMs_"e�b��S��g�ɞ�#;���~���n��|u�m��pt���۪*D���[mD�2˂(�R.�)��I�����n�{/�k�Eei����}<��p|�[�X���(-Q��j�;a�T�窉v����`�8��%v��U3�����F�*��V�QLP$+<H�%Ӎ5���+*�*J�tڝ�*�H�/D��\|���+�&`��� ��~!T�)���s�ܑ<矌�(r���*�mӧ�R/ƞ)��y*���|����k�|�p���|���>���I����E��*�����5cN��<i7p��g�F���QE�����'�Ӿ���Ţ����4��?T�2)��I��"�����~�YW�Z����u)��h�k�f�;0P�g$��-a�0r�$�E���a�$�D����By����3�'^�/�#�>$�>�uE�d��`Qc0l�׃o����:�q+�
�-�4�s�?��e�/0+ˉ�|V/�u�]6E�tRcy�Wv��1��<�d�m�Z�C��%]�Ɲ�����*4 �%��Z'yC�B�eW%j:Ɔ,����]mX�~�ʴ-�ց���a9l�dX͆�\�q���� ��g L�!W~�E�\�y��ѻ
��J�b�@�?���R|`a���o��Q2�9��,����>i�Lڬ���7^qPf1p&�K����.O�IC��J�9 ϑ@;�o*J��i���h���H��@!2ݢ�@�Y�Y��@����4�����ì���Xi���c��FNji���!�E��f��P�E��6C���!`�A�A�1� �n��\��%��#o���������a(��[�u\��+�t9��pv4��s?/�cI�?�'m��:��4�D-8�<C)+�<X�8���*t��U@�������[�,
VBJ�m�j�Ie���֟��O��E�����3���p�M�Х"U�h��t�mr��&׬Whd��}�>��*��㛆Y}�=�Љr
;P"��`�@�����S��fܗ��h��UwN#��k���M�2�a����i��i���yK�.Z)9�&.ж�$E {9'�`O �E0���B������Z����z�>�}=�������8�+���Б���:�8Y�3T�jЏ_L�%Ky�Խigʅ�P�Nԟ�����}�cJ��yO��������S�⼴
�^�� /$���4��k[Eq�㟹�k��Q�ȡSɔ�RF�����)�ۧ)��/Y�sU�(�$E�V��03]mX0�4D'���{��N�?�D��ul�U�R�4jV�yo{����u���j��kg���;��U{�B
Hy�3���_�ƤBBt֬%/C�f����/�ʢH���x��
Up��
���
�J��B:y@�څ�m��u�]5x7��CI�֋��	�Vb c�5��	P�=/��XJl�gI)�����j
|5R��0�ݖ��j�lfAA�r���%x� �%4��b��b��� 8M6��&�#.�1��S���*_A�.�y*���|=��G9���n��RB�q��Ui׿	�xṠ�L;���X��X�bvl�A�lwu�=�Q1?���r!��!���8M w��w4D7�N::�CVM�E	/`�0(f��@���$&�a�2��q��A�q3�O��([��A�B�C��S>�>�QKs=�0nO�'9�c;�8^��T�d��J;d���#�U�*"Dx#��4D&�l��i;�d�|�3��J�D�;��];)����5@�엪�t1�N�Ы\�ϐ+�GYO-���*�͓5���Z�~��C���w3%�b���68/�-����&��	'�����V�
T��9�cX�b9��7d����=��L�[
`N%B�A���J����-Ϩ�7t�L��e7�_l����p<"�J���������D�B�܏��F�$z��,/x"`��Άo慩�����2������&��׆�Jְ%M���{2��H�����7�=6��k9����o��(p'��	���)Ep�(�Z�:!>E�Ҩ��2���"20�Fᆳ:c��!�L3����ߚǩ�eL����2G�oT��ߏd�++���bw��'�����L�R�P�Hަ`���S���x��x��0��g@�y��h�ֈdK;�+\��E�_�[{P]���72c�գ,~v�cR�0KwcL��*U���~�r��̒@�֕m���",����Xsv�eW�boe�����g�C�/��W��ϣׯ�]��e�#0��l�+&w��;ĵ�����Ћ��4�%,=0�L����2�z��':����2��v�e�cd�z,����|᪬�~�~�ꅜ"i��c� �LtG��aco������3X6mX�d�_�F.��e����}�7�����1lػ�ǎ[�䤴�4��b����?��j�6Re*;.�,MG��O	D+2��k"�/��d��}�&�Y���4��+�ԀIL���*�4v��#>W!�lԶ_��b�����;#��\C�Mp+��+����ޑKF!ςT֜�ι
���#�F|��������J1��s9����?�ƶ*�Z/=b�$��Iq@�LF
�{��c2��Lh!)�@��iV�d�w���KC��c�j�����^u�iz�ݶ�&��ֻ/q������&(]q�Y����*`����H��es8�q��h�t��W��{���<�X��T�YY�lJ_��o;�@�����V�n{w��¬ǳ�=@m��b#���������,�oB�FZ�����C�Ԧ�i����k��@�/��xs��ez��(#�lޏ|�4cc���oq{Y�ru�~1u���yTV{�����PF-C9B*]��')��/L���k��HUe��	�G@�.)׫�ݪ�F��\$�J����$p6�ĺ��9ʆ
����Į�:r�mf�����פѱ������G��Zv��q0ӻ�����;����"M�x7ke�R[t�&k��3y�v<���(?^�`��\������iӻ�D��;��Xlj�:�����H[_Cɑ:D���?��S!�K��bx|�)_���� �}Mn�7|+��u
W'elA1�<3|���8E�8h n׭�������Q9�l[��D���ɡ!r���˘Om��y���޲S�#��Sl�� ���c�?���8��[�!�K�;��4r$ v;X���6��N�ëoZ�
g����z�4���l��4�o�t�lk����tn�)KHK�ɮ�,�j�bC<�)����p��1�֟�VDq�5aϣ$&�5�@�%��O�d�jî������$s}��{�n_��q�������@ό���TB�j��=�T,I�ߗ�W�;)�'z8�;�|����.n��φ���fJZ]d}_�./�n<? =,vS[Ӛ�Npk ~rV^3��*׮5J\��7��9������4��9����y��*ȡ�q7K�2Zr��6^75%R�Edi;D$km��FN�a�7ʪ�j������%;3o�3�X��s20=:d�`�T|L��|���j������xy�ᙶ@�*�S�����Y�`I��p�5�t�|An�qܴ�#� ���
Q��ҥ`T�(������E��~�o_xx���z[�ye0҃ESͨ�����u�P����,\�2r�AM]��\��c8K�f�����뇆��ہ����P%�R��I����">Y��44��ֵ�_觍��Ր�2����O(͓��ː �HК7�!b��:�V@�Y��Kc=��3ό�8��(��`E����[�C��b�,L���<��E�*�!"�N��H�0AY�u��y�~?�}#	�o+��z�E$!���%ÓX��ʨy4��~rc�ǔO,�d��3�h��'~�1�*_��|f�,w1�0�1�&3t��fÔN����&Uy�Zб������(��0%E����ݩ�s;}�Q�6&���g�9/�"f��u]�r9��U�_�^}��L
8(#���Z:��D���@ueT�C�+�\D�(MG�-¾��̄Z�$Y!ĉ]k�Q@����$��)/L�|w`����Nr���D�L�#�:����x=�/��ï�[Δ#���S���*�X|+t��ᅡ1S�Kq�+���ncr��y���f|�5r���/t�/�H�G?哺�\S^�%q���Z��2�K������]����5yQV{�(�߹�>�e��خy 1r�hݹB���r11s{C,h!�|��s8���J"���.:.$��K�Ʊ�����/��-w���"��4�y#^�C�5J����o�s�<��D�#�N�l��u5�qЄ���	a���lz):�(�m�ǅ�=Ea��R'#������j��V��Hı�ȓ�L/u��X�\�]��͠O���(�n�n��@��h����GV�B�)�Q�ȋf���@��*Tَ�Ekە*�����Ћ��k�>X��.mPhx����~W���3��
���Z��E ���8��y�W�A64('nJ��o��AP����)SV�؋��9���K	������O#jx�(�(�}�?>شł���v�*#�6��dK�i���F�r�e��#Y,�H�bO9�F&��Ԛ���-��.�Q>a��D���v��ʽO�\u��x����q����#<���~7��P���EZ��h�߄
կLˑnR�kFO��m�>R$�Eb����nef�jI���:�=�MUOw�v���e�KN��R��s�v��|���S��,����|�D��]}�������.�W�yX�(�EjnT\yK)q�-ʘA����*��l9�b�PƤ�"��2Fm���ژ)��b�K��SȢ=��?�A��!�i�����NJgr���Xk�h�6�� ��~�5�S�>jU����\%��8g��z'�46}U1H��-+���6Ǒ�m���D�j���JY���o! �UD��vG����(ܲ�E��&"���_��H��.{�j׭nk#V�������qx%���m�9�Ab,�@��&�`�y�=3�!H���.n�7F�u��s`T+��@#�I��]ӗ���pM�BgS
n��23�勭�J�M�G�h���\׊��}3���z��ԺB��_�N�@\ف.a��<��� /�(�>�0��[�����n�T�[�d����p����SDO�V�,���e��A~�F�^S�s�bw��,�MGF���[������ಕ<e���=jTJ����[/Z=J��*|�Ǿ�6�ř�l�~��2�i�t4���q�z�a��@ }��oBf��LWe�ҟQ4(y�O������?RG�/D�:�_듏����*Y�Y*�~�=\���� -h1rP=ĵҦR�Ԑ��sxdf���_���_/��w:Riu� �w�G/�����hP9vvΟ�6G$�,�y�Z~��0�O2i��6GU����܄	������<E��V;�{����I��~;x�'�I9<�	q@L[��lt��+U[J$�O;U��^h�NĈ%"�t�����3h�Xp�w�q�y�%�6��t���w�
�~,Z��&�a����]p �21���f�TE0����;�|�EG��ɵq�Q�BM�ᠬT��ޫFG��c.���` 3G�ʧ�� ��ܢ�,C�y�!�7En�	ؗ��P%0��Rf���Mh8��Z��cޖ&����9)�6u¯������򹲟������;Ef�VN��e�=@oKq蚎�n`I0-'Y���*�sɪ�uapyl^�3+gw���F�؏و&[�pG�g@uF�����O��*�E���F�i��wo��4�i��Z�w�&��/��`G<7�\6W�TR9��%!���>�!C�6�xF�D���o��n��rS�+�F�$��e�Y��J�Pu�yn��(`�KrbC�&P�ãD� ����G���M���_�b�ߢ�
���^"a��p�vr�m���(��*9E�?а>�L�ϡ�V�n� ۾�ah0L
��*�ɣ��Q�u$( S�%Z?BEr
e��c&�3P�-��󵏞q�W�(�c�Mɑ��屶�Q�l#���B !/#�_�pb����4h�j�� ��;9׽���Eo�hw�J�qF޶��^u�qO�]����BbrkN��پ�R�S3��2IN�dB5��~_���!���,ل���ĕF=4�P�DßZ�be�ކ�H�ee��l�7�2 �E��UL�3���n�pȁ]Q-`np⦈q���"���r�?zEiԃ��h`b�13�u;(�?���,�bNv�z>��0��IF���G�7��I<�Yd�S�w��ya��y�*_D��1���XfYf�1B䕌��́��'�)��Z\	g�iA���Q�bT걇�n��0�T������;�Q��'Ȯhn
G@�h�#�@��A��c��ovto|R�0_�m螀���5A�H��o��|�UH\` f@�_�^:�E"�ͱ�[  ��2v']��p3���]� J��G�i����۞O�>>��$4��3�xai,R:���J������\Z�;oy�\#10I5�R��Vu;ԋ��u��]��k#>�������������e*f����%���'�e�}k�n�bh�D�\�0���=QD���Y D�Ñ�w�v��W j�{;�!R��Vp��u�C�}�ҞA<@ �����I�z�V�=^&�&k�Ү(sݻ���"a��������j~���T��)�ڐ�aA�)�s͈���?�,YQ��pWd��z�S�V*���t*>�Jd�Ӳ��Y��}�k
�}K?�4���:��
���uN���a4F���m�Ttwn��������^�Q�P%���R�lEP�>�b0�c�$�������n"��W�ۥC�/h�g���Io׺/�G�6�7`N,e�M��K���`*���7�X��AHP�<�,��ہ����M���$g������6}Hː��!|C� �VɃ	�4[�t[X�����ϋ3��s,��셲1����D����%��P5f�>M�R���.��E0��ft�G����M��?V�������*GU�Yf�*����=v>��W���e7����l/�_�)'���; w���"c�t�8e^��)4��,삂�[��c��_����A{
Z�I��f�N�P��L� � 9=�KR��
+��v�l��0T7��8^踩{q�~{�<�v�c*=ݟB�RTL� �H5 ��4�v8�ɝ�j��p�f���A���z��QK��C�� �����*ve`�������ˡ�8��]�g��hV��E{����CY�p��\O��kZ����%�a$��1���������^�'?�X�B���ުhExP�aE�@�v�Z�)����7�5�!���W�"�p�V|��c�"w�����nU��ғL.�)�-�F)#�wz�Aw5 ��QA1<c
�ÈAQ��Z��g���򜦽���`I�R��YH\z�uʐp�xo�T�\NCM���U"�ʢ�%[:��oX���f'�b���go�+ڢm��n�4vc7��ƶ��I�Nc['hl��>9щ�r߻������{r���q���TB�,��W�0Cw����d{�)`�3��6�#k�F^]_3��R������T�#_��������N��[*�H�H\KDצ��/a����-qR*���9����ԉ
t�^��S <_�uF�y�=�u;p��C����c��i{x�N�2����6$��D��H�ջ��yPR�������w�WJ����ʍ-Ψ�ԻI��*>�'َ�/���](8���ߡ���[���D��P�X�ɲ�g�Y��]��t�W"G�Q�>�2a��>�k���ϭѮ�]ӿ��$���P�{�R]Q�A���n�#�}��^j1�R軯��a�Lam�bƲ�a���.�|�'X�ق(Ep"�a$��~��G[��g��w���c�NM�R�����B?X�`���: `����-��Jl+�Z'���H�97�uȥw�d�4t4E��1%:�F!�#Q�&z�����F4n�店4^���]�����i
&;��w��W##��B� Om^�M�
gM���`m,9��������� �� ��[P+�"�|�#�7�3kG�VD߄�M�޽o��vG�1�ʃ�9�{"�^�_|�)�g���Y���m���7��:� �I��?@]�
ԏ����T:|u:�TS������R��lQ�o����OH���v5
��T���kK�`��������K��j%�T���\S�r��Q��'ƫ��'H'�0q�J�_h6�Ve\qp�Ig���r=��Y�.���H������Yk�t�����F���bZ}-xf���0�U���*+�2_&R(��Zpd�pF�UKy,�����J�m��ת�i���X��b�Z�ߦ����~҈�EI�EG���יFlc��*���^4A�#z�j��tn6����ϐ�����&w�?�w�����+GR�F͟��O�76amD��U�7�S��YQ�gM����[�Q�k�Ϊ�׻�x-3,���Jg��rM<`����ᓪ��]���<Z�O���R�O/�mǋ�'�F�9�8_ٺ�n�m�t~ܼa�CM���q�ڟM���c2K�8ѳF?:?���5O�_������!�������W"�u��J�;�+��Y��v����rL�q����{oi��؂���N�s������ub!�"@:�UW���o|�G���C9���Rf��[��?�.'�eA�_���&���wEPa塋���]�PCm|�R�nOԯ,�VO S��/�.t�f`�?�1�7��P�DY�dz�$�:_�,��p���~G�o�e����:c��^	/�ö�������'���و��Ozp����Խ�!	`��l��:n�(�?�Kd�H���&�=��G���p��

�/34���_�i�h�����<�|l�^�r�+W��m3)gIH�TW��f�tD��,6�D�xۊ��gNS���bU��M�Y�������qWD�/jY��c�%(��BiH�cz\�I�;A�_6dL�o�Ƥh�4��p�|��j썀K`Ǫ�.C�	]zHiD۷l�gc	���̉�;�2i������o�ے��8��:�����"�v�8^8��v93�6�A*BuF�h�5ڒ�	0/����/,��V���g�� �U�B�+2�P�LX墥pa�2��)�̢U�7�� ���%&�_a^U��!�g�A;�Baִ�١(Ez|�5!��GN�ͬC*j��["��5:�i�c�=�J�e�]�X��"-�ϛ~#�)WVH��ڊK��H���� �݇ ��71A�}rRAgiI�[��,�.	E��w �T����*���L)����7���9��A��'v�O����ѧR��BS��>�:���@=�!ve�5^�2���SƚC���-�7�m��T�t�+h���A��U4�B"͂�r�Q����<:}=� A�H�������SR�����Wd·Z�<�K8/4F�'�>��"!�������$*ݣ��ز��������,��p��5�;���������~�,"\s�~� b�c��P0�$�+��ܬ>���؎�f��E�E=A�I�x�2r�?��.�������ZP������,�Bxi�짯M�BA�o�0��2ȁ$�k��� Vb�Fɋ-W�#�¶@��S���?�B[
u����UU+��~!�%Z(�	����
]5�zڂ�U�@;F�Q��9���&���U��b�v����&im���6]��r�a{�
��:�*R͝���9m)&m���"աo��Z���Ԭ{�:����$)�CA�	� R�J����9h��;������*`�'�4Uw�dV�b�@���C[�a�9�7`d?�1���0[��}1t��X��k"_�U�M]
�$Q�F�3���:It������d�28mK0����u��d���VcVJ�K������k��[��~�H��'l��Rl�����BF�H.b�J�V�����n��wH:s)W-��c%���V%�ma�*�;5@�$���yEI�k�|��(B��|�mUȤ:~7*���<؝��!�� ��_��::Q$�>di�;1,=}���W��	?��C׍_qN�s��P�L����	-���2��`n�W����)�\�=���!��_H�~�ȥ�<^��#S�8`����G�n?��%?c�����f�@�͘�o�'oɪ��i�v�n�[���)uw�����0�й9�z�t/3|��ى���ٽ��!M%o��r2��g�����:�53`F�o����*uiO��_9p��@�o{l6����p(OD:pJ��<�7Y[?��v�hL�v�[��l�#��gF�k��249�ƃ��z��
����@�I�@�֝�AԤ�_��~� ���?�%��H��V�p�����/8p��1lM�c�H��1�̴� ���>^v�v�lk���=o�g�[�ƙU�g@��!q;խ�qܛ���]7S!�:.�{�F	�|�UF�����S�����W}г�����*��ᑮS�R�2
a���GS^'%i�w�5w����[�tԡ�B��f�����o��
�%�@EBa�U�X�b��}��Ͻ���h[P�F˶�0�E]c��-(�vgo�B�M�㶆(�~��g��E�n�����(���4待��붽M��7J)eq)���l���z�-80��AF�^sP��;J�!�s��h���� ,��waD�������GBvJ�֨�V������ao$I��ܴ��ޞ���P']��	� ��n��Ǡp��kj��)	~����~�(@OO��!\���@�*���H�����Q�B����;+E:�l�����wo��y�ԣ19��{�FX��f�a����X�r���.WiGbAA|�8��E|{���MZ����C��!�)��Ԩ2KV��y�����Q2E�6䓜E��7���n�ݷ�;�I���;n
�Ǔ�z�qz
��z�H{e\�n��|�9���7O�+��8���/I7璌'Z7=&>ezy��1�3!��}I�����ܦ�g��7�6F3��ȱ�$s7�GS�����PB悄笠�_��F�&n��&F����1�3���r��C<��l�چ�1�7qDD��[�[`�z�t��B��WQ4�eo�G)�w(
>��ĂR;��}9mL�mʒ	3l��h9|��G�^q�(U���]!q{� y����l�Ċ?d�����Z�� S	�3�����	4�����MZ���z�� ��r
�1n�7���j��F�J�Mu�w�$���76��!칀��(��[Ȍ匶X*�Ķ��N����I{�r���*��+�L&GO懎m	m�X�	甯\f��Gqìf���	�nd�������9�F��"�q$p\��y��s-}�fm0s��Ҍ���[)���nO�l�G����j��fp/�����		��!i���`U�f1��¢�VN+�v���6��n�˞g����.;��b�^:���Y91�3�ܙ��'Q���C���a��W���D��_Բ@�� ��j$�\�lo���$9Ů���Y���I�i��PQ5	z��,�����2���e��&�ʝ1����R7(��������7i��1�B�p!o��� jE�H��3K�r�����ړw���= Ki{��7��q}�ypq�����z�)�hX�UG�ɩVt[�Yk-��ҚZe��^�7��x3�!j�� �΢���Z�Lt�����[KL�b�ƕY3P�����nyܩ�)j^v9/���Z!X���5	t����뾶�����H����$���u���BXQ�yi9���F xъ�x�|����}ݾCQlvU;'�'�R�͈/ג�_�M�5fȦ�0Z�\_K� ��^�r7�g� �ٛJ�{��J�g��V���ragl��k�&��@Q���F������Ǵ1�v�*��"��ٺɨ�VsF����ߝ�>�����h��jz/1��*z{K�TNQ4�_QLj�Mݪ��2���W�:T%\��b�|#�0�R(x[����=^~1Ձ��i���� a��sy�]����]�٥CZ�2/�Ƶ?#V���ø��5 ��;1EIbG�I�--�g䣞� �)=��d-Zi�۩�A�{s��t�l���#�=�6��\���ZE��DY�b��Ә�~���
��IY�n�Qn��L����6���]b~ٍN ��w�3����pB!�
-�����+~��F��\�Ao��%��*+��љ���(�9�*ʽ)+d��U�Y��L�l�	;ߒ#�z�x��.��g�'��6-K#�Ud?�|D�M��c��n�����KipFw���-)�a�'�+�%�f���ڍT� O+2C^r�ƽW��=���5��u�6^�hS���?�z���o��ҹ��G}�
����J�NP���NB�U�.ӯ���~?�?YL�|=P�ll�IE�i�hc��nU�+y�T>�����?7�F~Yu?[Z�� f��N�
>�j
?���)¹��ؽ6ρMe%['/��CS��J8������Y��݇�-�r��3h���pr��[s�+��}�8n���@cR*h:�:#yB`�d�}w��RI������7Qmm��#�Mh<�9��� �yF��]q�8�Io���# #���dÒ3-2��Kʺ7��Ɓ;�7���0�i�w$"
���O)��	r��O��g����F�ˍ�&��5I��q�@�]�TsU�=z"PTR���[?�ki1>�h�e�}��0���]���6B�='�2t��*���z{���@�һ]0u�?$��@���&_��ggy����X�2���wR� u��63�HA�A&�gQ����gF֨�N�o�M��'�
����$������Y��W~�Lv�IK��a��$J<�_�h;�ow?=H8�2Yu�qcVz8���dX�vcx��2o���[fE^��O���J"]����ha���k�����[܈d%�^�v�|3a�H�i��R��P�P�;�)�����<�;���r�Y������s޸o<�#��)
��EVh�x<}��^�I���.������2#������3
S�4�d���в����7ME7���i!=�F��e���V*gF�z��?ʙ�un����ڍ�uwb��=��=C��*߇>������}��u��ݿ��E�}��ۃ)����}��q��I�Y���Ƽ����yoߊre��K�Ͱ�Z��-Q�=xg[^g��?������k�Z����g��8	(�5�e[�J�����<aV���a�q��;q׺Ք��
}�����9h�-�����wGV�d� �x���h�0YN�6��:� ��>-�� �)@uh��QQIK�ݗ:ҋɷ�2�����9��R]HGu���E�ފi���3#S��{&�
����`%�1�vQ5��|���/���e��X�Ԛ� O)�bLY>�*��Z��΁������Cq�� L�?�gR��5-���p��ZC����}P���SV9��/l&���ę����� �{٤�Y[�~0 ���7n҅$��>�)X`�ě��D���y��k�ݒ��8S���w����m��e;�=�QX�0���e�GT�2<&�/����ܸ%��+X����!U��3��t��ES�a(���vK�QK�	����FO�:�!ΜΔ�`�/`�����ǫ�3 <����G �K�;����BIM_y�ؙ�5�sn����s�ēt�Cߜcls��6���H��|��z�\Kr,�Do�B6}�Dd������q��S��He9kb-�S<{�ޤ�4���z��K+��	ʼ�H��c���o��H����H!l����iYϞ��I�$+�c�3-�����l���0��1d>����C�N籀�J����%����孖@q4�r7~v��b	14���)����	�����έj�j���ꐢ>��J~ȡo^����`d����'��Q!�t-���������Kvk�<9���z|�!M:�Dt��|�S�gv��s�6�\�u�}���V��&��dq��Az4>��Ӡ���f/+��Ok���䑪l��s`q�)�z&G\ C����t`���!�P�۟��Dx���_��r��nJf,��o]H�&"s�e����`��f�kd���s���Uj�(��Z��ߕ��q�ԟC��D��#�Dъ�Q��	[����M�j{��Ћ�����=3��D�����^4uE'�G����a��As���R6#J¯M�nv�fY%���<
�CIBr����MM�%o�^�*�g�j^��@%�$���=s���(̏�����ҫ���$�ͳ�N�:F�R�@/���X*���}?`̪�d�#ޭCS�YB�+��r�Q���(jN�x��E�&?듼N��.�i���U�%~c(n�~�֓��Z��-�q�xm�VN��jb%��D]WZ�_�%��D5`J�)��l�b|"�p�a�k4uS�$c�0�BY]�/k�n
�O-n�?�kkM�HaS �9j��6Ӭ�n��hT�COb(mk�.�s
Q"!j#��D����P�k��Ma�Su��<�U\�3 I8p�3�����1������ԉ�EK�Ê�!,�.q�؊��x&�k��������O�ꨬ�.u-m���}�{a�M>>c#��+#,5XӅ_�RC��^!DB��w��H�6+QŬ��0RU�����B�b��V[��UޙOJP�t%m����+j����݋��c���~�>�D,/�2o��rfƖa���$LN���⇺���A0@H�i1�M'��d�CD���;�Y��}qa�E5 ,5�ܺF:�'���1���M@�"i���i�UN<3�ښ�`KQ�Q��ܭϧG,f��}H����ըc3��8ѐ�n ���сH?�e��I)��8�d(+�5,��ː;��K�Se�Ma�鮤���"+�F/�*�������S��KA�n}!���͆��rP�/r������0��|�g�aH��資(��;��g��}Wbp�����Q�5�>:��:64�#��Ӵg�;e��T_9_N�W}��&l��˔�����2�5�1邥���?��Rsje|��X�Yǒ���x�ʉ��>��:^ˏ$i;K��Z1�b���c���(���Ed�~,�u?$M�8J6!sgj�א�w����D0$�f:.A��g�-��_K�􏵠�R!GbH���Y��:Ӄ����
�f�a*-U���\�����P�}bd���.�K�=�.������|��PV�N'��3Uq=}hiՐ;���Nt�]ծ���|.�G����i� �i``��׶#!�N����0C���fYs�g�V�B7���Ê��"�h�����n��->.t�)Do�����o�4P�-�-��r�.����t5*P��X���c�T�,ؓ6I���X�����Y�,F�jr�Ҙ�*���yh�ʁ���^8�?N����P��յ�lKUX?=`�б�l/��`z��u0!����Y�۔�x���-6S������%&���y�P+?ڂ}���(q�+�-(�K��y�`s֙!f|1v5��/U0%�tV����J 1�W}M��.�����|@�"T�@�	�sf���e4��lc�Wɪ�Z���B4���zMa]�1�'Pd�n@�?�9�P�i�@�5�Az$^�;�/3V�-�V|H`8�RF�Gs��)3[���S!�����oľ~��0������t״IeA�s3�+{R��K���4�N��|\ϗ���6�� ��%dU<_��7� y;����0n�}��7���,I��
M/ߠ)5Ɓ=W�M�k����4�DQ������$�a-�R�����%i�7r���=���3UZ��>����-b�$��o%I��7�k�	��l��7�㋟}3a�5�h��.^�1!u$���EV�<�뙘�հ'�.��D$��㌙�]~n��M�4��=����v���[�Z���<�Nʓ��qe��ݻ�M��=��nw9X���D����<θ���au)��/&��6�$��a8gE�5��H��������ȕ�ҽ��#��EWQP�	�W�t{���)r��ex;�q�\�N��9���1�<���*a��B�w�I�����QC�,�]�>>z���$�.�a�=w��� #�����{b���S�5a\��:oqK�����'�un��;lu��s��,����%�GTԊx����]:D{;h)=�]1��8|��d׼���v�W�PȜq���͕bkO���.�9��Sk�'�����-����LK�	R՟�|�˭+")��Dj���4��06��È9m�'�I-aiv}.�����y⣞U��/�y��~��,�n��;4����bF��~��{:lPU�e+�������4��T Ё��0eUIc���J���:��:������9r���$ ������S\�[��]	�#;�)F����O�18D;<��^�#�5�]ŝBxE0�b��x��!$�5̟ ��CS����҉�d�1�/���{��Ǚ\m�K�ռ����0*ʬ������~�!'uvV:�L��(��e\�f�Ԡ޽嗚,w��ڏ���d��':qV��E���r�)!'F�eO���9�B�տ�i{�_�dH����tx��i�X�}�&h�,�9�yM����P�%+���x���Q��#����Կ�G&�ݎG�*}���]�,kώ7����w.���A�	M�7�����;��#���ԓh~̿���Gv�par�/ ���.�&�v�cv�����|uƃpL��
��r���t��H}��'q$$�..Gn�@܎�
�,�j����⚑��Rq�ա���xp���(!�ch��U>�8��!�Fu{�=��%�J�u��Q��u��~�I��L;�Ȳ�t$����b�N֐$��nW�_#J��(��t'�ġHt�_�w�Z;M󊃰���* �J�#��#z	9��39��i?Z�~�7����κ�8ϓ��E$e�g�_�-n2O��ir"�Й>�d���I�}����{e���h�ʸ#��!<�<���.���Ɛe�H"��+ۃ��QP�����I~���m&�pLm��i L�aF�
q�E��5��zx�}���E���+�_�3�?��w����(uM�$�쿯��v͹�]��({��&G��̬��U������:����.g��g%��.-u�mM��^Ъ�|?� *�:��R.w�]�cc��v�	_�C@��  ^c���A>��|ud1:d��ߎ�V��ztzt�ﵙ!h��7!�}%��'�����K�g�v�vv�:d2�`�j)����Gwt�L�Si���՝�פ��f�i�ͭ��o��q۹�a���ۿ�e��RY�f�Ñwe��G̀�����*�ֲ�u��8����g`i�`V�0}<��h���<�Dާ�"�*ن�\��oS===䎿���Ì^vq�\6�$3Y,�S������X�ޤ���$M6�~�]��0$�Bq�U���pq�%�y3_V;�쉬��8�`��i���Ym�F�r����˓X�C^�-�PW9֊,V��֭�'>gh���GRy�jaH���)ʴE w�Hl��Dx'�G�FόZ$�j���h��6�"�4"�i��?j�0&*!|�X�P�`N2�EZ?� :�[L��7'��M봪5#���6&*ϙ\�12�%'$C���12]���ek�������#��;L�h?��Ǝڧ�,�K��ܢ��Y���J�O�O>S��^�&D��=���J�D��z����x��l��usCW��`$ݕn��0̮�V�E�ו"���Pj����]�,���{&A/�[ϛ����ݾX������o���%�s�%�6���b�TL,jU�_����X{����8o��k�i�$u���X��)T}Y.�楒�&���T�F�F]l�BRFb�V��?�V�e�c�c��T0rx7��r\��}%mR����B�E0^Mͻ$���p�����䑘�U���,�k���!{^��&��`(ʮ�PѮ�m7��s��ws�9
>ҁ��B�]1�"��g���\�e.8��с��\���b4ȇ��ETζ8�xF=�ݟ��Oe�#I
����.S��=�s�џ��l���ɶ���N�X1YbN�3w"��ּ�n���������ޑ�����Y?_��l�v��������blWӈt]�z�v8L�Q<���f��pI����"'��c�y��Y�E�1f`4��O�ޭhHfJ�fjE+��{��W����B�AK^�RƷ�{_wVA�,���Qz��l�#^�G���A|G�A���o ����	ӂ���'�ܭ�i�?��H�t��^���yv��s��k <�	m(��|A�ІEj�-�6�����4�{��%-&����}��j�פ�Nܾ0A�*jq��D��P�:�L��q�(��|yK��a����uw�6��г��j���ܫ�(^�/���З��z�A�d������+İ��AD緷���wB���8���E[8j����=�7�%�9zo�����G��A\^�S����%�]_v���/5/4���4�Eϫ�"�g|�l�[ k@v�Y��(��o���M���T��D�����Qrs�+y�t��U��ہ�lHH�vo���]���~qp]s]I�.V�I59���|!A�J����pd᧨9^a�L��&��������:ǝٞ�A��JD& ��/'�H`�5�٠
=TT�u��s�xx|�wÝ#NiKc��}���'�.�ͳ0/>��{���Y���wե���0ssc�{�漙#3���V����b�9��Q���]e`d��%�2���u�gq�n��M���1�<�Tq���O�z��M�f=�z?��mE�x�g84�Hnč��$7/v|��|�6z�Kk�}Ox@�8��)�F�Mbyl���P��و� ���+��%m�J��}	s�P3�\�d?�J�Id��z��|��g=1�A-6|-׶����C{�S>˩���h�U�&���S� ����a�J��ݝ��	�d��J��x�����8)F�K�H��#�u��u����)._��r�X��ƫ�(�k�Z�9��+N��4�x��xX��O��	t;I=��X�7Ub���3�����?�ޯZ�V����a���p>g5��*ؿ:
E�1z�r���t��}��7��T=r>��o7J���/Z�P1;x~�j*�1�.�{[2T!͸� U�V��Yҗ��7X`�5�Y]�n�~�2�.0FȈ��Ld^\�:`����-e�f|���2�r�У�7�^�8zA+
��"l�)FkG[<��՝r؈� &�>w8�'���N�&I�\�'�"N����w����a�/g֤��	V����߄����:K[1�X�O䚛T���fe�5&>����@+#Bᯐ-R�<���a������l�<��¹�b��0�,�ӱ�)�!nҥB6>3�{:S@�Ka��b�R?�Vۋ�ન�P�%ъJ�N�Ba��ܑ�`0RS�d�W�^��m��/�ӕ���6�0�N ,�]��UXz1�D��6V῜d��I���Z|�l���o!���r��{�r����9��O��]Lu9�#M�Ia�|}��:��vVpI_-?���7À��dGɖ�8�%g�}O����Yn�v�PՅ�?�\Q���vr@~4�|�dD^�A�ݍ���Kbf�kצ�7���k�+�ǻ��{��a>8]�ވ ��ѯ�xf��^��%%�HΈ2�JyіNi�ރ��r�[`<C��6����չ�WAfq����`brN/c��W�Oh�;�!��Ǜٱ��.p�#�6ப��_'��f����tg���|�>e��e����l�Ua�?v�����&ݬk��j��,��Пl��!����s���k�_J|15 �X	����'�g�q��Q�ٝ�3
�cp���W�̳�M��,�;ϛ�����Ղ�i��&8�1Ǭ�w�6��r}�D~J�Y<,C^�V(�\�B(���C�����	2גkO�9�\�Z�=1�<3��S��݈�q���5�q�VK�i�66[�[�ـR_���y.�X���������$��R�?�yz�z7\6�5�eJ7x� p����>Q�:�fM�2lw��E��#h���.��������a�3;��S�R��O���I��}�Y�d��@L���F���*�+���G���?`��������pCz��zO�|&�F�x�9�����~]��nx�C6"4s�YB�v:q�������+�<CER����m����ƳV[:u��{�Uǝ�'r���'���C�:Oqn�R�Pn�hS�e*�L�(��W�c0hΔ�@��\�;4��A�m�y}�W(�I�X?��wS�
��b��:�AZQ=<g��e=�i��Z8t���f��G:����a��2#�S��`2�� Gku�n�I�9��P�>~0	����:3��Pp�D3��~�2b.n�4%������뙑T��[��B�2�/n2^��5�1��]n�O�����]�������e���=a�"��d�\d�~��^ ���+]�'��gnJ#���+�gg��	�6�&
(I�	j
��¯��]Ugk����U��hD�m*�!�D.aٙm�NG[y�z�!X�_H����������oh��7kf��־S  ��ul{��X�b��F~Š��y
(Rc�`�7c�	���LGk�����]^�&�]Ϳx6���$<F{��l�crynE�;u���G_/ӌR03��Ǭ>�ށ�|���j�;���<�y�ng�[=3������y��bz������:5�1�g����['�H�+3@q��G���u�s�4�)��(��P��}�E�m,&/��ы4�[�t�f�pa��Eh��rOǹh0�vhg�{7��"]M���@V��ϕ�ܓQ����VѦIƒHloa-Q����7L�g�rr�q_=`{�-�P��;��iǹ�z��ݖ���C]v�����`h�&���j*����]�'Y�Z��f���.�V����t����)b\�ǚ��s��ݐ�'g�W�b8� V�i,lY+�fxi���S�o��m�K�_*��fv$�Q�,�%F��Z����6��&:]K\yz����|\�Go,kޭ��~��%ˠ���ٲ��*֚[�WϖQ�Dihr��BqeLѝ�Ϳ�)�zv�yu��t�=V�#
4x)��l��(���
Z�nB�.��X0�/ :Q���[;GH|���F&�/{���p���-�M��.>f.�.�^|/���ۂq�+��xr�RQ�ߡ�Ճ�$Vb=۴�s	;����S:-$&p���|��Q�H,]W�혱�Q�l�Mq<���#~���x� ����U�ɇčpoF�0��%0`����)�ʙr�y��Mc�t���#����xe��z>ƈ׮�����{�>An{�j2�Ӿ�䝗�@�&K	g��"�'�?�E*H���l��wx��J:<-v��Taa�CgN��[�[k))Q�&1	t��|'�^^��W�&Ȥ�X�IGxh~z�\���F���F"b��aZM��o����(fOg�Gj�GH��rj�D[�A�5���V�'ɱ�Iǀƚ{Q�ؔ<�Xr���u���T���%ܪ#k����C?��Hx&��Ṩp�F=k��v�pD2��� 0�����Ϫ��!��)W���%޽5�T$�Y��#d{���^��`~��&@�LÇ��9��4�	Xy�^���u^�Ѽ��~�#��N@�s��L���O ����ӊ���j"�TO5��E�c���/\%m���,x��7%8s*J���r�z�B�y�����t��M��L�݈M�}�%nu&v�,��q\b�1�p<|��<�`��>��5�n�M}<��}d\9ر|��0ii���^ӝ��P��tn_!���KS�
���{\/�Z}��e':��4	Ȃۍ��S܋�0#�b^&������C�ݦ�����8�z%x�M[�2N�D��� ��6±���%�r����|����LPu	-�]/|������H�s�&�m��H �T���Ű��C���n^�J����T����g�J<���s�)`�jR4�fY~Ci��
$�o����\�i
 �/�--\���[��䶡�cS��ڦ)S��{|]��K��yplf�ْA���zҴ����q_�1MRI�j�|{�Ұ�����/�H�V���-?�&��h��XC��(;yڪ� � �͆W���9٬{-����C�0���؝��9���l"Mj������F(��� �1n&��^�Zn���R���~�ȬC�W\���<fG����xO�KUC�đ*Gl�b�#yu.O*��5=�����Nj�Q���i/䮭ֿ���u&#�Z��n���b�'Z��M��턦(�u.�X��e��_o�!�b�wߘ������՘D�(kT���e�
� �n4��TL�_=?Xe)"x���S�wQ�w24�ּRF�x���% ��ena0¿�V�<�;Q���'���v�!��r�?Vj4;���;�,�w>#��(С<r;�'T�KVO_rз&��A�P9W��lW7RAy@���q,�<�A��m�#C�+�Mz����qDԯ�X�̰�cB��uZ��[䣷o<�;���#N�.��凨5�}*��M����H��"%8�%4V�B��S��ϯ�n/1���qD�Q��b�T�-^~�\yD��&;lpb��@��;cQJ��aN��bU/U3gU���ry�}s�"����	m��KG������﫹k�ܛ^E8��$~h����~�!k/��������kom�9�.GɸINp�-����6�7�$>����-��"K`�#( ��<f	|D������g��\/(v�-�acZ��_1�/Y5����Ǌ 񱒣f�f\����9��i'�[��i~��xu�i��;�x��r���ն+� ��n80��':�#�6��7'�� �4W�Gfc�59sdu[$��),ԗ�4f�����"���<)����aTC~=E-�}O(����Ѝ5.
�����8�z�*�aJX<�s��2�1��$#i�D.M�~Ka��eV�t1!BO�nL�g��<�h�o\j�t`�d�' 7m�,o�V7}�����_f��/�(�й��@ aQ���S���i�3�k�D���,ʅ�������7�Em�1���z��O�𻱉����/���]7���;`%>/�ɚ#�����P�<	��^��CH�~�T"�#u��{O{�7�JQ ,��u���m?p߯�=]Y��ً���q`?/�ub�"j��<��C>C� 9�vl�`#j�r�ȍ����KR�Txk��z�E5.ƭ��)F�V���T�	X��N��/��iW��6<��Cy��p̝�8��_��v~�*��0����o���Q~���`��x��\���Ovm�}��9�.���*v�ɦ�{�%�@29m���"]�s:��R�J��j�¶���&����������5i�j�9�D��Ic�u�������a��p9ic�� ?���w��G�p炊G�L����2wD��F�AO�UQ������� 1W����!�:[�J�x8/��Y��y����	�]z�%��5&P�ƚB�n�8_�5[aK9�nSY(�&ݤ�!WI���8�����Q7����I�@��+��8�M����H�~�����ʸ���m��N�a E��C�kh�n����k�B���_�������4��{����>V�"�f������ewja-W��e=呇+թju�٥WQ���"x�*_�p�}%T.���m�xM�L`�S2�AP���T�HYF��+�r��W.�N�����VU�������I�����׫�p!��s-쇆-�D�Q�`���e�{u���a��~��5vNۃH�T�� ��+ɆeA|\���� iW-���.L���+�?0�΋����τq�!0Z���(ێ��_��}��Ą�.��>�H?�G��?��\�?�H�Tp�o.��ݨ���^�'��-�����3&E����:2���6����1��Q���?�nS�N{�C>0fX0�P��`I�P�����698]��ji�Y�G�jÐ��?���ق#I�\3��I�����م��@�� �Ǝ�w���<(�r;��MF��/2�PF W�kq����9��ɘj��s#�7��'.Y�:a��/�:������3d�r�x۰嘺���c�| :��V�h"�*�ZhQch����/�*�(��~�Y��'�~����]h�ڹ�z5n_��������k�IIރ@٣Sׄ�������=j�D�U���^��ǌ]ol���{��E�_�ܯ����������@����k=�CH��k&�%X[Ӧ~$�-��`�G�Q����n	�\�]o)��S�\d��O�4ҫf��I�0��i¬P���f?������ :�v��Y�⡷>�ڸڨ��b���$�91�c/�+lI 9������;�4�86Xs��#v&/�C�B�1��׬#	͞�i��s�rbk��W�'�5@��[֤�}k��C�����΋^M#r�c���}.��D��;U:^� ���3�]I��-��f�m��^���/��3Ó�M�d�ܟ��޲Q�f���^b�!�q����{}A��� �������Cϥ['��PV_$b�����g+�3iw?�G;&��!!"���^� �iv���r��N����gK�/��җ�˻��|���޻���(�*U6q�󉚜��3VXs��@	$Gt$�K�6�H�#��iذ�б�e�>؝\c�9��G��bh�!�1&������$�+�d��ZU_
/���@O7��d�&�n(1|�{ëRP~�>�ӳ�afJ�C�t��:<FtF}��+�7����np^�yV�o����:IF�`���gk��N��6%���a�磩8���q���`�`_;��S
qUI^oc��?��l|����	Iw���{.?���f��M��N�~�`��2<d��ɶ��0�B�se�^ɹKPW����B��z9�v�o���b�C�ow��;��Q
y5�v[�(yx~b���`p��ZQ���!��Ev)����7Ϥ�{I,��Ovd�$�z���2 2]Ƴ��l�/~Z�ȝ���?��]�c�O*�כ�&ŐG��*���Y�9)����-j���|m;�.d}��`��r��]j�i����n����atN��E��oPo�'��X��jUhf��,*x��������
xʅ�P�z���t�y�VQ[���	�|�Y�J���\�ѓ���Y����MW�t$��o�X��{]t�)!0�����}��-���48Y����۬Y2f�9 ����Zet�ǸYܶ����ɞ1���0�tX�p�uO.��^-�).
��ؘwE���I�G>�^䝩IY��.wjE�zO���i�[�)r�V[>n�s�C���p3|e$��=n�*����#E	��l���NluY�n��å����ERYʙ���������1� ��do�]8�rWH:�i{�̶���[���@7�?Cć�p?D��}U�K|wCbQC�)�2��R^��`u�d�����u�D�J6��w�	�;��=��B�tw�t@��_}�奏�%��}�����������[�)6}� "p��`���J����8ꥴ��J���.4�0j�g��mA�=�r�->�:��Ӌ�������_=Q*�w�\A������G%���$=�'�mzu�ݕ��J�g�50�+�p]\�����м㰰��N��;��Y�Ë��t�˨��\���ڎ�"�1ٯ8��x�0]���	�t���t�3������xkF�(K'��9OI����ըß����2�ۯ�qɝ�J�١yF?��	�Ȱ�l�[��<�����7k���P-�;�8ITxZCL?-�p�M�ےT���/���Y�%��>FNt�ɤA7��d>CҊ���П����Z�"��?X�ٛ�r�ȖN��/@4�q:�탦�֙CS�C>����|���%���9��G�q�{KV�f�if�f�Z���Z����ehɊH�ʸ�މ�z����}[F���_��S~�@��ļџ=���	"���Ԙ+1���;?"�����:ΰ��n��f��
	�{0�5�.P�����6ٯKx_��}���Ȱ/(�d�mNe����Q3x��n�dc d���mqlu�¨l���R5r�C�I�~p����%�-ב�U��.�{d�Q�g�ݶu/�f(���~[S��2B��Vi˥�����҉#�/\�w�X�O�:���D�ѵ�ea@Ҿ�II�1(�c:���VY�Bpkm~(v_ߗ6���%����#��u3f�+�c�>�t-dZ@>}��2��E��k�(��T5C�(��j��F�A��5 ����U���BV�.�����x���Wn;�Cϥ;��O���w�}u���_	8��`'
�ى��DX�N�$:���i��@�+%	LdOӦ'��0D�,f>����9{�~'�:�w�O��_��RBA2TYdO���L�����6i>;B~��J���	È/~�$jS�"�k�H�M�9�
.������!�
���9@�"�V�lǼ��7����>M��Mj_xb-�^����1>�׿����W����=[����4�&�UҚ�畦�F|�$�������)��c�7��C�U�E�^���I$iPn>}�{ے}��z@<�u�A���q��)
!�=��M���7$)�O�sw�Ň�ࢺS�Y�Ƚ�o�K��9�~��
�:zn�L��B��-�<�v�sf��okktcS���ĥz+���Cֶ͜[�PXu�UF�i2rOYUš����%ո?L�f���Ŧ�jx�o�[ۚ��������hv<.O5a?>�[`�Ω�!�]x���?�֍� O"ZUWGlkk۸���n��jV�԰=�n����h[2���}ߤ�m�&�>z�ζp�v��!�C*�tLy�5�ҩ��W�DTQ��ȃ�;��:��vr���c��3 ���wcO��a6���+L
��S��׸�����B5�칵��BO���3]ݫ\%0~�-��nl��{�t9�����+���z��e➥k� ����6П��qf�Sک�����mï�Iм��}';pH����&�N�S�-h��}�!�B��AȔ��R�ǂ��~����	6^섳�Fm�2M��ducU[��f�s{���-U�ir8<��^by����u�w�D��#����=�e��5?�_
S20��v�.��T���Q~���?�t�����N��4�*`qm�a����Y{���O���z̑��\渲7^��Z����U+904F쾱fœa����vn�`[)�"��I�s�{=�4���C7��PP��U���s����h�Ŵ~�p�
�+��s͎�ަ)�>�1��0�8M�{�T]ǰfT�o�o�m�.���u����Zz��֖|i�M�?�N�`�%k�']ѭ	���c���C�����9�ա�\,��vTX�G��jeA�ƙ�F !�������}^�.�~9e�:�!�q�W�)q-�*@Y���]�����<m8���U.o�#�q}
�e���!�s�����2�R�9��?��>�o�#s�}�.��2ތ�3z���{�zJ��p���H�*����3��ڱC''�׸����%��[_@b91P�kB����ȱYX�{��[J/Rj��>]�(��lA��g�&Z,�S�'j�ĺ�z�qa������/>0��.�?w ��$��_�O���\��Hŧ�ch"��8BL=��|o%p���d(�U(�u�i��uz�|�̻��څ19��qr��wB*��0��T���S���a�f���+��� ��yM����πm��Fw����<�pq��^y����ܾ�_c@P;����.��p�o��f;�T�;��*&ϟK��Q߲�FGE�������vJ|�=�-�f?�}�T��fN��0" VV�:��k|���%�3��s9�g��V1��?�i�ΗU� ge�q`�)��ԁ�=�t���9��|h����2��'Jx΅15�g"�t�:zz���uB1�q|F%Hk.�i��[QY�Vɘ��f�5�x�����9��ǧ��2�0�HN$g�Q��y�32�z�&��y"i8��Kf^��[��U��z�id��ch&v_�AƹO��:5��ַ���X��P$��#�9⨿��G�	�\qi�4��!�Y[� g"��>�c��'��u
�W|�#%��jE��e��<-���m;E?�qN��;�@3d�L�q)��'x�n���W[s�,kxp����k���9ѥ�|&�Ȏ1�V�6K:t�d;l������Ǔ�F�p���<��9:�灞��LS����r�	�@*����޴�o����L4�[�?'���e�H��,jg��f�x;���$���&��8F���2� �j+[hW=c�:��!����ӯs�v���F#�ʧ��Ĥr5�<TM&́�0������+)Xݷ�"�y-�9��8`L��=ߣ����sy���1�55�j?�6�.	�@�q��#��_�6�Xm��n�4�������P::|�(��%'��Wt���'��Z��L���G�@~W��W�
h0�.c��?�b�7��EE��~g^Rص�ɝG� TG6/�4TzB�iEГ�nb�FU�C˶pҜ�#�'W �Ⱦ����g���1 �(�t�`a�5Z`��"J�Y)�LR�����4�x�«�F���I�\m���fU��SwI����`�x:'�.�]��O�$���`���K(te�&G�LA�^�#�s)$��u^���;��b�Yl��jh�����C��8Ơ�D�.HԶ?�>�XI�T�xuY�����������d4�����Ϸ��:+��Ы+�����Yҡ�"x���g+<�u���;�A�vGC�/�[~��3M4�$�ZO]j}��x�G
xշ��M�q�Ax�����nF�kxT��s�N�%���ڶ)��1#5��Rί�wX3�C���٠���!�F8e�Ҧ����uN����|q|�fG��E2`=����X)�b��Y{^�؃���-�Νj�9c?�颪�j�jYh[�J|�����N@f���y,=!�˳�S\� ��ű�{y�sP��_�
����e."2BX��0!:����F���u�¬o,+�\�r�
�CYfHI�_�,N�Ǧ���,�5ۗ�~B]�r,Xhr^7���Ӳ౪���j=���A��p=��7�:/�t��wz.~y���A���C#�::��9z���n��z5��ٛ�w�%M��w�C��D��g|?)�y����ƴD��3$�CO���P�7�;d�mR�^��@�F����TV)���.A�}���w�1��o�S�ŽUC+�g�v��y=�>>�R�򁦭�i�0h��>�E�j�S�7�7�4����W��̒P�Z1�>�TLı?Y��MwL��˻����n�]���*��l����'�_�f@ ./���������Y��$2����'�'�������Gt��L��;�<�%�<|��KoD��:�@���J�Q|@Ra�ct�3�!4*>��~1���6�O�����V��XP:�������ǔ"�1.4 ���@1�ϗ������'��n�TV.�e;&��7/2���#t�N���!U��.vZ��0���Yo�}Y��\|)ܒwb"Y2%��%n�,�C��B�\ݾ���W�K��f��:�"���ӛm�Y�h����(�Ѱ�2��Jyc��N���k6@�N.x�}B�Ϝ���\eCd32�H	Vh�2Ӹu6P�&ۍ��Xw]�7�T��|(U���Q6Rg葤 ���̈́�VYDU����ٽ�n�� �Ҫ�'�0iB��Pt�)*��[�=Џ�lҵh��7�gJ'����U$:X;O�$Y�}�_�S�g����~���|?Ps��UP0@�I��l�?{�v�V{�ٔ�p�,�	��tj��D�T� �I��$e��a��K��,bI0A^c�:[�a��v�j������w�V:��g�p��n0n<Ǚ�t (@������hTR�H���$���)J�K6Q!bU�Ui"�����o�U�~o]�.ȰE��èZ�v<[r���vxE�Y2�a��fk�MU�j��70�:�j�F����6p��	�n~>%�骹dp�Q�`ֶ�=W�t=�>��о�	Çd�OM֝��ʎl_���9�i(5:�c�FI�`��F#���x]��(��v�<��c��OHhE�#6�G�#�yr2 و��������8�W�Џ�8���<�w�j����Jd�>���m_~DZ�����C����2D�|Q��P_�^�c1�t2��|��C���C�� I
|�Z�@ΰ�a��B�L�`�6�x��a��rV�CE�Bd�D��
���[�SpR������%��*���(�]��I��3Wf�@ue��Y:�"��
#�)|�ۂ׭�Z�ЀB#~����ʕ�`\�&��e�-�� �l%1�E�̄�y�<hhA����ҭ�/z����x��ZT؆����7ń���n��$QA���'��4Y�p��f��QV~d��z����L�B�NԏK�+j���k�<V����gwa�鳨�	f����I�����+eL)���f��C�?�YK�j������R����g�e����)����Ğ�j�bY����E>�����9��`�-Jm�,�������m�]����+᣹�����Q�����4��?W�*�Yh���+>��뎻8�"���x	 i�����c)x�5ܘ��V�&m� _<yҴ�l�գ)���0�U���A
�F�NT0���s�|�����Kx��g2����6ĸ&]�S0O����T�j롉�;��@2�P:�^[���~����d��W\�m|Ҡ!����bki�ib����C5Ӌ��
Z@�Z�NP������o�f����0��6ϘxsR&�~����0���	��r�!YhRGZ���@1=�,�v�D�'����v$�Z�^2�a�e-HE���c��(���ϝd�+}�B{?�`�]iXO�*'+�KjVW�HZ�ձ��d�Q�q;)r�mq��y]/���Cy�7a1�V�E�:1����4c�����(�z���X��L& 8̶��z挃��U@q�]ҞoH�6��r@�\��"�i��2̢A)�G����"Zrr	���$�fO`g�j'�����B���YA 5i��y$�'��/�qQ�Brj΁ƾ���(���ʲ�W9Aގ6���)�GHrM�/4�Č�����lw����KJ+�<{�u�޼���Hه��eb`D������48N
2Dr9z�bWf9f@��e���lG�uņ��pf�	(��]LyTZ	mH'��]6�I)�m^���G�۱G�gְ}=��[%(ە�¢�;��dW�9a��.�I�i^�� �?9�ۙ��ǋW�_���q�"C�XA�9 F[�P�������f�** 
�a�7o�I"rY����K��2D=�¿�߱ͮ�޷���c�տ�G�W��r2*���S(G�^��:��av�ڋp&��=�;�,Q\�!g�+oUa�b��.wT�yb|�|ݿ*yn����B�*�Y�Rـ6��5��^��O�اb���h�.�T6A)�ץ?_��
�Z����������MW��мܹ̚(*�X���r�aE��u��5�6��n8����L2�V'c��N���|�|�y�I+B�2�P�Y�A��Rf���6��[kq�x��j��1�9r��L-p�iX�/t]Ϡ5}$}���(��♯���]�7��C��w�*
u��5Ѫ��Ap��+!<���#���r�=]�L�}��a���]��9{V���q{/0��;Q��tg�%�-�J$L��$V|^�� 7�N\�F�*ʙq���p^|��� �~�s�r�YqX|���@}�M�M`�\|E��������럩�c�_� ?�,�Ӳ����[�%�Rvj���,�^�-�p��ߴAC{w�)ݯ�Q+p<�u�G,/7�jz�1+���a_�W{z �l��i?��Wy�;�;@[:*RQ��UK�|�'+_VaS�b��N=I΢4쩼�G��j�R�Z0�1D-�ϣ�K/^�q�{�L��Q��- �H.=7:�OYD�_�gJ婢YeW�t$i!-���ijk�X���V�J�V_�� �x���hk�%A�U�� ,�9������F�ˡ��6�Ԍl�������x&4<E�hG�@A\�$g�E��Զ��9Q����||$]ޏ�wѫ�/����`_���߲�,�^�O�m7�׶�}O ;�=� c��Bx��@q��v/ݢ��(�8T=ݢq]Y]�s�$����������&|Wヾ!���)�e�^���e�D�x"mb�t�d�܇����s
��͋$8���ʏ+��G.]�U񌃧7Cƌ��d�@��Aʠ�O�)E��gnu'>w�ۏyr�
�b>Wx<봺���"
o5�"�ׁ�j�:�q�>�W�&O�ۀ��$����җ�k�	����P����uq}�@��wj��i��vg}F&��<7�M���'�-W�V,ZW-��+GbԶ`R �� G���K���4���c�N��OŤ�]����B�*u�$Q�C@=��:2�<�xFhD~��J;{���[,���)�jV����Nw������3��oHj�pZ��6>��Q��j��<�S@����T\�e:LT�%H� ��șN�8��eП�i��S���f��=�cWcW�O��B@F�%�a�x��yd��(YBUf ��A�#�[�Mxi�f�!�$�ݱ)�B5#�7� v�/[��b��<-9k`�G�ju|�J���˒���m�򍠆1,蔧{�!��ǝ���x�72.�8�ֆZ"��6�8,���k�g'B��un%��a�k�!�tQj�6>����`�T����"x��b2�z�FP <x�;���f�?��s�9-��ȸ�K�&�&ռk� ��t5WvB�����L���R�vZ0�p��s>���4�O����+�AjM���������������YG�S�[��U0��3��Č��^���?@�N���ZN1�>5<z�p��n�ޕ%�j�V�(�rcD�oۨx�����w��.b�/�yϰs>����|_��x[yR��9\�j~��2�. �ĲF^��n�-m-c3���D+�35�{J��'/L�3m�lw�<1��S���Q'���q�1X�>$-6��m�y�4���=��T���z��S�ڸ[�E�����qh�[�g�8L /��=�iU���m�U1@��hɢŔP��:ܔ���"fw(�ךȵ�R�ٺ�]W�0rBz~N@�
��s
-��������p�����3��:���V�AO	c��
�B��rw��]�F=fj�W+AӸ�6���r���x��`a���25{�:ޟ�jB1vT]���1)�7��\	b���z=���C�:a��9\�b�ti-hK���y�,
��83a��z�Z�o|�m��p!��~-��`�.��;�N'K;].j�&��
��'2�}���M�|�#Ud~�0��J,O��[�)m��H����j����������J���gT���e��7��K	s̤ȷ�����̭�.��U�p�h��hU`3�.T���l��.�Q	��f^�}a2߶
�_� 6�M'l��[�8�":�,����ib����q=��4Z�&�w�M7�`�j���u�#J#t
I*שEϺ�(8�sO�?���(��"�~}�AB�3!���t.�1�e�K�����~���T���-Z���
�����\2G#*GJV�k��+�%��&@�.o5�?tbF�WaZ���PY�t��`��']d������o�;�c����X��@?�igG�Z��]�֗5�P����L���%�͈���w�B�t�k���סs��oT��?#U6���e�ֱ(5�7�,L�n(�?N2H�����b덢I=8"��S����i&��$0�a����G: ��4�q�޲}�:�E+xwF��k�xynh����1��ʃ�#�iz���#����d���P�~G�+c%f3��D����J�R�6�$����0����9nV^G�be������6�oVK�Y�1�9yo���N[��z]�����8�-o�<��n��� ����L�U��������u�����|��x��X�h�P�X��o��q��cV��E�(я�ʊ�������Gb#��ǲ�����Q(!��.�۩wp�X��L�VnF`Y����,Ay����ay5�;�{�O%�*R���&�e=�����A��Qd�;�۹iĭ�M�og��A�I�{�Y�
�K᭨$������!�+�w�RzﳴS^hu��T}�0�m�����3�ʴ�æ�ƚt��TN�y4�������G��-Jl��:~��K���vr����+�9{z
F�<�v��7�n��5���I�����5A�{RfF�Z�Ё`�����ϋ�������_`��2�A����|t�c�.�m�,K=k�%Ź^ؗ���5X>Ja�^JQ��D�����i43:5����G��%�aZU��0��xҐ��kʫE�^�KE��=���닺6�"�E���a�T�Ή91���! $5/�������ž�Ԗ`�����L�L��l��>ި�W=�ޣd��>����zҝ�4E`ˇ�*צ5O��p5Ǒ�T��xSH�,��qّ<<�xY��cu��Z�m�C~x�r�ɦ3t�ESȒ�쁊��#47PͩR�)����MPI�
�l��_B���k#L�3����L�N��Ж�'D�w�܊BZ��.$�9-uk5x<��#o�Z<<ۦ�K�L�62Wt\�Y=/����$aӪx�~���W���")�b���W`it�Vi,�3�������c�e3�?g�Jm�]�g��$����UBy�?�J����� ߺ�j"���T��E��v�m�1����0�#���%��o�ɫ��.��+)p4����~���h�f:S`�4�h.x}Vw ��b��@?�x�ZUV����,�u�H���
Й�����]u�EXyC�� ޽a���[7����<�x�%z�r���S=��uu�N(B�L��[��8�D�5�-x����6��d��67$�?�No������3�E�ɟ��nFBj�p�i�jzz��ۅt��O\u޺�
c�z�y�Y��Ņ�|�蕄�%fݎ8ќQ��/hq��?���o:H��cc�1sd�6�li�/X�e8���J�܉/���g���J���}����^�׸l!�;�v�O�'�>S
�J
�>���s~��@d�.�֛�w��D�$&d��e̪�����FR�0Aⵉp�}y��݊��ˮӉa7�}#QA����ǟ�mm�E��w� ��n��m>�v���.��[����(q���xLqK�l����J.y<�c��D�˺�[ܬxm��z�A�W&:����h��3�VJ�H=���1�F�P_�ӹ��`1��y�c�'�M��;����M$�5���c
�
A\����!�_Otڦ�uu�Hp��&"�����vƔ���o
����9�C��bUj��,u�՗�_W� �~,�^�Ee��t� {hS�� �P�e�or\�S>�O�K�ڷ6��s�c�zX䪇�5�d0���L��ѥZ�.$K�QS�5p�R��o��M�n�VlipL�i�bTJ�nT���`�d5�y���[P=\�ʼ��7/@�\�����%�"���/�:Lw��A9�l\*�-2=8o�ϙ���:&k^�j�3X8������C����Ee[J�	i��J���S������;\{�Ó2���?+�1�0y�
k���%��Jh��0�'�&"q��^���,�\8n�G�Gw�F�]��?q��z���t�n�w�P[�0�1�z�b���|}��ݏt��ۥ�>zN�R���\��o�-:~�ۚEuBRb�<�5ጥY�G
�aU6�&��&-�����d	��*�w��Iz�t޾K1zKR�-y���~LS�D�!�����1c}br��A��;]!6 Q�%,�yh&��CU��x0,&���"ҁ`/UJ�� :K��˨��C�O��f�O��Es.:��N
�s˓��%�''L���w0eا�6�-�3&�v7�f��ݞ�hW~�A8{�r�s��B��ӛu�x�j١�z�݀�C����>e<N����D}�oqpy$çJQ�
�i �&S+t?n+i"�j�!�����'�r!��Wh��#���)�V��B���5 ��͔%�{r���M��6кW#Q�͇�����r�(�M�?/YV#�dq��7�[3-
$����W��DwV35�s�(~3�4����aՏK��nױ�kG�{���A����_俜{��j\��'=�#R�,�yF�(2���<���dā;CH1%�5�{/� e��y禶
y����4KN45��Z���S�2��P�/��r�D���vx.�3#||��5>��6���O[�M� .���>u�>5�O:ЂI �CZx�N�C�|�F�lB�RN̚�p��!����n�nct=f�.����Y�����A�/~��$=D��OU<W+���	m�r����Bă߀�cL�{n�c�>���`2����Y�"�ܿn��ݣ������i	_<I�{��CPa,�piX���͢�U�ƚ�qr�de��@����Mdh������?@6�Ekn��M�	/	��;���Q8r����tj�k�`�7g��8�yeA�q��>���Nح"�?<U;�\����:��B_�F�gKj�"W��g��рE�N	�]��'�ǟ�k'g6����_)�W_����l�����]�q�����C���Vءoa6�q*k!!څI�I�Â�B�;�������$�ϐ��ʉk���������o������9a�7C6��k"��e�G���sr�򷻊�	D<%o�@qg��$��H{�c~WIwM9T���~��Dz�;1,N�yZ84�F��{��cT�sf5�j�4w+=hRc������ՊŌ�/z�4?#���j����3�GK�r$X�I ��7��492ϸ���N�prxLK���9��u�����֮u��Vf3솟����rcDH��6y��\[��܃>�ǳ�W��ܩG)&�F}H����5�M�b���k	?���M�G'b5|��$G��||�+,��n^�Z��Q.^��w��]ս���������%˳h�<"�_�;����D<u���ƙ�C�bd(��}\�x[�ن���\�p���ܫA�0��w�
���hE%�h�ZK�EǰJ�~O�ć��U�5ql��>�@ �K�S�}���'���c��$�1�k�¾G:v���Ob�����P�5Θ~�u�T���x����Z;^�l%�s��#������Sោ;�`h����fzP=@?}�R�	�Uy��cƣ!j�ʻyd�)���{�C����F1����oɇZ�N�iE]�=�<(��/��˺��0���h�qt�3m��p)��w�g�e�>f�']Y$T�M"6��>|���*Dl��A��b�#��۸�nc�T�u�=J�$ݵ�ʌ���Bv�XT/�l,膜�:)y^j��=2��yhG�޶N�����lVa�����_�pE[:�_�B�t
�#L�6i�w
V��^h}�j��3+��Ni$��	ݒg(h!��B��}�3֦��4N7�vY�ͯW�|/���ʪ�~�)�∣΢����i�)�T�	*���_ӆW5���E���CF�K�)��^��L�b�r�-�}�>��N��d�94�ěnq���\4|�y��</�ܓ]I����@8�my�d�J�3��FY)���T,�ڢ;��W��7����_�g����	8w��v��w��Cms�0i��)�V�Z����K?��כ~Y�t��"]�l��;���J�!�q�f�O�R�r��ϯ��\z����~(8���:и����)B,��?�=<~�a�x�h�����p�p�c8�O<�m2t��,o��|��Wd�(w\��Gl����Loqe��m���E����P���������N�t�Lp���,"�����R�	��p�cY����ì���X�S˥M���a��zD��m�V�S�v�	O��/�(�_].� ��hnD���\LPgK���H[���W�V�����8�T���?'o�l�Q}�EƷ�: ��T������.i�~�t�#��(�%!����A4|���Vϩ
�:g�=cK(�~��������Q)<���n]_����	ó�/��!��YA#iN��~��V�<�'*3/6C
��Es`�C�Ŏ��\��ẔO꼭8KNsy�@��w�l���t��l�����i�����T�@A��ś�"�bQ%t/WG�=i�@݃�_�g-���vYu:��l�F7�rY]
�r�m�];Ï�d |^k�s�M%�Up�����G��6�nB7Uc��P��;_����������`O�Bt�me���ňF?�D��!UJF��7u�%�s���8Z�Nۡ��a���m����F�ÚTJ66,�F]� �N��$&�����m�Y]�b��]DOU�ҘyW��� �'�1��L0�%�Eǟ��h��?=�=d�M��%*1�X�3C���]�Y7ʝ��}?bH�n��Q���~����hӵO���U$?��m��%F/:����ʠ�3����4ܰ{����Ȳ��(f�'B� }�L��sʈҩ1�9/�i�-���6oe��{˽Ak��v��ۃ&��R��@��]X�zA�c��ݹ������`O�鷵,ێ����7DLpk}N�������ξ�Q�G�ֱ�p��R~��}��Ү��ʞ�5*C5�,J1��$p\�vu��G��4�iU�M�I��)�͍=�����n�X��^��<��\XHeHE�z�ob�1��Q�lC> �!Y�N��RE�����
ɆnB����*IcO\��-����ͱ2	�[j��4�:���®#G#A���^O|�ѼV��R�s���f���8�y�W��7�<ϗ�pI��V��kj"c�ʇ/۝���IH��>� �����vn�ɺ�/��d�|��ӽ�b��Ƈ�>�ї������d?�b�vG�r���'�:���Wl�����Ոsz�:���GM��45���{o��<W�
�cm!��R��=;�xoo����(T��w�Ç�����&6@��U��3gx��tm��b��ŷ�XE=��pY6%5�o?�}�h-�e�B=m��:��:Ũ�% �,��OJ�Z����{Y&��@W��{��2����O-��%Q���F���_�v)�\o���'���*]_Z���,�pv~f��X#�e�t�oT�:�:3�3'k�!�C��"1B=l�6�,���崦X��={���y���ٮ^EO�P5/Ud"���ZhI�fz�n���q�Ļ�<1������陵�z=Ӭ�thm����~�RY�ܶFq��u#����~Z3��vh�̓�x`��P���Ty;Y�S�r9���~����[��ۗc���¸8�ԧo�H�k���S8ʯC�c�<��gޙ�OH�Zp���[���0߳��!��N>e��G����h^�w�Qu����n�Ű$����J��;���}Vݗ>^\7W� �T��R�J╽q��/���V��O��3B��
�8j�xa���F���� �$�$/�x�W m��\>P(�	��4���ǳ�|�g�P�ֲt6���ٜ���.����P���a�	����6��T	}���K�b�%�Y\���婫�C��A���#*��O^9�6+����s�n=rzQ�ϼ}�_�o~�r�F��f�D;��:G�q�8���-���\W>�)�"��R%�"s>�D+wa��F�d���R�n�I"�Oi�N1f���?����@�M�y��v��M�񶆰 ��H��k�h�0n�����$�}ck��N��ox����am�˺Y�\L���t�=W~e��%��}u�JaS��E'o�c�p�	K�X^��� ���}�/\�Z�m�9�X�-�^a�uce��M�g�f�����|C(��s{o�'���5��LY�b*4q�l�?��2 ʮ��
Hw��tK�� ݝJ7,��t��tw�twww-��������<w�83s��e�rȉ���z��h��(��]��hQ������6�H?�=�G�$#��BW���н��hU�9�:7�w� �����y]q}5����>G�����5����g3�q�.�%[1��H玩z����Jum���Se��lp���J�F����0`����!�5���(�Xv����?8� �D�#�Y{���f��[i��W�����Z0Z6?��~� 2;ұi3��Y��a-}�-c��l�m��й���|˭G'���9�����	�v�F	��{<m �h>*3J�����a������O�9�=[3��gr���:��ܸ�Y�ɿ�ݧ-���0�,���X�����<P�����.�=,��>�/.�gz�(b�(Pu�K���ڼ�V��Zӗ�^��%q�ʟ���3��ĽA!X��^���99DJ�$���Z�K#\ېw���ل���eA�-��}��կ�D7��3'1D���m�Y�Jp�l�Q�߭�bl3I`�nG�t��E��g�f��bQ��ƘbP���0m4�եd�"�D�~��_!]��Y ^-2&!p�BIJJ��+ݪ�f�K�J�8yp�2n��Y7�+{yޢi�Ll�O� U̬P�O'�ϊ
!˞��M�>��c��K���;��Ib*���O�W���Cܻ��ϸ���n<z�����������_(ᡳ3�7ȯ;2��0V
��~A�S����Ձ���guk����/[��՜�Ä�/�>S�I��B��y&V:��6�	��]����]djuU�w�Y�������$��v�2!9����z��y�1Y
��'[�V�Xp�|�g����e@�J���>lT1�N�P��<��Q�Ȟ��g��:�� .���s%����v+>�B����K��E����	7x�F�"��7�y�����p��-�[��Xcf�� T~���d\8��K������b�l>с%r�/�����A��?t��h�!FL-��^�_OW4�YC��7:XĊu��׷�}W��!�Ť��D���7��[L!B&(3#M�J�p=��ME~?�0t�|7 ���~+�H�j:����C*�f+anA��d��v['�� M������]gM���56H�GM���Z����cR��T�=�����_ߤ��K�uE���0s��5����IP����hED<���W��nx=D��4=H������gm��Akq�FYU�)����~�����4�*�I�h����v{��k{��^G��Oe9z���������]��wP|�rL��8�t�S'���Xp�2N�)	َa�g��b�<M�ߛ�� ;9$|��[��d����>�uSr�^c �Hl`��GN.Z�M�@Y��kX��h��6�-[����P�L�p����_!OXzϥ-�)t��˾�w�<sdԲ�(�u��Tv�IH�z� �Ş|�mu�q1�����oΤ��C���h�FY�ݮ7^["0�N�/̄F����2�� ��=�8B�쇤��B��P]�(�ʉ`����9i/y) y���6pW��"O���{n�ɲ�O�w���}S�w�"�'q��oLY 	��=,[|���z�w{����aD�UR*Lo�a����b���t���ayƘ݄��\�ߵ�q���~�"�'N�V��5{�y2X�X�H�aQ)�������Izjr���(��������5����!x6[��_�ȐBx�����$���tW���Ol�W)�\�d�*�2[?�����"	9�5�	y�.Ŏ�h��]�)��'�'Q&э���&���DK/�~􋽅'���J� �q���lz��V��1gg�3�6S3K},�������ń���r]��,X�6�N�0^Ȍߨw����V���b�<y}."6������<�����y���:��sUo;���	�>x$�3������Z>rcy�M����!�I��d<�?� Rʑ�e$��ɑl��͟�j�����Ќmݣ�(q)�<�,ʛߝh)L�Ua�'`g����x�=�lm�ޮ�.e��.X�>����-���l~��G�g���"&��Es����qE7�e�H_5��2�����`0���a��4�m�d�^�m�u=?��>��6�U�a�Ry�斉��c'e�꒪t����U��.�e���t=�������VH�E|�� �����1�R�5�=@ˌ���wޘim�r���A��Ĺ@K�.c�Ú3tsV����q���o����!��mI�Tj���n5� ]��*M*���I���A�-�����;�y����Oڜ��䖕�v^��������r^�cv�y{�m���;r�<׼�`T7�#��ˌ�� �u[
n}V����h�fY?�p/Dl|l��牣=�<�tm�d���o��[�Bc�v�̒��2�LRT�Z���^�|%�{�Њ�p����[<�b�[{�Z�J4Kn����	`�MZ����V55�0n/NP `���z�����s���~.Z�',����l�4�Sy���x�	�t8������̖������y�_htw��~��'.�gB2T��9����ǱҀ�Z6�+�t�E�����E�ʶ�T�#��ۮ�ތ�X����>��AC�^*s@���i����8c�K�<�Do��N�Wj/&��~)7E\�Գs%c�ik<VT��ʢi����"��d�]! s�:���ȁLo��&�~*�v��o�I\|?3��QA��e]h+v�c����@/���bJ^�lf�&�� ���筎7'��1Np�Ȼ��|}���-�_T�__�{�2���l����ZwȢ>�tpTA@�Ӫ�R���q)�_cC*T��i�|U��w�y���{�_�����6��Q�[K�9f��ʒ����3c�Ey������Hy��,jܮUz��qл��#]�.��Ԋ�����>O�"�O��,e�����T+�p?Ҁ�ƍO�ɼ�;q�N�ɴ�(��L���Eɾ�N#F!��s�y@��/'DDr �[辝�𤳚8Q�nn7��p�D���d��oDǦ=����WG�z\�f�ە�ɏ7?|Q���;̍%L��b�o��sK�f�����m5���ɇ�8�v�S�{�s���aس=QXE��kF�l͍TG[Tb��3V�(hS��rjh��J��o��ݮ_g����Y�R���ؤ�AJ$I� ɜ���)t�v'N4)�>��{��]�4��'���|����674�_�6ť�d��o\��x\� ��$�n���Y��D�q�l�8-����S64��
�K��1�����Zȝ���=_�5f��t`��V��v��Ǭh?TE�*��9Tw۬�%�.���f_e����3*�%��z��#�L5���Z��1�^&��X*sC؅:���L��]�s��ls[T��g"W2FVmBz���O���������J-yQ���� �jnY@}cwL�����x7���j����O�����S���.�\���;1��6���4]5�ϳ\� ���X���T�\������y���:����\{M0Đ�
�W�n���_��G��:�4�e ��$e��Ѥ1�Y��5����(���;���t���գ�a^t��� o��$�-�C��)C,;�уɔ�@�������fW 2�?�,��/{��L�])*�@/J��&1w�5�����*�;�?�o�#��9<2����Y��"�p�s���ïk2����V�?*��q_3=�&S��x�W;�$�y��hI���ϲ�'��$H�5�O ��)E��ayH�p 2ʯ|�j�ϐl� �����\����Os�r�X,��T�<DӇ;a��8 �a�x+�ٗ�y��;	��{�B�za�n9"�_�{���m��(��'&�l~�b~��
l�ym!�r8�n��Uu��	,���ߋ>��i�3"��x�MM��%.=M�|�������XMQª�1�e>@׮���io\Ĵ�|ia���N��$�b6�mVE�
mOP�7�IR�t���kt`t��f�:����r��=�&2U�����$�>'��j�޶�x.��4�N�Z��ϲ��[ I���^��(!����c�_5�P =���yR���o����چ:�P�=�x���y�l�KC��N��i��:y)=�|։IY6Ӹb�(�g���6Sl��a��YUE�X�fK�.�m�}~��*�M�T��|SN�h��t���%��[4��!����8����&/�
��נ��#V¢����T@��~뇅�[�����FT�&\U%���A�b����W�B�E�1O=�U��L�<�S'�"#�}ʌ�k-)�ᢊ���q���&��\�.Ǫ����/!��H�����ゎ��/P�7]�&�\D�8�b��G������Sq�CG�b����'|6������V��#
K�z�����4�Ό���M��8F�$��ҕ�w�x�J� >�K�rq�����v����o څ@�#s��F��_FP��r��ĺ�B׏D��7:e"�
zO%E�C�ܪ�z?f�?�i(T~8��>�9��Ϝ�Qq�r?�m���E��_��;�!�ǹ��/���=�=� (�R�)O��_��a1M�<��;Jt�k�L�
hUc����2=��^�����j4",
�1�����]��_'o��E`)�)��h�U�m}�����8յ�����B;�.�UA��{	�m�i�x�9LoN�����I!c��|X$씀A�?��}�RYp�K�S!;.d��T(}6��..�\4�q��G�Q?�\;��T�m�5���ZPfC.@��!��
�_)��jq��\m���F��4�t,l�.��ܹ��K3SoQ෽��S��YR9-���T�2.h�}�����?g������֓��Eه	3�׿���vm�zW�4��1��|�H�u�	��Nۦ�A.X+��e#e�1�&Pƹ��e����$`��c�\�	D*�b�E�S�h6�7v��sZ������U�% ׄ�a���3~��g+a�D�M�gρ�����-��W�^yL��Ԅ,�9����zm��0�lu)��EYL����Z܊ swXƔ�\���7�J��Y���&�����\�o���*�PW%E�T~�F��$}xI=�Ñ�Lz��m���r�2�B�_�Z������W�`0�P3m�����kA�F�1��i���62_ݧ# Fg�shO�S�KnH�����t�>RUNa����ʨ�a�9E&�0f`���|�v��e�DL,���=�@��Tg���(Fp�Bð�h���H~t�̀ǩ�%r�<�cֶ���GTX�ɛ�.f�X��ѹN�6
@�X�#!Q���ɛH���&8zo�Mp&h�ˤ�o���rx��~�4��Y���CIE�1N��*��(U���Cf�;���I=LdA��,s|A��Y��Sq���G�mn:D�׷�魜��6�:C�:�~x�En����j�k�:�5��il䨾�Op���`�ze�k>��P�]�L1T�_�C��#�J��b��'ȻP�N��Fw?�88�6m����+��(������W~�^2ȧ��&v�_	e讒��bSc�����}��l�?�P�&:��ko��M.F� ��n���= �����s�V�ht�a��G�v�����$��}{��Hx�a�b��kB$�zjk�����v���bх��s���u��S�q�0oۍL��"F`v�
�IPs�(�gC�(-�Y�Us�s��S�'��-����Q��²���㲛Z�9j�3�F��F�'Z��>���U97�m�������ը���-��=l��3���%��o=�y�l�C=_����1�=[g��K�� {��Tf/��w�6 fnf�4#�%`9V�%J��'� �@��g�5�{йw�����擵'��
�z=0sZ̋[uEH#�]��|e.Lb^twg��wK��.ǟ��X��pd�*�$��V���)�0��a{�&h����(��	�-//�NvW����n�^�x�z��T`�`�ߪZ2B�ַQ<<+�-z�l������:�WL�D�t/�B��Eg��j��ls8�0�L�L�����b?���x�'���mW�U�Q<�b+�X���v�o$;`�<2{p��p����6G�G���jʩN2 �me�
��*�l�?�N?���S~�ۤV�����ˣ��mg&gx��9Z?6^�}���6��loc5��(@7�x�d(�e�kl��}g��X�|�۟Y˙΢�̎=��^��n�k�¹c�����0F�|���c��0��@Gu!�G��X��	L�� �H���s��W ��D=2L�����? V�E�s�|<ЧY��}P�~b��\22�Q�+�;��ؒ�AB[W�$�,W�跼�nvxƹ��[�=F��1>WT��f履���ߪF�N����i�i�)<��-�k��������3�}�eO�T�v����_eSFr��%S�U8vy���.��>��Psϯ &��k�6�~"��y���=ȗ	�U$'1?��(4Oo���k.<_��U���gMS"�������d�^�'�QEm�� �a� �Ģ������d�?���T���	�����>V��Q��
q!�ɚ�ݷ.[mu�#�!|��d�.�7ˑ���h��E��0�־i7���9���c����p����~Nϕ7��}��?��!�2�\�Q,�ہ/��=��zU<Voܙ9�j-�:��P`:�G2O�3��"$��,u��GKY��L�8G7�Q�U���ut�/��G[q8�M)k�F��e�f]���[F��;2�恂wG��������	�0��߿��Ð�'U�Hn07�Z�U���#O9�r��k��)�+�[��i$�d.�9'8ۦïNԳ���
I]I(M>$탪B�)��y_��|ۘ�a��nO�WL���6��a�F�:]-��A��ܮ5�b%+��������g��C���Vu%���nk����K2� C0���jk���V`>v���&��2�W&<��O,GyT}*x�!#�
�ĸ!�J�J�[mx�g���c��j�K�,�<���s#�*�u��Fo���}~��D,ڃ���(�41�!�xzy��5(��װ%��~t�8ˋ�!���3��asuSn���y�����HtAԂp����|f"W����2��3��J^����
:��س������c��n(�ޞ�u�7��4i��=K�i�û�S1A�c�CMs�M���S����B�8dl�瀽ڻ�hTx�]���F\1�]9�p�tIL�[ ���y���0ө���c�Rsu~>0:��<^���K5�j�B�U_�N\j��Ƨh��v]zo����MClUOD<r����t3���-m���xZ(G�z@���E2����;�)������	o;�c���iM��_��R~�''5�ZƂ�Ϲ�;����HZ+ =rZfC�Σۯ���:Q56�sTd�KPi��ʽC�\2�2)L
~���>Q'�����Vt3��,��j0e�"53��agm�������\M��fN{�桲_BP��F2��o�GW|FJ�k9,Hu���[�QH�P������;�o����Q;dӦ�qP^�o���ӵ@o�l-@x��!�5��B.Gj6xb�|&2"J�`$�S���n�BaP�i2�lHI{`��F!s�Eq�*g�L�\���������h]n3�
D9��u�s��z!A^�]v+��ҙ���]�d�fY�U�{���;Z�麜/�$��a|ۯ����:?U���]�1�+m�M�l��G�����t��V��9�<�f]O
|������,Kj�| �#��8'ܱ�J#Hid�o���|�0 k�h�t�e�����[��������qo2�pZ�a�N��OL��/F=�<!Z<[�1b	����x.�|�E��4lB3�a%�l�1^��L0kn�됎��\����ں�b�l�SS�Bw+?�n`hoI?�]��r�%��3Be�-�~�S6E{Kﴲ�|�
��Y�kQ�A�rsQ-�zdj��hiB�(�7p�b\���]0�ծ�+&�U{��K��"]����o�t7y�7�;���a`<��KS��e_c���g;��g��o��=����j!����O��U���j��D�p
c_U�cq}l�����1}kn��TJ��fDM<�@U^�׎c}0��~�Uw4�G�2 ����/����
SS�0�m���5����x���z�eT˟��Uv�J�6?�5��W�
����&�(�'���p��Z�������E��l�
���	S�^
����ޒ!��o�F�p��z��q�^(d|���p5u!�1mĮ���S;ǔd�ve�w���ڻ'�"�=3B�z�J#�}T�DJ���N�������B\9�^3���͖������-1NF(�ξL-'gí&2*^!�͞�YIo�p�\����^�������: V��G��4�����t��^'����`�`S�ұQ�c�(�0ϗ��8>�3��0y:�9x}"�In ��W�����Z�s��6�B�>��2��7oR�>� ���[f���Y�MO#����Fo�7T�Ƀ��%7af�X'R,	����I{�̷iC��=ĉ���=�{5�H�m}\�a�?	�Q)�����mm�s��NJx��"��Ժ�۝���cv�_"���:��,�+c���YP�I'
`@qժ�ys�)j�!�{xo��k8��Mq;I|?[�������o&�'[��^PF�p��b
EZPZT��&�5�u�e_YV2�ܻ�tA�\G|��[a��Ag��$�q���-�7�;8D�߆�CjfY�)����e���S�1�ō̜�N|1�{�*A���.iȏ�1�P��_�x:�x�z��W�o��F�{�j�veG3�Z�`��<���
��
6 mU�}��[�^Qͻ�J
�3{3�v�E��֩�I8w���t��K#��Ȳ��Mg�4����u��h�ᝢ�Wj�B��f��ι�"��Q��V�Xy� �:��ߚ�V�&�Zu�.J>�z?77q�K�Є��9H�&) �"sp�Q>��CY�i�ǥ�'�WV =�/c����s��Z��|H9�����ñC�Y��w�w��@��V��0߆��Q����1c��V�a�O���G��3\^^�ck�����
nG�vuҼ�͠~�6w�/��Ƥ�Nm4U�����_e�X� 8�h�h�akѺ���9ִ�<:��o�n<$�M4U�����ȃ��1gV_��8����ց�,mWӘ��7\...W��H���G|>�O?8ap@֌_�qˣ��sZ ���\��G ORR
2�R�_��XwF�7�P��x��3��S�g�9��|&���!�|����]�R����6�&�N��Ŕ��r����x��%y�?�F90�YQ0ML3���`�nx�y�������iq�������%a�9�<'�+?=lܠ�Oɻ=�A̢5�B����{�#,L���m
B1���)�x��X�H,
*��r��[7��3�z�9�hTV�<�27�f�m"�-[�2�V�������C��/eBm�<��_�HB[�)�`�E�T�aT��Ѿ�̼�������@[����Za���lc�Ѽ�h̷c������otO����H-�qD��V��*:v�"�E�o=��C�U������D��~'d�N	o(Zb�\FY���]s#���-4����{���l��;p_fܶZFc�"�Y⯲H���n�Ӧ��s'��gk2 � ��ǻ��jV]j���߈)��L�8~�3���%�Ԟ�q�!��#�*l��:�:ݲ���%�Of_o�x8Ζ]�Y�P�2��1��}UPS"�!w�q�6�HcJ��S�LХR{�Z5��Uv�xi�J��Q�%�s��b�]2ZV�RcU4m�d���m~'���}�Ns]�<�3� �Fc�������{y��sb�])eޮ�a�TZغ�Ȗ���������io�J�\ �J8�5D���`�p�{�E��G�
~����x[�&��WF�]�Wl ���v׋_9���-�۶f��5��M4�E]q����mo�Po���i����N��[|�u���4�H���ww ��Z�9���3q����|J<y�9O{�����;^_�L��+�,��r�'6���Z�iz�U�{m�e?���C��b���?�UyVz�X�\�j||��8�aK��,S��D�x�Ȼ����UxB��|΋��(�����b�h�Un/��b���">�4~�!$%���Rd�cßӲ�&|M�+
����9#�ϭ�4xn��k߾�!
����z�O���l�2sKXINR{%�W|��:_��%�r�ù�Jb���A P��rb�*F�?���
��#�i1���[�}g���J6.K(�讯A�sHt|��˖�3oP�"|�7#\�;�|�xu�=7쑉M#G��6�c��A�5��9���J��he��3�uT�O_�iZ����{�WE_z��/Ҁ�+��9�J� ;�w�B�W%�����XG�#&1�M�h'k���9)�6%>���/��Y��wU�����*�N��P��R�b_��������'�+��6�믨�m�Q�ᷖ6���^�w���0�wˍ�l#6��3�{E��2��O����h����GC�UI��}hs���ͯ1>DJ�ǚqr}>;����:{�G�H���6(��J�|?�.��M*0�jc���D��Z`&GyE�/��Ч��)"�܀�3�O��/N�㭙�\��i$ƥ|��s'c��M�xi�y��c��6�������䄄��3N}A�nM�٪ƪ��d�75�z��S���i�6g�A�,@>
��р/��Y� ��LNȇ�󝝋�1��te��/+���ѯ�`��]~e��ŀT��89���nk�g!G��3��.眣��+���Dx}W��uBڍҀ ��Z-8��~2�|$Ij�\;@�HI����:�_�8�ahs��;[�eT�4ϩ�ڭ����i_�2���({�͙3�`�~��+��IT�l��*爚	O%�c��>�����享u��������j��G\�"kcrk��w[!�'�vU��}�P����2yab�{��2��RhTP*�vb��be"=;h��@Au�ҥ�KQ&��a֑ͬ���*�W�۟����/�߽5��6�����Q���e(�Y���5��*M��ї4;_n��2<��^�6�'��	��9T���h	�9�d�۹��M	;�t6}� k���JI�@f��p�������aｔ����Jڢ}�E���c��`��'I��A��1{�["���Q��3]& �Ƿw2���Xf�\ں#�ۘ<����v�1�5��h{]���k�ʨ��-�ڼK��� 7����PYvOq�m�盕�!�ԫ0�3M�;�-C�-8���2N�3�-V_B_�A�0\�Ҍ���l�c�2�W��ħ{֏U�E���e�@�Mz̅	�: r�`�;�^^�������� Zx��]�E��Svs��H�Ӣ ���y3�+n`��x-��M�E���Ƌ��^��F��2�|^�
����qw��{�gy@�na����byN��k4ZI�64��x�,ئ��� u7���s�vN��X��_q����"#�X+¡��<~�xIok��D��-ld'e��y ��n�Y�M����u`�@��
���G�5ȪNe�q������1�[�����K#��}��߱!!A��gaF���H<�~~�S��v1̈�Gڐ��Q��B�W�:¾�M�xL(�rH�4�
�i��`��
-����<9;T�O�DN�bog�k\�[Vt�Τ�Vc�$��۪��A���H2ĭh�A�H'AD>�\�T����
��I��W���'�����������&��+�~��K������(��6�Oa����&��&t�$bc��
`y�L��K4��;��qk�z�eQ3�_�j�0����4;�G�7����/�LWl�N�j���IHFϭ����a�΂h�Z�o�{*J�l�&����t7���?���i����pP�,.�Xe��vʅm����D��!ɔiqGS0_�W�iJ���uS�R��"E��X���ԓ���)A�q�2���R��l/�@��:u!Fl���dFCgZ��M5���sy(	;���`�3����a(#��g�g�������8�kY$Aݧ��~?~�4ڌ@��W�MA=�Ӷ����)�YS�u��lv�vx�OA�<�H�a�#x��a�X/1�z�_��W6�H�ō\���,��M]K��9�az_"�V��[���n�8Z�^V�@zz:�mfL�܃;��͒9�K2�6a�g��m�cH�]�W�L�9f� I2?�;$Q>�"� 1U�a�.��L����'d\��������ZU��ۑ����欧��B8�0�l�`��0��wYC�-E�`C C0r�����,K�b�"�<�G�"��_�nq;K;��r��������|V�xc$��[r�=C����q����5�����S�~����Z���[�V2��U�i���e'�k7��\��FQ}�����%��N �)�`�톯/�e�xD�|���+ȋ���2u#�_�1��y����;�x��;�l]sXE��N�fK��v�b6�9��q���^��1Z0�_��hS#;⟗M���X���H>#�P���їc��( m� �E��\ ��%��#,�3�����г=X�Z�;��L�НU����2���F��#P����u?T�<�궫�Q��hׅ���Mf�.c�����~̈́_�u���ZǞM7�'/N\>dl~n����HTG�D�9J���q����_����]`��dF�@d섷�+�Ч����Y>߱�gg�uê��-�(�W���i]%W4���=�&�1)IɊ��|f_��m ׇ�w+t����݅��l`1�,���[���ш wM�|͈�%��jo'KDɟf}��鈬:�����M���`�(})�����t��(-qzV]���٥���{���������d���e���՝ȩu��"��V�4i�|aR�\��*��q' �k8t�J�Iׯ�WWri�+�e-t0���]	�$���IG4�"��	�V����|c��~E�J���<b���--��3�����L�9����wE6�yqT~�c����|��	-B��7[3���{��gO
*�A�_]���YL���g0*��n��`��"
�I�����j$is��r�丛��FZ�M2d<�SŎH�}��njF�4e���I��e��O6M}j'�cL6B檣kVض���p�'Z����)�d��$�3�m������v�/���H�X�7���sZ�z'^��4�G�%u[�f%����+Q�]�Me��4����%ό�����cO�牣2���ί>E�$=�P�3���b�z/���K�L5�F���n��(�x��q����y!���.�@�����Xs�IݓP�����DךJ�~L>*Q57���c�̋�u���p3��﵀�z�43Q���r���m^�i7�iH��"���=jO}�t	��6����8>������xb�%[C�5�s�~�s��nq\�0d��K���$C�l�U�'	6�u?�e��x2;�gA�Ȝ��@���N椼I荍S���`%�9�X����z��$�0n�V� c<��>`(N ��#�B'(�3���XksK��uDO�"�cHm�Bӓ�?hi�IՌ�K�x1��g�*�Ұ?�!��y��g濜����#��8�P�	)RuXQ�ۇic	w]���YT�)_A�����&���Ͽ��lH7�Op:T}�ׇ�2q�k�Y�۟��w��} ��bR����ZXXXI�l�,U����k���]��?:���8Uq�ؖ����aV�[����^��\�ޖf��BE�Lz4�T��߈ʶ���=|
��mɗ�k/��'��J�fJ�f�&BX�헦�E��]�vd,Cxo��f�8@�i��Sx�2��A����vh����*&B*�Մx��ɜ"L��'��c�ס���{H4��WJA���a��p>�L�9N��d�[`줯ݚ.}A�x�!�����_N��pԯ�I������7��x[8�^�^`ύ��� B�DV����\�(Ql���I��ߒ���������g��U�0���_�\5_V�7���6u�^"݌e͑*���`|
�$ν=�s3����y���CRi����>���+�f��Ǔ[�8�U�~8�nT̛�2X�pᵿQ��D28|��)���Q�\�����գ1Կ��Ww�1F�5�q|K�����[t�)3'�o��`[N"�Q����%�w����<ӿ��N�neSdڔ��X����۶���--|�9m�"�欮Y�^hA��<�Z�v%��|�m�E|���t��:�5�HD�4z{�)�(>�?�Ȍ��W-g�GQc~_���u+�h�� D+�~Y!!q8��R鋎��s�����HϔG��C�X�,X�&�\�:�5�r2�{�/��N|1���6�7Nw}��n���P9:d�hq4>�D}�d4sa^�J:a�V��1r�d8?X.�ʭ�X����;ȶaUM#��������cYO����I�2DEE/>OfԄ����s�{iB�b�\�����yl
�7�������Ty�q0�����I���%����`I�#\^r��u�AvNǿgD
�����(/I�mME��qiƇ�?s"N�?��.K�5����*S�8�኷�u�B@���4!��X:��E[=�R��O���x([W����}��=��N���Kw<F`�Oȕ�������MY��_��[�c����Q��|���f��o��%L&N�±H��sKH
�����P\����*�떷3&���@�Mj���G��tg�E]	��ҙ���m�F�&���&���]��y�"v=�'?�Ț�뗬���ѧ?gZ�5e�g����8 .1լdk�r��;@���?�S�.>�Y���.;�,ˤ�{���K��ph��_�&�qP%��n&nA�/:���.g��.؝�I�z,��r[b]��Ո��{���>3Q��X�����Z�0G).�fvO�gJ��3s���s�ϡ�d.��2l榔�ӆÜ&�ok���GJ�X/[Z�h�^3~�@��~���x;>G��9J0S^sJ�_�"wj5=t�-=�x]$����Cȩ�t��6-s(��v\?&�&����(��c�X�s���kaK?w0�_�ݨ�ԣOLߪ�vא|����`Z �7X�fI�4R]�U4@!�(uThQí�9x��6{��M12z|(���i�v��1���TM�B��n4CHWSt�8��6�[}��d�\��+.���i��_�H���d�nD���ǳ�c�86H�s�!��9��tw����]Fτ��2S� ��xIF��2��Su�8�K�
�"1;�w�W^���B4�~��-y�y�����vM��]��~���x��3�A�No:�u�����\�N��֌&� ���9SH�?� ����9����s=%4�w���x��H�u	fSV�$cV툑��m�섣��BpW�CV 禕W�>������_$�4FOצ�{�e�LC��&ԕ��k��Ԋ<��sx�Th*�쒤��Vu\�,Š�.���Ȫd�:�Xү��h��xw�B�c�v w��x���42y��?Xl@������f���b���@�wd����.��N�k@�+�J1]O2G���:�8ZE)j9� j��)��k��X,DQ.Q�#J[���[D��x��	�2Z��ǌ�x���(���X�p��D�`�L�hƊW!��5ʎ G������u�Lo��K>�=��HBmِ���Z��}mĶjIB{b���A*އ�\
�r��PB�t�	v��*5��M�5]���}˳�c,tѦ��^�#����\��0�	����.��s�@�J��Dg҇!��	��,�]��Q��1���<;(�m\]�ѷZ_w^�*�
��.$}�ĥ����;������&2K;�/g�u�S�Ik�_x���5, ���|���7����R�E�n�y�6�La��ʔ��dn�tp�z{�m�n�P�[j�^��LGЄ���KoGd|�ٶ�ʶ1Ʃ)��ll��������G}��A��sVF����H�[ݔ�ۀ`�X�?���!�_q|�w��h?b�M����<��^Y������ཬ`/��"�84����k�J�#uE���ر���,!��5)M�/n\�Η�=�n�0�L��2R�E����`�����?�@���\�=as���	��f�K�K������}y��*)v�i�é=�v�i�Yy���G/�>���ŊȌ�T�vB(�G����!�s��B�m�*�ũ	�?��=!\evd.��1���u=��?ܦ�դ�ո�m۶m5�m5�Nl�<�m���ϫ���}�s�=3kf�s��g=��a�T�Y+�ea,z�z|}�7$�5�+�pB�9�F�~�E�@��i|��3�ǂ�dz^����C�R� 	�6LB�wv�V��s�g:��������~<pc�GH,``�����#���o�Ǯs`p�N�E�S��� �A���ƿtQ���~9c�c )U05�}5�×ܕT��Ӣ�n�,E,ڦ�l��޶ax��z�K�Q?4�2��[A�����P+�6��i�vT�7�5X����]��u������I�����`A���[N�W<S��o��"q/�n�J��;��Viǰg���8mp��X�7<��3sOnwi�ZP;��l�8�6h!+�'�YN;R��Q�z~Y��ˀln	�\Hv釕�s�f��n�T�S�&�t���d�+�	�3d��%�n�+���?�Qns�m�r�7B���b$��m�,�6��D�MO/��k�"���޾��E�!��,��r�f(m���~ę�1%CZ.߲��79� �Z���k��L���T5��wC�&��s�l�f	E)���.����wNily��l�����Af��>��P;�!l�N�*$CR�n;���F
wm�)*wr�mNҤm�3�z���
�0FԱ�\���d�(;��7�*�}%�_�Z�\�EfA�O�k`��
�&���e�ܳ��ݨ��2�g���H_Β?��?��-����e/h����z�S��:F97��S��8}`�L$��#Onu^�ћv�$n_�^�!OH�b���!���s�z ������S�'��@��͕�Q�:#�K���MS
j�El`�,��.5�I��
���a�e���	c��ھK̠��ʕ�C����[�Ad�f$L  �(��ƈ�y��z����0��8�AB����5��HR~H���F|���ֶRUIk�4�1���Sr���=3J	M�^q?���IHҀU&�y�b,��`����6����#Y�C�����hځ�s?n6��������O�2|mX���Nyy\Vu��oy�G"Qm:M��rZ�)�P�f����6�qKe���9���:򪢭�w�H��b�|m��l��4ْ�X�vW8�(�#���S�R����6X�X���
RQfB�#E���
��� [�׈Z���?j�2�[e���t ��|Myi���b�5D�BM�<�RCrC�C�E'GIQ��RtF��姾������9rs�2�H�j��݈O�d���_�H
�2�Op�vH�̱���ͭ$������.D�F!��_޳L�3u����|;��QϵJ.dYs����Rs&j�A��i(Ɔ+@ ��bv��ز?�T�$8 >��4ck!$-_�D��0@����U��Bm�hj������3�������"4����nn�-���J��)A����?]��%9g�F���`� �a���ɖ��G?=�2��(�ǫ�(V&�9b�l�i����=��7J$����w_A����������\�T^K��/;*���#_"���f�f�>՝d^Po��EPL��P��Hm�&�V��<qgE���U4��& �tN�>r�����{�m�� ��2?� �g~����M��حo;��+rF�q�)�zgDjr\�R}h4G_��� kTg0�T�B���zf�+W���ь���H�}�Sn�����1�5N�z�[2�&i��S��z�F˸���2��1�`j=���HE��5l���ѥ���&/Z_�]/�����ɧ�/��)��"��X3B��q��4���Q��q�6��J����V���I?9ewj��=�d{�^v�S{��`r����7g$�4���u��Z�G7<-=H�>���J�ps��m$cL:�J�ktm����?�v���yg��o�muhBg!+ϊ���$�B����G�����1��"��������㺫3�/O�˴��q�ؙ���>�i5��7)�L؞���:T$-�����zXD�9�Z!�w;�~;����z�eD
n:�4p��c��5"�A��۔*�ʪQ�
�\��k=�ፏY�{���VX�^1Z��'z>���Į|A3t��-Um/��s#C�+��de�$�xT3�]O;l����AL����y?��������q|�ҳ٧��h�G'�;�Uh��UB�7���B~��F#�.�AX��x}�B��'�� �V���R͘����L�o�\�t��^x���K>D����γ�X�b��w~k�O-�J#]�����7l�M���-t'��A�Ly��[?/�r������� ]5t!W�>�H�3�D	�vx-'Z1"ը���;#��(�Ih@�U%�Q��5tŲ}�0G:�(�D�@KLK�EK��K|Yi�K1�����U%Ij�������
���2�� �?nI׀NwV��7M��W6NV�O�����hA �<$(�8d�˷B���R��&�&�c����Le�ab���\�������a��UD��H�j���yKU-F�D��3k(G�57�$4��d�V��<5J�.T���uݧ}��l% 
h.�n��w��R�"�XԱlluDG�����v��v,)h�����%>�T#+���?�(�䋼Qftj�e6M�XܞЍX�W[�G���%�W�@�lW`-42
�s�"̃�7�0C	]��(�N��7�Sx�qP$m\�\��
���p��K3$��N�~���'a�h{�U6���!
ж�%�*��Z���o�j�A��$*��6;|&B_��\8��������B�B52Q'�?�$��0�[���l�	i�oS�����ǒlQ�:m�8�: 9��[6�*�UE��q��8�`9͑���QZ��W�#������m��<��`��J�?b��U7�:��ǂ�~�@���e9�#zPŲe}�]EM1�9k%*�I�P�!��?��!r������L�Py�d�A�i��*s�\�楔X#�2���ܓgH���gk�	�ݠSk՜ ���X}�����f^\A��v�y�G����"��f$�PC�YG���ɝ5���P���ɝ9�4����b��v��B:yL��`��cّ��i�v�V54Ѩ�s{䴢#��h$	��;�{�j���!.�f*ϯ���W�\�!�,� w���|l~ε&�7d�0B�T�Q��+�t��>�f����
n�v���)D]�ưo��m�D�P�3b����tנ�z<�-N��j��D�C^�(W���I�թ��/��h�[���?��Cxd�Gh�#8>U^�7/�r�%���
����Qh�Ū*-A�V0�R%���NƄ>�{/�M<rS,A�z
W�qnO��E+4�)�L�N1K�x����[��ssȡ	�Z$�d��>Pzsؿ�ҨG��TxO@p�/2�^P�7�0�<��C��`�b�f�M�6e�����m�o�����VKa�#���ʧ�6X�Z���.lk����)���u�hG<���)X6�`��,�e�E�a�B�Js�2�iRZF��=7d,Gi}w�+�'6���s����g��z�ag ,P5mT\ޔ�.����	����J�)I ��=����f_	��5�B&Y*d�ݠ�e�����N�8�/���m@��w�l40����������M뭡�dd�(�`-�����s��+������L�n:�lDk���饔�mdo��q�C�H��^�V��,�@��n�&��g �Ӻ���$���	�Q������ʝ$�h� ��b�}��Hu�2��������ہ*�	u1���r�%�%�V���x�b�P�!,a��"jH84Q�Uf���f��&qO���5r�b/ⅠH��$��UdC�(FH���ʹ��s��|�pϰ��!�� ��<�?D��к�z
��g���d����}EE��ڋS�nv^��"'��R��/�R��:b�4}�w=��A3'=,�C��gC23��\��B�t���qD���¥���&��T�V�<�.�Cyq��1�}�֕[����+)DZ��;��$�_�To�`p�^úSk�ħ�h���Zp�˰8.s_��a��~��D��rY�Q�I���;D�~ ڞ�3H��BTꅰ�ێ2�a�3�笋���*���#���圄�p�[ [��]q&�}@�r8[��P!�D�w���}�}*�R�ߟ���ףʕ:F�%�c���Rn$=Z�y�'�΄��m��ߧ~<i&��B	u�	�	��p�9���ٝ�������!F�THT=[9�� qCen��5�;�.û��71Z]n�=(���QO�`I�D�~T^�R�E�DV�N��[̜��b�G��3��/Z2���;B�^����ծ�e��:��]�o#�����=hޅ ��%.���YA�3�{>e/�ZL��ړk�L��e{*.�,@'X�+�,�f)��*�0:� fP��o,I����n�ujqs��|ffy��rq~t��۔yޮ�r���{��3���&jIĖ' �v��7%W�a����s�6��u���$������.�*�a�XJr+�0��5�w����$�ڢ��H��I���;M�uzgR��-�B	a��8����/�m�m�����c'}VP,Ĵ�S	��B���[����t��NE[+3XB��V�ɠb���
��Ev^�F�i͑�0W9$g&Vd�E�U��=H�_��m5�NM1W����,,���
�T��]�V���G�!��@^[��a��T�CC�董$b���	�P���إH&lU���.�h4�ڭ2�u������Wt��b~E#�c�!��8rC��#�+i���@��ϑ��:oRu����pѡAȉ60�m�Pru$�S�>I�M�1��Ε��C.J�{)�*&3&FAM�I,��Օ�p(��!�A��R9-��8DXq�~{C��L�	��	�$�ymL<��'����۔�^N�m�������lF�E�����G����~�	kP��RM�$�^%\t�Ȕ����b�C����mR�f��2O����⇘���k}q�:,�4&�w���i<����~����&�@� s�]�0���n�A	��/���1a��9������·����F�Q= �W����*���i �q����H��"G���
�^�44��Z�0��<��l-Z:+����E��h|;�1�y�(G����a\?éx�(��:�k"��ujq!Ty��
<v��9���nhj٫s���<����C�eH�(���?�ጷ]w�DI��!A��p���3�8�x�P�wd��º�D��\�yyʨT'akiYTW):�t�o+Q�\�)�����11|��<��RHiִ�{r�<�xm(�$����i�`����n��ϑS�X�?�R�N�%�_����(�c��y�b�Mc�|�$��!�bn���A�V9��Al0I��ͬHnÆ3��H`|9A0�l�/�^��H�blc
0�������]�0~�d1 ����%0��#����P�6���ʎ�ؼ�o�)
%2�gj`��Rd�[c1���I1پ�Dc�_�i�=����Dwk�����Q��.���N�K.�u]�� �~T�ir�۲w�5��p��E�E"���[yړ�Z���ʩ�5b4k�Jw�,0;ੵm��J��ړ��_�簷"��V�ƪ���ԏ�[��s��nu���	^k����ϕ����3&��2��%t-d��x'܂Y�f��幭V�޹HV��[Ȍ��֛���n��N�a�7+Z����0X)2i��������t�D��29���!xm4	�^���-bd������05�V�`.:r�Io}[5���u7�{��=�����7�dn(���������%��-E��3���e����`�Sl����4Ɏ�U�$G�2�����?� @4y��]u��ږ��yr��@(�?y�Az��U T/�.+����k�#.� �rʐKs
|΍���8�!�]s��w��8�EѴ?���f���;L�8�֞(@�J�}��8�o�"�s�u�U��
ϛ*\j 7���k�H�G���B��@|&R]��&;�獥�p2?(���-%�ެ�l:�:'?�k�x�Z+͈ G�ҧ�0?%J�Ԝ
�|ÞBK����P�)�%�"/�k��jH9nD ����z�g�|�X#ݟ4lH+��Rc�Qvz`j��,��mW�v�Q� v�$ �h*t���ͧI,�̝u��N��A2�6��l��o��D;rP�"bLT�.()�|�������Q_F_|��KϽ]p�+�O[�%v���'B����V��%=ska�3����E�6I#a9���㥨���YU�e��o�`�a��p�Y�Ӯ�UB��p�}�0I[�Y#��ɨ�����lP�q���k�+e�,4`'��bd��uJi�Kؿ��_�e˺ns
}�FBgA�ް���AM-�L��CD p���n�*Zr^༞����,�[���V�q�~p��<�]6F��G�F#̍��D����n!����_��n�g�b�m.���F��3͏���h��6�O��gaA���|ND���oP��^ۻ�o�Jw��=���*�Z
Ȟ�
L��BѸ��d����s�l<Y'�	Z��y�����Q�!��h+��z�I��

[geCg�\z�M���Z&ַ<d�lS��G����
!T���qMV����+F�����P� �Rbe�ؿ>��fu\T�۾$�W�G ���Ɩ��ǒ�g�CG<(!o�(@�وNӨ��V�q�D�uun�䑡u}9��8˼�7����@Z�E��'��_1-�CLc7cl�� �	�.��*V�u���Ip���s����G��/�"��,>[��&�l�B����1��"��8��G1������$���1>��1�1rS���xQ��uTP���P�*b;�����S�8�dq����a'-sI��]�a;�A��v�8oa�*N��r|s�	��a2��i�rC����˵��k)���efR%Y֟�l����W�R�d[^B�H~�9ii�#�7	�8v���R�۽�g<�Z{՛��i��.���+��l�댄sY�Ó�X"s�W�^��Z��"ٞM��^���?4J��uk9}&1�
R�Y3Rv?8�B⌤�d�lr\���|��ʒ�\�`�U�frd�6��S�����@�/�Zq�.q��&e�p�{7 N]m��tY� �N�nE4(3�4��'$�@�T�YN�6��e6�_cW}z�����8�$ǽ�YY������g��"��V�w��XZ<��߾k���2	�@f/�m(%C��l�)��jx��V��^}Q��!n�N᫪p(����-kk��[N�����i4��a��+,̞���Ft��Q�px�r�2ҿ�j@C���GLD*� M��?��o��Q��]� ��{%��-\�6�JL��E��^��`Û�jn�L�2��[|<�{ȏ�C��S!H8��_<�}��pӤX���5'Mlb&3�Voh7S�.�,>oS�O�d<iP�%��y]�KUrdE���zt�LTp�mK�<c��[�8�A �����x�Y�cX����8IR���yA;쓖hW什d�	>���uLz� o�eşBG�i��s++�xRRRİ��Q�bwww-���)c���練��iv�@�Ƃ\����,QbGK�O�to�vw&�ޯRlN�������+rh}��5D#�kLd�"$�Ѕ��۝㳁��`_�������J ����T��ꒋ�R{9_*������u��T��,	a��Z��K�?d�YG��������[N�����딃�v	���{�o���ҫ���p��<�}�u/.+��6����X_h�.>%<�ך�M��«���:��w���|�%���8x�6
�e�R���|s��8�|�����j�o5��-�~0�!DQSv��8�����b=g��*�gNy��[{�9���e��n�b��]V�!��h��V0^!�Dҡ��x�ZPP�}��W�[�ps��3�M2���B��R�v.[��5G�*��r�L�Ac�,h_p���P~,�B̢�70�j%�Qex��DI���bQ��d:��O���a�X�����N:���WK`�B�F��Ǎ1�ú-�Ӝ�sa�s�(���N�_���c/��K�W�v��G-�5�3����GxP4R��팿�}�i��m:�H#�x޿uԸN�$8zLr���5,j����E�gu��N_x?p�$Y���8�������`�T��s�q^<�8Of�r�t�>�\�}��������� �=�՝f�g���������E���,��E��nN�oT��^�d_� .|+ +a�UG���!X����B0���pߒ�}�7��0;=<.�Y��:m.n6��x�̆��לgÿ��pڬs����Mb��Od,s�obn{^6�����_��_,I"9M���y�a���)r����'��%�e�4o�r<���^�S����x,%SF��~c�����z[�稏������ՉMe) f��ͬ���6W\FNg *���"�d�J��褳�^�|��=rF3��|�2t�?R$�����.o�v��0/��Cߞ��X�'B�צ(�,��7�d-g3���ܾ@6�=�!�{��q�>��i)Ur�?64�G���px�m������A&��o�����ѸR�Y��"�j�� ~w��6纙`�gn��S�Q�������l��T�磢ٛI�`l{�Nl��C燖�K�W�w�� �z�k������,��G[�ʶk�7�㒢۷�*[���4e��V�;��lxvQZ:��A�[�62¶�*�����b�J� ���B���!f��D�G�|��1IB.�{�V����Bd��<���1�"��i���9.�"0���3��ƽ�3�����'��j.w�ҰS���B��:�C��.>������w2_'%	=��	vk\��o`c��s3^��踝���x	*��xY�0������Q���|�'9#2��8�Wx����Bq�,cY8:�me �{ ks���by��y=B�h������
��F5m]�X�di�1����s�fQ�+Aۮ�,�ؽ�c���ɈvV)����B�n��g1U)��/3�n����͢l.�_L=;6�=D��j�,k�ê��*Ia6��6��޳*�]�̑ldG�۹�*Ys�5��O�]��yn0�9���Af7�~�B��)���ޅ�y��X	('���0�pb@#�i]��J�yp��@U[�y>�1�h%OU���\��T��G���M6qUs���L�l2���a<�K�$)�����έNbXm�Zu��1����l����T2ޔbj����4���D��!~�4����%���C�=�C��q=�n�Z�[���0'�����x�.��������vUaK5�h4Ew"O�;�4��߱y�A2�ה�;Oz�����Y�>~']h��:S���cv)T�Iud�:�*�r���T��2�ګ���0��>�:~�����xO]Ձ�/�n�TI[�QըM��m[��Z{Re�%B�QM;Q���EoL���
vo[W=Y"��+P1��h�42I�[� {���u�o����Wi��rwҝ*~���-�OaIBD��{~�V�t��rZ^a���U�غcM�=}dκ�	�P�:���|0�0�]Mv�ײR�dؽ6>/�{1��S�i�rs��A2������?�/cb)"Qqw��~�-��$~B�}�������/�/����lws
w�����g<��r�`���U���V);]��Q��j���I֯�Co#�x���xdE��>�5�4�M�7�s��F�[������V���iV��2�?�G	�R��6��ERk���=��_E�$�j]�/E �M�wk:n{mz�ˢ�q�Mz	��P6�h>]�3��#�ō�]t
=���)-�q�-B��3����Me���8�i ��bf"�|b�`�iNU+��s�d�Xc�{�n|+}v���͚�44|��J���`�G����6�Ƽ��MP��Yܽ�<���W����z�<�^�4n+w�}dp��f����4똥E�C��x�,SG%� j�SR3�ğJ��n��B߽UR�0�Z �ԾQ%DĴ��q԰G�jE~욕��ڞ{J��A��/��A\�.����$�S m[�+y�cz �3�����I���KW�{�PG�#6�, E��������`k���)Tڒ�8�KC�!*���Si�ڭ��d�]b�
AΤ��{Ғcs|�7vN[5�-l��������e�?�f�ߒya�D��Ս�<t;yLr=��lWL�d��{&v\�F?���^��^��A�7du2���봗�pT*�?Ń�j2�Ȟ ��.'�j��v�A�:�=�����,ծ,�:ĠC��'
�I}�DvBakR�ɮ7��(tQ���̔�'�$a���J@��X]�,GV������_rZ����L��;4�x:dE?��^*H�L�4�3��S	��H��pf�b�tS�^?�|�WO׍?�k��(�;K�P�"*)��t��oi��n����oϩ��v'�&�l�-u�D��v�bv4S �	����$ދ�~	Ѳ'��
��M���W��v�C�k�M۸�co�ݭ?��Mi:{�[�"��e�M�W�8�o�)�(W�H��v�4�����C�L�}���?���+�f�_?���f�������H~7�ny����Ř]�"�.�V��.ٝ~Xh�k�N�w{�J8$�j��f���]�k䄢�����yՓ����̴u�ʋ�2�:�o�S_J�ő��{��ǧKc*�)k���r�չ	�&�q�߄�XѤV�<j�@���u�6��4�c@��w���%*�)AP��C�~��i�D21�f&����h��n�|4u)��Е�9t�G�a�\��lE�^^^b�P�����:M{3�ch���H����CW�į�i����ٳ�2�O�Ǖ���<�u�x�wĊ9�H�����',)��e�A�.�.���;�N�
�1U�Z	F�^�Nl��W������/�-C:�$x4��Zm�%�M�xc�-9 w=d%�GM7_� "��/z���AW!���	=u�|V���5�¨��4�2P㆕u�s�u�m�˗�X�W��{�;�s�k�����>�������<1�W|��A�8���fr¶���"J*s�&�����ΓEK1T3�&�}e�����!�U��~!��V�3�� $���bp9��I��0������K^���q���4~�#�K�n�àOu\v~�t�*-K���TE@�����x�뇮�et���Oh��' EGoZ��>��cl��Z�tѫ��Յ�u�i��UU��A�����-����s5�G��[V�R�{�s`���[z�˹u������1Mm��-<���E�}#��J�R"�SOU4�",�eN�8')�*�P��{��V�M�"e�nZh��(Y�{�~P�L	a�N)R�v��C����t�=.����;ܒ�-T3�zX�ineUh�00�q���$���'8�M���e�~�� �đ��Vז�6"�CU�R��f�O"�������)L��w5����g(vk_��t�ɮ)��yӇ�����x�5��ͻځ��<�Tͺt����$`?��������@�����Z��񫻊
��vJz���ѯ+�����_DfC+���f2I����ec�-���6C���gl�&�ڊ�-G:��ކ�âi��引QV��O��ac��q��ac��'��7�	�B�\�Qv�e,tO����1-��߶Sɴ(�iz߿\0�8��z��@�ՄP^#��13G6U��O4e%+��{4�tÏ|��F��wƌ��;.���QBH�*���(��������ȹ��l�#B����y��
�bP��> �cђ^���Uو�]��Lfur�VS�og��u�ѷ��-�|vf� l�����q��k2�A]���nr��"<�HP�`+`�����zB4L�T�./t;y�����.�.��`�H��_a<�Vph�j,�_��Ą�X�ֈ0V��zM񻜄D��uK��F��l�G{"�
>v����.U�϶���� �`Ͱ$
�*=���NM>W��+5��Z���ܞ]��Jq�*��l/Ѹ,o��P�w��3zI�n����(����z�:-���{p���8?��*v�1��~��3-U��s��[��Il�^�T7�(��w��Bڲ�`�ϰK*4�C�8*Lg���Q�F�6�;�6���֭~���/(( z�o�*��{��o��o	;���&���	��� ���5m�^T��*��F!�W��"�c�C�G�al���!E�T�/^�._K87�v�7���c7�^��y�4�xg��K��&��K�D �fP���x{ ���k��N˙T>U��ǒFPV�8N�,4���� ��q�5�y3�v,�Mݺ�'����e�a�}�鈒�cIy#B�c�U�Q�f(6S��DnFzz7S$_��Z1�\��`P�z�?:�Rd$b���Q]*xV8���oO�kP�ed��s5�tc�qM����q�ktT�q�@��ڑ�m�L�G�3�g�lڦ�\j���}G	�TE�xF!�H��h$�*h��PK�Eշ:�M�aH��YʞFl��_玳�r�Q�!��=P+L}�P�i�fp���Ͷ<O�֠�h��=��(W���"�b�{�	쓡��x��@�LC����s������S���ot�'��Q����t��U3~N�
u�em(n�2]��G&S̮��α#�t����l7�8��i\�647�o,�ч҄�s�m��t�X=�X;f(��4[���qo?'U�P�e<��
������=�$��8x��Kd����z��y��u   �*"��C�ҥ��[��b��Dq�֙�/�K� �X"1�i|٥�m~<E��;���6��bz�hZOk��o����F��j��	�5�?�3"��a����4Q�ʣ
v�s/��4W�<�a���g��N�N?�YWhlD|P:�ϡ�J$��.u�\����1�[ �I�^�{H�h��ec&c.9�=�6O%W�&7�(�$k��X���B�o�M��=\��U�eQ������CL�Oq3�R<Ed���ٮ�����H��Z�ú
��]ǳ�}9�4�%��y;������5k E[�d�B �P��/�����/�8�4�ࢂ�0$�j!��#-g�k�F-��߲���*#dU�3�g�2ކ�i;D�֕b��aX��ؑۘ���~;5�d%��tp��L<u�r���I"t��+��K��_OY��A&/yZ "k��w�>5�d�z^�3�wI����ʳ�q�A|��8�B��J�%�s��|,D�X��-�Y6,SP�7ϩh�>TE������EE����0?Z�������O���}�� Z������`�Z�f�B��K�c6�a	6Gl��m&��K �������G���y^g*R:����`{>����7�t���v��R�FK���]���ņ����I|(����?�Lf�#D7�zaSټ�I���V�'���+������/�[��4h0�/�O		���-�l��1����1��p���g��P.�Eٝ������o�щ�}��z���yJ��J�?�n{�a�K��L��y�Y+��R�9�"�"��m�=��/�_�"t����J�X{hd�_ $a�0��g��x)��)v����a�Uh~���If��K�g��m���4�n@ ?�I'Ċ7� �ՠ�!�d�g`��bQE-q]_�!��Km��̓��m	%rD]�D\F�d�V��	ౝ���s��7t���OU��5rژ������⑿���Δ�����0�\!q5z��IkuB)�A99��nN wkR�iD*�:��	���z�[n�<�hϼ��
�[o`�2�֒�!�_dZ���Y�XD��Y�p��e����X 4I�.Y�^�Bq�nOW�b�*m�'̟��)����~R�2���*b�o��XL.0n'���;�62�$	���E��[�xK�+xj�~#c�ᐶ��Lh��qÞ���m}#�vӶ�k掊�S"�M��X��D�ouH��l�_eT]�m��<��0�^���0��\����4W�ӜG������O��+�O�l`�5��3�޾�-�i����Ο]�ٸ��DX��ѫL��w#|(z��<iHѽl����a�TIA�XlHg�c�n���m��L��#�ϖ�9��߃�9�Å�Sm�m��T�n���뼬,2��t~�X�d����U6���$��}<�Ns������%&�qƨ��.����Ro��RM�+�ܳ	��8��:�8�=u���A0v��S	d���!��*v��d6�K��o{�)��m����B��S�=_�:=�y����y���M|.�Ҝh��2�I@����\�S[��2iD�{�r�a�^YZR��$�"r1��5D~U���#��pXj�-��q9I���l0�	��'�T"�`���t~�3V���/�̭�=�0���ל�_&\:f�j'	�>Cr�p�cr��wN��w�dM�E-�5c�UD�d���{��j�a^� ��L��o��h�K�L�UH"��@��7��$6�� �ǺM監4B�*�4:�5��z���i����0�;���V��^~��m>nE��ZħC�۾Mp=h�Ũ�iޭ�P�K�h�.���Q;�{�F126e��
��A�R�d$��58����3Si�y��N�'��!��������A1��&��z[q'WeY�F�²>D�pp`Xs݉T��\�����LY�ԢT�È��۱�GQj2| �˭5B���yn�/��:R�~V�Zb��fQ	��ŏzd��Z�=�1O��tL�Z{���>��P�X�=�,�j��o��Ρ&Z����Jj�#'���D�Atv�t�i��m���g�+D�s���9��Y6$5@���T�.'}�o�]��n6�ط�?#'bE�g"p*0�A�zI�$�z=�F ���SVEY��Ԝ�ˬ�k<�������,�Y��x�x�l���M��6�Y9����T���-Jj������5�k� �q�D~I!�D��72�eb�R��$C���%c��c"��'TK� Tkq,A�6Ʊ����X��Nz�^x�[X �#V���H�:��ɵ���c�����f%���>/�ͨ��+�I�%Zj�Тj��<�@��PVY~�P��
�^rXs�X���+��>�/�RݗF?�e�,*�s�9^��wkD �xn�[;xb��!���׀.t�s��|Y�p\�����m��~I��p�n{!+ �kW<�F&�\^UF%2�:f.�\$�֙7��?���'���$�k] m�Xi!��Q�vAG��\��dG�<)��3=t�	M.���������0��}|��Y�+���ǥj��j� $d"��O��G��Oq@�&M!A����b���c܂�3����g��ó�Ǥ��dL1�	��N'��[���i�F쉎�������[F��SP�'����`�y^�|$��6u\P3q24δA��z�������P�S��7�Ay�k2�B�h�ι�������S��oQ^�PdNY��q��$��
�.[����:x�`��j�B��Z���5�#�}�>L�].�=��O��VwY������.f|�Qg�e��Q_ʯ�D��4�B&���0ĭ��@V���7�4��g	r��kAtC
=w+Z<���@�UBO�%�]fy�bQi�-з10�Y��4�t۝����"� ���f�G��T>
��ӓ���dɁÀK7@!%m:T"�,v'�k���J��*�g���2i۳�q[�C��RLmh���~�ڋ���vf�ҪID���d� k�������H�iKČb�+�p(T��k,
�[��1��+��"�m����D�ڀ�bI3���j���=��&�)���_m���n���p�fBY�����L���򩢋c՚�xX^���v����Ie�
�L�p��u�UO���;�D2l��c�����&����|Rˆ^�����lɵ�,z�}Ȧs)�a��3j[3I$Ԑ_j݁&����9�Wř�}��GYxb�0�����V���)��7�G߆�b�Ĳ3�
D��q�e��:�kf�u�u�z��'������#�h��Ҕ�"�7�������R�lz`i��G�t,�ǣ}a�[�y��t��g�����������:LsjB�:i�Ngy����#F8<����]�-�=�/��^�}aݣ=��4MLS|<6a��QQ���`�â�)m5Թ�� �ܗl�t��r�(�h<�YT���o[#7CP�	�C%W�N
;��ĝ�z2(�W;5we��i��5���.�Z$[e�f�{�i՘˻��m����C^̐pK}�
H�j��� �Zq�G�	݇	�����Au�$��M9�]��K���x�ea:����:�6��*T"B���?�_]A]:Y-/��f�*�����;0f�4m��m۶m۶m۶1�Ķ�+�ض'��{���������]]�����N�>-U�~����߽�~�F/���$!�=n�hR&���>`�u�@|ǹZ3 e���}!܂�Ņ�*����q��,BI(��ez"�D�f'|z����X�U�p}��q7��I&���$e�pcAH��^��u�����^/��m����ݍ�~��}��uF�B��j��B�vP%�4�+�pRe��3�W8ü�������q�j�8r;v�~�)@��+D�5����8��Cy�xS��qB��n�#�]�pF��C���\��X,(�^�|5�PĶJh4D��/<��@X��Tga�,�HI��6*�e�:r�,�mZ8�w���aD���~�sF<ʄ1���z"9��NE�^��+�#**=�!ϩl�Hi[�j�pk�����p.��9&{��,<���1)SA-���-�O�\0۷=6�ҺP� �V�ɭGPc���:��U��gX�3qc�/�~	]�pR���.~e=E�KZ����=<�@Vp�Dq�S��l.�����G����>��ypMwh�J0���Hez�m�ӕ�S2�|0��oɔ�#NK��"���Y���IV��X���!ۯ�#�H®SƘ6Y�4MK�[rJ�e,cdD�3�Mh��V�Y���R;T�� ��E���Ql�4?����hZ9�E�rZ^E��� t��}�g�"�=.�EX��|{���pv��G�;���gN��q�E�Un	�PXƞ��~a\<v5H�������{/#��/5��=��)V�b΂�{�=���햀����cƖY���0G�*�0��A��yɧ_Ƿ�:�2�{�+�~H��*+z��u�_WW׷.�i̮���q/#$z[�`�n�s��2�1�p|o���X�l��J+u^P��+���6s:n�tţfZN�R�!�m��������x�`��cˡ��Lh���k2��.뉣/*�j�Z�`�g�G.Ճ˴�a�Ғ��z�~�񰀋�ND����b�ͥ;�t]�g�2Ը]��{X`���J�g��X pk�t �!V�g�=�H�oL�z
ɰ7������W��uth!�	�y����iD�߽ ��	�$���3p:�W9�~⮵#[���N����Im���GX�̃���~� e	�w��3�d6T�IL�v�ߓ�SӬ�T�5��)�F�qJ��F����ΠcL310SYG�����!By^{��{aBd������<��W����a�V.@*�]5�<�5��T�'�-{u�S�A9�(�Zf�rn0[�m�-�9|H=�;A�P�f��c�.��a?QyȾO(��:�@	A'S-7����La��w������ ɽޛ���r��8��l�p\)�n�:��X7�D��u D��c8�@;�y>�^�:� ���΋_���z��'�T5�����C�A<!+�*5��;5q{u���4w����<��������m�k؋���.�����LH���7!F����~��e� "���9��]C�7,�ݫ����k�\�0�k�Q^^��4��k	ֶ!Ε��ب�uL%i��)��XA�01�A.�L� �%��E���0%�L���_���T+�]z�.�E��↧�/�xY�7�xe�I9��۝�L/��β�0���2D��/jT��#fm�mDo a�y�ʟ�����L�����J��-U�}ҩ󏫆���&��vu}o6����~��6]�z����z"ܖ@5[��5���M�<ϰ-E���4 D��Ď̓����-�1����'���ޖ�cs6�Y�{FO��a�1�s�S�V?��L�̲aaH'V,Xױ�=�c��cڔ��	�`=�mN�l����z^�{]DM H4D�	��r"*+� *�-�n`�zp�iX��6��s�?�jAbJ�:��ce�i�	���K�N�D�0�׺eu9�ǌ��;�0w�����5��O������Y���(�թ�wST20㰶�m9j��
�����7["!s�FNa��rh�����U^"��[�����E�E���0G$������btG��� d�.�f)�W� ���XB0 ���|ex.�|��#�ɮ�)~�؋�P
�1B�;�P���4`xV4n��O�*�*��>b��:����`l�n�7d�=WH5/�y8�ҋ@�p0ځ�,U��N\�a�U2��uwr5�3%�3��;�?���Y���b���*K��ӹCbɴ$U2�����uGZxh�Z�*�*�PvVC��K�n��RٺՍ%�eo�&���J���X0�V��r��Z>�
8(×!���).���$g\���=.e T������jd$(F�e����gG�WQ�����-W<J���;��l: �+�[�Vm�@@1�^�"�
]����`�~��^h8)]�O�`�����e;�3J�g�-�a�>H���{Ϭ�$n>�OI�~NQ��#��`����N�VN�3������B�|��q�Q�)z���z�ȢLy�E�&������1�9bO������6��f�u�}�{?ϼ	�\�����ƑS��jF'3��Gnm"T���Õ�����ߛR�!��s�����/��Q��j#�u[C�4 \CC�����xDwPw�"e�Q��L ��ٳ-c9+�rZ��>�ww�h��t'�@�o`!�_�]��lm�l�WRY~�2�ݬ��J��� (
$����$�	ƾ�b��=���9�6y �'�{�$�P�����\�V�V���w2�iW{fү����i����{B|ՙWݵEH�A�Q�<�(���υ�	X4i��b��V�7\H�M3V��&����O5���6�rnu�H%q���˔����ї���1+��A����@5�:��wZ�o���ʒ�r;MM0���^��9��{^�����8  $[| �t�5(v�l�,&n�&�%)���a�߻͸���;dxz��z�)	x���.V��*�øj�YgA0�}`�,�v���ƀ'�6�!� ��f���9��Z��~�;��,Ν�+4:�_6�e�������}�qDo#��82���wD���`�r�C$�>
��h. ��z����4���E+���|����+�2K*|�:u3�9�f���)�Z��1g�y&f��n��5�r&q�>_�f��5�W+RKE��u8o����{��Z��|I�P誙CkYV���mKF���(��1��`��ٿl�V�5g�xRs`�^L[ߓR���RyF)��Ie>U
��X�@ U�	i��x�bi��U��jQ�_M �g�-�?�5<7"6��.��W�D������2��a����p�7����ΐ�Ú��cu�WW�����{(lB�y�}U~F�k�բ0-�b7�o�H����`����@�
l3��pҗ��{iw8v��Akd�ް�9�q
\���D�ט6�e�'�t�UD<��RQ�[��G�-@�A�w�Ou4��;;�s����q}{[+�n�
�혂>O&�l�T���eK�_.W�^|��S՞�6������#��	e�
��9jd���z�k-t��M�L��5.�T�d�
�s��:�&lY�5v�$}E�U��C�ƨQ/��Q;|��{~Gy�������1068��]l۾�z(�d�j���uN_ӳfF�t�x�W�{ h9Tg]�	 '���C������m��.sL��������������j�/�D
�I��1l�Û�#?91�T�EqN	��05����jw�'`�BԎ��=�8i��慡��ÿ�Y���e�ղ�� ��WJ�$��)֋�ʒ�\�J�@"�B�J�خ�������cm8�1��N�_�
�z��Z{�;,�sc-���Н�J��1c��`Y�!oa�׫��� $�Ү��u��_^�-����8���ޅ�\����"eh�J��)���ֹV�����q���׮�q���kt N�*���wʻ;����
<��dPҲ�l7 6�U�h���%��e6���^�q`��u���u6Р��u����2���BqT�Sޚ
:���o�pK���D��XӞ2�2��ئ�z��ap�;���	LoC0f-`u�e
 �
�����B��a�ɬ��V �A^�b�s����,|Ap�4f����s��O�/F]���`��5��Z/�L�+��cH�K�D�ݝD���!�-�5��t�-
�F
8p�%��>�����E�(p��?�l�#�+T/�AT��g��������98M���b��v�u��P$KF�>������ɩ����a	/�.�!���P̰�z�+�O��/8Y�>����K���D���ɇG#B���f����o}�ϧt�X܎���2e��>�y8ԟ�x��xgU�"� ) �/4�b��f��	������S���5)���*��Џ_��7����)���e䇫)Ji&ܒ�-��B��DƓa�����P[��温Dm/��m`^���G1���}qt�$ ��pX�6K�X��󈳠����03[����]����TP<�MvV�CK���Xm�T�����Dx��g�q�G,��c�g����z౟O��T�V�����`�+�Af�=N�
���k�����\"�C�i�}p^ʰWx��Z~4?��^�#V@��C4�������w� �x@lfƝid�����zm����2!�m�M	C���u���e7,N&����zd��oO�+���#��Z�1�lEU%(t�)�!_<��oy4i�(z�o��rYGFŃ�����&ewG��6�~��C�E<�~��I�Qx��<�Q��,݌�������O��cs�z���������/��w	=Gq`X�Ǻ�<%���Uh�7�=���jEG>^�e\����F�3H�B����<��;���d���%p�4>mh ���}��ylXWX'b��1�9�vpM�a�N�Q�E��4����2t��:1�2wD߇/��6.�;�)ː�������jb��dad� Q�U(yS�5�u*|X�n��~N^���p����<�{� ������M.nĽD����#˘������ϖ�$�� )��-$��t�տ�I��'��;3�7r"�;�7�CS�^�Y�y�2�k��;gI��t�`�:�.������/ݑ�Y	<�z8����Zu��>�M'�β;f�Cϰ����t�m�v���|Dt�	s�E�iܿ��_���=0���e�M���IJq���PÙ�s�M$'pᭈ�1�iY�'���E<[p��ϟY�	E�����bf�������?��	Z�t�T�3%��$��	�`�nn�,$�(���s��$��E�����;�Ԯr՗�z=w�4m�n�x��.�?�z;��ǎnCbh����Κ�-�+�#��""X��O�K�N�� '�w�jz��|N�`/�G���j���ƣ�������s�q�1�@`n!/qI�2�����:˸���|!��}'k	���(�`��˴3���NȄ_�Wֿ��aH.�
f�u��y�f�k�fgccc�m�~M�f�� ��:�N�	J��wf{��a?M=�1��$ ��FX�V�8� 	k�f@�/C�X���J^lkw+��UA�������(hkݬR1���mj���=��ӕS����+�i��hEmӡt�h4*���o<��=��_l��(k�2)m5����"j7=r��?��ذ��J�5Z���
=s43�Ƀ�adi6(�`�N���T}���?dׇ��O��[E��w�tNgP�Ѥ��/w���fJ1��?E����1ھ�n��6�E�^��%�|-�i	v��
]~Q��c������F�L'Q興��U ���r�:}\/�ݻ�L��'w{\�|~�R"����af�S1+��>�-wq���tN�<�b�ǝ�,,��N/�<��q�E�5���ec�4[='�v��~w](�*l���7v�����W��aV�^����:>歸u4E�E=˺��9��+
��}_�Jw}eHrӡog�(  �[-e��
u\�q�J*>�20�U�Ee�p�*�p��N�7>^,���:���Gۦ��=Gr%v�H����h�"տ�Q����wc�7�m���^V�T�w4C�pkjc��������
=?��6��.c�>�-ܽ��k��^�������tW��5�\{�w޻�[�P� �6]��gN"8�M������L}���gBhhe��0L��ߐ���c^^���g������!Z�V�PE�~S�Tq~.=h�܏z�i� U�6ԧ��g8�0mzM��t�q�lǘ��F�z:Um�9�^H(�����[���	�d�CQ�c��~�l���D
���%�y'tډ�)�A��,m����u��<�G��rZG�T|2�����x��;�A:> `5D�X�z���p��C��aVݥ5u�Ox��2 {X>����6He0Nc-c��/�N���c�Ͷ$������B-��@ES��H�������x(�Bf`C>��!��PD�@��L�=���+�e
����w��[�;b�u�%�
-�D�]ZR�W]�WuO�����M���k:x!��v0�{���2t�� �����{3yF�,׸!˾�Z�sf�5������u�f�l�!�M-;����h*�m�T��\'j(�2L2���r;ﻝ� @hZ�R5|��҂�������+:}:;�����A�l�m{�x��u9��Hm�x�F�?�8�,tΧR��?&�p	��ţ/��]�q��V4t��j��C��`&F�99���5��O�\&ǜ�zo���s�~A^o����{��������6�
�D!2�oI���d�I�����r�'ᇖ�azS��D~��s������b�N���2����j�"�\�����R4(��h�_�Ak����ʕ���<���G��E��,] �� h� B˰���A�����-���5[�+@�T/RH�E�N=�'k�>�u3��OЇv6�6�O�P���x�a��V�����b�YHjy�nK4>J�'�L9��D�n$ ����H�����>���
IGCM1M�����l�������ec��f�����2	�O�Y��TLHP+�mv�5�_b֗�(��{<&�3�A_r�9%H?�~��	 �9?�--�`X�15�ev�#N�R��`�s�.�k��������=�{�Z��Ss�;`&�W�-/�EeB�z�U6��%�l2{�GL]��-"lî���x����Umv�1�hݲp�a4����M#���grcK&���&Y�M�v�e �L:���ݽC!�m��m�G2�Y�gҝ��������K�Z���5%��t�.{�/���i��y*	;slm=5)xpJa�B�2~���D�B"�����W�|6f���fe;���Z7$�
h$>��w�*f$��<�Dwz;=~P���V��m���U
�<�]� �^���-��('��8P���c�^�����2�����q1Y!
���!�,	�t0�b�ɒԯm���g�d�?�̺����1V�Za�Yw����û�>g[|���1YH�y��;�F��a�M�/�h�@���,>\��1.�r�P���%���v��	6O����c�+Y���X��(/a�7���wBLǆH��\�{�@���S�ޖ�=ns��t�$-/�Gź!��R<��#�Gn����n�"|	�9ʹ��e��Ezܿ��cj�m48�����e��-(۝�Uu��1�!���h��:�ڭD�:x"�z:h%SCO�[��U���Je"sd>皩�ʺ��}Z�a����i�1���Zedw�]$�b�y����8(n�"�]+]"g�O^�� ��|d�dA�2���-�d�m�d4�y1�G�ƙ��y�/S�書;0q�$}�݋��WJ'ׯ�B�B����J�o��������[��%"8pX.�%��sn5ĭHݹ���2��v��U����"������|8:ϯޤp{�(F�6���C�������O�0/N�c0��g�^�D�!S��|kl�.b�g�_��mӆ���
��غ!H�˦�ޗE��>�V�EүJ�Y5X���z��� x�jU�6Q�
��Bo��$郴���֝��'`q���m:_{���<�z9+!_H�Ra����L��DKh�~s
L��S��ʑ�i5�JGGG��݇��`�tG�����:n��p8�0�$û���N������b]��2�=�'Pf�AA�hk�".�-��T�rA��!�< � �G�/�a�~���?�d3�&�����W�Jd˳cO���g;�r�	"�!S�+d�M�c1;�r��]�5|�&_����FV�\|���~�i�E[��1�}1��ڇ��,����>?��K��酣L�}�{������G+��F���R���Ҽ���؁�d ��u�窞��=�z�j�������l��A*�F���
�i4��׾��BT�6��[3,�����_�c��Vު��QeGV����jo�̀�k���E-g������A:���Q����
??+Itx~0�!��[���r
��4���m#K��7?���0,t_��I�>S�k0�l0�I�����%_���*��'�0>|=J女j�2�"�
sC��%Sa\!�&�QǺ��#����E�j:���et�9�#�zkɧ�'�(���c,��+��P�m�5�#�o{C�]iP���,��F�0g�x������ݚ�ON�mA"z-�Cm3���B"����B� g��U�m��[��
Ҍ�@J	�l���.��_�哽)H�\(<
P4����~��w�'�����w��Δ�l��<y��PQH��x��R�4�0��<��YT`eQ�4�	qYX�v��7�o��K�K�q)�YH�nն��ӝ��g4��IǞ��.w���<n?��m��)�$^�
�
ٴ�z����	��=�vz���G��|�Ǯ���V���s�k 2h0�k���q���B>����ۡ��&�28k+w�q� j�M���^ൻ^��t�D�=�`va5�F4�6~$���:`��3��a�[��|z�g�O���{"����,�+����&�!����9J-W���m���$���R(���-��^�q����	�56y�O�ofy��E.��(�J�����U�g��)i֫뷢m$g��<�,���Z�M�����6DU"\|�,P�?�}��G��x���S�g@������ܟ�GX�ڴ08� 4yC�Nbi7�N�T���[��i+������T���ɂ�^�zb'�<)٫�bz��1:�X�.�KN��Wͬӗ��q`E�N9�OÔ����7��d4g��.�q�?yc�>�N?�lW�0^�SB$\�5�i��Ի06����_���C�?��a|�*v��*>�@�Z�1Z�/�}�	V�E֤�����0I�s�)ˍ����t4-�?:A��IVA��N��F�yw5�-�? L��r3�vO���2���h�u8T��M��PO��J�Þ2�(��^?!�����T��t��������%E����3
��es���9����o�?�h}�zv�VtcJF�����--a�f�:��L��{�(�+3+����慍��p�����2�IuP�.��^Ii�M��G�@Vm-�k �iT���d��ߘp�i�m�G��=8�6L�ܶr�D�-|h���
�j�&@z���\5r��@{Yċ?�C�3��!�ǎ;��.�	�"�q
e����\�'�Y���帤���7>�9���0'������~�h��y�Ua������AiE1�Q6��+_{���u��y\�R���7��a�G����H!��y�����t@YT 6^FݠPF����眜����w~�l�QO�:TA���w�ݯ
RO'�mi�($C�<R����*�ۙE�kC-DEN#��5�}��0/����0 Υ>� qKT
@5�X���CN��P���S-��A=]Y�!�U�C�l.�5Yr

"�*6�ùTI_��t>�K����C"���2Q���/iz��Z��Ȑo�O�u�Λ��e������6�o}�]�3e�`�a[�"��!v=�s�(>m6?�s�>�:���S�������k�m�(מ��<���g�%i�����ur�s.�?d�E翗8'fE�|i��*|du�E��&ޣ�8,U�׮��#&����Q��c3FN��tȱ���qDB\���H*ޝ�)�Y�td*��\~��d���C��씈����&�vӪ�|d/~�F	Ʀk������c�K��.�5��]��ְ�0s�]�����x���n���-�3�Sk��d�nw`�"з�i%+6�'�B�	~n�]�H����ς�����⛶чYq�b�u���H�L�d�X#�L�]� cTB�~v<.�z�����B���MĒ!�R^��|�L*��$��Ԯ�&��[k?�W�F����Z����*�~��3��#i��;����[�@��H�p#��Bsr�D�������>�?N����MB�̐��Pw��Ÿf%2@���c���|�ύ��4�h�W)s{�l�h�%����b�%�X`b�m�RM��Ó�4�g~6��N	C�<Uv����_Gm/@i�H<��ÿa=YZO��hk�{8�a�Kr�¹�n&%��OVhWuj{{�V]ݪ���PP2��%��]>�5���s�h���
a�~���t��,���,�?�0��ٙ[�sN!���)L^tf�?ܠk#]���?�?:'zS�;��5�K�*h�����$��t���f�M[U��o2�Y)[�|> �<ͭ�y�������l} �����v];4Xs���)@��V�P8鋷��
.\�[�<�o��&��$��ZTg���.s�ʼwҚ^������)�I&�"��I��`�]���`��	�v]U�_����ē$NQ�i����m�3m��O���.2}V)r�u�y���ەgh��O D��x����x�D��8�FiU�2q�g�#��(���� ����2���Nh��tkK��<0�}\R�6��i�GS�r�T��/:"�2z�_u`�(�������$-�C�'�xx�s��A��Ὣ��b~�"}�����c/v ����o�G��`����@��v��� G��d% �&(�����'O$XK�eC��"��'ߝ��$lsS~=I*1.�ЛK(�\Q�&����>~�r&����33�"���?�Z��^K��p���s�O������O
@�Ŏ_2��Ax6�Ȳ�����U<���������:͉�%.���^���YF���o�'6�x����9N]�JsW����!K���N`�T�����Ȫx���AS׮����-�a�JO3��栛aQ~<��]�)1?\(�^r]�@F<�V1���x�}��q���F.�l�9N���_d�m�H�8?�uP�/S����<��QF7�=��J�0����/�B%��V��t޷.ަd�*�t*[�u�������_>j�-��yl��!w�C��95�
n9AV�d��M�\�.�V�.�� ��ή����z���J\�4R����#�W���
'jo;�݄+�p��ݔq^֢�n������_oz[V�9�;'�he���t�����I��ȉ,��<���6-�� NYIY�r�g��,(HT� �ċ�K	���Z!C��W~��q���c�H���W@;S({��ն?ﺿ�@���ɖ��bF���K���&S"�p;#湟[mo��D(T�O�>I�`���"�\5Ԃ���S7�B�v�7�'�ˣ;��^�K�w��"�۪0��.8�m�ſN�sh���he��(i}�؄����E$�P��7�w���nO�9c�؉SC��M�����%,:�\�?�+8!�>B�J�e^��6���u��[��(���M�\0�;��HaJ6�S�?ԯr�}�> �#YrY�.�����l����I���#�f�u��aN��������\�;�����<�M&肑&������h�����H+�O�?��B��T>�FNa�W-��dA�Ѯj8�}�e_�gFn�fw|���dre��p2%u����T�?�KN����E�	�0�.°`A���Z;���L��d)�;�R��ǯ����-x��w{�����g"=(���;���m�� �	g:�Ҭ�&�6!���s�Xi��,�!&�N�6���B��oI�6��>�1���Ӹ"��Z�N�힂�U�H�鹭˓�-ߣ�hԎ���>`��Q���o��#9�6�+���K�r�%bᕔ���*��}*B��� B�L2�t��ޠ�b�{�����ۚ3��s�ʴ�|�_������-+L�L'i%��>�͌�ÄE��H�1����m���%2�4lg�z�w�C�?.(l�9��M�-q�~��=��qc|(����s'�̏zj��9����@D�S}V	1}´���v�Uw�{&\�Gb4z���eu��a�_*=�81>�A=��eH������s�}@���X��9T	�ן��hM��m�k'Q�@�o��:t4��o�P[(/P$�I�@�[�S	>�|�x|�H �7@L�����7	�
:�ѦY� ����dD�"0�R���O2Q�G:
���(�U�?�ȹ\�k���gE�g_D��?�s�-�g&����1�Q��t�>G9EӁO�Њ���ʫf�0��}��x�SO���)��X�������C��T��KaTY���+��-���Ǟtk�/n�B�8��7��266=Mμ/�N�`�5
�ε���5w�[��:u��r۟���53��C��F[�np|�D"=
Y$����~��;���D���v��T��8I�u��� aV	}(�;���5��p��>Dfz�ʙ���DXl�׬n��bv�۵#�p]z�S�"�U�3"Rw�k)��V��  �?�B��o����kT�j��5���Bz���A��͌v���}&}ppj8E�ؿ��C�_��b�z�UaQeI�)��V�0bhYx���Cq�h44������Q��!x1e�xx� �L���.㜬�8�x�HN�՗$%�ws/'��[�n4�s^՜��t	Z���NîC��z�w������M����m�-|�>R�x���r��h.�DP���\�Z�Ŀ��ܺ�����,�H|�Ɇl������*��o��o�E����΃�<�E����~��J鋖��0�BWA}��Z��,��eP豥��.@7,4@���ٶ��#�D�0BvȪ"w�(�1�Ju!��8��?Mz�����%��IPȴ?�˱5��l�#r�#\&q�	9��4*�f�j�2���~���ޡ�~�	?���x8�dM��z�J�ɸj�G�x����/�5ʠ��N��M��X>b�<0?��F�˷��b?�G$!!��(���s}���Q�0���1��9����{ֶF���o�a?顷]c*���IF��I
īM�0Ձ����̟�G?�Gn�;� 2:c:���6��?3��?� ��2W���!�4�P�����¸i�O��J&�%�IaG/�c�uwvsXzO��_W�]
?��\��`2��E8�Ҕ��m�}-�+{+;;1��q-�z��U����� &��׾�o�L�����Ŧ�w�'���}π��ď;���Ycol���}rj�Ma��]�鳒����bڬܹ�<ݒ`6.����7�o����@����d���I!>' G4'iL@��g��z�Q~��0�^Sf�lf>�զ�,Y�t�]�y���2����"q�!T���>"��iv�F`��#.�Xc�_�T%�[���UţI\lȰ��z�I���)�M x<���kf�ݸ���y����1;����}�N�b-�8�O~(e���$;a����t9v��wl`YE���O�p�Kq�`�B�b�Ǜo�}�׀J��g�B��#�e��b<����x���a�?|�x�fY-\�KK�������GrzZA���ĕZ!��ƴ����(߈<�r�Uqv�&j8�O���4^��\A���������0���M�A�,�.|X��p���U1Q廉:�y�̪���-B-��x��g+HO�K'c�����l��eO�x��Z0��� 2+���g�0��WF���-w��ۛ+ۀ�j&.rH>�Ն�|�b�AY�E��\�m�O\6'��[+�am�}G��ӫ3WA~�$��Jߔ	w�k���*��m���jD������b���j�%���j[����qzB�cH��Ȃ`埭���������&���K��׻r�LWN�tK�;�b%�04��9���\6)��id��@�V]��L��<�((��,L,�{�+�i���w�,�fS��+0��/�DT�B����Bi��B�����&���V����Oۃ	Lñms���4�ՓB�B;�<�B4�(�Gc=Y�_�&r��,�ե�i�w0#:�\uJg��B�{����`�	�(OE<����۩%��)pb����^�\���f��j�)]!��Iژ�'na��;іd$�R�i�����r�m��h8!�5�?��5m��� `�k'��o&m�7%<̦&����V����hڔ8�\�^r{�_:OF]+X+32�:�8lH�s��nטvMq�x/��sZ�f�a�vlCK����?LlX����.]�������C[�q���
I��GL��ܓ���\�Z�i[e���@Ivj��--�N�鬜�C�X Z֮�k|T�j�^�.f���)���q�A����R���L���2D>��51���\i���Y�DߤH)���*%]<���>������Ncm�խ7(��Cl�!h٘V����D/��:r��5&v��;6I��9x�UuW[n���r��Yz��݇^�։l����N(����{�5����H濲��߁�B1QX�`��/`��
C������[���g���%B�����G:=��c��l�X'a����ZebDHD~�6��� ԛf�����&s�^ɣ�F�5�l�减!@�6&AT@ZD�\��(J
�<�.I��,����k'���w����)��p ��-���C�lm�n"�nxؑ�t�*
2v]�T��4�̄�N��f���p#?�E�K	�ix9J���G�G%]�mӈ2�~?�^ }Z��,_����q'��/a���RM�>�~~�eg�g��):
!N�UR�YN1�P�đ۱�ަ�
ʅ���>�Y��[��3��oJ����&����m�P�.�ꇬ<�jhi+RgVh�!.�yq�(��6�G4�X�q�Ԥq�0�m��fzl��8�p���\#� >�y�n*�׫>+y8�O+��>;�mb�I��>�ϚXEA�^]�y��۷��pJ�9����q^z%��$��%5nϮy�T[(�Є��C}�ҦZ�Xe2��M�,�tu�{tAq[�a@��~�rbr/#]"��^�ٲV)w����*2��MN���.VR:����)ݯ��{{�Q��R���������klL�˨����Ҋ|�I������B�s\S�J&k�=�T�]4?����FŅ�}�Dc(�lA�1R���9x�͕��1�ᴮi2�#����R���Nф����O��--������W��.��^�@���#����� B.���t�#;���k�?Z��o�W~�vwclx��dY'T�Te\XK�������i�Y�:�]@�I5�9�жA^�W Z�UX�Wi��$��B���� ����8�T�k�L4�)��8�ŭ�?�����	���
6U�9\?�C�Q��3���z!H=ZNK��g(*B]�:@FH���k��H�s!����#X��VBr^+��@��:Q+��fn�K�VU�I���^Tg:�����i�'G?��,Wߝ�b�N2ߕ0�Q�t�lx�q�Z����D�*��8�o)�Y'��2r���M� ګ�uk�7J�1�Ae���E�lKj�.&�,/�OC4F���y.����;��uO/+��0�/X�	��4�yX�Mڑ7 �:n9^q��2P��D��'T�^� R�����y-%� �-�h�Z$'%.�D��.]�d]��[yy��.���,=��a\<X|�플_+0�<}�i�������� J�!�\�eeޝ��y���)e5<_���l!a�F�m�­5К�@�^�C�)�l��;�R���;Zf���Q�O�#�.뚀���?����f�j������ 곁?��T�AG��p�?#�.�%����>@��������1R�Q��!l�)��Iƾ���ĸA����ͺ��ٓ�ev�+���M]Ӭ�C\�$��5l?y���ɮh]S>L��#~퀾-������*N��>Z49@XN�ir;f��0"�Gu�Wt>�����<_B�,��1�k#���6R���k"L�d����ox�YZ��D=7\�/D�/>�8v�G�n���6�>u,��fڑ�3��z�x˴�g4���8vw�{��"Ɨa:ר�v�.v��&p��D��"��&fW�`dIU����I�ÈDKUnm��v]4�~*����([z�tJ�Q��@� ꖡ��8�0NCW9b|��j���T���@`��Ҕණ�;�g�W?�6�2q��ov�9pl����x���4FCuJ��#?�)��ưOk�͛Vq�
�)羒(H�;h�찰��a��V�˅�Xh�$xS+�#xZ}3̱��#MRD�ױ��(���z5z�����˯�;��"��7oX��=��1b�u�ҿ>��4�s=�7�hAE�g�!LÂ��U
�oNi⨑�M�ؾ:3G6�lC�AF߃�&�B%�y���`༖�b�-���,N������C�Ԙ�p�c;
!��,�p�ݩ��R���%�����U*���^9jA-7'�����_��}�"B|���N����.:�����Gs�5?`��%�smZ�R~N�D�a��6�}w� �>�9�r$����4rX�r���]��Z�v-��UU= ��l�D4�b$Jd� p���>	��eQ��i�u]���ĔѮN���39gQ�r�l�E�F9���/�ò@��?Ώe��V�E�hyZ����]W�KFݏ�oM� |��߫���g��i��X���I=w��֘Ll7�b�1<�19�	9;:�g��6�B��M��6���)8:�I��/%aQ�u:X̳iEA��h\��M�2I����
o7�;m�6�`w�-h�F*d]�	���'�+
�!�2�օz���Ӽye[�E��l����9�C˃�*^��`�x�m^���!�ׂ�־��=�E늙sԉ��SBb=���s;��C�2Q^�:l4u��ͱ��Г�UF���,s�\��.a���H*��
�qDk�Ǜ[	�~<�E�ָ�&�|�%�>J/�iW�Pd~5f4��韶M^���%�,�،LUV��B$���?l��&�퇛�އ_����7���p86���ׄ�o���	֗F���ށ6���ؑب�U�	9W��̺(W��AW'��G����K1t.�9��*��B��Q;��$�s�"�"�&v�,�J�"������sp�1;��Sq٨�!_7?�{+|�5��*U�&LϠ[L��f=�s���#W?��p���W��Ϣ�����{ʡ�l�uVGj��G����6�X�aN���Ba�b�C��'��M,x�kx��M6��7Pm�E�Mv���`<��d�x�9��V�,��Cw��#�A��X�R�WJ%t�rx�jmH�^�՘J{#ћr������9Kk@h�8W�W�o�vD�~��p�E���s�T���Y���3�\�B���v�iF��:�Mn�������?�CX�0�}�y���S�e�\
��%��s�3Q�JjS���j��8m���h��˟BX("Ŀ|4��Ig�v��k�9W��u��ж)����Y�ZÀ�8:j�ڹ��#p��nP��·;I���G�� �a��m/�!91���/�"˅�b�G���8�ф\TO�/�<V),��:�s�}O���O�*�V���ɊU4DA�����|��e 5��D�O*L��L� ��y8"	�s�~��^�$�y���s����1t�f�꼻����'��vO�4x�:eVݻ�����F��y��E4��N�8��Hb=R�5���tC�&a��AUO��C-S'w��:��x��BD�sN�0mKE�p	a�j�n!Hc4��j����`�i�հʠ�8����*����(���8�.�V��J^�e�P"�ĉ�|2���h.R�ddO><�Vt-#W��:#�:�x皠��I0p�Ǝ�s���&\����rq��'�;�Dte��+��!3i}"��sX���9���v��V��\"I�82��s@�݄$��B}�v�Q(Hi=�>d+q���L���ﺔ^2R-w����p���1��{~���)X�J��BXr\� ? ����U��䶠F�gSc�_�=���_r�-Î҅���Y�	Z�Th����-r>�J권z�x�����ޒ���� �nd���(|
�r�T�U̙7m�UDa����N4HD�$܋��B4x%*K��k}&9K��ng��� 1���E!
s���a��d�~1�T#xn��V�q����\��zSQ��R��8���D�BZV��^B-!;0�>ۃA¡�D��7�Uǩ�����}^��M�\mvqǉ�~��涢��]�tgb�M۱��XD�^-hh(�s�+[��g�|ڞ��`� �,�4�)|�D�]�v�_��x���W��a������_�q�l^	K�{y0]{��1��E�7@�l#%[��f��@Eq�C����2���c��B�C"�l˶Q������^K��ҺRƼy�h/w�/@ǉ��T��nA�~�T�o�崞�q O'a�Jx�I�>vFj1���B��Osh����MQ���Q6>�v0N�í�D�e�����;cЊ%d>�5�Hh^֤ [���i�\0Wm�r�͛��ɯҘR��K!���Ày����sox��f\�C����Pq�0�'�Ј<JQ�k*�2���������~��^y_
l}K�����Ŋ}L��󙹨�19GB?���S��ih�S��0mWG�/k!�{ç��I\|8m&f̜�����g�M]t]>����-�t���a�k`�A}���~�㤞_KO���%�:�`a�'(�ա��\[>��*
��s��F#	�ۮ8��3>��K^��%ر�ީ�.:��,���j>�HP;�E��EX���&��Bb�PU�y����i��fVC	r���̙�0��xi���8C�S�k~IYs���n0�n8+��U�D���:&�m��FY�E�P&�Xѱ�F��痊� T!�����u-�-���/N�Aĸ�e8�j@��ʁp-�4�+�ӥ���y%בI��v�ZkT~���}��^14�s�N?���̹����x���xmrGT����6dѧ��p6�`uЂ�+�R�j}qIpǑߪ	o*��h!��	�N��к���h��Xep#���p��Q�8�o���fĚ4�GT	Q�[4 8�!�-���zj�B�B���[n�)��/��s ��_��%��k����q���*y^X��賰��+��٨Tj��J����eXܯ�2?�gG<��U����p�ؔ�0�L+�VyZ�^Ip�bfX��$*�^'��C�G99�%L�p6&O��kn{Z�f-�O��Bɭ�_�<������v^�[��<�i 	��4�q���������U���m�<ٌ�Gn�(d��t�~μ�VL��*>��uK���Ht��e�	Pt��ɉW-���o����ָ�������Un?6m��3e*F��uZ�[.�_�[�^�҄�Ս5��?������Xs�!��CJ�s�]G�'�*��~� ��XS�k���q�f9F��7]y$~v�u�D�K���q�i���l��5b�4>��I�Ҽ���Z_l�v�Uc��\�v�)m$��$������w>�ݏ�E}�v1Y��Hs�q���Y�Yï���2V�����z=��9�<�\�
J�C�=�HqP�R�^	z2�͸����Q��V"��������� �4� B��Tkmh(�G{{���e}���>�]�	P���/C���3��_a����� �!qn9�n�$���m��G��[0d�]$|�q�9��\�ˠE����v	~�)����q��n������_��M%r�3a��I<���Ud9W/�b4ݚ��h�O����
#uItT��g���x��K�[������G&�U瞸�[k(��|D1MG���H�pU\>%��tC�T�nJ�Rb��Of��.ん�ž,. �g�%�͝W��5\�3�KꄏT8G��-W���a@s�A��H�i�fk�,o�?���/|�i�c.���߅]�QA�ܿ�8h7��
�s�7���Y�(/ �ld�Vh�\�Va�i��ŵp��?�A��ElE�ʨ9��S�$A"�=4O�6O̡�P-��'���"Ӳz�Ĕ]TQ�ֆ�?ι��z_�����������8p�-����h���g�����z{AD�U�}���8��*I'��!��p�!8��[T(�����W�s���R=�Tf�FQm�����K�c��r4�� ����{�� ,"ėn:��Q�����?�
��4)��Ļ�5�_5r���>��!��Vh1q�A��U}R��o ^�.?���ԫ�jY�rX;�,*e$	l�	A�N�܄����I�<�p�L�����~տ;װ=��{���E��Շ�F�A7r�Y��z�z�;��rH-ș��-�T�������p��� |�^n��0��d�K뀎 �ILhd�����r�NO�#dY�"	�8k%g���
q�9A��B�x�<�y�M*��3�ŀ�6\�?!� a�9�Z
�6;�i�(&�qw�J%\s����i�dN�d07_�+�V�9��zZ��$�3��*��p�Aͅ�Ӹ#���蠒�a�{�8�ռ�u�/�����3�����C���CwE���F� ���1��E��?ǵUtX���a5���+�jhnvp�Y���ȁ�7��G���kD��U�H��	�i��#2�kh�33U�Hh%�~��������/6"ĻF�\�w?��8d@q#�x�ӠGI�*Ъԣ(�+
K�ONk��)	�-6^/M�qo���V"��EUG?rPT�[YG1�z�����Ri�*�ϙ3�U/�DkË�>��<�TW���n�V#�������vMe�\L'�Eõ���O�����Z5$;uH ���_p(�<�F�-,l/��qZJ���#CU�7�����-�lr�I�$-2��*<U3Z��?_�]��ƝsU�=O�s��~;m���ݘ���[I�$q��"S�h��m���pM�z��}p�E� �v����Ah����՝$�u�U�9\W#XEC9�q�#�r�������������Թ8���p��������cr纗��ުҵlÂ��cv3�P;y��59��:N����u��9B�z�(����-7]��N~,���gy�Xd��IV��7�a��JWs2=\��؈��
|x�y}�W�r�ޖ�F\�9�UDn@9)Y��{�K��q+�6my��7���w��Z}]�b�������&G�[�uV�U�o�W�)y�!���B_���Y����ݤ�B�����h�y�C<3�j\t�O��jP+��D�#��
\��P�i��j���$@rz���G�\#}ƅE����}6��~L�����i4�:lbn���A����c�8g�%̘5G�{���
��nl<�|l�t����܂j櫖L,��{>�dqğ���������&��H����2/_�I���-4�r�j�,���P���fo�s�VN��x�) Mm����c}��FZ^���wխOb�?CSK!��yj�`���!���V�S�lMUVOC��a����i�u��3oJ}��	�J8���(�ZǱT9�z��������IY�0mZ�I��i'�sÿPI�Q�!�u��m�K����N�[���$�ȩ1��F���J#�Tڛu����P3��5�$�͸��?G��/ҟ�k�[���V@R��i���|J�)�Ua���3R���,0�q��-[�˹�S.�;�9x{l��z�H�� �pB�+Ts��8!a�թ3��>Jf�
[�x�հ����k˪",�z��~�`&5h�I´Hs�����l���|�LvdZ��5��1\������b�f�s�Y������ [kA���I�z�r���N��{�	n"f͕n5���t����ƫ�J��2��2?E���U��j����h��dK�=1	����
E_��G�z~�>Xg���jm$ ]xܒ5	�y�j+2膥���0Gq�c�o�Ǟ~S�w�x���?��M¢�d�@�,�UX:��׸�,w��D�w�(�R��ڞxf"���C�R��!�t�s���m��U����̒�9��ZCCj�vh�a�1�aB��c�^�%�S𫃷��<a��Kҍ���CϊH�q�r��p�����-眂zS��k�����G����o{S?���%�5M-M�[)�Vj�� �U๽�z$ɳ q� L��x��� B\�_��]~����WB{�l�Q�f���BC�F�Dx���8�A5���&ি=�e1(��3�xG���4��jJ��I%�$�:��(!���|\|�8踫�^��	|��]HU�Ϳ�:�����=���X��4,)���n�Ǟ}����r�E���#���t1w�\�A��ň����^�.��aME��pv�(u&,x���л�k��������A98��%�%�y.���%G�æn�ϛt�]��M͆�!�t��m�i���.=�o�����1���a�rj�E��dU�DD1-ږ��GËc��շ�CX:��ÍP�RX������	;�:c:��d��U�5�����Ƨ�,ù���y� ���� �����l$����TlBf���Cw=8�������?�.!���߱���o�Ĩ�d3�j)�����2��<���r�n���xw>��eߛ���w�A��Ӷ��؄�V�<,��8�	�1��� �!�'�#\<�Q�s���Ek
�Q��z#	mn3Y���W��B�d?m�������Ij_V�����~}؎1|u��
��i�L�C"X����ǩOkk	�����qc���q�#���m�w�GJ~b�c̨�j2M�^�UU���q��;�X]R�&���u���$�~��A�ʈ_z����i3fOZig��}���y����w�\'�6j����=	�̆��8��`�_]�배�e��TT#3P�͇��Вzz��ķBC	�Jo��.��,�#��+S��r��O��%#@Q�P��+O,z	(ǀϡ�Z+lZ�K��< E�f��Kȭ�l/�n��jH�PA5�I���z���|%էV��!4y��ţO��;~y�8K�^8��$�|��y�:�S��ix��w%Hhn��\Ps�uW� �7�{{���FMjQM|Q!�Ɏ:��qU�_7Q��p�#O��祈�:�Op٨��#sl<|%��N␿�H6��ؠ�Њ��'�`���ָ���r0%,��|��_���r-�-��k"�H�K5IJ��-�J�	����hy���gN����{�e�P�Ad.=x}��g���]>t��g-IZ55���3*��n�İ��D�J�q�7[M��
���"{�Mx�c���W�B���^r�^(�r��Hr�i��H�gZ�=��A�mr�-T��<��^����������w1h�A�n�es�h-�����;�۱�E��&nv��s����J�d�7_r<?q���Y($�<F�ۈ4&	T3M辏�*bܛ㖿��\�!������>�1b�i�Mș�`Ҝ�gܺɡ��W护�B��/<��|+���嚳�א������X��=�kH�8O��}H�V���S1��)�UD!�_�8�����J/�� zFs 	��ʐ�U��M�:�5 �kЄ��贽��������p0��W�jcТy���7\�:���{�"�L��Z2�B~�@��Y4��od�E����jA���>��'�eS A�K�å����g����փV���A����0�NG�΁��������Ĺ�O�']0Z��%��� G{>l�C�8��8�A�i�J<�Zk*�ƘS�p�e�ay�+D�p�0�#�X���,FC���JYU�傀y���戹Hݏ2��ޙ	��CB��p����3Um�[ٞ�0�M�WH&�a��-�0_���9?�/}������aC�!�ˀS�a���ˍ���i	\��(z�1�e}�u�XQET�4���ɱw�*�ʵ8�*#an�s�JLEI;&}P��w?�\���g_|/����ѻ!�Ev��J�r=ZK޸����H�~���hV��p�N�Wmn�Eӱ�ZP�a��KNa*��F򋪴�Us�*�����/�K^�[;�%F���g�{����{�2�����zf�%Z�i��'��{頻!V_�7v�f|z��/U�~ -f�4������m�Q�P��(�-(5�m��}�(,�� ե�����A�]��p�)$g)KR$i�D��9f���%���ݰߑ�6O�pۥG¶S�| �ITXm�����Дn���f�ԋn\���^N��ݸ�cQ�jG����3���ކBҨq���q�eG���г������G�4���Tj@���[I<q6/o踰Uw��/�g��g�֏��M��H���لa�y"�?���iD�gp����g��ξ���������a�51t��t�c䙥��bуI:YW���}D�ڏ�p�J���ԟך����1��K>��%D�/}�)��;ힾw^���<8}iR�:�0�'�Γp	K�:)���o��?�
'��3Z!,>�_<x`3��F.���P�yg�D���i�-�RĦ�g�N��[�%����y �����j��ʌ��v<�o�%$�m�2�C4��j��B�\h$�`��+	�	]�i�X�]��0 g0AHs�i;���Ov{���O��{mK�)�˧M$�uOՀ�fVZ=wT!�B!�}-�B��b	��!�TQtm��$$B��m��j�
��ShEME_t�ٕ��c����[G	D�l&�?�t5���M�G@��,��q������q��۩N:F�)A�G�L�#M��"9"45�C[��8��r9��l�1g��(���%���Ed�~=���&N����ڃ����eTM	q��T�0���l�\7��E��T�i�&�c�9�!
E5r�t���K�@B���+z��sc\��e�B�W��?œ/��-F��4hS�ߖi�����%>�̣*=�㜓~����~�l�#|����@b4�%D6	qr�R�ʠ��ު�m^	�f��I���'w���ȳoaӑ�`�����%����-j	,��"��.���ʳ�1���g³�N: y�C7H�Ӛ��/��:�)WM�p]/�1���{l��͏��Y���4�/°�����]g��X�H�����G����?����!�"��Ƃ�KO�9]/Q5DC�ޣ=׹�]oI�H�tW�r�ķ�R��Wf��`��L�t<Y��t�.#B��%��3.=���]���VM���8�y2��Eۄ%$6ai1��(�9n��0��� R��Q��7\��EL�/��Xȳz
E��X�`�y �؄Q���]�+nz��hCh���T���sSS=O��	.�OP�5�#=�E���&0ԉK�W�i�j��'[�ł�]�E�lg^�p���<��{��'@����Z˸O��ۢV��G!Z������fY���bRrɁ'/�O�u�S��3�-��9�'�bO�F���ne-9��}`N?�@Z_Rh$��,�5�P�u�@�su�8�F��\�ń+��p������QC�W=�^�hlq�pME�A�N�D�����m��r<��KF����	xZ*���(�}��_|��7?���&��F�i�j������K�f�Z�BIC�x���N�']x�,h_ �(r��&�ջ��vZ�,�&�uy�����Z�x�#L�2�>����b���Q��������r��<!��2�`��Gb�=/A�yl5rU��<ph� E�F��Ӧi�����"�${I���2�7>��u����@�q²�omDH��vt��i!��du<��=�?{�h38��j���"��v�\�(h�pH��^O�4�[Z˄I31i�4_mED�
�o�e�(����]�>@�C��O�%����=�?��Z�[�Mu�F[�|�<d)G��\����*�LXrr�Q6��Q,μ��'!m��@�RC����)m�?���l�֚�[�
�b�wg~8WMg.9�]'&��Z@X���dH"kX�1�������Iձ��I�V��Vn#�M"T�����J�Q�pm������n{���[�~�źВ��D-�������u���&ݳ�͖k�/��,�=]3q��[�Ou4�sҮ���	8��q��L�<��BwK����]�����K�C�(s������ҬH*D�%4��Pp#�ώx����~�,س��v�">C��?�h�X�TA�Y��7J��)���ItGx�x�/`�?VsCL�(��k��m4�D&�����_�ߜs/�oY8��V:6�"�J�>�(4�>]����"�/��,,!	y=i�W�N������Mzu.t)!B��%���G�7��F��B\�dDj�,��U3�4�fN �D�%4�)�&����94SG��y�������� s��� �0t��� I`�ñ�c���1эû��q�����7����!�Ͻ�Fn��C�9��[2�s��8����<8NVlq0s~ ��P�sxEi� �a;b��6V�,@iЊ$Q����a�}�T��!ޚ�6X�zVo��6�[	,CٌnVItXh.�t��#�b�I�����ڑ;��BYFs��r�-�P�j�S���X���k��?�ԙ��
%D&���Mv3��-��N���	/6�+�&_&������믄����,�Q���}��\��P�]m%�a��胥��*�6���9]�qm����� ����ǟ�X@��b���K4ۧ�hlXb4j�%1��i;1$����A�Q,i�f�����9��̗������s�ٙ��e�����<�9�9�2�D��凭j�'���_��oyih��;BFĻ�`�x��[���(��/�B����u�a�<�#PVq��W�H���c��P_���9 K�>���.E6-��S_@L�P������_D�h��=���0i�I�k.1�l9�q��ći��F��rC<��[�P;X{h?����ǆ�L�B�r&�)�X_�����Sѓ�{��w?��J� �x-� x���/��Q(0|h̘9j[n�نB6��`k�䡕̄s_�k��IBD��)��gaH�M�^�RP,o9�e�x�(���D���w����+�!�:�{�c~E��Y8�tξd'���%�
y�,�x���W
`��8J-��)̠�OCF¿sdD�����>8����{`u_3Ir~@�Q W��9÷��h2��0-��۱4�Zې�������߄���o�	����N���3���<n{h
z6�;s�6�ЧQ�������d�N��CWM$Q��w�
���T�`�=�&*��bg"ԄG�$2��s����0�c�t<;�#���]`��B����⣝b����EF�kr��I���X�PI�-yq�j�,k���?����Ǧᠽ�A(�<��E0,*F�G�!���� �cb�Qឿ��+�����ׇ°<��A��"J�2�8��u��'�C�zHh�ꆎ��1�e�w��,�}62|�Ȉ��.�{�/�<9��~6�D��K~�(X�$;`ZUȾ{ՐA�����r�T���k������ޖ�0�����Tʊ��I�W&�>_T�����i�F���aa��<����)�i���`Q0E�.�N�kL3Gl0F�Q@�ˑ.�b�u�*��A�BSޜY5N��?�5���G>_A�R���4E����Y-�#(��T�ѷ���>i,�'�>t]��Ę�?�S�"���x�WX{�`b�8�z��V(t�8v�D���I�L��w����F�L-ܙ�7x��O�!	ۡ�6�|oœL��y��j�|���}��V*��$;ml,���f����]6�Uz��Ȳ�]���X2{^�^�`�]�2��S.�LU(~Zs��[�P5�a ��a�-�"ؖ!Bҫ���Cq�e"smd���{��!�h� ����r}:g>j�����/��V�1Mx����S�T+�r��`a�8��M�]�	����t%���jI� pI)�65�Jz7֣������=��~���鋕Gs��t�.�PJ��#PO����	����#R��$Q�DF��H����_��Q�$�̜���|)2��|?�Ϫ�T�VbE�o��e��/je'��������*�(�FTh�ᢾ�A�V&����
xlkD���ۨ�m��Y���HXE���	o�4�.I_�]���`���v�KFl����ꬍu�p�*��+�8 4�8�R�W�����|΄\�4�<��!pꑻ��;_�y�뺼N�P �����$ᝣ�:?��苚�[�N��3�w���|έ��b�%��cgx�+�H�<�n̈x��wZ���Ô8���1)7�'W 2^B��7&O�� �^{�{��r�M�S2�r��J�^�d/y"�-���ѷW���0yN6��[�t�\i�z���6cN��&x��y�7�i�x�۴~�
�*�ߡ=�����/�X�Zۂ�L�q�NX{p��8���y"�����\SYM�*"Ѡ�T���x�`������E�Z߽����ӻةe��.BFĿ_�r��-��<�w��?.���9��YƗ��!}�r9��Y�-�:9[RC��Ců�su�-�l�����L���0�	�E
B�G�*�"[�2Ҁ)�Է�V�	��ͭh�'rt�PB�M<�,� ����"�����⭏�#C����*4"�Q� Jt��M-@�B���PC[[+�^Z;"K��V �|s�1o�7��wf>MՔc ����g_eD�0tp_9�D�
��
�l�"!�Xܐ[�-kF\CL�w�P;�}Ä���ۑ3x��8j���aˉ|pU�D���~��F�c��y��D�m��/ o�,�HX53���U�H"Ī.m��K�-%X���0s_�������}���.EFĿ,���W���[��ڻ��ݤ �HV&mƼ)�C�,G�^�@��]�v��
m49I>�:l�[Kxe�g5ۃջW=݋"""�/
2:�8������o�u<�琲�(����g\N1�jB��@�~��=Yb�:�,ڵۑ�vb9���/{��-A��z���I�;�i)1�п�������1x`�΀���w�n�c15^����kO��RiCN#"�x�mK�\���k��x>]!�*s����7�������ˇ56Â����^�}�� AQ�r�rE������{��i��{�޲�����ǯ��k��#6\�W�224�"���i��f?�aq�-�ɪ�g��uڏy�(P,`j����
�:=UX��R�/��!.�3?_Z�d|큽��*���t�J�
B�2�����E�BC���~�AD�I���iBO|�?�2�6�5���".<'�v@$##$
��kG�a֗m�~� ���Y���	�Ԙ��B�
6ڄG�������Tȳ�D8�*Z$�������k����9l�AfK�G��r����S��P��a�൷���$|��^8������Ss\�O�,��Ēj�1'�h��H�w��"��;�� 1��R�s��=D_�i[m�.DF�W(�Ǵ[�}r�'������t%1�<�8�i(r�a�d7�5rn^����Mp�)���3�&��j��7�d�B!O����SӖv
����Qk��0����5��7M~��d�t�K����N�����Ϝ�s=��f)��d�����"3�)�j��C��@���В�1;�#V&N����/����������a��}��Z��+T��~q  ��{F���� �)�;�(Q��7���$Z�o!�*5�Ȉ��/�%��7o�������r���m9�#^؆��X��P�AL�o۰�����J���)��鳍�4'���z�����x)���|̈́�Ʌ�4b�Tj�G�\�,W�EGۼ�y		8u�e�*��^�u2@���[��o�e��aP{���ˑ�V4E�&�v#�	�A��W�zd�����P�y�>����*U�K���/|pŇU��w�*�G�qby���9І��A��Yb��jCKJ��upyl^���:p��≯~1��fOFZ������[}�����M|y���	ԤW��jF�Uz�KE� (:}�NW,&d����b��W�M�B������#p��wה��C�h���C�bZ1�U�fpϐ���d����OWse��&����
����F:U���L��C�c&�(��xy�H�R_xg������
�ZAZQŶa�ZHm$!_��+*�dFܯ�
�����C�T�P���ȷ9�F-�W�5��k���}��"�D��fpr*��R&����������H������^�(�y�ʿ=��³�['ƒ!y�T�e�6f�ͧ�-��P2|{�hEW�CC��Ҧc d�%�k&�i��_��_3;��R��+�^�t����d�'�L :��gI�.�D�?O]X�Օ�"f�,�K2����O��rV�E-����_�!���f�A��e-
ܐ��X(��f�K����	�IޠW[��{C��W?���}fR߽wq��(N+J&0i{�>IF�U ��*��%�x]�-��Cϗ�B��3�����\Mdƹ<�ga��]~%%�r0�q3q�x�t�nWTQ2d��,C,�Z%^����1eyz'�5��1���k��"i�O�?_��>�˵;���J��Γ�>����ÏM�����O���������fj������w����E��^��""�e�(	37ۥ�C#15��s�5��/���jo��jFF�W?��|��N}r�]�޵�6�/a �����lZE�D�}�!,˂�+�<q������;m���[���~=mm%r���~�� IIT)��
�h�����%���o�ז��'�����PhmmG���V����g�G,t���$�7�}�*�a��@��p|������ �<�"(Ԡ�%� ����Vt�������p�>�c�mG������~����1�+�13t�r[Y���?AO� ���{DFĻ*�������e�ky~y=MU�L�̭�G|U 8�K;��� ���f�Pun�R����:�a�A�cޒfL�6=�-e�	g�ih(����,���>^�~[k�,��D\H�7�'(=�62���2�m� �+g� �dv��XV�q�f���*�JG�zzP��F��Ғ�A�\�i��\^���8��uQ����6�Z�7�\��9�!�x�̅��O,�ź����Q?��H�t[๪]h��UH\�vg�u�cГ�G�_t��>h���}����t���fuk�X�#݌�dI���S�0��kϙ�7В�/� @�X�!Okg�E=����!�!~=f_,�f}�s�d�.\�@	a'�اk���={�@D��|���ڱ:��]oAIbZdWV%t?
� :��AA�����P��p	�[{0,�������i����("4"�J"��u��k�`�l��@;��lDdW�:��"��v��d�|��È��I����D�%ɲt���=��S{�ٹԖ��߄ب��5�"������4�{�Y.=�a�%��6�	g�3��/h�r�,��H��%�H���������vx�?[N�Bfl�����ks��i_x�b7BFĻd����{a�=��/�4�ITg��"��e��ڑ��eY�'<h�
d=�>��T�0M1m�����o��a'_+��{"/ik�(�o'x��m�鈮ۚ��_Oמ�� �t�~p�05YR)���b���60A3h?�� ��}ږ9Z2�@GO{:�6�����!��+�WO�}�I��1�2d�̞�6�`}�A$ER�-:#�#�Ⳳ�li��5Pk��Oo���i%D�����.c�c�89,"�s����8���S��^�X�Д��#ސX��G���x��W�~���92�6dD��A �~}�-}o����;�~��*:D� V@���n8΁�T�Ԍ�BA��ا���4�(�H��;�T����=2LX�\JG�Pp��+�W^ 	�������f�X{ؚ�K!켆6"W�,�M�bY���G��ϿF��������6���7�B�C���XST��5�g�P,%	���	�TΖ�
*fdD�V0�˅�w� ���g}6U�h�`?KdS��1h��%\���#2���!ha]֯1�Fh/�,D�cE��\1���c�	5>jO��k �&�h䶊����r,��;�_|�c�m����~��{������5���F��%�&EL��1q9�9�H��"��<܊�2�lSQA�Ѐ��=	G�z]���[<)��O�W8B99N�!��#7_���4��XgH�*�M �#����a7u�'�EJ�XdXK��C3xo��k�Z�ZU�D�uZ#q��`gǭ���7g�����v�b����IµA�N%��_m�e=�Xd��X��a��Ri���<�����8:�������&̜����.E�zrX��
���!�:6�EN�Pm�m=/S�$�αG�28I�H�dD�K%(�;"�h�� ���翽������g�W�a�"#�����p֒���]����C�H8q�����RaV$����4�#u2���4��gݲ��{�/)w]��-�}�w�;G�rC�*Rw)8v= o��ىkH
�`E��:C�B-���V����S`�a`@3�u�x� +��\=a�cᒌX�
��`U�D�	)t,'h�o�ʆ�u�h��x��x�ߕ�7��˳߼o�*�R��X���:���<b��_c��v躃�w�j�<��3^#���9�\l��0|2w�����ts�&�Vm�V�y��7o!�b�Q��Cs�P�=	L���(4jE$\��m���w%t3A���h��f��Ͼ����ůї�!kn]�Ȉx����:���������+��:��I"��T�6�4Q�x���~�ò5��E,�Y�>}���w��kN�1��=�5*x��9�f�5� `��/W�������k�ǉG=}��!m��r=D���@Q�ȷ&����8��Gk) jq�`��V���p	�M
�)<q�+%D�P`h*F���)��M������E�3Έ���˯�@���a9ZK��;��u+*��z$m�Xw���r+V��b�P�~@�[�C�x����uCKL96�c�wߟӣn	�w]u�<t �:�_��c>��ٺ��u�����؏�ʉ�O���s_�L��I�Վ��w_,�y�/���5�>���~�W.�i�8z�I�2|;p��6�F^�ƕ/֣yY+]�C�,W���p̙7��]�Ͼ8[l�x�����+g��q>g`����Oѓ�Y�u����R��;D�"�8���G�S��"0e�{�I�R���[�0q�<d;"��3�"k�9��}X�.W�Dd}�M�䫞]n;|P/4֥*زM��1ْϕ�x%����������x�m3��B���N]1����4#��V�s��5v�j8�/`?�<�|J�%�\�O{��2��Ԅ�=ƿ�_��k����Kq%����&'�2z�����`��KP�(�3λ�A��)��Rd�Ȉx���K,�<5y��{�Öy�P��-)<�yy�RV�d'��.*������'�R�g�	�-v��U WTq��18��[z���9�k��V����;�<p۱�&�a�����G�3|�GѲ�W�irv��w�u��DO0a�d�-���Lq�62{�&6���2V/�ˠ�:4��^;m�O�y�G˶�� g�bmyi�T|&"��-A~j�;��dGW5��&N�N[�n�1LS�1:ub!`�:|�c�7>��=w�l����v(I��+!���I��C��'3�>���=G􎫉�'���l�"C��*�F-ȇ|=D�.Wo�Z��m�_�t�¥�c�*�g%�����hf�_���-Gna�Q�Q�M7�8�e�󩪙�f�w��3+�,��C�cS���<4ۃN���i�?�ν��w�@�h�,4&m�m.+?�t"�m���c�M��lpO���u�� K�dWBW)x r�Yq��-8���q><|���Θ�𯱸5 �!T
�3��`p<�}A�'*�,��v9���RO.��u�����AX�T�"�=�L��O��6��۲`��0w~��F��zG[�5��!�5�U#���D�`�MBː$�p�<��f�7�`*�`j�!WD=��Ҧ��Wp�eG�hZ�n�r�VȘ\� �|�	�@Q�I��++,Kj�(<"������[�.(So���H3�=� �������1��7���/';��7���m��;0�����)�ԤXWS�:���18��[ ��W2�|���pҡ��u���PG�a�)=�@��豎��쎱����>^����B!�HW&�2���2{�Q ��|EL����T�*��g�V�������Zg��a"!;Q�W\I�`���c��>4����l/��dD��b�B9� PI�x*�s��p��x�շ�ؿ����a֜yXg�"S�k��J:�,���N�(@]��9�=�>z�J���{I�����"�xRg6�R�%l������4S�`��?�>�&�{f��]	]S(TQ��V*⬓m�����U*e/p�<���=Jo�R�����!#�ՁV��&_w��N>b���$\���m�Zі���w%¸�B#=�P.�B��ލ&�9�H���;��������؃v�f:`AM.��R�Jœ��N�S�^;o=&"��%��]v�D�����prf��md��Pf�ӆ�1��g�������;^���� �S5�D�YqA�u$��jF~��Fn��z g�ƝF'��x0�\J��D(B�`@��U��"n}�e�Dr��?��o��9\�����f5VM��+M�`�2ˀ��k���x$�l/�o=j�Ӱ�j"ף���a���q�2<��&�y�#T3�Z毗�~����)*2t���(��q�p���M��&�����&L"sd��l�j7DFī_N|�I���l�C�5����4tE0s�xx��OYh��^AC}������5q텇㗿��j�Ί/i.�O�:p�M]Ι,4�d�)T�Q0�෿��x���t�f�v��}7E�<4ႍI�@��H�D�%�6�KQ#��l̚�j^�ka�y���
"
|������DBCDa��b/��������Rg�'�K�O:bE��u°�~D�v����t���C�{�+>ܰ��*3�
��oCB�3Q5�%�c e�*���G�(�}���f������
�ӏٍ��3ܱ���!�]Uc�+B�v9��'��El+�[�Ρ�5����@,��o�B�xx�"���nr�c�D�UZ[�xx����e���Ƨ��_"C�DFī\N��c��������E�b(z��ѥ0�:���Bє�����q�y��K�R2�෗ݏ��>����k��&Jn�����6y�!\
$�6[O�z�{��K�B%֤����@C MW��)L\:�#6;V��d6��?@�	3������$�:i�E�I�&�X����14�P����v����:z
8�ݖ?�����B(1O���K	B����(&Ê4��6>���?�f
�g"�U�\�w�oĬ�`:Px�vE�w��<�6z
����)�ښ��D>o�b�M(���kȫ6*�/ۡν�^�jk�\s�Aִ�R�b�!d9~���mp�(��S�t�"D����x�yiIz&&�M�����L<��7����#�&5����3"ޕ�rK5� �*,�z��P5`��F\q�h�����Ѕ&h)��6���.XJ}E�rm�h�,eg�����NT;�<�����x��OB� �Kk#"XI�87E���ϱ��ݏOˈEM#��w��F1��/-(�����D�s�J;t`�cp��oA�����C�S��Wd?x�ƒ���#�)ڶ
?��'&�xw2�2���[�w�]`r��Bm:+q���=�TyBID�!�BQ��/<�Ǹh�U����rژ���*+ȋ@3,�'���ת�\J�!QĲ�����z���a�^}�D8�>h�T��z2�ѕ`�+�G�����xE׋A�:sF���K�-oٜ���B���3|����g��t1����e�K�����l.��Hx	y� ����f/\y��8��:2�������y��--m�su�,]�)P�T��	E+Ӧ��W��9�����TՆJ�����F`�͇�ko�i����J�L��I,ئ�2���ޞ��;h��]����O����lG�d�5W���H�'҃Q�au��T�p����תv�W��N�fN��� "reBc"A�3�\�·��	�d��A��7��;o�"����͖_���&d?<�=p��66�p0�s<<�-��Z�̀ߜ�7��ҡ��A>�s�(1Ӂ���D����;ը�{���폡k�*���2�D��A��L����2-
(5/A���R�����W?��L-��##p��k�~���m8l���=��B�.����B>��!��AQ#�C
6=�ZfʑVk�a��F㬋�:w���_�U-��P	8p"�>g�˭�l��S�������{n�G�0X�r�5�����vCTYJ�`^�����9r�J"O�'Q�QU	���)d�����7p�>#�ly˶~�����B.2���#�L��)>���ϘM�U��h���6�=w=�`�xQ��%��J!"T�/�1��A�����Ӑ!�[��6���-RS�ӱf���A3Uh\}�8�Ga��s0wᲪ�#a{9p����F�a�
�mm���^�oE(C3�TP�-���G5��s�оCa$.���vU�k"42*ޕ�X��`��J�]��WK�<���\�΂6�yh7GFī\���W=����Ϩ�o/�QQ�}4݁�ñM
���Ҍ���Ⱥ���"mRwD�r
#g�bT���b O���>\s�h�qIu���
9��1�c��L�E��T��m�3}*D�Q�@��z��p���ዯ�`��˪�\(�]�Eg��SFR"�QC�D�C߅i�8���)f�eV<��q«�Ha��n�w2�;lw��/�C�u*��0�%T��x�'ρ���#v��seV�Z��'شѝ����r"݇c��<}&7��AX���"_�q�Ƶw=�,���	^/M}{�64�#���0��o�D�\MV���EB��4���p�Y����i������C������'h��-	Q��-**��_��6T�{�X�����~}�Q���R %D�-�[&�3����>��;�x,�j�v�&�R���������z�1�V�߯�^�CFī����_9�7W����?�-�p���>�	9z����M�.�ʁE~�G��������#p�%w#�"���`޼v�������i�#��O�ª��(�����q���g�U��-�!����з���%Kѫ�3	90�<�0�>j"J*rΫ����{&!C�����O0z�=Q��^�r\��)���1�+%�9���@�(�*n��w���Ū�3db?Qq�O${��/(�uQ����8&"N��֊���t�}�ղ���gȐae�x�d��fS�q�9r�m��"��
r�<|�lS��b��.�ϻ��+�=QU�&����9�81����£�ܫ��dx�{C��u��ª�0���X�R]:Z�׻���1��d��]�����"��)�ǭ������"��/�����O��Y�����U2"^�h&�5��g�}��CU�e`§����l0!BS��ebn]	�z0��B�r;4GA�&W��S�u�2���AD'~s��x��s�+�hm[
�鍐'�s���k�r��R[�\���q�uO�Otۃ��yz��8
��QVѫ�*A3�ź|�B&�e�&\�)�r��ݘe�2��s�8�s�q�� Ǡh;���Z<���JR�d?�K8uw^}�;�V��趇WL*����Ǡ>��u[Q_$�T��|���H������% r��:���!+���`{9��[p+����]Ψj�����u�9֋��e0�hA����ʣ��3o���nj.r����ܓAA�%�l��#oX���XF��ި�C�Q�<x8�;�ƿ(�C��MkBOJ�̞.��h2�,���9�=q�$j�/{����e�J�֌U���W?f=�������{�M�-"�
"WQ5a��TTd$�k�3Q����6�4K�Ё���W�q�PDq�}O�g�:9h\p�D=N���\.Mr\QC>�oO��r�x~�G�n�{?�_�u(��H�J�Id�Ȓaip��׀IQ���#'tma|��b,m�!ÿBB���3�b�6�BDm�FD�w�E�\ZGZ(�k��=�5�㦫��������c_��-6�_��#��2<"�R��c�B�|=*e�XTL��F~&�t�^�2Gfh2&��_�����a�����0̢Tgb�����!נ����&7t�5'��?݇/�w��+&��n�.ƌ��l���iB�5g-�أ�i�Udu�*J�t��q��S���*�%��Qpͅ���"��	I3t�@2Iƙ��:$<f�?�6���O���4��2T2"^����W\���C~�Z��ػY������Y��x�TCCM���	O��eh<�,�t�@�F�^z$N�ݝ��D�ܳ��������bКy��$��x��צiȒZ>ɷ��ǮC���G�5��p��S)��.х��������Y�k����r g�#1d6�4��)G�hzH��O���c��'ÿE��w��6d��'!bD��B?���v�����\>���7'��ǿ��_�����w���tw�^+���b�(�|��$'I�,�4U"����D.���۟C7��2�F0�>��p�e' ���T�Vد�uE_7��'�}��c�;͈p��G��{^�s�}�m����m�~4
�hC�s�5�|���5G��u#�	�@Q�P[a8u�=w1�?�>��^R�I��`,��x�=gA��g�2(����w���3���t��W.���ӗ�CV�^uȈx�@m��|��w?x����-ٰή/�>{�*C�AcQ/
DC!��AWmz� �*t�Y���<g\tJ���d�E����]��OǣO�zD~Z���8o�IAF�u�Gq/yj���!����j��8������X=+g��N>j/��p�£߄�/*=n� /&�d�XE���r&}=����(���n�@��+2�6pi��݅�ǎA��!��8�t�P�j�UI1������7���]u���`�0\��Vs�"�.�Ձ�n?D���<+A{�+�^�\�<�+WxN�!�1JLvo��mN��NTO�O��>�<�q����=�Z29ۧ ��"��#�"~��'G�<�Dt�;r6\ ��<a����/ב������ލ��6���R9D}!�
ٹE,\���⯤:�X�P� ����X�{�I�Mc/=�f�Hyx�ͣ�NC�����HA$c0��l���Z����'�s�]dW|�ۂU����4S@����xb�S�گN+k�b$1��Ⱥx�<)��E1dY�'��=獓���4u���	���oAs[��cU^1'��&�z����8�#���|��'�p]7`�,�n󛑣�_��}m�z����I���d���y��{�۶�q�����
��Ce%t��e�&�e���:!�@YD�ځ?��l��d�"���$����v�/�'��OC�M�{,Lť�\���y���P���%l�a_<0������+!O�M�=G����#���=P�#�a¶uy}Q!J"�r�JDd#����s�L+G2{����xn����8l���,B�?�rl��ijp�e��$���X[o67��<^�:�{�Xb�r�n㈃w";ue�^g_9w�(�5�5U������0���$T�/λ�*yy�U�q��A�Y�"�_am�P������WP��d�oq�ű�e9�+(U�_�:~���	��«�9`kmy��O�����w9�N���u���it)�؅�;B��!����[�����cY����c������f��;0^;��qx��12�%R<W�ҙ�~����H,E]C9萮_��"q��8���1��xe�G]�sX��ƃp�{����Ѓ��ð
��`(�J�'��Gl6B���B��:c������+�Y��� �����8�]`�gu�2T�HDP�E��*�����mBd���q9��j��ѻ��v���<��f�������m7[�<bg��5�HD Ŵ�*6�1��^3X""UJ�-���-?�~��������7s!�{���&"���+ۺ4]��L�5g=��.�򘈮���(��S����o���L�����ſ���8�g?���P�
���F"E=YTĶb4�Yއ���OZ�>�e�6'�}�}�p�h��c�Ň"�7�׆�� f}����cF@{��M��R$b��#Ά���뢵�uћo}4��I��Qe</<���Y`C|�o�O����������]n}��I�´T�%���y8Z���� R,)f�����\��*݉R�O$�;��[�p�q8����{��p���קp��P��r�����y2Pt�AD�.��Y��ђ�\"�:r;���q��I���l|��݊�����6����$�YD����׃o>�.�%U1d��=�ߝ�3c��#2L�6}&��ob63<��o}~��h�]��5�� 
Ц��U��-Q�A�5� �m�셈G��ç�8���%8���ԣM�r��d/s��F�.Q��n��8��8�kh#&r�Dd�,tA�_��L�\ݦ=��p����f�>N���^������kZ47<4E���[mBk�#��&��<��$��!�ъ�T!G�1)���L_"�������'a��s���6��Woa�M~�cF�Ava�\B˹ٚŇd�ZB1�"kc��K�U��o���P��Ki���=���[Y�z�~��K���j��������Hx�ç�%��S9T?BR�J_,^��5��� �e:2^�Ȉx��Q���W?�p�5��E��w�,S� ��1�&�.H�o�$C�!U��y㬨�S�a������m�bA�38�����j��8��}Pp4$~3*-y�������ƀ�pS����5�����m�~v�8�';a��f<��T̚��T���D��%�U41|H?�6jSl2b
|"8�eV�� ɴ(H�)�K�� ¥�.$Rns&��I�ERZl!��/V,���'w�K�8[�o�z�7`�������SZ�E<L�|��޲,=QJ���141��DvcV�.�p�O��	GY���<��t̜� �[��z}r.�o��aC��ߞ[a�֔�ݖn�\U�*̵E�	���(c �P�=�*4���b���D<��r$÷��+�x�k�[E\��:h�!�+0"�e��T�5���0�ǁ �*�Ug�ģv�Ϗ�3?[�'����>_�e��_�N\z޿������}w���%3�,������w�xr Q%O��ף�U��kA�`�-���i�'|���qw�Ǵ����C�M9\v��PY�&km\�ȩE9�/$���0�5;l��_=�O�>L_~	�zdD�g��ۦ�������1�m�e��RWm,���/�nG�Xd�BHNBa撡�`�����*䩦f
d.;�H\{�x��y���`i껟c��q��C�mX��DDzQ�n!��>|
���A������U��������.��cz��������p|�e�m�p�R���+����0lP��x���]�>�۰!�v9nL4���q&/9�ͽ�@���ɫ�PtG:55��[�WMLx�=���䌄gXe0����S�tY;�>|ԫKP*��^"׎T����:�2�Ui͆�L"!Z�re4��2<l4���;}���^�5w�|w�Ehi-�cŤ�t��N�Mcc�� l��0l8����(����]��~��G�i?8ك/�T,2��m|xH��V`�k���˒�p�}���Wgf�#V�玽�E��Q�{��ґ_Dxy�dx�MG
���JDv��/e=�2��>�ub���c�!�X��´my����E��9�l�<���DdwI������E�3�/��t8��%&�U����-�p��=@1���U"Nլ�<$	�L
r�����ߔ��	�����̞���F��+��x(~w��p�et}v6ug5#�i�[�l�s�B��Ϲ�����2��܊U����\,�jIi�w<����;��m�o$*3b�a�A���C��\f��F"���9νɲ؎��c�����������j��ͤ������kO��'@�Q��#�$[�D�X)��%�,��K�G��2!��Bd����@AК{lB�&���L=��Q6in�@+r��b��w@㹚��ǐ%���0����\ѐ+���K��u�[DL(L�}W]7�ޙ��2|W`����1i�'������.���u=�IF��m����3��0T#�C7T)�h)g%�KvH]��=d�z��$�LL8��">L�y�,pڍ�w�ko)�'/�ܹ�\#ZD�W����"�7�'X�$��g���;Z�~5��>��ѧ�C���d���\�&��?�y�<�_^�~��3bI|5̀e�R�C ��y��K�~T"�E9�R�x=����\l2<���A�yS���X�_4I�c�E�ׅ$�L��op�P������o�K޹��'��<��`�l��Qa{�\�X��s7�a�	�U���8`���}UxT)g�-dX}�-�g"�V*I���|��y�Z'ӗ��6������x��Oدi�=v�x�D���S�M�ձ,����t5
yrʾ67�����]�ɹs��A{m��MM���纽��n�#O�W_����HR3Lǐ=�,P��l�zY��sa�:�����@u�xDR�&"�}���I:��R1(�&ܓ�`�D�yff,�q
���6�H�RО���U���֔D@
�ͭe4���m�.{/rp�/ǢZ�����Jn���v�^|�?����Ϧ`"`�L�<�C��m+'gu'qZ&�\*N�5�2��}�&ۖ�J�IH;
E��UNڀ��,qgb�廚��c�(�ǜ*V��� �
���P��a ����6�^R��9��5���ⴱ2;����?���N�3n��h4�LZ�6���1���W�Z\1��/b��C����#�!�/l"��-d��⦂���?��p�J(�?��I'��#dr�E�\�.�o���.�LӸ��%� �%����=G�T:�����%�u�mU�_��9fOl��`���U塆p_>2�F�(���#/j_���������EV��c��V����S�2���Fj	�QYDD�^ڛ�u�t)X֗*�&
jYuܱly��D<o�0j�A���`�s��n�rU�>�#����-�ۘ�@�
J(���T���Y16ȹ+R��T^�������d8��o�2�HU\vM�l��5d���t���}��Ll9�=6�$�:�{IVx��F��'���h-���,4W|<�k\��2O�����Q�<�f�z���a�u���ՔPD�S�[����\����nK�&�a;�I���X �!� �$��؋8oå�Ҧb�#�4u�w�dѤ��Gf�� �t��4)8�{+W��&�>y�Gw׋���}��P��=�سn�E�����0S?A�g��9���ds�ةgR"�R��<���b������_G�p�EF9��}���{���F�=D��
C�d�����N��Hrq5:�r9I��q��U�:x⹩���Q`�}��~���u�IH�c��]�h2D!*Ȱ�@�t\.�[��o�q��Sn��f��w�x�a�"#�=l��/����rr�N�Z.r��A0ӱT��/O�eƊ��Q`���ڴ(`�p����C�1��Ʃ�����7b���'��)�ᒳ���|��]C#�L[g�ܠ�R\A��DB�;��<�`�~� &��8��S�PГĨ�,a,���S*N+I~��~#H�~C��y=k��#@�D8X�Zs
coyo~�EF'2|��������3p���1)��U�%�ɹ�\Ӟl����DK�Z�aݰ��(r�0��$�g$(CM̎�6	�3)�H��B�$;0Q(����9�q%N��)�W�D���ˤa"GC���.�^yf}ޒ�K����.���jD?�}�R�-
��C3UZ穆C�1f}��GB��q��&g�sKG��n%�/��}ĉ������B��qƛ�g�\$�.��'[
��&��)����
6�m�	.�������j ߎ.=u��"����gyK���n�)dX�H<����^����mȉ�z2"^�0��u�Mk\w��u��l�e6|b�w��f�:�V^v�\�F�Ĺ�M$1TN��݁I���&�]}�>�ƪ��~��ǉ�\��w�#�:g�/���2#ĺ��cR��P��3"LB��@�\�|8�s�9��A����T`��C����Y��"��^0�"���R\��ʽ����]��/���7���.n~p"��l�gX=���%8�?c�������4�Zm�P�$�|�%3ކ"{X�0�����3Ua �]�k;u"��b{I�nuYg���U�xLe��iH�ؤ�N���3�����A�� �"���x�ɸ��7�LeX�]z�_��ƘCFa����u�η�6.�$]�z����rn��>qA�m��:ҿ0�}��xZ5��q��Τ\��*���u���EvV&�m�%�\��R�-�`XL��롗���"���$�ƫ�D}����O�Oa�=��e����CVx���u��]��l	�Ȉx�`�6�%�������3�pS��IH$ч���%R��q��^;R,%÷G$k�ى�������;|�6��%�b���ۯ<G�yC��t�̣/~��^�?9p[�Ƕ�����'���p�2ې�6��2M�F$"����L"4&�)9��s&�,��(T:Uf,��~�,����&�� u�fy��2a��
bM�����SO��-Ȑau���ާ�c��w¾��p:b��i鴦�.X|*�S�����+F�$�[�?QK����X�q*J�9r�R��d=�ӲsE��^�azeDDD"��؈'&������Hf�R��>�տ=0	O�2����[�C��.�uE��D ��Ƀ��KLݠeK>V�#C;ES��Ȳ�N����:J�=J�t�3����r)� �J���Z�t�b�����������:����\؛�q�I(濠kl�1��Gⴟ�&�qF»Q��r(�Uz�A1��OMt�Pι�5�&�[� C�DF�k�͞��W/��蔆��x�~!JM����R �<2~�Y���Д`�,2VI��2t8�fa3��=غ�Ƽ�;Ǟ�ν���q����M�}��}��A?��R��P0L%&]c�ʵ��L� 1YZ���g>�mS:zaUI8r�:�I���=�<���V�EZ�D�5GE *еzL��&Lz��-B5Td�-,jvq�����g������� �C�Q�尿��A�$���P�,J�c�%%��;�6�H���4��ZDD��G���D�U��#�E�
x�ix��X��I���ҵ��������k�w���˨MP�ڑWڥ��m��i<�ۑ�[���_x�����y�/�М���l�t�V�yB����#F����u��������QMEV9��͗���Q���~8��C1g���+�ዅB���xlڳ�?w�m62q��������������i���(�mp���=�|ʫ�90�HjRԧ�g%���*���,� �BD�N`R�p�'����Ƅ)����H@���'�ၧ�aב�c�-�b�u~ �؀(�dƛqT)XEA �f��"p�@,�e�B��h-��LpY��19�e����
XN����4��ܥx�x��7��RE�Q�w���]E���3s�+��N��J�@��""RD����'���"Ho�;R!�Fh!	���!H��ʭs盹�A��P)a����۽���;���9烖6���4ܦǁ{���QC0r��z�srh#UfaɁc[�����=��T�"��y�l^S!�G����[���U;�弨T=LQ,�������w,�ęs�'��ٻ��]�D�����o��+�8p�-�Ϙ�1�_$�D�T�~K��1�M��T����}aK拺EU�I�2�2������쑖^�A�	����K0��E��Ԝ|a�����#p��{��ڶVM.�PлSI㊾���^�Q�$��IK�k�4���Wק�JI�ѐ�}��m��t�ċ�:x��>��N*�^�ע&�k���'��~^���u%\m��Շ2Փ���|�X����4B��L�b�xԞ9bm\z�Y�>�_�L��j>�<��M1|X#��fS4�b�h����<���ݾ=u=��IlR��ȃ4
��h���F��>ﾻ�>�
*��+���D�nT�[?v�sxp"��!�l���4a��7��Sc�D��Y����τ�#�<����U��kO�գ(�B����`<��,,\Ԇ�����;=-Dwb� Ο�����h(���-���&l3jc�&�<Z�D��Zn_�(�G�y~L-�j��\f����.�<�2�;�L�;�ӊq�g�H��(��"�)ڏ�m���V�N_؞�o��/&�ש��^���a#�#Lxmޒ��/���+��s`:�=�#����o��+|��U��Ⱙ��Z��v
����Z�� V/��k�^�W.#��<�.I�s��7m�"2;n��+���B�D2�My�%��g���}vXÆ4a`�2��K�׷�����}�)�#z4J47W�lY+�C����`q3^xe-i��7ѣ�:2���Ky��	h,a�-���5����o��W?;,��{;fG�=�JU?+-hn�`q�\,z���}Z�q����!z�Nn�%���;�ޓ���l�6jD��"�4�g����c_</Ο����`yK�J5ż�V����u��NB�{n���yg�����
�7_��D�z�`@t��eX��sZ����GϜ���.�o�
��cM�
�N����W���<�!���-�W���"�.����V�$΋3%a f�q*�BC�<���wj��0\��o��s�n���'���n���#O�w���#P�(��*R���������7�C��Gb�	��=�UL�U�p���Ms�)�뺰���+��h��$2SP�T{7��MZ~ST��v&
��&m�j}E�3�<�����z� ��{$�{/�o֢h�/~s���:�O��ij|����a�)�_�p��+�Z��Y��T*�{�R	2�q�hŰA��c��K������{w�����տ�� z3��P��,�����߈�u�4�ӿ���8�y�j�� �/������$�6�$ީȰ���DH_����h|r}�Z��"H���o}�ޱ������m;^7�(|=qK��:F��$2��e��e���<�jj���?�e�j��l����?;��3{j.@�6AA�=�l����j^�k���<�B����H�\�����i�2E������G&�9iμeS��� z$�	�)<������l?j���{�Jyl���8K�ӣ�T������I����q�v\<߻����˻B�7���c�q���L��D*8���#��q���AAD��o����VR��
B�ÁJڋ�9�!	M�6A"���I8��45[+(5�k+s`3�*��g�]<�·��
馐�)�e�'fV~����i�O��l�~_���n�G��4�y�g3����S���a6��i�X�0n�W�o�u�d,�[m�����.�����ww	������!�� �,N�,�z�����������[e�,��������P'E��G�ݰ�ʰ;<ā�ܺH7ڌ ����,�Sʁ�ft)Q�m���4Z���U��$�H�"��\�+�X��y�����;����=��^�*���r\��)ǯ��=ݼ�f�!�Չ�촸����q��R��L�Ϸ��-���Ŋ�POy�c��=Ӵ�k��v%�^�Wi��HY�"�0]j���~:p����#y�c��G�j����o�B�dyf.q-�ޙdC���o[ٝg�nf���ܤ��^B��&�L_���Bkv�C�?���@^��Յ��;�`�! �Fm��mtFji)�`� ���s'Qu�F��f��R��D���� ��a!�#�'�$����J�e�{�7�:8�}Q�t��L �Zu�����7v�F?�J���9�����g/���zE�HO�R�����ټ"m�8���,���!��Sq]��a�+�ۉ`��,l��GxJ����T
�ыן�A.�&��im�0��"ö��a��TV$2�!����2���n(���L�}O���oD�C���� 8�t�b�V�_'�ȸ��2B#��	 �)v��40� �Fw��BS�O��;8 �n\ʭ�O�+{g���
�$�ε�T�yƻ��;����@���?��Mn8\���.�|���ЛҀ�� �aj�R�|C�qwI�*��A����j!fN>�#�*b��^�S��߮�^�Ǒ�9nA\b��)_:�4fJ#�ԧ����6���]����OH�1|}�Q!�"�u3��+�����2��&��w���Ͱw�;ie~H�yݣ���a���狾�N�b���5m�O۪��x�NT3A�i��2�
sCҜ��DĲ�����9|��vz�E(c��O'`>�1C��B7<���l'�$�*ԧ�G{x�_��}$��c��������6�>�}]&)�=N�+˿}��zr7I Y���{L�y!�ɀ���L�٘��3�k��I���0�S�u�U_Q�����/~;;V��B��A��w�@Hl�#��㏌�ye)�^���j�WQf�F�n+��/�U��Ns9~]8��y�e���0���Iث�a{ʠ����~~^�䴻lA����o�@&g9R}�����*t��0����cP� S��5 �1���}��	$���69<#�2E}�`��+8���DX��[���3����8o|�g���0��7q
^M�"��T5����
��l�Xˀ�|O��S<�vBGY�bV�cL~� r�Hq=��q�O���D���6�0;ZZ�#��v��P�TE/�n� P�x]�������8of���|��{��%PiU����a�}K���,
Vǵ���Ԃ�chu�3���S�A��A+��ŭ��^�?���|��w��ȓ0ˡ�p��6q5��� DS��_����L�3B _����<���]r��"y_H�K��� �ߞ��ӟ����Y�N��n�v{
�����܅���4�����}i��p�̱�^�� �����4�@���](����0�f��k-$�A�aI(g��h��d��u�������J�6>O���Q2�~�u࿛o^0"�����F�gcj�E�i4?F���V!Z-�QG��oK��i�d�'(���ɞR�b@$�/��DcDLfD���w��L)�QOq�P`h0�J 	r&��JՓ���4�k��_�5�]=���+f�bn�`c_Ȱc�_cM����E�}�_�~��1�h�h����_-�B�ƛ�GC�u��JbT�H���	�
LwW�z���WX25��	e�&!�jX;YG6;��D
�,���Oӣ���5L�[sD)�|��{����%	�<`v&�B�o�vZI��b�'�$�G���uf�1�0q��"ʻX@t�a5�N<�v��?o�K�0�jnf�ɩGf�zc|��/�4�a�p��U�BeD���ʗ�)�s̨�7��b_��A8�7�(��2±2��/��9�����؃yq%�����f�v�^���Mv~����"|�AW���a��r\��D���B��K�Y[rE<w��\N�mxؾ]�;sHS��.�M�����E��)�=���DL݊�&砢�RY��6� @ 6��wy��H̗l?��vt8��}�=[On��<�"{�����s�u��v�JT��}ŗ霢��"��d��B_ Zu<���S!��2zB�|�o{;zj��5r�_�5�]�Ak�y��j, r�,�,GH�q�Im3�����T+*����"&a����7�-���P��r�8ʔ�C�����J��Y���A���0�軐�]o���p�=��wi��=���Fܙ8A�VëԻ�}����k�!����7���a�ݍ��c������88+�gٲa<<2u@��B������B�;)t��z��36ʬ\żJ��L�|D���MyO�%!����VwO�E�rTP�����o0�Ǵlz���xB'�K�]��ud�~�	̲��ڏ����͵�;���Wˢ����i�O�O��Z��Ē��j�O��h���O�i��q����˲p��*\���?@��j0b:H-.DqJ����������9��5!� 	��h|����a�W""�1�N�������3�KN��JP���?K��ox�w8��q�P���^��W#����F�rJ=� �"ƂɑW���@b�t��t?�-�\�]O����˦��V��	sg�@�x�+�ǧ� �%���S7L��4��8�:���f�v%(=0Q<����86��VtV4~(Y�OԘ	� ��?����ׄ���l�40�i/=P9k:���C��2�	]N�d%�\���i�_���yp�D#�y>�vcuV�G���qrT�1NI��,������詪BK�-{-1ZoB�H��]�ܶB��l�"w���
�!���|5�����a��w�$Ҁ���_�Zx��Q��A��f��Tx��u\P��v�s8&cB;�-�w	K������yh|���:w=��8����(kvUQz��{_�\L����]TŮ���-��&�܃qS�8��o]��vD)�1xo��˦54պ"�ȸ'pۃ�H[��'�/���%En�L��6-&� ���ϡ!h1yB�M���)�4B��͵�l1�y��j�eݶG�[P���I+�%��NK1A��	lP�M�&�O���n��"��Eڄb�8��vl�6�f�= �}:"��!\���Q)�f��y� <O=����H�O�����S��/^��y��d�e[Ql��K�^�;��^�Z����2��iΡ��0J^a�-�[,5�_��E>E���σK=��c4֕��k=�)�I���9���B����Q(����#�N��c����8bY�{t~�"U�i �՚�R�7��m>׊�*mmk˲��rW�՝�����K\EO{��,|��1=/CH�&���P2�A8�\(_�&����~��sݗ�#����<�5ܒ�V���T������ C;����&�=�j���ha�#	xj8����t��~[7�Dhj�/�1�����_!��ɋ���6[ӂ@;#>�(�c¹�1����� �z�����j��kŐ��n�Y7!����"����w����|s�Ӧ��u����šW����N4|~l+	�l�s��6#!�ì��'��o.zx4&l'[���\�c2+�!Z���V�3�j~
�7�%G�(��B�=��(Qf�n�Ɩ�rJ ׇT�֮`��l����=,&il��\�4�Rd�g������	� �Ʉ�H���@"�ͪ�f�^`d����~���C�;��5�#�������9�}/���t|�:���G�۞ľ�ܼ�uv�_Xfb��t)$�D�%������M���V~4!v��� �g`g��F�t��<�|�4�b�v2F��ᅬ �̗�D�E��t�j�UJ������8�����A�yp%�Sj��8��{`�m+
F�ش�xnIB���7� R����Ux"~"xޙg��L⎗�CQjV1BǏ��"f�Hh�5E��>/���u$��KWU%�)��v�|T��I�
Fx�2��`���c���6ylS�6v�XG�E� e{O�x{��Iߋ�
�щY&V9}�f�Ei0�VF������Ù�v����%��g�e���m���v}HEN�24c;<�M&5��0e���_��ⲱ��JU�斪��P�8���.}�6�<��W��~KUK�����l��JP)];�*�`�ػ^�Q�/:)ۺի����ʟ.�T��҉%[%�P�"Ew��p�}9�V�{���4D�. |�ɑr���M~x����)^h����!�J]�����-�'��c�V+P��$�8�٬������KN�p|��t]�g3f掄şR����v�
�A �}sY�����$�̞���I�[�������ď��tز�A�Q.���U�t�l���'d>p�y�!6g���<N0�6���Bv�\6:�q��ƽ}��%J��X��9�l�����fF��c��#Kݬ~O0�5�%��:���}~��:�s�}���[�^��Q��������������>�E�%���B�H�N�k��ͱ��]��=ӄ(�G���p(=�S�^j�,*��EJ�*��BM���o��_A�I��$�|���r~ǥApxr�g���ޱ`�I�o�V^�r~��)��ڭ��?>��Q�U�����ՠ�.������F#�v��&�n����>���S���C���M������}S���SQ�! Lk��k݅���2���Nh��o7��oH.�%�7������*�E�O�P�
�b�v=�t*�d8
D������Dƀ�i2��#��o�.y����qԀpV�)��"�sv͗�~U�9��J{��.��'�R`D��
Y
�L��f�9�/� �������e�Of��	?�.'<"��e���p�5`���W��ҵ�����c�ԃ"R�fx�|HE�h;u������	���EI�@��	уL߬�$�wԔ`��]�
Ʊ·�b��~7���Z'�R������{dI,F���e��� �7���~{X� ��@^$��حl2�0Qj���g%/�y�.�$��;�[�Dٯ�F��$2�x�K�U��^v�B7$J.?����O��ˬ$�.V�F�������	V\V����ӳ�1�n�*I�i4�b U��|[>޻�C�/w�������^`����vQ�
�	#�IJ�\Vw9�{���x���X|�\�4@A�j6�����Q���bR2�xn�#�R�WB�����T����������?�:���z�<�GO/��t\Ii#o0�RDչ�	
8ȫ�RQ�������x���g�X����k��-E�<����v�͎y�r�\��nؼ|�$9��'AS��|���>O��Oc�a�c���ѡ��X��u��I9�B��c�m���j�u���*��(=�\���e��*�uu 
X��d����܅\ɚXZW.-u]NL�Z��~,���˚a[ ��!�wQH����U	ͮ<\!�M1̺`��09̝u��d���m�fє\����������h"�9��[X�؞KuG�y�7�<�c`��5gO)%��m��@��瞉V���u�٦�t,�-}S����F�}���i�m�q^ѡ���wT�Ɲ�O�w�(�n�
�ƭTǉ��ETz�䖀�JIP&$qz�M:t(�R�+�.��vmV�:�����, Bţ������+[?E���l]h��T�y��R�P �d� �c�H��C��7�=�|��cy��RE��d�����Zq('��c�.m��P`�L��pYP�3�q�=�G���͓���?o1�[��tY�ٓqW�w�ERC��c�V�[��.R]�5/��|�_Va~b��t�	�.
���>J1��E�����["�
�������YXz�SZ}��8x؇9W��To}����O���Del�KB���flD��5L�/V(RX�ߎK�Gv�4p���Hg����~d����%-ZpܤT�B�j�V�^&�6r�L��O]�g` )";R�r`!"���=���O����7��ƪ�A�G���x�0Cb�������q�o��)�����r�1\�c�����mx>����qN*R*�m�[kt=,�D]f�o�t7�b:���_���:O1}�^�V�'��8�r�v�;�b�����t&��E�JO�B��ۇ'6Ĳ����%G^ݬy�g���,��p�K�(�m��p�~�ӗ��e��i�h��Y�6b)�1�?��Mk�[K�2C���Lb����b!��+��QmUE�F� �
�׿F>{�G���?���bl�p��u�?r��B�&��hKv����o���i�ƃ���5l}�E�!��p�����18����age���?�Z�H��W��2+�4i������8��ln�������<�}�ř���j������a��J.��i��8���CWOW���3[j���Bin���%��W�l�GQ��Иz\�����B��;�� U�@�����V��fKʤ��i������ʵJrU+�x���\�֋=0�i��?���;����@C�
J%�Y+a��Y� �M!ҢL1�o�� `�wuk������g������Me!V-z�S�N�&Y Y�V������#�d�Ȍ���z3�4�Ø*�(�s����y<b1+�Z@K R���m���x|��RR&Kv���i��m��a�!Kp�I�}���d���j�N~�ˮǯ`�M>�i��	%�RU4*1BO��cD<B�v����J��dkǐ�± ř�rd0��'���˻��ߌ��LJ��h�?U_��,HC1�>��V��%�U�v�q��k�@ڵV��qt5�~�w>Т� �����)���֨d���a����^o�8�g�+��n�Cb����a���+��w@����f'�"����� ��Vӝ�{Y39��ں�`5�
���z]i~�`ye5T�t#w�W�؁l�L�[��3'��>x��Y%,A�"�l�!��"�K� ����AoȉP�j����v6"Y�X��)��B�P�	jg����{��B�t��+��^������-�4^4�;�w���c�c�_�)�6B'ڝ-�
��{�<ҏ,���N+���m�b�y�������E�I���c�ὐ�������-�r5���L��q��~��ݶ�؉*:�d���N}������U-u�)�Ä�P>�c�^�l��`.�)y(ߜ���#�1�rR��ظ��D� ��l�����_q��'��i�x�?=�x�ҡ=��BdQ�I�NZ�9qi����?�K�y~�X���{d��G�5asL��K��Bi ]�[5�U7Gouh��Rz1��[�Զ��چK�];��ª��{�!�5���#8ÓI�I�yf�T�v_Ȉ�U����O6.H��E�*qw*� ���5@
fy�ב��*�>����h�����E&��s].m����� l����sϑ[w{�%��GZ(�0���x�f��8SXZA?�׮�ҹ�IY���2����"���itP�-��1E�aJ�ER��L-Ac�i
��lT�t�M���1��3�9��T�ة��&��輧B�wbV�T�>�y�(��Ӭ����aJO.Ŗ��� [��wi�Z
ͮPD�����CI1�F�JY������!�]�p��!�%�V1-�Fo���?�I�E�zc$�����\�#��	nq�^s�j�G�Ң���:�v����+���}����'�9��k�h��C���Q�݇���^�G_;��;5������=�ޡ����:V�D"�z��W���1�0l�+�5��5����<?�i`��'�kM���;��\�⅑�s�>�~-��2sdJi�wF����n�sW���ЊN�l������Rx�2�n�1�$���k����tD���r�+#�9}��4�=ο1��Y��nk�]Vr�����2H�ڤ��$r��-�"�[�b_X���[���V'Z���t���uϣ�m���n㲫�h�����2̤k9��m����H��V��_B�gGK��~�Ġb�����M�$f$��Yl$U�����D�$����cU��k�x���?�@�_v�Tl/��-S�{5C7:^R�nF񾄡��
\�:j'%Ҕ��F��M�����K07�c5pK��d�G���<��d[uI�#�i��0q��>��{_ܩWd��"�T�l߷���(�OM��]@�x�]SӚ|�o]�b%�w��d��긪�X��:�l&�?�{W�E��^��'7�4�	�!�|:+�z.*��o誶�o����,.�H� 6����<=�F�̚:�ܬ�cy(��bg�bs�g���a�(h�A������zb�&t��ē.>�\{s�C{���d=�s�b"�3Yc�jׄ�"�~-rS���OW7e�o=�;Se!�;[ꇗ�-� ύh��WE��<<��q}H�t�&ӇU��*<yG��ny�-�8Apf*���)_���M�V�̷)������c	�:��v�[z�&���g{E��RS2],����2�N�6�	G$��8�R��/��Wxo�}�f�j��
��J�"�`����h��ѵ�i7��%�;���G�3�Yt��Ys3������}z5���+�ܙ�wa�>%�� }��
�Q+i�����𴭕����rk=S��m�q�+�i��Φw��A���Z��W{�ڡ#J�?�9��Z�I� M���@�nY�������+���n��l'"�!�C,e�nT�{��eP��}�W_���B!��3Ee�~4�4���Ჷ�lO���7�f�}p���I�
�V�׷���.c��,�0�}�{"�u���vf!�"uu� �,zU�]1Mh��`a����27K0�B�G�`vc/1��b�_e��3�b�]u���4������ҧ%��T�s_��	�(f:TƎ5JHaZY��������f�jZ�ۛ:��7Z�i�Dh&����e}��VŮ�\+,���0��.�k�����^2^��<��1��vt��O˅p`����;�������:T����+=q:�8��m��Rkl����p[fJ��Ǉ^ޏ>��������0�Y���	F]��e[:�m2#��"�Ń��n��x��A��?���2@�k����r{�O�-���"D�XOr�=���⊿<gr��~I�k�&�T�H xoN��0Jv�x��H�~V.&o�pCzP�M(�_����%�w�`�����r��ȤbA�\����6\���k���Z��A�&��Y�������]�Lx���}�����
��[oQ�D�]����ԉ�E�|��Y���Q�̋A� ��0s��6�� I�~��p�Zd��i42mR����ui�c1~�bր�nl80��:��#z�U�~�k�ajy`�7^[�l��~9�͡��G��x/�资|��[��w[vc@;.(WO�f������Z���A�p��i�R����JC�N),Q�|!�����]���M��r��@��f��f{,_�g!��{K��ϗ�z�.G�������kƌ��Z��`��ES/��L������r� �K#�X:D#J9�+��B6�&.���Jy��ʧ�c���M��l@�it�	��<�~�~SB+
L�Я#�+ ����#�,g�X�k��M zh����}D"}T-����'�)��,�o��g]߉�O7	G��a
5�+�0��7ᐁ	�������:6��ǰR3�j�eɌchG.�	KԐ��5-��n�P9H�::niBY%��ps�e��`䳚�kۭ�$����o�F|	�x�R5�pˏ=��M� �Vf�N>���{G[i�4z��r�#_X���[��G�.٨���0����b��y��q�~Hlj���Y�yo��~V10�� �/N�49x�ޗ�L�^���=�,�M����c��D��YmR������z@��cQ����&�U:d��֣�H˳�����ǋJ�:�#hu����OL�&CmF����������{@��l����uE�f�v�Ԧ xt(y��@N�Ji�rj�-��`Z��fſC�|���nyg��ı�$V�}N��s��F�d�(�٥�tX�R��'f+�ʳn������T24i�%����P��o�[ɋ�0ML,����<����)t���QFvy����UCR�+�N]ƥ�.���)Q"�U���"�M2�P���/id��z��b00~~��xJm��`�#A���uy9��|��y>޷g�����.�� ul�JJ}�.�J��
�0"���;���a�:���>h���U	ᓺ��*����H�Y��c�	�{���܁���?3.�FG{>�y� }��;��;����z�d3
q���Řė���Ãy/.�v�M9�
A�I�������EE�\MI3�)H������'ɡ�E���O�/;�%�ϷA����YQ��i�G8���B� .�q3SU�G����F� �KХ���o��<�ZL�:��K�Q���~O8�oC���PI��ǉw:�����ɒ7zIf|LX��y)��G�#E�H����b�)��_�f� ��
V0�H�Q�WUt=_����f �@�ۮS�l�߱�����4�h�L�~]�[m-�P��yߘ�)�������Y��-v�A�*�&�(���6O��fh�ΐe�`nA'�/.��	݆����Z�텉�ב<bݤ(�mN�x��V�'(�'�� M~
�/����샺�q����m(� >\����l��J�To����n�wt�0"A��j��q�~DE?-AU��<��:�i��@Ԇ�l}�l����o�D�w��D�mu��UrXh�&��$���V�yP��\����R����5�~��~q+<���)�g/Ͽ�	67��s�L�mT�m�4�_V`1\8�7;O���RI�˶�"����qiR#����2,�a��g�ꏛ ܝ���÷�Ǭ��D"�6<�q�K�wD�>�}�i>������*����A2^���F�{iҰ���] Ó�����m�窈��j
!h�344�u�2KڏN�bz�L�F��o���lry@(@X@����t�i__L�?餒���Z�,J���z0�P���M(�����p�w�KiT����֤����$��X��s;ݐ���_oZ��k�j6�uwCk�))�!��x�cв=r���V���X"����ݓ?�V��&l�m�_�a�K��(#Wd�V�.;�S��[�q@"��~U_[V������ݰ͒&t�^��	�/�-s �h��L8���Ǒ�����e�em��X����2�؁h�������f���L�͐2V4hm�n������V"3Jl��y����Sʆ:�r��G��'Fg9�#�+\�S�+�����w�C]��H|FQ����jz9&�~�`N�.�������/���Nư������k�NU�c��1�p5�v��)����烳��i$b#�����L�츦����`��t����L�c��u>�:���%*���yy�]��X�^�O����ȢU�a�Қj[���o[C����q�׬�+��%�=dZ���I�?C�4�/e�4����n8,y��O�stf���)�c�wUlb����r9 �x�`n�m��'��۶���T6�D�)�CMz:(������!8Z���"��ʒ�)�7� kfg�,(�r����~�Mn�K���~��ʖp��ݥy�>�
����qP���Kt���=�.K�ȩ^���|~�ٶzܝ��l~l !���?�/�%m,���6��Z!�_��iU�n��F{��V��TN,�M]��F��9�F�CˤG_5������>wO��^&��e~��=�C�]2iMC�S	Q�f��ޭ>�jAS=�(�f.VQ�0�E�_Z,-V� !A��x6h�`�(d���*s6?���qM��4�/�SM����o���?����vx{��O�ɛ=�|~ه�m�O&��@lg Ǫ�?�j]�L����+�K«��򑜺�kw�p����l���P���fq�w'������}^/c}��E�F���w�ނ�CQ���]B�-+��������
L����t�.c?�d,�˽�LpunF�BuxH�q{�*'���6�4��tZ�i��in�.ܺ�sJ4�#���C;MF�SYHxm�{^�N2���E�l[k{T��	r#"��3���L��!I��|����k���[!�$3�;���!=V�!1p\0��
E�%�<났lAo2�"���H*�zg�_tU��~V&�-l�-{Î�M�:s�R%�ѡ�R��Z�b%�0KA�T����C�ȳ�3P�ޞ���%7-2��F�>����}W �I:t�����ߵ!�k��E���?�a�=�@P�&�e�c��eڐ�Y�)����PSsz���!#-uR�i� <�;�"FFn��膏�e�#��ҏ:
j�ϔr>�� [ ���囐��o�#�.N?�Ӽk��*���CW�p�t��[=��SB����VM���e-�G���Pf]��C�PYͰ]M%v�L:�~Q
,G;��˄���|�ވ�쑭(a���$�=��Kf:�n��eyYs��B%�^���w��0�i4�����^����^,V��γ\��
g�<��T�il��.�V;Y#9m!��$W�t�So�A e��G��J��c�*�Z��M��]�����uQ�?����Ӽ;biS+�,�/J��Ɛ��$Ԥ�e��U�!#���kJ!
�+"�?ЬP���n�'|b��@�(niχ���YuCy\\��;pU�$U�5XV�u#N��^\ L����N
��� g���jꡨ�.��a _�ȿ*��6���|YF{�5�KTۙd@w�v�Ź�>��*=�˻`� }Q1f��L���}��Uuo��҅t���sQ+� �_��M��ձ4�q���6�t3ޗ���n�6g;C|g;50��A !Zn�*��o�Iٵ�J���cm��Gڹɜs�!�l$4���0S���ꥰs���g��V�2� I[� �;z6]��T9��
�A6 ��Z�k��+u���i��1��܅3�w����,ZMjlW^��wc"�b�'-N����%��$��,ʆ<w�#hpf�9 D�O�x���\����_�ّfVl5sqxpW�縟�����?H��'&2fn��(s�4�FU7��7���:��?�/u)��nO��7f�;�L�����0t�� v����ô<ol����}��˔W�JkI�\��l��~�)o���_VA�y�Y�+�E)F��%B��ᅼq�:��,�-�4�� ���b�5u?�p���-ьgZD�+����A�K.��;%�-e�?���9W��P4���6y\�� �L~D
' �)M"9X��Έ� ���,��v��i���N>@�h�j�e�>3>�����|�[ӥXND��������檞����*���l��rj��:�UI����&�6��s֟@̙N���|�7��N�.Ⱦ�(��rfɪ����(}ȶ8�WA�)���}�<�?W��Y��g����lY��8�J��#�m�d"�_��U?n�����b�m�VO6�b�ଇ)��K2��~�7.�=T	�N��S�˥��*�\ND������n���/��;@��|�=��p�,��)R�G�|l閨���;�hČE�t��M��ǩE5eH�����Lْ�=��VK������XX��;e�=�j�:��SQ�<x}�1��Ļ�4��K[ �s�z~azӶQ��A#�i�$Ek�������W)��<�)q`�.ߤLta�l5l��W<oF�,/��$q	N/5�;$�ש�����eܬ������{�e���x�KN���̤=Պ�j~}ע�m�����s+�����Y�+T��[	���*r�2��B�
ҏ�q��`���v<�"H�R��DO�]'���G�B�Ⓑ|�)�Cb?��v�i��8�ݱͼ8�|�����\6�4<��lUR�q����$
����ڄf"LU����I�H�ܥ�	���;~`\ɓ�[�c<�v�:�ɜ�ov���1��$k�yE�ny��n�F�w���yŢm�u�xr�d���	����;�)_�.l��M����*�aR�}8���?.1�P%�V���b� �wH��)��=�d�e�@dEy/E��/���%�~T�b���H��ÅQ\�8��
_�?�X%\$�p&Xc�gD�0[ʫ'9U���L��!?>��A��ĕm����y�i�C�x��oA9��R��Ӣ)�E�U�/�G����,�O��A�p��^�����Tk;*VLh���3��	�U���[��Ղ)-��芏�3d�%��lsˊ+H��K�s��,�[���G�+�.�\ì.2��lx�-��k����u _����<�r3���r�����ܤ��W9���څ�,�L�B۠X��{�����3p׌JL5��DdU�D3�ǐ�)�q���83�Kt�ɫ _�Tyz��)����9ò�RR�<ڤ���tj�j�|�»�r���+�[M�/BD�'���Vj����8u�7>ϼ�6R.[�͑U�bI��H�'o���L�M�
Tk�F���	��(rH�L	࣎߳:�3��u���z��2L[t�0l,��k�(h���ͭ��?�σp��P���%V�|$1s��ܒ���-T�눟��8��V��6��&��'^�C�LI�>-�(�f����-����W=�#�A�{'���ͪ�G�_g�raꙈtd~g�:�m�n�dP������R
#�|����ڗ=ԗ�K�m8+�{��x���ɿ��1����9���>��"���c#z8X��A|:0�^J�7���/=���#�H���I�ˊ����O�P�P�\���##,��lT�W2�*%�a��؂��>j�'�^۷������*�!x��X��Е:�|�·6ㇷ6A����~!o32�][nc�W���3����%�~�W��jl�e�Nf�Z�X:gp��6|zW���A��y�{�)��}-�؈��&��m�vMT ����8xa\j�c���3�j�hk�+�E$�#_���H9���^
h��I�n�_�k`��̓�~�Ǖ�ٺ���g!�P�'OT�iVD���g(�"�1��t��c/�ѳ��-�X���Rg��'(ޖ�^:A���ڜfu���О������/��d���<���b�p�7�U�{���q>�moF�~W�mS�����h��K�!fs�:]��SW��/FǨ�f7M���a��k�t�����0�����yr>����}yW� 3���3��΢ӑ/_����Jv�$;�Z��kd��9�ٯ�ɣ�������
3/��)���ІQRR��r�sٌ��T�k���Y����,�U��%ž㤑��	���E&}���=���V�%�U'l`��R3"�2�+������c��1v��;Jī�ho�a�����4(V�*sP�۷}K��yhmw�f|��A�[������G����=7�$r+��~��Q����Y����(�W$�Q��bńg�]��%.{�f��ӷ�_fA�0��:ۘš�=��^�˩3�t	�eYs��Z�PM�
���Z;�]^y����T/�q���7�������u�\�hȫ$�@�h���������˅weX���	G���/���s9���e�u�n����P���J'���Hk0���𴳻d���O��я��O������Ā�d+�C�s�ե���t�J(9�un�~���/�q�V�P�{���~�*�C0��jUU�z�u�b0'�e�lyxA�Q�	��5d6M�~c�u{��E��e����NC!'o~X�ǳz�Ze}w�U?;��֏�xE Ї�?�J2h���g����g_y�Kٲ1�.���io�!9ٺ�����=�1VJ�W3�2^�ߒ%��/T���= �M(Q ��'��`��^�_�+�=Ae=�g�i� ��ChUhQb���a}!e��Ka���L����e><���������(\*�F|�ͤ{S��@��̫ �ͳ4�~�L��Zo	x���m�� �g��N^��ADQƹw�d7v0q�n���4���Ϥ�re�8��_�����E���Eѡd�`GU����iG�h<]��
�_�[OZ�@1ݞS(��B�tKwA��ə�ԑ��A�3��u��DR\�,�m���j6���{s�v��23�l�(�if�uD�4����f�_����v���i����g&� ��u��z�C�>�u�y�_)W����DD@	AB�C	�F��Ke��t�#�i�Q�f H���{��l������v]۳��}�s���5Ǳ-�'Z�-p��������"������\3��wy�o����ṙ�lM���#��q�6�1Z��	�ǔQ��ɝN�P�J3��ȸm�d-3A���J:���)f5;km}���l�K �'���?�Q0�싞i7�	o�
������弽�m;r9>�;B]��<��t-��*����W�ˬ��	i-������k8"�^�h����t�0c�/�3�Rd���\
��x���J%���텺]�f�ńh���p�T1p��G������u�IN§\��*�7cu��q�jq\i̒�eQp�1��M����xJs(�	�tpt2۽�XH/�3&:����c�x���i�v�l�^�A���W<%3�r�ۧ�ՖL�vJS^Q�T�LO#�N�G�W��W���)HF���_	S���=�kp��8��^��r�.���ch��WPI�켓�C��x�{��:/�MH�斄j�э�,z.�^įA�6�F�f����B-)"a��s�I��F/}��(�|��(�-��u��q?Y�Q�Đe���AB��]O��C�5Z/UpiO
���eૼ]"�Z��S\��Ќ�u�==���n#~������lY�)��S��l���������"7?^���K�^4����,�L:J�o����av��
��  ���!���'	�Y��`�5�5����b�/�i�+�"�A_�w�+����>����~K�&����?~��u�k��nwo��!}��9 �9.�4y\��8��sV{jR�j�hr����7'�{?\Г	 �z6�9��z��(�_�2vi#�"��Ƣ����w�>��Op��?۰v�6�󵚊���G¨�x�煙�2d�ڗ��C�xm��.�����Ȉ��������ɭf�78ʈ&X� ��9�)�yI��	�+i����I��Vu�Ɏ�I��K�SG}�CaO)v�/_cOtxU;	ڈ?み�Ty-V���^Y����qE��'�ٿ&%�c�|����wIJ��%��ޅ�]�&M	�0�zū䅡�d~����s�5ǻP�%�sa.�'@��7����bI=� ��GP���ˇ�PN�s}M��IXk�9������&#^0���g�D�Mn�t�/����LbF��lw����0���I�I*F������Z�g��v�>�=�l\[�ȡ���%��7�t,�/\��pG��� �\�<�zhjd*�/��bԘ2�!���g9�'���*���.@1�7��ugdk�B���O��QY���:�y�>��?���
��y�������s�v;k��"v7��������\j{��8�{}b<�\6�"k��XK܊����a�gk�Du�<�Ŕ]�$ �:��_�	{�L�1mm�L��'Ɔ7����0+��R��R?�)v���ײ�X�a_`�7\._r=���V����'��� �@���s�|�!!
��. y��SN��nchF�he0�-���WjrΡ�R�_�[i	
�Zp	6��t܂;���_�ӻ��s��
���9|lW�H=A��T�-��<$���}�:�2���R�d�O&^꼸;�l�=�F)���zH�e��'�"���M�N�\7�V��9&+E�tf�@7��L=������/��\���.�F�HC���7I+�r<��P���dLRY����|;!�,�y��<aw!FMkL��<����𢎢/��~��$��]O�Z$Bv�y1�mi�l�i�([l�5���X ���&M����{����-ӠqK��߶)�4���������	��N�>T��Q�F$�R��qm&�	v���_M�V;8��z]Vf��x�c�B�X�'�B�~o�؛W̟�������Z^���
Xپ��Z~`�!�SPw,U�}�F��|g}/���``�'i�Q� �
u���aI�,��v&z/x��j ����Bj�chJ��ha;S����9��U�gz2�q�bD刃�l��0yy ��M�<ڈS��~���}�Z��-��.�8����+�Y��9��]W�p����0��c�As~����_!��.��*fZO8��ӟ|���~;S^��W�)�ez�Fj	���r�&�����;��M0pvJ6�l��4�Gk�����8xo���vL\M��HV���V�+]�C���3]�â^Z�+x��il���T��4�?�}� �(4?��nZ~�l���ut�e^��_R4��T�oR�8N����쮱2)H�DR����p 䇖���o��@�$������J��2Q'����Qy�>���g�0M�� �s89�a�+_��|�)V���Q1 �#`,+�Z��*R���g�U�`rn��Y�̮֠�&`���b�V�Ɇ��ɴ>�D��YӾ�R���zc45WBS"��S�2O ?�B�T�
�9ة�ˌ�u���\�Og����or6Z�Vo�0Z�f6O
.���c�?�&|���\�py,�3~u�s�51ߠu�9��mEO9�8�N��V�������5¶;5u\��V��ҋJg�^K8� u�^Ó8��>6ݤ^o�h��'�'<2>?��<�lZ_��/kǍn�;_�x��y]}왎�Oi�v��<]�2K��jb����#�O!τ�5��z9�Ѽ����T�c"�_��X�{���A �"�36�1��-Vaٷ|�Fh������;5�}��?��5����ad+;�r�n�W����e����a�	�#�n��O�원!z���hL�J{��& �y�Q��7x�P_XV�}M��"��{�+ڿ�A0g�O1����p��5㩘~��s�2�hBr�ə�[m�7+°�(:%�g! �Bk�dV�z7<�:�l�ڟ��Y�^1�m��Ŝq��)b�z�9B�W	?\lkd	e/'����N!�f�?\�>�M�A�&���G�WE���
ו��b7��#w�h~�25!�t8G�H_��a�u��`��I���e Q���ٚ��ӧ���ءփ�	� �F��w�e�m��EYd�/��N���=Ax���3����_2܂��hӸ&�;�UUY���s�A����C,�ѹc.�����ş�d��k�zRj&ڜ���'.��'�y"���0;��?/w� ���"�֌r�a?k�zi�{!����?���򧌜7�y��r�ot@4x��4�1�9�6��1�љ�n���'g<��Ȏq5��#�Z����JW���!��[ʨ��V7�q?��vMC��ܠ��M�����3��r����qj1O4�B�3UrPT�#�7��Uj��:�����l4y�uW�H�W���E���塸�A��񥨏N.���wfw�B]���1)�����.,g�Xо��Ry<�A������Ga~яnZ�k]H/�9Rw�51�R-8E�#3ţNN�SY�:�+���$���}����K-<LJ�FS�����3�21�F����3���[�o,����=2�q%�mقE6=xj�3���`QD�w	��0v�<U��m�~�[��6�e{m�����Lur�H�7<u'�爠�|P��)����=A-��_�ډ��!6EO8�Q�I�%s�	u���d����z���=�����9��s'��j'��<1OX�/��+�5����F�V"�x7����l�h�/��*d\C뿼��Q���0wE<>/V3	$��e�X��������Y�ۦ1�"��I
�S+~����C�E���=��}���ov��,'�FYI�ƃ7/@�W ��F�0u
�ܵ���bA5\U���@��7`EoO'���3Ž�S&,%�m����A��?bqt�� �J,%dE8$?���"�)
�/���CyP�k�5���c�}���ѮtH������a�`�4c�d�4�e���-���n�Ή�W�j�@�-��U�]���ci���w�T[1k�!Z��.�q��9��(�W��Z�W�߿��'�z�����?��w�Y$)��61k�MAs~��ч�=�t#�ĥ[K|% ����1����=��cg����d�L]AǙa�`+jȽA�Hb��Na�P�!�Hg�ڟ������u�Yx~��2WNՎ���� ���f�0M��<�hxMb ~>*��]U���{_N|.`4|��s�o;�&�k�VH]o����H��ۡ���#ePF`��3/�ƀ]Q�O�/��ăv�N���òr��f���h���Lv��@֣ܯ��i%�M�uٍo@�i�&d���l�;\�5��Υ\�=���҈�;^�[?�g�z6 �����&�S��9����}�%b�����S��n�U��ņ$�����QcӲq�U�;r��ɹc�ȓ'ߗ�)���1%��I��T��JO&<o�<+<Av�Jv�5�����-��ƚ3_�� �C�1?���i�uc>�ׁ���f ��DZ�	>5�,��h�Ɂ�(j<@��}|M���*o��։N@K�UWbS���T��sX2W�K�M�cPU��l��`�q��;�Z���S��䭁�t�S��x/͠��p�<�ou�?G<�=��;����g��.��و7���ڗ�/�K4����ȩ�渵�樶a���_7�W{QFZ뾳��W^�/��f��t���Բ�f9��z[���D���8�e-C�m6���{~�~�r��B����ͽ3�����.F`a0�'��ɨ�J���Mo���l򇱥j<Zj֮n���u�z��T��p����X�T¯�#]�#�?��X\��N{�.�7�͡]��gg|��?�>����j% �F���˭%�pS5<�,��ř`0�Wߛ1����^Zlsu� M$��w�iH�����x����w�L�t�f_vB�% ]ӛ���g9��1V�p�dM��f�lC���㵓q�Y�Z��h"�7�t߸�
Z��%ގ�]UZT���t�r�b����g�7L���7�8r��$�O�y��t�$��_���m �`~��n4*R(�s�o7z�<��((�J9��h��]]��V+�k�Q�.��ͮ�T�fji�pҹSk�	�Zi@C'��d�/$c�P!+:�}$��d(s�hd���+��?��%R[Y���P9x�+V?=��]]�Ѕ����9��v�t�5�(�*��c�yK�Cu��{��y�6�V�Rw��r:b�u���^�q�}Y��q�-S�?�������R�t�GX]׸�Gl�Ei�ͯ���5C`��|9^'f����ôC.��\��	���G?����dG���B�M�U�d��3��&3�Q3�	R"7�OZ<�X� .���G���}=�;aN�O��5��m�����4@«"���w����'�;����g�Oj�+�Qk���=^��}Q�N�Z����n��q���쪕��f:�(���Y���t��c��ƫ1-.^��5I�S�g�s�?+�*��H�3�2�	Ok��z�����n����-��W0Hm���#x�s��,ݞ�P:6�'/n��$�d��qR]��\k���碞!f��v5�9m�a�M?C�RH���F����Ϻ?Q�FLff����3fW����@ְT����K�LM3�Lo�׭p�!2�N�lQ�e/����Yit��	9_�2��"׬�rkz���]و��!�W07�q��$���9w3�jl��m�4x�#M�r���+�X���ȯӂ#o}l��H��8�y�\1{����h�ּ���t(Urq[Y�F�T�ɪ���g����"e�	��i�T��6u۟J}t��亴+~	�rS��ʪY�~K��UZx�E���O���<�#��M/�ýˌ�m7��� ���z�f���&���#D������՟-�Q?�����.]����b�%�Ծr�l��{�Uc<'^���&�e���\f�W�pLK��Ҕ#.}� �B	b��l��B+ƴ-33��v��T���1��xx�����B��.`q���*����;�4sWy��Agy�5E:iǰt~�é��Li���>\��Dˬς�q��ͽ.�U��-�,����q(}Q6��X����,Eٶu�<G��/4��W`�k	]YD��~њ�L��$��1z��w!x�ǌW���E�KX\�n]*6C@q���S���|7TR����c;/�پ>����h������y����L6�v�m'��O �ׂ�)x��D{�͹RZ�N�Qi�d\��7������i|�,�j�î�F��3�����,w���5:��W0�|-�p��|�O?���.���8~�ő����L�HI�BdT�`�,F`�Dޑ>ў�9�����U��ݩ[�<�s��c�h�;W��U#>�q���C�����v��5e���|`��Ϣ �?�<�W��'���Y�m'�bՑ*s�g��"Y$�Bv��Ͼ����������1��E�������tyS��B��o�:Q`���ώ�Dg�\�NܡG%j�S��u,�Q�P[�< ��Ï߶^��ڢ1i���-q$py~�����*=�q�o��p�N�8}��#ہ2kae�]��qTH�^n){��j������w=��,����b����b-K&���G	ų�cX��N��pv�|p�����.TL��s��=���^�B����&kb���
�4���MK���9���HJ�m�E>�����z#�==�[���W�.��h#ѷ�t 2":�}6��,"�ۍu����؍�XL��Y6�ɭ�.���?���8&��[Hp�W?pS�d1��^�k�:��ap �	O7��$(	e��Y*���k#"��+���u႒�ZL�T+�}�ڐFʓ���ְ^�M���-�[��_��6}v<8�\B��j�gM�b�t�*hI�g-SL˃�2o���@��"4i�(��9]Cųۀ�#~F s��Ŵ�I���m�Zϻ�����G�u��h3�!���u�_��I:���;-	>��N�"��y����~�{zMv��$OQ1�C
�F��g|]~�B(��%}���MYu��R}'�|��j4���������$�r�c@��qK�F�������	�J�Ꞣ���+Rq�O�o���������>EO-��!�ٯe���v��h3�w!�
^���T}��y�w�^��c,Z�&o��ڏt�n׾��7F��e{�`O]E���c?D����e-��>RL�y���6,͊SB+I�Fl�O��/u�qU���"���Ϯ>9�M߲��)�i��l��7���a�^�G2���)�'��G/���u�����0�H��ũM7O)&-�j�^�#�g���h���<ٰRqgţo�V9��3�a�w�C��sJ�2���	���[�=�u��3*��Wϗ.�j�c��Xz�{�|8`��:��)r� Ȃ7��������g�}}!�&2������YJ;1��.���p�kz�����y�%B�a���;�ĭ=�HeP�,��{]QE뜴�s�p�[[ �_<�ʩ��)I=/4Cg<a*`Q�+��,�%�v�"�z��7��V��E	 ��F�����K�~�$�H7`e�q�M;6h9�df��{��
����nE0�A�h��դ�9�v��N�t<4C>�h䍸��>-��	4�B��f�r�_�i#~V�@�?���o����`3�X�Ξ�te�͐J{n�ڔ���(P7#��8��Z6���$k7��	-�%���xG�=�5l����8vPP�l�ۓJ�c+��Ǻg�F�{W5���z\�]b���H�e�����E�>��ݯ����qI�s#:ul��Ϋ�m~"���zL�0��UU��Xn]�U�M�b'UF��M_���ٽ����.L$��y�X<Mq3p��I��$o�)�^ʌ��A��� �D��h��@�Bqd��6-����>�?HL?[47:�G--�.��	 �Ю�$�� W�6���R,vL��<�6�nGU>�����vkt1Q�0���S�E0�Iy'I"�����:Pm��D��sFn9"0C8NB4Y3ɓ��|�b����עY�ݻ}o�SEӤ���ФҨ������]�P��e���g]�7ۯ~]ʾ1}FA��D�����g9WE��]��B�u'��~�N�i�8o1Z���Tv��W��p�.Wʃ\�1kGo�&O�/;O�^����>�׭f{��~����ޅ�~~-)H�:R�g���;�o@��F�m���R����.����_aLH�QZ�)}J�u�K�Àl�ƙf�,�Z�e�Qȃ"�TIj��!����a�Q�;����z!���{�7���ɩD.�J����,��쀧v�S�e?����oZf�C��V0�*�Lڬ�;�I�;���;v���BS�M�z��������.c�d9�c͊�~��h������ U�f�Ze�|n��ȇ�һH�o�n뮵�H����_���o��b���11��-ǲ���{�5����Ѥ��S�3Ł|M���0nÕ���]���U�9�{a�ȅyu�Ȯ��7��-J���.��o��	s��p�1�*����~�_�ȍ�1fQ���Eh2�M�f�_odk�$����_X'��H�D�]$�û���m��U;Oc�m�)��otAK�^��.���j[y<��&{zN�-]W������^�t3�|�|Bۅt��k�g�SG����Oߟ�r�G�&��>y��SrP1�+?jg�V���ii�H*�3�2i��N���vt�]0T��]���4t_Q'���2r:姇:�O���oI�tR�:��.y�m;wQB�Vnr��D�2�_/�V\�o.~����G|� ��r��ȿ��nA�US��sG/s��ן�<���_$�����v���8�27$`?d�Λ_��Gh���2W�2`�KG���>���	Kى��D�䉶.ǐ@,7�8�FV�k��#i4���h�Nt�W���T�^��JC@��=bGb̂��ؽ�[�.w<�ek��溰�+~Id����IZE�^��B�!���͔FM%y��5�g*&������~�����lrY]����^l�6�Ɉb�dGk5�*�����㣉íc�Rf�c�uC3���f�`H�T9�q����t�4��<�x l���id�j�Iܞ�P����AC���pE��I��I��߉\.�\��H�,��y�c���5�ET5E��Y�%�jg�k����"��9��i�TH��<����>��Q�ɾ��yw��n�}Q�`�����,�H"�n*^ߩ������ޕ\<�B�wݾ7m3'���D߿��a�Ĝ�ssV�0_��\�jhƙ)i0�/ �|�,�p���C��5k��_�B>%؄dL훛�z�p1��4���e��l0��oٜ�)쟒�P]>�3H�U�b_9�t��	"�^|��WS�*�ij���+a;��d��mB|+��7�0���]�><�[�9�����Ʉ�
�"',��l�U����}?�l9)c��-a���в�|�\3��ޒI�,r�^�N�b ��l����p��v�����ֱZ����l[�z}#1��3��$��{�*+p
Ik��W^�+�ſ�*���g���Ji���{���쇲_k$XV��*�=8n�i�y�B�+��v��Zw$�����/�B�&&��1M�	�-����pk��N�O|�5IH��`z��j.e\ہ��>�!��I��7�ۊ�+%�'��1f���SAj)�y��
�%g��i�YAP�Y�V�ꈈ��U��{ �`m��H2v�H����E��~�X>$垚��}�?1����"m'g9��W5����k���/���F��Lnl�N�.$Px�W��cM*Y�.�xQ������6ыq���P^6o�� Ěߩ���e^~?�����m
dX�)/�5��P��H�wL����ކڬ#:�2�����i�IG9��|��>!S�yX��C	%���N�coŇ�� ���zm]����%�4�@����474�e�IK���B����j�	CG��R��v~����1���t1�[dh*����`�(#q۞��k����m�8��0�*�j}���/Խ߃ܠ��o��'N��^�'Mt~[~)��Mn�|�%�A��b}�}��`>����?[jp�X��4sD�S����k�yk_?f�����C�hi��21�i�Sœ�RV��l񔖾ᢨt�<W�V��l�Ԡ��:�B��|���/y�|��G4^19�){TO�\e��|�1����ټ*Jo>���i�,Vd�7ަ�%3�����=�!��l���c�PYV��Ü�s��h��O0�d��ʖ�@�d��(]s�'b��]�����S�/h���^f��$���xK9����҇�O�o&����y.t�XG#}% �8����,�2����T���$g2��-ˉ5&"���'"t%�b���0�>���7
� *��}���)�޵��Z���:�ɅQ����b���|�A��"=9�������C���'�����)��Z\�8X�ױ���4�D�Y��b2pK��ۏg��=_
,׸s��<����H���Ά�	7�VC#�����S�{[�j6�x��3~u��*����k��js����N�#O��~�t]��N[������H'hL�F��4:;)���(���~��]���)�@;~��ͽv|Z׿��:���zJ���\�1^����,�}�Y�����>�z}w�h����(V���Ǹ�6y�ZCEG�h�� PK   (}OX�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   (}OX��n�% �, /   images/c1d4a215-2c3d-48ac-b15d-f6239b4c4b94.pngĻW[]5Z��/��w
/�xq+���^,8(R�)R���w��������;F�8$#cﵗ�9�	�J
R�(�(o޼A�������&��EB�~�=�.��"%��b�d��LT^�͛߱�����vҚ�o�`t�^0}� c臔Nߜ�L�,lm( �&o���9����ٸ(���?q�s��*_˿y��&�E�w���Gҗ��Qj������DB��i�Q�|8\�VU7���IW�Kj�o� F�VOL�� E>����0����a<l����6-�g����)H���(���/D�tY�d@��� 
$���������~��2�]�4)L�ׂI��������� ƒÿ�`oBo]v}�]y����C@�7�����u�aM�gz&»o�^5��s��G�i��%���bQ�@�A{�&��P!k�p]T6��a��V����k_3���2?�T/9�������Tu�X[��I�H�4��-X��\­�����Y �dO_#V��;\�|�)S���-b�\tQ�g�%�{���UQ.<�-FSq��#=��Q���M2���ʇ�����.�	�`���6;M�t�{V	��E��Y܂=`�$����vO���8h�Q�s�����7���� �Y�ǬL����1$�q�aw�L��T���@��_s�k���5����u�B���j�ً��mcs�%�"'@ջl1����������cQP�WSGX�������|�7������n�d�dtW�cJ��kh5�E���Fp�nwY�><����`������7��a8�9�TjjhBj��!����d�^n;�Xgvu?��`s��8�I�Yg�R�6{Ր���9w���}S8WR����M4�j1���+U�o�0r��k����O�y�6V�5�FXfׁ���zcH��9��mh�"T�	'��[DP),Z*� �T���(�ni��tt&�{�w��(U�{��P�6��mWx����`iX�Pp�� D3n#�O�}sGn�3!��WN}��B�=!Ǌ������"k�\�N�'��	�"�z�>Q�qYǍյ�ҟ��r�֝�8�����t,��#VS���e�9S����1��}�"	bX��!�,ѷI��{������4 ����8���������V��`p�|�l�D����ٷ�ldZ�*a�d�Md^��5�,=al��Q�/
Bл�oYT�6r!�?�罵{�+�nQZ�`�Ze�P�\�u�m//�~ Y(����C���bm~�tA�/a�i<�@&%��j��JK�l���rf��A������\��T����jmڊn�2�b�`���a)�:��v�	�!�K��ζ�*�� ���_c��ABίP� ���z�ߒ�L��t)�?�h�����{�<C������)��@�3l+��U�Dcؤ����=�� Jq�X�L�n'��av�I�b�ATܳ���bl�Xh	�}#���^��Es1p��^�v��j8��IG����I�9� �d�dMč�.�ފ���~�L	��Tׯ$�Y�ޓ{iS�1�������t�
9W�x��Cx�x��s���>�_� \������8�)�H2�����剗�kY?���L��˪Y�W���{`�VQ���l�F��:pGQ��c+%�\��r(枖?��T�<����:���eϰ���B,^&Ki� �ʚm�	!��%����uX�.[�T![��As�vD+�Z��V�����¤83��6p�B��
ˌ7@�-�;-�.>�����F�ޅ_;�'��0�i3ナ�KZ�ʅ�/��������*���C�����ֽ��@�>����C��qA�|Zwh[���Q�3�Mv��%R�ߟ�Ҷz�g�N6���}� Υ��߀k�z�u6�����\�1n?�qd6x��w�)p�k�G��\BZ�ì�γ)ЏQ����5K7BJ��p������ �Sy�%j[�2�x���>;ѱ+W����m,lb�M��SnY��!ǎxyP<zK���kn�M�@��R�Lֻ!�����	��BE˔�9���Q�t*K��>�j�˚jwVw�}�~�$��(��������|����c�i�	T��(��W�G:$]�J�"��Ц`�6�[[]��QV'���eWԗ;9��ذf�XVٲ�/�^���a����$�҆i\��Pi��H�A��[��7Fw���^bV�P���݉���m����q;FK�|F�5G��vW |�c��4g�^�c��"�H�s�=U�Q�y�tǜ
_�S�zr���+�u|,�フ����kPE�`Q��� �>c[��$�Q�C,m�����㘔���y��_��Ʊ�s���ɳ��{��k*nVg2�u��1�k��<�q�go^Z���m}g �f��د�&�ab��	,u�iv&�����O���L���P2�V'��P5���2��ύ81q�3ZV��̗$*m��c{p��A<�q��e>w"�I���(�.�@�L��t�sϿ�W�p'Ki+��p�of{�ӻ=��R�������P�Ly�8�'̊�-����/����N�R�Cy��e�r~Һ�m��-�60�������<�|~*D3��x��bF:&9��PM�����r�d�OV0��d���e��-p���C�jq�� ���Ȏ��� ^�ī0�"  ^��!ݘN�II��n�Q�|'WQz��Lr��>r=`�_��������Z �������.~�zσvX<��Mޯ��.�IP�GL�n-N��ia�	�9��6�I&�K�N������0�O�()�g���\��0�P��j�Z�K��q$ǭs� ��2�7dK{Ֆ���u����3 ��;��r�b{� �$RiӜ0]��p��- �M��������}6�*wl|��_C4m|y��s	*�����/u5�f��{W丟ge���0�#�I��S���P�CR���w�g���"œط@5�M"e�ڷ��i7��ȳ�U'��&)H�,>�%�� 㤃I�R}7�i�@��|V�""��\	��G쓂�內$��r��di
x�X��Uo��B��I���b!�A�C�&��H�������+��h�� ��qmwR&x%��2�gzl-:L$Tʾ�Z!t:�{��!�tr`�������`��b��2��9�q:}v���f{=�=uHy�+و��t��rΐ����W}Q'��z5~@ʺ�/;�d���¶�.����v�=]�Ҍg�r^���}_C����B�� ��;�@{�źO�O������<"_�nYȊ��o�+E�@�(���g(�.e�^��8��.�B�dG3]��DZ#��ѳj7̞�c��;�h܅��|T������8�nai�ߝ�����gO��1�r���̾KY�@-�K���矚D��%�1U���;���>C:�_��:�Cſ�Aѓ�6���(�}s؛������^��Q�t�ͨJ!ѼX,���	;w�5�ۈ�2||��=+��;3��I�T����|{K�����E��b���m�$+����w�7$�?n@����.1�����FQ�iX����G����e3���d>�mc�m�H���w� '�<�q�%^� 1#6���[r�v�E�Qo��V����^{ǩ]ҫ���9ۇi_G�Ȏ����򨳝��v[���/*��o4�㰧�y��;^�a���6B��F�x#�lf�x9�D��ws'L��R���u�-+��\>���J��\��֬��c��<zk�`��sa�!�-M�/w@0o�w�[
�=�{{"���=����33�4����8�"s+r�K�h��B!�����k���P�Ǔ�І��`�����b��?<;	~�Ũ��H�f �����F�?{"*i9���P1�.�Y�N�,3 DSՀԖ��9����N����e"�j해��Q�HA7��z�>�q���Sj�� Q��2' �*DN�/d^�[�X0h?���t��Y7ouf�I,��Ƅ#l�Ϟ�A�b��Փ��1�\��������υ�>_�fL�?Z�Q7I�`��ﶯj��z}�r���\����zV�T�������5v$�}e-q2�H�R�R��'s~Ķ-$?������ց��2�M����UV��fg��	;��­F��F��s�]W�G����d�W"�\�1��ʝzp�*�5��I%��%�f}�v�ҵ��?L�lGM#I�Ez
ا�1��&K-�$9�k��i��-M7I5�*�ђ����;f��|�z/���N���?@c�<��������/������})�$�-P���{E!�Š
"�^g��茤�+g������Ձ��I,���Los��'B�d���G�#8p�BVƸ�����3�ȯ#wiz��nB8����
l<<ּx���m�u����H���t۷B�hQg���({��s4=B�� ��
	�P���= ˸O���n��uw�b�v����<A�#�uo� ��"��:�$q4!���8���Sv\�S-Wץ<�,�uJ��(m~�c��p�$�"�_ �w@f�)Z&��ๆ��qE�2�Ϣ捁:m�
�����,�����1$��V��-	u�c�?=�vR��뽖��~�&�j��JQ ������h͹P2�;�H�Wb
��_$�갡I-�eL%�u�i#�ߛ����k�t-�M�Ȣ�ܣ����%B�>ZqH�-������r��" jt\u{��$N����ѝ��٢�ʴ�B��S�W�`[���d�%�6�(��r"��F`A\a#���������JH���F3�56�L��1β�\+���0���1�X�}�Z���#mJ҄*���w:h?��ɺ��et)#CMJl�b����9��AR�XUn��q�Xewkd�umL@y��E)��I+�7�̇v���p^�ӇR�T(̼!u��ȝ���_r��-r�
��@��v[�*춯t�nk�$%HD�_�_0*�b��%��\�)=Y~
�
�f>z�f��DҜ�[%��+7�±��;W	Gm��F=�Pȵ�${�6�F:��E��;�j�4�KR�7a��SI'�2�I"�	�)�r�F�ct��a�<��<�(;q�UfȌ�}���Ȫw��@K�䄀o�������s�H�Q��k��u���t{'Pwm�JƎ	ƚ����V�s�p�99�_��q0��0{5�+8�����y�d��,�B���R5uZ�B{l�ل��T��K�$�o��%">>��Y|��M����>�����Ȑm�C�U,���S�Dq<x�*�
$1Ԙ�^�4GE�P�ц��m�ǈ<"��:)�E&�^P�87�^Fw̱s-�)�o�?שS�����`�����g����ȧм���8���j:�O.�*��@+�� 3{���N��}3N�@��w\G����Q:/�����=�Y~�uo��Hr��Yc�q��Y;s�wb�UB7U��+L�5��b��o�����˹���|�F�J��:����P��C,kP@r����[�D��`�cj,eȆ6�#�Ͷ,�a!���qfB�fs�E��\P�G��[�S��T�m?�K��V��傢�u �*��ޤf^�hW�l4ä�1���U��
eǵ�ʋiw~GAT��9@��� ݜ�����s��Lq�!?���2�T���$C+�p�3�m���.�s��]�IM�;��Y�NtWDj��ty��h}o��[�@q���4����/����G ���wu��^U3�i6�ٲzO��R���M�J9�hx����P��~���?:���"�6ۻ�p���g~��d�G�(�S�>E3���Մn"��4k��������LU��.z�
���,�1aL���(B��Ne��-�؊�c�@��m���Ǽ�9%d=�S��vV�����ى��f�r���;w�L�����0̷hW�1'&�۳����6h�\<˗��ُ�!&e�=�*t��Y�1_t��}��v����V�ߒ&_���a~c߉���}��=^��5Ar�]IN��Mh���PpI�Me�^�MS�{�v�C#,-�ա=m߬�6:�6޵�y�<Ip=����uH�cG����J�n/�؂I�F?l�?���� �xK<������u�b��ngD8̪��}��Q�x����ǃ������������UP4(�^�q��{wH�oF�?m�80�eA��Xj�zw'��O'�kM�v����s[��Ў���	Y��o~�%�X�����\xh�sz_XFI_K�����9��g�`�o�g3��:g�)t�i2�6�M����I)�N��}�����ďo�^1'��g�ƞ���O����7>۞7\����}v=�R,H]q�L_�f�o�����d��M�(�W~�/޵7
��莗O-BSd��E�:61�YR>F��As"N�;j	�Kb9<j�����BI;f�t5���_����-�3X�?Bo��U}�k������?��|��t;ρ; T�E���Kb�H��Fshߘ//h�<=H�|�-҅,�^��Z�����\l��i����!����,!���Ji�����#�+E?�#3��%W9*��j 2B�UO(�;��/����>99��]�:��|$G�m�^��&�x�J �<��^:�%^}���t���%f���[��3Q2T�D���r$^[�8�I���V�H#�e����ڒ;�s��ǹ��+^ylP�P�JE��3�(��,iŉ�����~�q���7:�%x�@EZ�N�괪{3]�m�Yv��Dq������_kd�f5Y'�ߔ@�7�N�9�;QAU?O��	ݢH��1���w�s��Q}{
�l~m6���ה�a
4�;g��k�́Y��R�2���-k�`�5�&5�&l�%�:wh5Q��_��L��,���I���T�ƫȵ��9�!�,���ͯ����v=0���X��0�'���͂{���.�(d���-[��X���#�������ēh���Ah�i4$�S������xVd�K���w��iu���*�(����u�Nؖ��T[z���Nܴ?�L�z��!3�y�C
Y�Ҙ��l����O�
~�9`��7%�9(�v�!���.ZU�<Yĕ�)���Wb�2��++�^��ϧ�$�����T,P?���m�8;r�9{�~�=��WC���&tWl�~hβ�Uo�@Ic�(oD3"��:�~��O���й�6����5�%iQ�m�@�:�v}�\�f'W��:|�<�i��yH�lψV0y��|D|�Lߠ�V��B�H�+v*v��/1V���'F �th/�.xzf�K3E�*6����J|�r�)�ME��p��4>e���q1� y{{s��9��k$�� I4�	��^*�#z�|�5E��o��4=<T�]���N`]z�2�3�4���i�z��e�d���q��!�9�\��+Ӵ�����w�1"ޠ��d�|قB<���'�2P��;�A:UZ�+Yy@tO���Q
_���Nl�0�e�E�J@Hc3�E)f�_-�� _�(�t�~�ֺ�u��m��ɘ�3�����Y�!5`�6JNNn�b��/��dP��0��X��5۩��OQ���NH�_��l%���:�|������M�[�X#]���(����L�PB�&��|�a���۞����E/�O~�]D4�9a}�I2�ꪑ|E����eǘf=
$��OL��x���rTn�ޱ������M]�m{��;�C5�,V��v/	����W��s�R�'u?9~_q��H`�P$�e^�;=���]k�s>�.F��j�8~+��^T�<б��Y$@�w�i�����ekڬP����G�_E�4F�\l�{�m��'CI]�sQ1м}M�m��_Jʚ�/&�C�Q��׆	K�U ����ٖ9��S��ߐ1X,~�ǫ�������8�ʨ(V�B�`9��@w��W�`8V��j`7�w�.�9�[-3��C5����_x����oS�H�iI�Q��~PǲH���)	M~d��%��k�'�8q~�N�/o��$��k^�X�Ɬd���y÷��Q I���o@�q�1<��|iV��1��8�2��Z
�ҥ�O\j�z����+o�K�;��0�'C�<(7�(���﨡�T��d�8:�ߒ�>���~�d̈́8�ܼٍ��u��{~�h�Q ��H>cB!e�P3~c�֋��*4�n��Q������mWg�j"�1Õ�JP2��nb�2���$:�}�����!�`OՍRHJbޡ��α�?A,�8�%��I�j}Ƭ\
A9\���f�(�`W����<��@y�<n�CA�$+Ǘ����і���Oo���hF�c+q�����*�r�ԗ�J��� Eq1z�/�B׾Sr7k-e垊ڠ���\��u�l�m�&�*��C�Y�2ҡ
���g^�nփ�k��MLFN�f	iFY�!9��J-�ź�Ͼ�����E��X�,�GU�]�t�h��oe).K�_c%���4��:�_�;��vUޤ�ݑ��9��w���D�N��t������+i��~?�
M!8TTW�}��ӯ�Ν�ts������n֘�mrq���Z�#�f:��CVMG�z��>��策Qᗨ�k>F�߀�A��ϼ�hH���b�04�]�U������fX�`m��΁�<!\�����ǝo5���e��M2�6� ��}���=��|���W�7�<QG�,c�u��Ӵ�I�G�ߡ�BZ{h�I!�EG��u�_-2��z��xl��A<�$�ޢj<߯M�me�쇪`ٞ |���N�nB���J��g[������獃>�5KR�z��0��&��lv���"�hW�Hz���/M�(!Tj�Ճ�3��6��ܒ�og{ĥ��� �N ���~%4�jB��8<�z��}/��� ���Nִ���*���S��
,m1B^hi+A��&_Y���X�LB_nF�(V�T���0��ʠ��8���B��bS5�rHb���"Jɘ^>�:����:��y�Ϙ����b��O�.0�uf I��3g"�zM�!��&�� 6%�zld{�YZ4�Ҝ�X�)�pR��>T��$�Y�|Z�_>V/�8p����$r�{�{\a-�Oz��Uu?�*YK�����g$ݶV�����ȼ�q -.�׍.b�� �{ܻ����/��6����-W���t�
6$6Ie҂բyML��i�&5���(��nӊ�#�-��}l���W~i@�W:�uG&fȋ'�$�YE	)���G��s���f��&h7���
U��~�Ķ��ؚ �0�O:��<��p$der����^�������b���q^������0�n��B��'��уRd�_���E�j\���}��ө�}�C�Q�ʛZ_�P'b0xf�o�g��o&�N:�W\e��^�
Sz����Rîʎ{IܦVˢCcC��A���TG��M��S?+H}M:�d-�͑�[E�"d��z0\�y�L��4�/GIu�]-��(�8*�,����~�CbD<2���f��,�.nӄd��*CG�^ke�h�$ ���5f!w�IDو9��U�{w<��e��|�V���Iv�����Y_���?������̓'F̦]S�Fj���_K���E����,n����%��4�p�n��A���o��-5) 7�)���c:�v�X]<�˒'ӂPV� T�2B��&6A�Q�z��fJ�bY���-�5y��mﾱtN�������t'����^���b����I��3��������)ڶ����^����n[�S�+\�uX$��9�G��F�#��C�1z,PL8ϩ4��O�V�������Z5>�&�!d�������]XRL?D	��2v�u��O}/?��M3_]�0H�I��8�4d��I�H5��>�I�6觪اƳ�'���Y�o'�+^�\�.��b��*Trm�1C�����Mi��ny͊H��'�ď*@�v5����ӠXp���U����a_,�Mi�Y�i�h�*Q�����NU�jX���Q9�0�f��8<h��
C'W��ufצ@�"����G����X����=�|<���Wu�Gf��l�y�����s/�6T_�B�Vש�F'��������Q^�XM�P��tS�J�9gҠ,�&)��wy���ʡ�p~�C�X�N �����G�u���Z;�Z���e�����V�(�A[������OA�y<�����^�r���U+�����g��{ޠ�	_��Ũj���/
�^���w�����d��޸��)p�k�2�OK�C(�?]�e�ҖUյ�����k=bd?$�J�`n�ږ2�]v]�2��=Ycz
(n�ټ��.���?��[�������K�M��_3E�{��k�J�<-E���n$YO%ځ����$���x�`-����yQ���G�	���X�\IEj/%R 	���~���e�y�b�2S���ҩ��3���d((�mZ�Z�?E�������5��iI�|]sܝn
=j���)�����f���L�f���<Y���l����D©Y��Q��*����u?Vʨ��� �6f�`������q���y���٥鎮�{��b���j<E�����
CZf�F8�Z��p����<[��!^V�cd�H%'��⑟�xO�Ϩ��[��"�p-`�-v�N%��A�	�]�b��L�f�5�_��lk�����JW�%��(��{��:�&4�[�B[;�����9��g�k�c�w�ʱ���D�U�
�!,���Q�b@3���C~���0_�I�w�]�,�m5<e��ln�u�����g��I��������N��P�H�pZ���u
<F��x���D� *���e��ɈL���t�����y����	ٖ� h#����q�e'�QL83Ӹ��4�<�"ק�9.�!QL*d��Xw�X��=e�:]�@���*�-RIT~��{=�A�J>�	�葛�B��e͟s&��i�*���:Հ�F.�1�!��D�A����/�oI_	4�f�4݈W5���/)�ԟV�B����ic X�(Ť^�yD�����=K��ͨH$Q�ϯ���Z��(�Ң��!t�a���`~X�/�fS��$����6�(� ��t�L�uex>�x�]X�]n�@I=�t��ҕ	�(HA��F��{[3�Z|ݢ�5�O�]^?o��x�q.��o���[�B��ԃ�ٶlM�����؉�3����&l���m*[g7Iŧ>RǏ���3�c�l�*Ɣ>&���~���I<��>�2�-e4	�J=���1A� �������%R�m��y[,�E7����
�!��
���d޴H�{�N�(������nӱ��앢c�n�%���}���ӹe��'�m�f��]}Q�]o:��)��iD1�/^�؞�3GV_�uf�|h�����q���p�V6sO��ao�����pM,�����[���7��x�b�%��i�]b��ҍ9�.��&(,��x��P�[�=�ݓ�#!�Vs��Ng��9M�����v6�h3�k���)��S�A2�SAq�����A�ĺڐ��R�?��M���u��E[�{�&�;	�g�a�~�k����n��R�K<Eڳz��*� �.w��z������cև�C��w�&s�;ye,���Y�3��#a��Hp��M6V���	�� ��o��<u8{f!*j*c#�F��v��I�a��Z�����:���I+]X�an3�&� W3.�LLZ��f�����;�ײϜ��������H"Ukp�L�Ja���OGX^�O)L��qA�۞;���si)���>wi��í�k)���<@1#��43�\Y��.8w1A^�2n��ɣy���b���X�(�2�r�d${���?'n/edx[�{m^t4>��*j �]���VxA+�� �m|�.�?�k��3�1��,]�h1\�'�z���$�󀛳"�`ecD�|�+����=�O]+Ɏ
�M9p Ța���9?%�J�w�#��\�=^/�����^I�f߸U�2�΂�K1�ʄ�t5���x0h±�������}T)e�	'��L]�z5��8ȟ�C3>TB�.���\)�ʸu���3��p`�[G90�-$����D��p�[S��,���ٙvX�ci�Gi�6ex�Ү��,!�$JH��z���2ѩ;�/[�!6�� ��_�hq2�,*ћK���MGԥ��X��i�h7{��@sFB��K9�s��-�p�._��ʰ;���H8Tw.�;s0Q�ry��n�b��s�5V�&�Ϙ�H�V�d]9k�"��Nl��s/�g����}&C��r�x�18����X��������RA1��Pb�t�Pr�D��}��"�wv��E�~�����{�Pd�1���@Qy`@qI��jn����"G}7D鲜���닽=����i$�P�IHZ *F�X��x#w��8�$~��x8�$�U�N#��B�\sk���Z!���i���dj�N@��ݩ�����m�q}����o�-ML*��5C�uh��2�	q֦1TpNI����yS#�Jw�Ut?�	��x�����g��&�_a$N:q�g�R+oW|�
�� ����xQ��WԂ���{�a�~�� �Sv%\Y:vP�خ��:���yW�c�:�O�&��Ny���V�-�p!��~�s3����;dH+���[�%T���sf��s"�^�į�TU#O�<u(Id\���(J��w�6��C�wF�la�d�������.H[��2��vi��K�7'���'k�}� i:�'�(��*Ͻ��:���B1�W#���˸�φ������[�VAT�P��C�N&���%r`-r������~8�a���5!��<�$�f�@6��#��AA �t���h�eM�'x��V]i���_5&)��|Ǖ\�L�efܢ�[�i�u��`.�mg%��
���!dOc�>:%���u�xO���-����8�N������U�քE�3G]�C���l�/gF����o'ȕ������އ9�i�6�f�"Q�NhZ��ʴ.��)T)y��MƐUE�D��nd��h!��g*㷁����q�nRw����lAb9���P&Q 빃IB0�4{)?2��L*A��w�D�E\���Ŭ�Md��uKG����t���V̲B�
���u���IJ�������}����-&K1�6-�%�+�ػIGT�le�VH@Ihۍ<��Bwƺ8~$�T�L�@�I{�U�5���^&,u��w1�8�f�}����kvpy X�݇(S&��?���$@�jN��@+*�4����-�,!^s�,�}���	?��gO������Z�	��0��s��'�,��8�#k��Z�9*����+�r$ن�z<ab�$A�T"�p�k���X�Q��j쪖=%��[�
�����S��{�-�?���3g�xD��|TB�/�E61�ck��v�#��i3Үb�8�9�!�_�z��Yq��?PgM1��~֣g���l2To$����ʺ�-)���~�7 
��R7ۼ�����%W���O�����Y�7�p0����+r���wa#C������#��?��C��A��zw
Sh���%�J��l��JxW4��d�{M�p�LI���ߢ�Ut��W^�߿�1�>־�)�����v����a��K�X����R@�;�Ee�TX�z�y��鶱�;��:刱������>�g1�R��|��z���X��CM��������ZFf���U��m8�d��ک�	&���U0.�?9�`1VmY��Uz,�/�����2�7������:�#��?��x����S�"��.M%��z���f��p�9��p+�_ք*õX(L�=#�y�jJe�ONp(��`��p�_�s�"�$���*�i�Ae��,��C���8��vc�u��ug�;,R�D�U
#j�e��/;�P�]��܎pa&{�A%�f���4Eg���sR ����y��@�&�sE[gs�r9�K��,�"�\Bf�T��=�;)})���~�F��1W�W+Pҳ�@��:T�N b�o[�����a���z�Dm0�q|�΃*C��R��������2RWM���"q�^0�r��Y����qX�)����a��]����qlr�j�93R�;��^;���Odo�Z��̢���{ѝ\������4���l����#?1�/)YTR�p��Hr�j�܏��������V���UG������.�W�(�SJV�V��ೱ��m!��QP*-�,��R���� ��AO>/DѲ\.޼`Qj`�-�=ZEZ?�g�R�r�!*�o��R���IV��}ƌ$�&!���؃��v�2����J�*ڔ�C(JS��w���|���.gr7?~v��(>��w��Ug�R���m���x#�>��G,6��h��9F���p�*r�W����[�Xǡk�fT���C�2n��	��6xy�U��Y��p.���X�����'EW�[����Ӻ�J�f�n��쮍:0Y_��I�]�̠D��2V��6�81�"����SVF7^�6���,}O޼cE�{���E�\�M���� �蟵��9?��k6�m�`9(���h���'�6�|�F7Z�Hd�dF��E�kM$�%��&� J2G䌚�I�D
���/�ңmVϿ�xU����z��_%�PZ��D`;��%gw�y1�e��.�bQ�X�_��/iaϩ������~	�����F|����L�D;�9fZ�~P<��쫊$�jk�:
qq��)oL����Kێ֟�K�N?�dp�^���􆣐�R�y�Wrt����OTO��yTcro��B����ߕ�v��"�������#J�w����<o�뛭��T���􆷢҈N�ɼ����0��f�������t�f~��2)�2���Q������Q�3�@|��'N�`;�x��T�[��R.6N-e�HH۵F�Z;#V*@�t��]J����8��q�]�Z�����+�����7���}��~���&`�%ݽ�vR�8��l�ak(�4OǗWU�����}�3�?�@�K����&�\d��+yv;*��3A���F2���<�=c���
�@�0���v��Y�Q�Ul"}����a@ߺU2�����{�+,A���#��!<@6�!���C���Ê�2#��sh����Q�]�u�r�a ���x��;M(�T�ˑנ�ݟ��v�>��������}
�,�V�oH�L��Ş,���/D�$@�0E�V�<�>�{x�h$��uJ���+휚�͢��Y��̅iƪ<)F��0��d<d�X�����I���	�Lߥ�������	cP\
(U٨:i�˰}�&�V-����� ���E��w���4�"f��r����1���Qŷz�� �{�ڍˍ��9����Bn���?("܂3�Spi�>�/�{��eJ��V��.����	?6��tZbJ`�)Z�$�?���0,.�S�cߒ�E>�p'������uG���
�K�T7P6�cHFI��w$	X޵��?X9���=L �&�<�+���}�x�d��󮘴��U�B�}]ӄ̮G��!�&�'��\O��$�NMܠ�p��z�eF_��G����1�?_E٫��G�n���5`�r8����l�<+X8��2WA,A�(>]��Il�i� ^��I�����[F���T�~?=�`a���������1�_-�L&�@�~����ڵ ��7ܥ�.��M�XͣD��ԧ_����d~W��1�ט&Bw�Q|H���BD��RD��|�xy�U��N��_��l�&m+��" ���q$���N(T�w_V[�7.N��9zl�A�>��vĻ-��p�S�/>��h����sf�����U�鶙|��UE����.��uz�?i�(r���j?����~�gkn1��yr�1��7�|e��$��z�H�����f�w\��BM�Oc�Ղ�-�����h�ܲy�a�DM�]X��登�z��#L�ơY`�SZ3�=�6>��ܔ���8�J��J�iw��r	y�Y�%��nG�����Gl����鰤L��"����O�l�N��&600�Dc��C6�\�DB�>� ����I{ʈ�R8$n��el���)�ϒ�Qړc~�O�~G�^��r�YDʣ6�kc�u��న���i�[�q�� �Qo╲����h�P��	W�dg�)J���ǭ�k�5�P`�8�BN�l�� ߢx]i�Eն�}o�}_�׍����+9=h���z^,��!R�ϡ�w���Y�ٍx�Z ���h�V?��$�!qvZ�|d��d��_CJ�j�v�.�y�j�9﷉��sx*�O46���p�2U2�E	e�By�|91����7S�$}qG'�)��Ub	��F�Ұi���6& -�\�R��2�g�Q�����_�u��5��?l>X���m�ʷ���t�!�z4��Ӳi��L��GJ��doP�m�XMzz�A�z�vT`v�-��xr����#ci&*5�;��Z�d�,���Х062�c5��Έ���08�B_����96�p�rt�굵碷��?4]c\$���l�f۵����6�f�&�6k��Ͷ���d7qr���|�w���չg���J�A�:��[�;�n�!	�W�l��f�3awԸ�W|v:�u��$�(�zV�
T��CK�ۚ;:?�@���C|"�a�2q�2nf���8��,r��P�,q����J��O��5S�o���_M�����,�/I{y�� ��_�Ƙ4��Ȫ.����o[ZU����)d��V�|���ͶG�︙j���K=�),��Zʉ��U(�!/W�3U���qF�FT)�#��a9g����Pi���&���jh�!4(�M�qnGB@&+��'{V����ɶ3����5�p�yJ��KK�yڔi�t*����%�d���uƯ�C����zE��jY$T�')���H�2>?��`����`���I� ^$�P����ڽ���]�aV=c��y|@����󄶓�'4�h)2�#
@�Tݢ�X*��B35����O�7:*в�]� Jk�m5@2T'mH��d?�M�ܿ�/ p��[�{������9I
g��~��\¼a�V�4�Bc��5��X�b\Q;�.���6�+Q�	3,�4�F�zD�<[��3�k_u���t˿��9&�=�=�_�0�g+u}��&�U�3��Q���L��j�i����� �9"���/���0��P7A�9JG�)pU��~���z#�XS�$�>`*��(�FŹ��0B��6���a�Ͽ���tQ	�k��D6"�����Mu���H�%J=a�\&�h����p��1X�g�4���Q:� ���(�����0 R�A�h�i��O˳/���_3��L2�O��5Y����+�����9���T�C����:�"��B�_s�n'�^����o�����ϕ�SO�����K���������5��B�����e$���qp&�W���x%����Жp����S�ha3�?j������T���C��P�6I�~�G�� M�
z(k��/�'{9��[�i!�݊Bqή�,�P
�t�u���%\[/�~����}��D$�l����u����������a;�� �G�}u��_�%���:&)�@�B�L��'{}�c��ܯ�����s�j�v�+��P�X�d�z�Ʈ�c+������$�BR=���;H0)��JayOQ�;i̷T⛮�.�)U�ˮK��r/���|�V�v�w�U@�1�������i�mw�K����ә����M$��m�hp���t��q��0�,�~V*|^IY�}ԅ�T�L�r�+*��#o�,Hӊ��$p��S-�NiC4��|�~ny}[�r�R�xΎ"K��1��25,��6!�ҀS��
���ތ�G�K�UI�Åy'~:���Q�q^�V6o�� R������f�_:�$��F���ӿ��Q�%��j��� q例��Jp��M�H�8��U�o�R��3�Cmq>|�\\�^�x�i''�����"�om���8��qU-�0��|
�r�	���B�F�UD�{<as@Y��</�� �J'H�-Np�7�/Ť8\f髡�n�s�Pi`}>2�s���]zO�ԗ��%6
�C7j�Cʕ�'@)�O���y�MYeϖ.����y�FVg&��e���}a�����f�-' �|��Ma.�"��7��%$�k�=L��"�~_���2}w�x^zZ�!!��*��)��&հ�w(EH�xK��l�ÈH�RO�Va!����>;��렉�������b$*d}T�}a�.'���Y�q�{c*�t�ע�R6������.�d��2���Z�sz�ʋIvǫ�˛k�*;��6¾�+?:�{?d�ڱ6%�,]PXy�>��
������������jdt�Y��IG�zS�h�7���=j)]��/��}w�R�J?U媝���S�L>�������ih�w�0sR�N{SCCUV{�:����JP%~\)/c�����|�䓉*X	�%xELg�Q�.0uQP��<���ٽSaʹQ_�5b�Ω��sw�9v�B�
ǎS�:��I;�$��֑!	u*֓����;O�����q��B�(B��K�_�<
=�r+f�*"�26i�X�M�ľ��`��3\q�՜�2���)��x�:ǟ�6�X�:���"�52��!��;H̽�K4���� ,̓��>{\A�D�g�$� �<���"��lh[qc�.'N.[�*�aa�w9�����\��6�����[~�v>��P|��c/ +,W��i�3���(2��&�:���]^���X�����u#X�>q,�����	�ڽ����4�r>�-J�u�A�]BpKR�-0�s�-{B�֤���Ϳ�s �������Å�;w����1���49�8�x:W��ɡ�/0M��:�L��)��z;O��"�r�8
wƙ�r�"["�6/����q�g^��n��}O��P�����.ƪ��Mc��.z���T�	�,��3�[����V�,D���_q3y�~:�}���ڛ�X.�x��C�3'�;S��ڲ�};YP	�ƉB�lJ���� �p~�U0�ڬ!q]�1%� �:��I��vB�ؓ�"���	�#��Pu�t�*\=mg>�H��(Ӕ �:������Z�7ZE�?�&��I��X[�n������G�	Q~��D��}$�%�漯��f��$�ήO?��ć[����fΈ�L�m����fm�����;C��.��*�9�:��`\��G���Ӑ�Zy�ƴtJK�Sz<`B3rwX�8�p�R�m$�����KM+�%�%	�.Y' tu�늶���!��/#����K������G_|˴od8�����T^:�C%wq�Wke\�o��o�=�,0d�Yk�B�Uб��	�i��˗=D�Z[V�W����֧LY��;7#tSH�����6抱k*~�F���g,�#[_�t�&��y����	����P/�*��Z��6>���}ih��B�(�L`�9U��1Z'��8��$�t0�ϼq�Uϊ�v�6���=���n(�7R�����x�#�͏mk�/G�[��.Bu��x���۹6��`���y���PZO���K!۬Rnc�(��y�y�H:��͠a�-y|	ɤz�Y���rm���s���^�n��!��]������)��U�ހ�p�s����+�h���{�W�V\����l�v���l�r_����^��?����͛wGn�G�\�0F�f�q�W�>K���
��"�%I��}^4�p�z���"��_ܻx�ɥ�b�YaE�1��T0S�a�V?�k���M�b�$凒?�ᾄ���g{{"L��s�!������9���^�g>���"Q��n��$�EFh�hB��(�L�+���Ֆ�K&JX�DV]���DIk��缃��k� ���5���}��8W��,@�xT�[�c��fB��%A�w�{?��{ծZ�AU�?�����R�J辝�x�w��s�,�[v�h����&���bNf�)So�D|L �#+��eҵ:5(�"�������0��D��N�.B���T�l�#H?�h�Ă����L�|�tqG�@�&~b�N?o�F���P_�F4�KK+Y,�B���uo�=������[���ҍi+�i���w!0�Jkg��9ŋ/�I,�%�@T�
�K�[�����G��-��3�U�~��SoG�7k�Gu������g����{`�
窠1'G�*	�=���b�lsg8���F��*;�#n����nd�
:�͠m�h�|D�����P��#�r�2��_��yK�j)QJ����n<��vJ7��̲	�7q�~�@����@�������WO���f�m������{m��2�ݩ��"�. Ioc;�L�I��fR_o]��@��$�'=DLs�Ʊ���DD3:���i�&�)9	V�E9��)���m���"o��׸�w�;u\���(����]7*u��.��b���sڷ��Pq�ҋ��hm��x��`��A���R{����n=\T�64ƿf�^����`�9*��2����w]�s�+W>H-[T/����q�Q�"��R�u�סWɧ����LnMFl7�bU`�$I;��Q[zc9����gYA���%�A��!��zb�G���B�TD�ILP��zZ��eFC݊����I�xɢ��
�H��n��[�U�!m�]��D%���Cb������ЏK�K�^��s'2��AܵY���<�����LtԠ]��X���{�����/.Ӷ���DP;pi��F��N!c$�I��X�3��N; �w��1l>}���doGv?ld�m��Xr�a�
E��.�'ߋ�s�k����8r��8=�oW|�5-P��H�k��h(���T/ma3�0"��y<����D�?�n{':�}nkK�7�eOK���y~�GA�L=�VZ�(�����}>[�
��-Ls�t^'�S�@���{@���kE���*������C"p����&sb:����!��(����O]�υM���^'�S�w-2����nrh���E^D!-�G�J8�� ��b)�Q��ؗV����F)���v#�D<�3���!TcHK1�ۑ]/@%�j���T#nf���锼��T�N��a��2[��C��S0���ܿ
1F��52��gO��5��d3a_�}/�PT3DN�F�X!�j��'Hk�93��ru�\秮�B�F�-[�a��)����o�q��,s���p$0��M����gv5������YQ9�i��ҨUI���&���mb�e����Uu��p�B�=�_2L��&v��4�w��mI2��PsJ7�uɕ�O��RIƛ�=L�^Ld�M�?��q6Icݍ���Q�FW�q
��}�@L;8M�f�N�f6L��3N\�ΐ3�g1&���P�[��q��
�p<� (�D�iǦ6;�	�A�Vl_}�]�� ������1u����6&�1^��
��'��ʓ��AlhH�S�=�fm�P��=�I�k���0���W��`�
aI\�5j&�b��'w��l��<�X6dg��qQ��I巏c��p��^2�7_{Q��)"���/���[{�m��C5�Z������C��W�A�������W<]G�w�I��.f������%�^ǌ.�ۓ*d�ĳ�K�԰�3gtдȣ6�
yy�cUM�����EE�DDb9ɉaK�"+I��;�:y�ƴ��r�m�)�d����c�S����]Ϋ���;L3V��6 �U��GH�A�"D���e�/û���=b�Dfiw���p�-{}H`"+.�-ǐ��+�[8F����sE�1��dndˬ[r}u�bF�Ȋ��ȞqF��OU!Yae�s��������/��oP�T&ľ���\����^��θfK��筣�>��[c���G=I�!g�g�)�6b!q´]1�L<��!);,l�_ �`�N�����K{�T���
��:� 0|T[��jeh�d�H�/�yԚӂv�̂��ċ�lJ��r3��5Q��<�W1��^.K�Jg��������O(�`��[��u�j7ӵ'!��)c4�G�����D>��4�>ơ��@;��u�"�����wse���P��FԔ�����e���<��ek����YX��u)�b�
h�M~�7 3d��$�=d��I��a��05�K�up��"̕�r7o4օ�8|����&��,Al~o�r�CB����P������8H��qw���u��������g{���·�1g=��ɫř��C�.8o�?�~ gi#��`���@7=3�,~�'vۋ�����ɦG�
�׍��9��"$ݹD������.�����TKK�k ���{��yZ��oM��k�s�L�^�ώLM�}ɱ���M��҅�������,�a�|o#3�r��O�n���2	g��z~x5X4���j@l�^�^69��_E�1hg��/�:w͘w<;�O��H#�ã�z��q�F)M���*lq�,sG"J�!�R�o�s�	M�l�J�:Y'�F*Ȓ�O��NtĈ<&D��r�ɴ27r�(+J'+�p�El���4,85i������&�!�qk6����V�$�nC�	Yg�Nu5��.�ͬaf03L�'A1��H~��F�2�}h*��lG�]��3k�l�$D��By�M�~�1|��LD�UT��r�2p�5����r�mՅ�
w@�`Bp�1���%7?�+�y�����4sG�����]�pTK-q�}��a��J���I��AJ���< .`B9��^��sqz�=#�6�&6����h�R�5�%���&�1O���V����*y����)^
N�e�X�M0�řE� P�G0S�
��8�]�VǦ���[=�?�ʭ�i�,�R�[Sy2���j��T����&\�����(<��V./��B���D�s�嵿����+�!W�v�\J�l�*# ;�xr�Z<=�X�Ļ���-C��¦7��eE��f��Ϙ�2�uOi{}������9�7���t��h]����n�d�W,�:�մ�
 ;�:\DJ&caZ�!�򢋰,u�`!/������Jc��w��%1�;|>z��k�0n���#�O��d�qH�Zu�o"TM�r�`|��o&v� »>I�<֘�y�
oʱ k���4����j=|_n~����^f�/"B�X��X��>�%��:�a�֗��i%�X�J�����3���c��^d��7K�EcT�A(]"���%��eh�+��!}"!�����1H+y�j����{�+r�ҋb�iȨ���P�y2�;�K�q� �Mru��l�&ҿ��za���j��s��{g�	�|\rs��{[>����??�s���tzi��~�#�%��< �ٍ�pmha��B�l,��+�<|:�>w���v�D��Vס8�Q��n�њ��t�؍�9-Ćb,䣏��?�����_J������sH��R?N�9S��h��^�#S:iI���oy�R"dz��!M�1h�R��`6����3�f�N�9�F�a��?W.�$�&��H�)�F�*�0���MB�K]��5;�w~�� ��7>���ƒ"�@??�j�n_��'����N/�S���&]��#M�x���|2�������7V-|�l�łȸQZ��j^�2���_4���֐��6�J���j�ԕ<���Q<{.:�D	tW�R:,�L��1{����g�1z�Ǩ�&O����B#�%7O��WLu4�+P�g*O<�7Pӄ�u)�q*��	�7�-?�4]&^SktZBq�BÑ��y��7�g�-7[M�����3�fޫ߬h��b�J� )�� ��#GU�8J���m�yk@>ۯ�ɉ�ܠ>tG�������h�K��K���u���hy*~v�x��ȟ�tEݷ�*�"�!�xB^����&�q��p�~xE�do#P�F×�1�����:Ċ3�g�t�/�}j��d���ƎiWe)���<g;�h&�#^��\��ߟɅ�$�?��o������\]�{2au��6] ¹���R�V�c��ϗ���RtXZ26���_�Q��k�����<6�^��1���_}���@��un��u��i6�w�z�L�;��d?�Ǩ�o�ϐ ɶ�'*v���#�/��ؘxl��"�@�(T�,j�&D4�4R�Arj��g7��J�^S�0��.�ȣ�5�^�X�>�Bൕ�>"A��90eߢp��Ͻ���쥈��N�W�r�O/�#a��ʢK}4����%���Md^+�{�a��u=�P�ͅ��x�`e����l���\Mc^��oǮ�n!z6��Go~�K�$^ψ
��&L�P�K#(w�YS(��z�*,ը��	X��.�u������SЄ��~�b�1�Y�Fjr�A��+�A���~d38���#;);�k����ʕ�X8�>��t�60}Ta�BY=�O�ٯ	��HXf=�ک��2x�hBKeEg�Ygf��부�^̩�Ѷ�e��1� wE�$�_T����`�Z�^Sͭ0%�+�}A,��țñ8��U*3ҐKs��������P�J��3�4��)�y:��M{6�*��b�9u��lcձo&,�y��rd$Y["��T�A#�J�po���}�zkݴ��Ĳ�޻(I,����Z��f�귱��>uE���8�4��\�>�Wl� �{��V���tt���!mW�)(.������\��tb[h@��u�[V�^��Ŭ+��Yp��ą-�V�x6xkb}��X�Vbc�E�Gl�۷5f�<�"���{�#��im_�hѤzvE֋13G%�'��[�AV�!t�����R��G�`�z��GZ���!g�XY�Ѥ�p��}v�C�?ͧ����oM�����5����"�*�
�}����k��f�4�u���9��)�#����b���6��ݼ&�cN��$�	(�]O�3E����o�$P�߇�H�Ԝt02���oY��ja �I�t�z_yi���o8�H=�Ww�
���@�q��qiu��iA��d:Okx���)]��1���A<�Λj���F".kꑞO����ŉ�)�?��W�~h��OP��l�?�»����[���}j.�A��%)N�I�Q��6����ӎ��ʩ\�\��m����Z�)��ݑ�p���_�n��<o��E�D*�f�u��ǁEo#�I/ ��d�k�ݡ"��l5�WY�{2n��h=������[�4?��:��%O���p!��9߲$�� u���c�zU�pQF�Q@�N���������������H>�P�G�׏6F�b�꫉V�җ���o���}=@u��s��޺���%��Y��%.�}N��Rk{������>�#h ڿb}c�"���>��<P�2햰�74��=��T:�ҡ���*0�+E<���Xz���
=f����/.
7[�10p�}�KIY��%�P���Wp.=Ӫ3�n:9F�� L7*�KWv�(=��[m�o���W������H��_���9����l�/�'��u8���&�� ��a:7EO�s:.���� /���|;!(��]��6F`���S	�L�Ea@��n����-�`k{�;��FJl!#��#�Ö���خ��'����VP���-j�}icrA��@o�&��7��pӒ�e6��M��CG����{g���w "�
�vk64f�Kl�{��\:*J���O���J��U-̐Q8?����
:���Q���Ҝ\F���Ε�Ƙ
�B)�6VQ�A��Y��,Q#b	�Ŀ��َ��+�m�t�D>��]Kf����MOŴٛu��W�-d���J�T��R��P��)o��Iހ0:��5)3��K1 �0��w�ã!�9��.&Pㄳy��?�F�_4Q9�"�tq&���سL|�K�!f��yZ1=`��A�z��� �4��1�J�%���5?����D�j.?t�a�U�u��⠁���|׫�zG�-Qu���)��BV���l�m��� r�0[P&Z5�v��z(���A����R��A��?�h3�s:�+A@�������J��U"C�S>�4��dh���y�=&�zBB%����N����.�����;���݅�C5f����\	kTm(�ۥ��g	v؝f`L��+Ώ+B���7����~4����x�ڨ�z���jOM�8�	���>��$�CQI�w���o?#�y�Q+4?,���]�k��t��7j���R28���\�<������O�ZXz%�=7F�(�?A��׾�ƪ�]�Z{*��ȫ�ы�����a���?za]�FZ��FBԂ~5"�ѩB�?Q�"�K�-ZheD���մ�#YJ�D���]_/�����!Y1)���
#�T��nҳ��o*8÷�������Z�с�s�t�	>Ф��%��a�[�͠�K�����?��i�$�`�u?L6'�>Fa#3�aP�	ă�B(�a�Ǝ7`���PE��P���"�z��4��}������S�b �XԴM�!0����V<��<R�fv����r����a0��_8ޯjy��F��˙�v���ա�u"�ć@�����xL�{�讹��>yiZ�������ii�Se�?��>��o�ܭy3�5�*!Z�瘏h�M�Q����hw��Sr���"�TA{����U3��|Z� �z���I�?a3�9��d|�P	f)�`� _���NwYb� �Uւ��W�K��U2�IE�6�鳂���ȱJ�!� V�S�Gp��8��N�0~7�e����Y�h�OK�^L]��2 7�Ӕ��2BD��op��m���R����W�*=)���6��<W�@�k���{�$q=CϤ6�!^u�G����=W���a���B-2D�6ꁛq
���&7���V������Z�e��>�ǞVN�ᐃ��R�FD{r�@�3���6'�F"��62�B.�0R���gdVW*����5\�����{{{bI�YH)�����Ǜ�s�l8�B�	�D��"U��RJ*���]Q?�el#���-�v�"ˠ����P4)]��Jڞ�[�6��9��>���xm�,~1����!�ɨ�TNGN�O�Q6��wp��v�\��� �;O�.+�d�!4�%��6�P^�)�F(������lc6�U�|6��mGϷC�:�&)J�����|mVX�� ~��(ģdm��~w��C���8�d`��[��"b1��1\x�@��*Wl�x�]{�義׸���c�H���O��!�p�]��)[oule�� +�l�0�,!A4,���j+���_� ̦Pa����Q��Y4�"{���絾�����GwB;9|?��bB�R6�Ã����|� j���0�=��v�zz��� C'�!��7��h�.#iF�ݰ�i���Se����VP�XR�w
��ߖi�L,h�|X�L�ƫ��O���L�J��y�/V4��f�Yż�8�C���Pӳ��Q�\?��+[��k����G�ۜ���ׯ�n����0�%�Fe�!�0}L���nP�:�{��վ�.��CU�u&%�Я����$��q=�0��xQå��XҊЏ���飀	�ؙ���+s��m�s#-�D�������|�"=����*뽿s:`�9���$�GF�,�љf{D��̿�� .��W�|Y��>�a��e�Z�<�e����&�'�O�V���RԗG6�D��S��5��ӵ�����(R}�����w�̤�	A[\�mۑwOsE<_*xt���~�����UK¶L�tz^����IGU�Lb���T��t�y�m�`^?{�k���d�,|[�B�����1`�/ F��DV�{Je�mۗW��ZM�R1�-yx�v�a2��]����u-n�L!꽇���Z�%��:�5ǔ�O�5*��ޒG@�1D���1L�ͥ~u�=�xU���yD�XM�Y��M,�N�|���]��-d�j41��e�L�H1���ۜ�?�+uEN<et�	(0��G��kK֒	=凵 ΡH��P)��x(�.̑������sIC]Ͱ�T��ό��U]p�\�E9�_��k�fx�@E<�ӯ8��[΅�·�W�5�:{¾ߦ�DZ[���̦�8qn�ZL��N�0N~ﳍ$y$�Cʮ�m�N���BHo;����z�Qs�r�z��N����t�#;���,S5��'`/h�Z^�ҹ�=1�y�V�ӊ���2�j��I�l��0��ft1�L��5{���Y*6r�Wd�%/��+�}����z;^F5��XPL����-�%|	ļ����Dw�ʋ��k)t���i~���R�2eq�`�$��BBB�̔h��b$�z�T�CP�C|�a�x��ވl�j��Xo����ɱ��T�nJ�F ��4�:,�3Kf�� 6ҁ|�9�:X�LJ=g�*9�H]U��&I+����=���:M�u&m�۴���ʢ��c���,� ������Goi�4�I��u�ywg���-����m[*>�*�ݛ�!�-z�eq�Y[�Jb�$��K���E����i�Z��p8eӋ=�)jt:�#��˄<M����:#\��=7��I�d�]9+7�$�#P��nW�����bP],�8�-�	QK�˩f�xd"sc�����_��y���b������� �����q��w.��Ίn�*55�A@?Ñ��2%��#1W^�%8;�-�_�\��K�bA�$�?���s�`>@�bb1M#�(��H�z��b�l��G�k������� �-��Q;N���K�ٓ�~j��J<���8Y�V���]��ޮ��6�l��X���݄�,�%;c.�A؍���	3��`�
�H��=fg��b*���8 ܰ�Q�]K-R"
�޺��4�oR�}S�l�[N}�iu��S�"m�1o�n��-�����ڀ�����i���w��&��=v%���n�4|I�l��BNx6��aaP:�.ƥ�E��ƻ؛U^���?���4��6�yTJJz*���r�G�CC���p^)��۰���2�Tŝ��F�A���W��`	�ٟ��a/cxC�%�xB��\#�������LN��D���^\�m#���8�K:�G��9�J%*-�0N�/�4�^�Gk�9���-KA>��$������>K��a�q?D9����PE|n+�����u!�v3ZE�e�a�۔��1��J��6з!�UOM'�X�����4�e"���.ޕ7U2����3�S�R��w�~�,sx������=��~X��0���|��.�Y���S����sA��m�i<ŉ�,M�x���9� �E�)��F�_�S�k��}�&`�xb�슓�'�(�����J�y�1�}���F�Q�c+�_��а>�&��e��e�^v
����k{��	��J�k�B�떦Dڥ��;����M�a�Y?��M�ql:�����i%ix��|�
��@��d��}s�5��T�HV�5�Sf��:p�ȃ.����&�d�K�:!I�/:�@h迸O��O$��E�ը�.,�,T����W'�I<�ಟM�aS/�N���$�ӂ7���?���b���U���0�!��2��C�Mܲo�w-Eܐ�i������.�v|�t"4֡U���m�aP^s����a�������$�cƕ\Y�����A���������S5W���K&U��L���e\�9�H:^��`�����A3�¤4��D�z$/���כ��vM�Q0����K��5��]�o�(��/4�庌�K�C�!@Xa�:��5=
�h�gf�6a��7�&۟d(_�P��.���i����jh��&mw�0'nh#�ޡ�4�������h�,o=	����	)$&<���C�H�fդU�&����wzX�Q��o'�W�< D�p�W�Ȳ	C��L����
m�pw7�C2��fҲ��N�p{���"�J��9.t�W}��D��(�L�kr��S��}�+rs
��/�K�U�*1�K �Z3Y�H֮2b��^�n���nNb
�Ɯ��j����PB�8N3fz�����4����~��ѧ�I���w�ӥ���2T!e��㉺TC�[��ޛR�����O�BsOһ4||_'��t#(UZ�H�u��:y.y��揞U�e7�l���ޚ:W�m���'�*u�w)c�u2�AS��Sx;��"�]'�bB�o7�Lюvj�H��c�Z��/"E�����k%�Okf�;� YNW��%�o����n(��D�r��t�z��C��C�g*��Pd!l?���?;�F��n>�}^*n��PM)켎ZBɩ��O5���8򭉞�� (���fݙ��%�HHX�du.��0��xP�M!=�b�<�I�oln
��}k��������D��\�u�0aJ�Zڸ7<��
>�'!}?'5�)�rS{]p�X��p.�C�jE���ҹ�����,m�'���
+ء���H��@Y�oȌ� �x�&�'�X_�%��Aӗ�Y�T�m�/�;��Á�"�(*�FW�4g���>%�R9c��|���']a��q�#_96go�g�wˠ�^�����eґ$�mG^� �ۛffd�Uh���&�ϝҦ��K��[74GSb�_�]����R�>��%�7�IkvAʴi"G�b1�:�$�d�#n���ǭN�8�������ԶTV�C��Ֆp���J�V`�ʃ��D���N��q;��7�P쩨���H�}���b;�1=$������Gk�e6yqVn�p-pAA�k�����-��{c�ô��e^/Ny
C�+�?�t�rɮ�9#�*iU�b�b��N��*g}��ڞ���j�gz�ފ̏����5��n�Wa��I�)@k�T7�T:�U/�=hSk�"�&H�i�tC�U������`S��U@���Ę�!XC똉S*�q��T]�Z�96&�������yO��䉊���-BL��Y֖��>Oz ����U~��l�Ҙ¼�5�d�萌iG��q��X���#�=�LՋ>n���נG_���s�)���W!��\�A�h�j��'��O�d�¥u���1f�P����.��H?�<-obi'+�����2h��&%[.e���;�c��(9ndt$ׇ/>�MjB�x$��z[/��]�rL���߼>�n��b�yӱq
�q��i�@[r�aF����ݮ�V%�^�V2$|�4����N�|A�8b���(����w�k��3��2][�&ΊB|����3���F֏F;k��� �P�<R�zR���S��HhMM7��Hh��8^T��	���w0	��U����w<"��1<�*��&�57눺;|�l��m8���;¿'"N���)��y����� �v��"��|7s�Su�(�7�ʉ��q�����$W�ʜ��9���&��8e��W�X�O���d*#	�7\�|;�Z�Iو��J�A�����/�}nw\'3?��!��I�>�$	�	����wX�h�Y�H1ڽ/\��ݤ������$�e��2V�U�dG����<w����ح��UУO=!��YY3߈�7O��t�Cn��h�ҏcXU�KuqP����g�y?#aD2]�ZB����(`��Up՞�;N���N�ߓQ�W���F�C���z�9�>Z�v�,��I?��8�`37jWGW���R�^e$�!�C�{徳a�!�LV�Ni�X���'d���"n�ճ���	`��F}ҁ.�>���`Ze��gr[��Pc@6���ሓ+����K�9�~�T&�Qq��n�]⩸8�+������x�L_cV�U^K���l��"ߔ?�������+s��1����^�L[�ˋX�e��k���w�9�N���	��P� *�{s��T���O�ZQ���p��<�*���&�.���0՞�)0@ޫW�ni@"<$Uf],e�߂Tw��~4���'
�R� 6�O9�Z�3��ޫ}/�[�����1�wT�)L�!��}y��CH�A�Qrۄՙ;���z���F�B<5�H'(Q:tT#[�aa.����s�����}�ļ��.����o��B��3�֊��/XpE�j���-�~|�qM^L�S�b0`ē�.�n�wR&���볰�19?�VY9T���D>������v���J0Ȣ�闫$����͗�,QPk����Y� ���<�\�O�<�N})�Y�	FR�s����e�2�UR`��x��!ΰސZ�ܡy�c���#���u�!R�s��v����y^��"F�)"�:>�В��|�Ա�H }��>��s4�^���޷R���g_ʦ�H{+-�: �%�OtO>�b�}d�Ȑ���9_,q��5��%�X�h�@ˑ��u�<�u�n%�������<�5SV2��\Q���/�H�qU�mz�%x�4$�(��j�N�x�ú�bm/Jf������ޯ��g;	I�9K(���q�0ۿ{r({�[f�@�xe.+߶�Ee_+X	��!=�n��ި�6�+�4U��V�.��vE�5����_3#��d*K){L�����@P�r��vY����X�k7̇�7����.uMv�V�Q3��ܢ�=C��5rծd���V�i�#��	�g
�dV�?�r��������%�����L������	9���o/쓳�-��X�ca�r��J�r�X,���<��|&�rz���D0⊥T]�+��&Ӛ�vHa����A��� �j��3g�wt'���s#=�=��ڗ�Cv�;k#0H�KNy���O���+��W*�7L;b������F�T
�j1L�htT�͹v�Z�5e�afB�ת?k����Tv'}[p�~w9�G1Yϕ�u��&;j���%����z��r�]�������;�?��kv��pL�Q���"�UN�5,n�F�Bd.�LuZ�&����_�
��.@ѿ�Ʒ�K�}����طw���\�=�o�����F��4"�EAw#�8=���Y�y��PUG�:j,ե���XG]p�ɛn��7_���_��8��P���
�QU��q�1�z���0I6�p�64"���op��$O��q�;��Sx���ȸ�x���p�7��{��#EÉ�W���8��%H��C�w+3��@�e��g��4���
�.^~h^x�����x��=�Ŗ�:~���}�e�X*A��=T� g��?�,��koz�<U�)\]��^��S�(r�|B��("2ʩo q��.�=^�ӆ�XP�@u��8���k�/_��m�k}�ndݖ^���w���K�A���Zԁf����D�p;����s�}��(Tj>�w~��CB\O�~�����m��k�D6ׯj�ZN�+:Op�s?��Nr^��r��_���勮���!pͦ^��қ�x�X0o.��z��V�o�6�c��<���g�+�8[��R��",�=7��ࠟ�rt_.�v}�a�P�)�)��:F�'��ӊ�"��8�dkߝ���4Qa`�fL�0��ok��S[�3%��E���n�q�Y�n3���*UIj��{~���<��Q���d|�!�Dc�=�o~�Ee.ӑ�S�\fi�/}��x͋���v2��:8M�(˜�y�0����X4��;����#*�yee��]ﳛ`��H�CJ���Uw��4R�Q/�<Ƥ��~�b������b)��A�he�W����np����aQ�d5�`5$\eH��L{d�vl�+�O��!n_���42�p��+p�!KKWtn#�� �p.,����Ԇ�}��N�Y�1~L�\������t|�gc��n:�����_���Y|s�3�f"q��N����х��x�?�~j����-X�=�>`)�� �ڰi�L%�VJ���4�U� ��9���P?0y�X�	�X�Ԧ��6x���~w�b�9�o���qH�-���x�?�*�[����l�(W�,It�hɢy�~z��k�>p��f�*a(!B|x0�n����_���>ƫV��)�;M��t��ID�.��kjNf)n����E'ϔo����>�ݝ� X�{�>��;OC{��;vs�V4�]ȩ���	�nU�sd�;ǹYI>��j�.��ۮ�w=����y����1-��4�H�g�V����Rh8�����q�a��m-w
�߀]���Ɠ�de>���w���ZA�ԑQ����Da��p���������}��R���wb��Q�0�:g�DP�����gv��{: )�`¤q�����F�_�?{"�=uD�F�шI��7��I��4{�qL�}�ët���ߋ���g�gy��>��w�����F��M��G�ځ^j�a{���2�ʱMB�[y���s��n����Xx��s�vӘ�C���Ҁ�YY�W�nٍ\�[�)�C4�-�WXԎ;f��K��g=��m"Ƈ"ć>U*K>��S^8{|�i��������Q���x�u��/d)���jx�ًNNu���
�4���\Tz�:ё��>r�{�r/}���ð�eh ��Ƈ�$�yw�,��5�Z��?vS��vKT���]�ܻR���Ʈ��W��@"���{�z�j`�v��p�id`ut�e����Ne��Ͻ��F{5�:R��U!C�q�AE!��}=����VW��+���s堬S�;�tǣh��c�h���[�­6�j���[E����b9�����K.�Cڊ�W�^�?>v�T�����Okҕk]�����Q�̎P~X�5!����q�%�w������ɣ0y�xp��z�����5�<qU�A��ԩ���8�}��v~�,\v����}�C���~ �7���6�74NҸ���cMx�1��̩��ö�m�rъ�֊�{̘��|�#��*m������P@���g�+N��ԣ��s�dR�:��ip�7\^�!ޟp�ȮC��K���4GX���w~�{#�(��q����7bt��C	�R g�r=�G�R��Fߝ"��r�t��O�<��������Gί[{	[�,��}.|h+��2���󽲋�*���G�%c�����$�{�Ф;Bh4;�3g�ǒ=�᚛W��{)�u���]�=s'�ѫ
���l�7`�
(��d�6D@��#C�m��٥�ỿ�eP�%���Y�4<j�fL@�D�����Nc�9�4�j�F�ڍ���'ᦻn}� ���g?�RtE5����MW/���q,�[�������1
�z���U��u�}�{�]�cܘ.L�9~DO�Lo�� �1�pI�-�+(�������\���A߃ˮ_�}��A[̓)8^����)�����Vs�K?�͉w8�5��yN�<y��Y߃+�>Mw�Ÿ0D�.B��c�g��8�sL"51�#e��11����B=m��9���?�f����H�F���.~����Ë�±����&�튌����B�Đ�)}W����CvG�'IX�G������OExL�{��ض}=���ۻ��u�b�8g#�o%`�G���~�(����vx�E����jh2���s�|��+�6A(�ƽ�ދ`�7��yT��3�Oר�Q_�S�a[����o��=�E�.�w��/���7܁��^��ә�r���R�B�xz	j�輁�Mou��ghL�0
�C���")ǅ<mm{hթV?�)E��/���ߊ��v�wd/�[�{���Ω
��'{;�o�����s�A�m�md��|ґ��*���O�k�����֛B���$�=�{�]�䎧���}�ӝ��$%�q'��:����?"�ޏN����A�ˡ	߷� �����}u��u(�n�v*���`2N�k&	=z(~�"7�I&BU��R�ix|M���[�0��9������-�7%Y���2�8\p�W����G���E[TAڤ�A��9��"�u��X�q;�X�w=�zbW~e���?�b�cqؾ{`�E���Qž{�+W]x�#1�e	��GZ�֊���x6��3�����W- H�hb�� ǎ4�+��!!���D��|�t(ȸ���Ku��[Y�ՖL'T�C�:��\�O}��!HP|��Sp��	��
L�LP[��!�4����/͑�qZ�k7�q�?�PډP½�7?���d�1E5��8�eHhL��XӋ�V8{=]P�����xu����~�C/ì)�9�b���b���RH5uT��PO�P�xr]��|ꧭɭ!�����.���4��v�*�whܤq5��V���ސ�$�e���ш7�}�4��Tn~����M�뿠�I}�mIzT����w������}$�������O�Jk��1��D���SIddR����A���O6��O�hD�|ܙ����q�1{C�w�"��4�C�#�#m�����R*�4H��S��΋@�&��Oo��O��׾}������^Y��|����#c����#��1O
E����{����пϓ�~Gg=d6G5$��)$�U	�?7$Vi��@��p��Ko@��e�27�Ou=�9�w�y�����>l���c�+SExp��G�Ô1P@�8��O�Y����-P�ik��������U��(X��|�=/��v�g��:�NYI�����B\���;JQ�Ȫm4�^�w���	n/���k0���p��k��J��&�َ�P��D}��y�����!�^��������S�"0	TQEn�*5��@��`�����b/vdΏ:6�xt�u�����y��U�m��}��fSI!!��[���&6�
����(v�w�V� �P�* �{o� u�����ϙ9a�黛�Μ~73s��{�=�}�y�{��9|�l&x�0��y����ö�޻o�oZ�'�mk2<O��PN�E�������O�Q�������8����x�#j/x���?h;dI���/F����������U�Xb�קK���m�Xo1�)���<��r������fKZ�&�W{p�O��k�Bfg=��Ǝj)
���֐:�?�#�R1��I*d�TRk*۹�F�<�o>|\�O��=���o��b���B�%�^����J>�ʾP��T���?}Έᄗ~���a��D��z~�8����4�%e(�JH�^�w9�*��}w�%Wqy[C;ö��_~\�B-�]Tb��|p9軾r��� ]es�W�ᯎ��*�����ǰ�>; q��4py�:��uRo��_b�=���;n�	���A��ȹs^�57?���1]�PpC��Q�"�]t�炭k����z�O,�ʂ��N)P�L!�W?�0\��0�,�Reo8x�Ãԛ�9��>�0`Xg�KMW�����^1$2$bhgn?փӿ���(i�5<��ǈG�_-E�["f-6u��"r���.$q,)�1ևJ��,Hp�#�����_���xi^��#�p��1W���t�8�K�O�/��S�!C���礦*y���Af��$��=@V��;(v�$���?Ė4�|ܒ3��-b4���.�ĸ��l�\6��P�z��Kn���E���-K�I9O� �㙔+%�mz��".tv ���ݱ�ޤ2�F��G�P���P��(�H�$�t�R熈� ��&��F2Y�ㅹ}����U����.��{v,*�$F1"v�u'�u��Yq����W<�����R���3�b����C
����G��0���g�[��pj9eL�L�pŌ��,���yg����ٙ��6\50��*v��Gġ��ŀkR����Hq��'���Ϝq�<����Ҷ�N�'O9�E/��c��
�V.Լ��
��)����_�bI��I�]X��ʙ��+n_�&����e�܏�c;0e�TQ)J�������"�RI�ޗ��>$r�Y,�K��R�Î�l��oz�iκ����T�Χ�A�^�#�j��<d�UQ�%���s-�0������[�#�������u�}�N��8S��"��ö#)F���dv�v+����`hG~��wI�{T�Z(y���~�ӻ�Әr���8�o7�� w��4���l����Q���#\�IX��{�C*��v#LYg<n��i��Ȫ/x����l��DL;q���)#�vެ3>������L�*:J\�?u��:tߝ���۟�ӸƸ��?L1#�#�]���c��{=�[V�VK�dZ���9��Z�T`�&���S/,�'d�qn�aI:|��ÐF!�:ƣ��k�&*�Y�*y3��c�;[e?�<�&H� 7��(N�ܯ��������������w�;����O�
��5���J��.O�*/+�	yN��y�b�Otq�;4]am�z�(F!p
p1~$�u�>����Õ��ǿ����֪��:�b)Ár�|_�#���R���s�1�c1m�hcd�1���� ���`���J*~GǙ�(NY^�B���ōo�R6�|��R&F)�Mw�,��#�"���^�Hq}��fn;mĖ�r���%x������ܩ�3�4����YpľZH{��r��=�3����u�4M�l��)��9lt�.[������/�^L�_�^�q�0TxE_�à+bd��v�xy^��}���""��<���q[c<��'�V扱�Z�p.�X"F��*ݻ1�rGo_?����o�P��چ�u����7���g��G�N=���(���XV������aY�{;p�8x���3�4{�0~ �u�*w^���8�(����Zq���G���[oy��^��-��Fd�`qjNF��2f
�\��m���9!��y��7��g�<lW�	=�,#�k"/X�H򅫄(fy���&W��P�K-;{���I<>�E)#,iW�A��=�Ql�I�#���z�F�x��7��9=U��631qG��A�J�WD�ܡ��-�
V���v��;�ݴ=�����07�t˃��=��X�m+�kRys��0l��k"Q�s�Q�q�/�ڃ���a!$�'�֟օ�/�k��=�D��{�CXv�4�F!�E��C%��9/�ݧ����3�:0�,�u�?񇋮C��)���t>*���u�`�bX�!�Ȱb<�E��<$չx�;���|aC�b�w���PB y��\ZՓZ��,���p�����.o|���~8����	:%��#�\���%0l)
��h\�;�`ch�!�L�p�*h!;�Ø��l�5Jy�p4�yő�c����*%\[�ҥW�W�LjG��TG.�h��G��RV|�?\���夑k��~O����FZ$"��	j��x�_S�1���E�[�~�q�ē��nr*��(�%ð´���>���9i?��f���܁��s����8Ͱ�$#��� ���Ĩf@1�.�Io/J��P��c��e.E4rˁ�y�������H�1�����N���W��4�#FG�ZR�q��\�epb�>��?_~~tޕ��1HE/QK���!���~���h��^�NI��<|��#F��dX���rA�u���s:+�_�x��"2`��>���<�諘3�u���j?x�	T�q-�ZR�-�s�]d��Zv����1�)Jl�m���Ei!�ꣾ�m���V���t���\�
w��XK�p͍w=�y��X��káM!7����$�
<���SF��9�)_�=������,u�:�z����H��GF������=IX�D��n�ZY
�#��+��{���Z����1U��o8Ķ�I������Ν�8�HwH�Q��f��c�+E�˫�ᠷB�K~��e����U�TR|�����-���~�/}�bL�"��6x}D�ђ]il-I�4�B��rFO!�;q�i?1)v�M��s/���T��9C�Z�^]��K�<�-y�X��7\�Y�-ǆ�'�|M�`{������4S#~�Y"��_���>P�Rs���I:���G8*���WufJ%�D6Z�:��>l�Ն�K��Bՙ�����u�]�:�p�-��}�K�[�|\�&z�T�U
�h�zy�B�G�^d\7��Ȇwr��?Ƽ��L��e�d�P�͘�EO�K���0�����_���N:n�#e�$��|�a�QqÛQ�O��s�Y���:麎c{mHE|���蚎�õLi@ƹ�""I�ѣG��TV��J����9�jx�g~�zۙ�gn��6�%�Z�e������1�j����z�hT�[��c?�C5>R����'�ǋ��.�gx1":��j��Z��M�]�t����^i�R�ަRmQ;`G�mm���ļ���<lW*�Z-B1(�ed,�_sw�[�˥�݇�J�TShQ|��.���}}��m8poy����Б���n�h���)n�����9�/7�a��Ă�5<\�Cr���T�M*m�/B}�ݶi|kd�v�O�}qEݳ������W�ݱ!������!#qb)x��i[���u�C֛Ե��6.��c3_����Ϟx��D�%�~��M��?,��?j�ZÀ(��8S�\�*t;���`�¹(�<�E��� �?�Ƕ�?�����$��O#��QC�C�TB���dP���8��K��<��/��6<��˪s��,\8�ʣQ,t�9~���v*qV�#���Pjh%(��r�r��,)y���U+(����V#�7��Ј��J,��^n�rfJ`�M�+E�۬������16���iSǩr�JICt�yDf>��'ۢUe���O� :����y�H�xp[y^)w2I�}v���-�{>z.z�*b�˅"���${Y2GW��P�X���*�0��v0�[_8�c�{'�L�L�8<�e���Ͼ�ȢS���¢cgV.b1I�+k6hl���[E�؁Z%D����9G��U�g�zx�'~�VXx���VXo������r?�ջ��r�+��$�F���x�|k��Q>�/��Wu/�#�/��H�=)�Q���*�8V��ް�N�bm1F�����vȈ ��c��$GWg�-X �����~��m!,�cO�P�����i��Ҡy����]�4�,�kH�������;it~�w�����ٍo�:6�����$��R�EזF%�Ԫ,L��ga�ѣ
�3�U`�p�G~���OlE�Cvz�$�Gc�P�#͖h׷b��`%����w�E}K��*������}g�Ŵ�ן:z�8�vf�e�ל�7b��ni�y��G��P��2ĸNDY���UƢJ�w��iH�Ŵ^6t�=d�-��#�SD7�3��C��ۜ*�:��+��_�p΅��sF2�F��7�E����7�\�i8�����\Q�+i"���G�����]BG���<�:C��@j�
J���n��uN�Ô�Q�P�ШC9�I�N劜ۈ�P���m�׉�6>�=&���gg�u�"Do��=F�iC<��K�|Ɩ1���;���"�m�T�!iZEw����2�����CZSAo��<CK��/�|Y��v�7\�{ϙ�M�[�%͆F�?ƌ����Io�/�©tE���Dj1}]ӥ��zc&Ū�5��!E��E۹�Ki�^B5vq��~Q�sۙ-6���pl��(-�c�F7�ƪ�!+C,�l��>���I�g^����<��^�ϼ_�8ׁ��M��mi�|T�I�c�m72�k���n�b�9RH��d�<F���F�!���9=j_;��k(e�P�SXթ)���k{j��u���Z��&H�_�a>�hk���ys��Ѷ ��w>�l7ǵP*w�Z�A*�V�<�:� tLw�yK��>z.���QnfZɡ���e�*@��{Oym�'N9r�1%{9�T�kS
�t��{_|�!E�f`��\��9�GŨ�Y��("����f�a`d�HmIyKҳ*BJ�B$���>|fCH.r��3��A�h�"8���q���Q�m[V�X�吏}��R�?_/b�/H�[I��$Q�:�3bv��}�7���v�.�2����uFI>A��JX���KĶᨸ�H�}P,�g�m|�M��=畹jJ����M��JM�44�S��E u%c�0��4�v�yA��EFx����h�&V*"����T�s��4W�u�
�(����,/��y�������{CW��#v�䫸!q��໖����C䔙��yCk#ć��ް�u��[��]FN�O*e�=ᣪ06ln��Q�2�eV�5,�D`�H-P��-�Q`��$D���+�.�Z.�G�:��%�mиbl0u��OqH�9�SC\�(��mɫ���.��g^���V�&���t5�4���A�ƒ�Rx��*!-�R.3K���æ�6���l��""��$뇛QT��z\K��F&�HO=_m|�M���ĳ���;�f5i�$5D�q�
#@+�t�,����&4�dhu��>�d����g$p�**a�q՗Z���ymV^�Gg�"�]�HŘȼ��G�Tl�W,ODy�aƴ��7Z�V�|�\�sց� u�%�,{ņ�Ħȃ���'u�a`��Z��*���""i������Q{�#���r�ٌ_K!><�Y����Gwԁ�x�;���\J
B5�GGGI�q��9�؆�s�_�TA>g�Ub�"���Ǚ?�s�7�m`�<⠙p84���2���D��;4|�K��{�������}P�K�6HV����E|�	
^A�����jSHRZ��Qj����G�4z�����>T��j�����Fz��Rs��^�e�����\E�Q���dqrcm��}U^x��u	_9�@|=����*�����_�����/�����(�ed�"iW���Y?�0�z��z�>�6X������c,����ÃNi����g�vLZ}y�<I��(�9p���{f#�b�lK6��@$�F����S�d�E��7��.Q\W�v�e1��$�X��>eJ$-}��W9p�hA���p�/���֊0���~XA�փ�{2��s~l��W2`��$IP*���M�[�m�CI��)ZϤِ��X�o'x���bK���̠vL�1��o���ϼ���i]�i.��ۯ�Z��Ϊ���;��>lc��n���߻�����&$���
�9��iXan)�0�����io}�h��䳩��F��}�|��G�zP��ێ.���8����ܑ
)�G�5�>GQ$b�)��G�4v��'�X.��ˈ�n��I����2hXIL�P����C��vj*���::��^�PD�ީ�h�r΅7�� oR1&�z ".�C#�K8���T^{��.�o\��aDS*���G{	�f�����X_s�����4 �Z��|p+w��gC��|�H}���A��r㔱v#I^_G�4���N�r�=V��q�-� b��"ì�+��ԧN�q�ah��$���.�[�x���/�(�f)�5��k��w�l�n���Ac;���eS�dy$"絆˰�� `@1�T� t\1d��}�%U8%�<1g�{�r�6�������/�g}MX�k�Z�ei�$��rI۟��ϖO���(KJxs�U���i,�*�}&�Ma@R��F:NCd6�	-45�s[>j����*
uC{М��/���گ��zci��}����:�˃w��s�l���jR�V�8k?�5��{v�����!3�����([{d�a�i�.��`珼��z66���f3b7G1�)r���a`p�N6pt�uP��Z12�Q�+�~�|���޼�vj��Q��Zp,&�W9O���q�"�<{�C�5:�Ry�E7I:�;�W�Yr4��gҲ!e�"�GwgMS%#�Z5R�X�l0=�g3Dt���bY� L7n�j��~�3�#^/�y�K����l7liGy�:Mө���q�Q���/�u	�y�C-��KÙ��١��5k��.�Ѧ��x؛$�w��fN��񵈘u;�x���m�$��r��J9�����D`�s�bÀ�E8����^E"m���x�����W�bD�r�1u4���$�!�Bձ!f�q1�(:�|?�vC{�c������Ҁk�3�#��l�F����r���}vݴ�=�H����)(�u����x�����$������	���5�Zz
�|�U5���S�->�7U�2�am3���TQ�!o���>IiS{{��-���'����@ZU�G��5�CK�Y���Nұ%g懎���bܰ�0B|��j�������4�J�n�v�(QC/�E}=5 ��������<^i�1�����N̛ۇ�|��Y�e��	������\��#��u�3ye@�~���'��3Mx^�F~�m��mL�P�狁i�k!�߆˘F2�z���\��1k�!�ڀ�� h?!�\I��V�0����J��F������uT鼠�_m���X^ʥ�*/�>����]vjYX(uN;r��砧';��DĸahadL*z8�=�]���̝����2.�k#������'�iw���cZ�V_�� )!NĸSKi��5:Q�����O�f�ˊ��g��g���5�3,���p��T�@�!�+�Dd� <b4pPΛ��77���x�?�F��`D�YŵO}F�ϸ��l��n?4yl��ԜW�sf�$��Q��������#�@�1R����2i| sM�z��Q��p�D��UG��O����C���+��]p��D'( �j�l�� �\�B;0�̲�^�e��>�D���8�( �=�R�g���N�Pyvμ�7��NJ[��_���^I��ޡ�jb'ӆ���R�@jṵ��Y(%�G,�TtP�L;��rD��a�$1>�!��aƞ���xx�M�����݆�"�
Ȣe1�I���yW���z�V0iy�l��DTh_��^3��y�c"0V��e-z��̳s����,�N����R_v��s�t�����d5z�z�z0=8Ң�s���>?W�7�>O=�<�W�`~�#�z�Nm�=S�pЭ���qc�փ|:��!�:�rvL����I���W���m��_X�_�w9��W��`�.�,@*�<aG�-y�5f���Z��s5p�$YgGGa��}�Arx�lf��cr�g�N�L���]�ܿ���B��a(�m�viR�88�/7�ƻf�l2cB���	k�Y�mA��ot�z任ʍw���/�Wr�Sr�\W��2�S^,w��Mb��)�>��S�Fu��?�������]]Ć΃}����kW�|f�<v^c��K��;h�I%��a��4��L�ХV�P���Y�I����z
�y�{��v$���ƻ���.�i������F{�<9'�$lZ�ްZГ���Bgp|O@2v��w�k�� ���ft�b����=K�t���L���	��X+rm��k���%\q����G+b�i+'��&#�]x�ig�lyt����EUd���Q>ƛ�c�N�4���BDW��U�9s�X-�o��w�~�8Q#|��j�Si��QX(&���5�ۅW�.�˖�!��>Z{Jpc�V*�*(��h����ڀ�fn��E}(uWj�9���O�*�%��\6/�pQ����ݙ��\~�}(u��z�&y�TL	F��,i���CE�0VC �+�;M�\��Q��ǽy���)�fFŇ#��L�-O}�>��l&5��XKy6�;�����G_��Ͽ��װ"�5'�[��\�~�h01����ܺ�a�2waK�T�C��r�OD�|�h0���Gѷ��f��7hF�>�n.B�1��y�b7���x�=��`y���¢�xy^���b/��x7@D;qv�v�khax�3��CP(��w!����M�%�e�^R91������ԥ��?ތy���x�H-k����\ջ���r��JH5����P,����1��>�����Ӷ��2C��k�ɛ�?v��w�nw'KI�۹�!��0���bQo_��_��<<ʥ/��v��U����s #�T���U$b8�'��%b-�uۄ�	�sml��$�7Z��6�M_<�IA^_Mᵥ��<S���W{7�Z��1c+�|��a$���
�X�2d�R�Rl��m�o��Ö���]�'���b0;�>wJo�H��?��s��h������:����`�,���tVە�L�v(���i��}��gKW|�A���bƘ=�T)�����5CA̵mO=��=����`�'���	�o:���޸��>���'êఛt%Pk��rύy~˥;)Z>�+��S=�,��h.�>v���G"��J.�|"6�2^��v���n7�usj]�S%�(Ƶ��M�#����ݣ����[n{@��k#��v��'��-7��Cm{��łܳ��	�	K��b�Xv�<�z���\q��F�7�����z�}�K�R�T�6���Î 8�s���\��M�q����g��w�����<�!���5Ô����3&u�,���\�$�"�Ւ8����g]ܼ|�a�㕜�ݦbs�� cR�7��>%�8�mq����ut�VBC�ˊp�~\���9|��Ŋ�;>G���z^8G�)��>�6�?�?\���m���ې��d�����q�n8�2Ճ�1�j��]o�K��v#=k�mԽ�9�%�������rP5*>�\��a1����?�<de5�.1+��Q��'RF�߶JO�ϥ(��Jv��Zy�i�=�}v��S�ɆA��M����9sQT�d{9"��v
�c�8ɜ�P�:�N�A"���_��?�J���S��ӗ�tĤ�]a�͑0�Թ���J��(2K9V���bl��`A�<k'A�v!��O�tG�Y�-Z�k��;���u��n��,�����I���)>\��Σ� g$^��U���z07C����"0��d��1�i,yD�K�{v���]v\�!Z��.�O�˵���� i e&
a�%��Q����9��CE���a3�������QPRuMYl�T�s)%mS؞|�����}���IZ1-�Tjn������g�SY�Ӎ��7���7�Ur���J�������l������f�q�<���a������z�5� �p�É=A���a���n������Յ2⥗�J:��Y�p�clYi+�Ӻj��MڍL�z�Ĳ�".q��`��y�;�~V�y,9���#�z��,u�s�bn#�|�뭜V׊X8��3Ւ���4��4R��,�c�Fρ0�q���ܺ�������#���]��
ަF¥�R~<��4�:�`�Y3�_lAN=�`�jU�q��/H�����rD�d>�Z*Y��؆�;ʶ�*$+˭�>����.�N'B�Oy�"	U=��QB�{�Fq�Ɨ�O&yԍm/����9�hٳ�l+dXiL6:hzw��-߱�F�gV*FK�ce"��٪1��fF
J5�!������|�W�G�~���vc��'%mW�����خ� �Dx���u{���NCr��Ѣ�~��(�s�}�
ܖe�`�c���eh���K~���euv�y+5��jp���������qA����-�GE|�����wWi�dCA�ֳ~s	l�C�Z��g�lGyN0o��&�����2���-i��rS�v�R�EF�v]q!�R5j�Z%���B�.�oW����ai�*9�������z@G���Y��=T�̘5��d�78�c#�3+��Q�����}�9Fvw�f��A���{���uP�L�(�^'�s���@���F��\�M:��w!������,�z~�2�qD��d[%�١���1�ڭV���&ʘ\ш��ް�aa�="�J�b�4a�9{X�J��h�f�>��Q���]W�?FR��w��B�Z/1�Y!p�
;%TzH;��N��=���m��/,��!j�a�t\���✗JQ�N�����*6���<hs��Z�����?<;���/�E����S�f!%�2ߏ�=��l��t�a*}�?��P���X͖J%���>�U�<5�>I�Ai�}���:Ǽa��d�N�Q�#ć֤S�u��-[�����E���Rk(�\8���NԢȜT����$�EC.j*U����ŧ9���9X�T�m��i���b@-?�"Ө3u� �>~z�?Q�:˗|_�x\z(Qe��S�������Y/D-��v�=kc�<i���T���2��������p��͟��[Ȇ��9���n�t�0J���;sٱ���MD��8������ߴ��c��c;�w�m�=*�#�;"lyÁ[ꍢ�#���c�8��MÊ`.9����[�jj��}5�U�5W���fCm~�V� O:�;^���6���G*����0���Q��b���==��<�zzzs��G���h��H�y��'���;:;�����._V��J�K�:D��MD�6�5�M��<�[١��v@��Q%F�v;��Q!pD��*���'�u��8B1`��ֶ%�����Q��	8�3Ǫ�����7>}���� I��[�V�C�y׳���Q�nZ��u��a�`���_oC�I��0X��>�wؖp�$֟��!~��,��F������_bx?���[8���"��{�hm�X�$M�" k���r�)/+K-��?�3����Wj��5�U(I�F.y׵��� ,d=ކ��[4��rx�l�м�U�|���g~��ǹY��42�rC�F�/�A�E5zB�����a xV�0��?\�W��kD,�,��q�\o����sC-;�<�曭�Oj_�CG���P�5F���餷��~����
Pd_r�=�Ľ(�<�r�&��yv�Z�?���p�(�|�>���G$����6�1Q�#BM͕�l.%T?��$�^a�۸�[UZ�恻�y^PW��P�R擀��99V�"���a��q���G.,/�=��I��B	��*�'J��{�� 5Gn]yMC|��˷�_Uh������:�T,KZ��C��""��ρ�W�I=�8@)2�兩څ���G_9�]��\wЈ�b�����y�~����YI��nf��Ӷ|T�k�8+�
R�f"�#3G|�"(O?;W��hc�a����+�����NJr��\7�21.Zac%�{?x��xbb���2�n���V�O��&9>Dh�5��yA����9�h�6
N{�-�e_���2���ܔ+m��(���}&���5���v�%�m|���|���Z��c��&��%r�V��&�9V�U�;t��ς;�{������|=t��ܳ��>���%UGp5���m��`�����_h|۰*�����G��SϣV��Cҙ��@�SÀ(G!L�[\��4��]w��\��;�	�I�.����%�����{���?�ꩮ��5���}��ʦ�cj��������V�ep�z��/ج���\�K�r�J����;U��}�R�AUO˲�Xn}����$J)�39�[W�R��D�mzVL����ڶ��:HtU�o��!���"�WO���G~m���+�)¢w�Ѻ�3�t��B@�H��Iu�z"~��9T�z��y��,~Y�r��؈L?�OK��k��R�נ�ϤqmG9�x������j�6��rL��lֻ�+�Vպ</O��5�a��Jqc�rȴ#��2B��q���͛�3m��4��/�Nӱ(�F~�l3��~$}�ѫ�|Q���ᤅȺ��v�,"q��~&B8�7@.��Zҍ1�)��d�w��mC7ag�Ԭ����\eXv,�U��2Ĵk�3mocUy�hnG9!L�Q���\���l���Q��"f�������&��y~&��b>ƺ���l�E�+����5L�:Ň�R{1����Jx��P�aѦT��"���ߔ����AM
ٳ�b����m�n�8�F
�>gY�f���7�Y]_/ۃ��ŏ��� S�r�ax��H{��n����Q#&��8��>����T`��0�'Em��bH���Z�Z�mB����ؽ�
i�I�Q̛3w����~���~*J^B+
`��r��4�󇽭���<X���J^�W*����;WSi��15e6:f��L0+��{�Hr��qV~r�I`���CI�TǅIO܆!"�kl���4�D�	0�N�d�N.6I�5�	�xF�)�Ԅ�)�������h~�ۄ_|C��ѹ����3�����e�*V�>_�~*E���3#��f��J�Z�"�}+�R#>����q
�Fe��������P��PF�'|sQ��:\���������0��-M��!܉��Y		��`3�i����Q����
d��V�'� ����H�9�����~��0�c�!��x\��/�X����\��
f��1��t<�v8�㵻lh3��'� �.zv�&zC؋����~!����W�?2��%l� d�_�{�ⰸ�yh=W-SG���#�xjU����]�Q�+U��>�^��{�Rk&[���9��YZ(!5���˃j����M����s��&���&Z��τ��b�ϲf���ޱ��
�D��$��ݡY�zq.�Vf�ZߐT��R 5~�&�� =V1��\u rq��|�U�m4���{Ujj�]�R�w��c��Y� �/�ux?q8��q�`�Zu��IGZ�j� ?��U�l���w.m�q�`f���d�E���y�Ԓ0^�yA`��	FK��z;<SȮ��9��* ;�n{�<��h}D�'�w�7q��?gb$��3��Ǒ�/��>@��R�а�j��/`e/�v��0����h��)GoQ�F�f�|<���)+�de�T����.amM�fPS�M���~������H.� �6<�4�/�	�F��H�+���as�
��][H�y�X�;_S�y5�ȿ.'*_~`~���V?9���o�t��p'�!�K����$�}}ۀ<g
x��3�Q���Èq&ls=0��+?6��b����D?���uY��y�Ű�R�1u��3#�����ߖɀo?|�J�j��ױ$�:�>��_N�o����e@�`��ͯh"��+=�����3��+T`tW�y���J��|�����9,S/��S�9��M
�*;�1*_D�G�����q��u���&@p+�<3���;�]\���P�[p�1�Y�U�������AI�å[7��J����v���9U��G/`�ZI��Võ�y�Kţ}�j����ǩ�E�2הR�U����*҈@������M��9�p������b	HN�D.?�>�u����Vٹ�K�	��!y���M��#]7�i�ߞ1T�>R��6�h׿L��uJ�H��/�2�
�,]vM��6��$2���g��z��P!������f(�y-DE���#�}#*83A�=-���%��)z�π��8���p �D�P\-[U�i�&���͏�%�����ac"�H`��[�wP�W���<~B1�6c|�.ń��-�=o��7UmСZ�	~�rld����9��L+��_�Nmq�%���x�U���<��h#�Q�9����U2��K'K�]��-�x�	�w�]]��8�o��6a����0�[� ����X�ҮQ�a� +�#?�-�H/Uz:��T�c;�W�!v>0���RZ�0z_$V��]�$��c9�t�\��:��UbV� '��-���%M�8njy��^ZG��lS^���*�y��&9�?�^����(�P�"�LϨU]s%o�}����ɔ 1S���Ѣ����L����
r�rf��W^����L��&��i�	f����2ii��T�g��[2��Q��������~�ϭ�0��p؆�߳�q�?u��������5��]�=�.���������C�Hv�螮	V���A)R��y�N�+d���G�}�;��4k���͌s���rP7�|��� K�	')_<lʁ�*�X�:[JI"ڻ�a 2_�����q��C�_G�po�0\�`��@���Mbt�I ��>���y�J�f=��>
�����2��*h�}��&��7R"oXv���`D��� �DBiK�IB.��Jr��"s�q�-��
ѹ�d4���Z��a���<vSM�n�RQ�)�6j'4LI;)��䤐.
|�S)�̚�>2ք���
�K�����z��E-z�N[�S(��n�J��hh��o У��M��T�4���2I�5�u���'�� ��K[��U��&V���~�b�j�L�W���|p����Q�� �}��5��z�P�|�6����$r���-��A����B��x�P��/�����~Dt�{9�j%Z'[*o��ϢX T�PZAɴ �.<��鑇�1m,�ǹ��ͷ�Y�6`.��O���M}�|�)���y�F�
:���@�m只L߉eE��W4.}h=o�����9���	���˞w�m�W�qqw���3�:�9SH�U�ԬɇK�#�tÉ������-�=Uq��Vz<r�_Z��F�H֤~��ѕ�)�>�K�ƞ��	W�c�G����&�s��U綈��~�~5N�{T7s��j泵�9�K�3��0�����QY0*�%Ә�e�0(�WwFN,R���-�om�����5;�C�;�Fd�7�a/0��̇��3e?��<��J�TQatZ�gR�Oa��fA�(�3!�y�Gm�hL#�|�>2��5�#���jՅ��f��o�Άu�M&��|�3V�{�qa��^szJ �{�-�2������3tL�jѯ��Ǔ�q���*�h��yޛq����ݡ	u#���7Ɯ|���3/��q�A1�T��֋+�2�ۘ�,Wٕ�����i�x(zd���������l��K=�8�I��*�8Ѕ���⪍Ӈ����2`���;X�<���j�oJ���4z���/��^��n�7��BcM�թ]Z~-;U�����Gw+�)�S}"mp 8�����l���w�{f���h4_��W��:�b�w��$�0C�	����h~��6e���c=S$�2H��]�By�Oy7.h-E����3'PB�6�Z7��I��-��Uh�NR�zF���m􌩋�"�F�$-��S�a�?t�{���߬���QH؞G0��9����~`q%���W��y�-���Gř������|y�sK��\	��Hի�u�V���brs_j'f�e��.�5�~,���c�n�ӽ�5\��l�c��<���(��Ia�0��u��h>�F]nF�!b�E�q��:��o���JҴ倞֗�C��|Y3�
f���XYX�z��|(j�q�=��P��zB�G�%J��v��^x��U��&�}d�W��+�!e�-jL�j5w������I�Xը�b}�%ض����W�UT%��ҧ�9 ����/�{�A�c�p����	}��;�
�$��T���9�ɴj�@���X�q�fJ2:�8��ߴ�~��	z�t��d֣�O��G|-��bRsO�H��1��As�w��З0� ��]��O�\�"��pլ��!NtTg_�k��2�M�6�B�;}�۞�_�w�sՍ�>#j�U�X�YФ3z!��ą�F|H����8Q� ��~茪�.XHW�g�Ny��@8k���Ϙ���\\��X(�AՋ F"/�'c��K����2��z�Jilq��I't�戥% �?���Њ��o��m��'Ғ�o8�?�(w� �__{
�A�Y�F���߾���G��*�UE)ey�ھ�y�'B��eX��CۅD;�����;��/��i���I�g�1�)��(i�V�@��,��9d{nr�q�\#����'B�WM�<�77b�Σ��XB�N�}L����_�����x�2{�b�^��])f@J�d��}���,�~
|zcu�����3c��:�?8`6��0V�f�'Wa��Sm�]�"����皃�N�^ٟ�8�ي�Dm�WW�b�DFo��R�?����GVo����9�>��z�}�X2p���ʡ��Z����ә6~\��x +}E�1r+Vd����i�w����pFo>p�c��c�Y�hCW/�	�G==U��gz���m���vP�tz�]�͂niM�f!����Ѳ�������c����czS+r6�?�9���Wr�w�x�IxO���N�<I�_��^���k6�jC�O�o�q'�.F�X�.濈 Z������b\䎜�E��]z��������U7r0kg�k��$X-R/F���g�חq=Po�+�h�x�2�!o������gw�x)pۻ��AFYr���3{��%ԡ��BpRdBe v�UۑRx��~W��,���Մ��u���ׁ���%Dʼ|�33���+ٵ"��]�i��(��;_�v�`�����r4���B��w����v����?����{��/��_�N���a)�C�$׈��t=��ޠ�Ve؊�W`Fư�g��~�Q ��d��9�����͸�#QO1�.�t�������#�!_�gb3����RF�V��뮔�T�������
�l���s�^zт\���k�@��65��������Ᏸ��Z�\b��T�` ��P��x�q�&�z� ���N���kC�{*绞���u�>؞���6+��s]|��F��&Im1�iW��"�#G��ht��s9�t����<�����3�#�nw�`�,y�C�
ɸ�$�녩WV&�S55l���O�?�O��A�Q0PdgF���q�2�6H�(�0f���a86R�X��%�&���˜[>nJ��{���I��=�z��'MR-ؖM�����bUC��mQ�šY�$�䱟2��>����E����~��(V1&�)�y#<�����m��쾧�I�5w�?��5���Nޱ�M����<W}��*$n")��"�rٶIl�L�n@��0U2���h��PIv��0�O�JE���0�<�N�];��$[)5�V
MU��NH��OH�Sz3h�@H�u�,����v� 8�<�;L���'�;%Z���&2%��V5�wĹy�W��e��W�ds�S9����22�C˩=�:2/5~�@@bH�������H���yLt��9:��9�H��5��{Q���I���l�L��r�䁳���_>V�To�������o��'0���+Iw�V�N�f˽P���*ֶ�N�@q1:���'��NqW��� ��ٚ��˳�~��'�u�4	M��~PC�������@��ýe�&���n�>����	,�����{�o\4�h	���T��u
�I�Ս-Q}jqR�Ɏ��g�f*�8d���qXB�zJ�=��i}�}F�_t���1l��rz\������^��а������*u{�H�?ݝ�`���Sƶס���5Z��Vo��y�5��Iɾ�Z�A�sS2zZ�:Ֆ�^��^��B@x ���cלѫ~�tl�͗8�7��z������L��p۫ek�"G�qY+����p�w~�p�N�;��tb����ζ�!��af���J�`��쾺�z�{��l�^�#6~)��M	�����8�):1O�ӥ����\�;D/r
�n���C�����a�u�Q��m�-�)a�Ce�Z`�s+f><YQ)��P�p�됗d��I�ܴ��Lr��I�M8��G�?q���+dn:0ۣ~�Ӹ~�*���Y|�=�C��f䍱�1��Q��I@�X�R��(L9#1F�n������r��3	\�V��$^Edf����Nβ���]��rK��X"�(�b�1��R\���;y�{����3^� �"@i�f��$��l������LE8�#�'�+Қ� � ��n5�v���ɋ���cn��Fe�/�d�Ա7$����"�C�Q���I�#��*ʎ��,�b�荔�C@HD�%�?�NճG6�R"*��֋9�xȊ�˹"�����`;4L=��m�&�c�.�K U��"z<�/Q��$dЕ��x�Mn���[�qŒ̛�Mڧ]C��âZ������=,N�(/���D��
ʻ��T�����;c��鼰��C����Yu��� �\U��Z{o$�{��7/����!{�x*��'�ۭz�����j�[�a�QŚ�P1�_��LM�������}f@�H�L�-�Y=��y/q��������y�:\�L����D��:�rކdh��@�+dKv� �S��%�ng���^�R���r�Kf0%,oS0�q�ѿab�M�A_5$��l�$D��fZ�Ly$K3Txsf�}"��M$	�}T ����:F��-�����=��+�l�WԷY<�,\�ݯ���B�ޘFQ�����{��p�,?�8�)Rg2����� ��9��4��D����bp�%U�"�}{��nD-�^]ݠ8C.q͠�t�W�*��	�q��螟��q��Tf%��)���H2I�e<X�.�%@2
�V�ȉZ���A=����K��J�p�}oy�B�*D܅��ʶ4�-�z�_������"�%d�7nkf��*��/��-�D�����JӮ~�:�XP�[�H�滎b��+_�H�a��~�%�B�O�Y�S?�2�I��K+r����U�_yە�0�&�##���� �� �w��*�z�s
f,uDPࣰ>�8�9n��m;��~p��������F�wEc'�\�Z-���7��H�!�G�w�gNmQ>=�#h�7�a��o�ɰj�Wp���sf�ܯ[����΃�#�����b4��J%�D���A=�K�<�����%.��}?��z�P*����T�R
@b���trD�s�Dpfj+�$�U����(��L,�Y�&){���.RZA�v��%rѯ�����!�%��%�s��OsD�e� ��`?<�UV�gwW'�x�5mD
V��	f�q�;��J_1�|g�g��Г�� ��n4�hDZ"�S�!2��k/~��ƔUR��@�홿�(CM.�:`�]�<��9���j�K[MP�+2�C�,r-��8�]��[�W�xNմQ�\�Pn�B)�fQ���4��g<�{��]U�s&�{��윬������<����a��c���q�s�8��	�
y��FP]� 
P�0i�jc�<(�|���^�������bM�a5��&��t��eWHe�Ll�6���W���_v���74-�α���d|�N����ٲ��Dz~(ۄ��ڵ�Ӡ��[x��6��z7e�����q����
+��^}1-�w����mm &-G���DAPb��˃�˽��W~�c���0R�C�f���F�����k��E�	N�<'�l�"��6�,���}���N��Vr_�hMy��k;���F;owk�*�l�Ng%���ח�'
�Y,�a�1���pZ|"A�x�aб��Ef��a�Pq�xm���ۃJz��t���ۿ��7Y�@�^�eJ+�4%�@ȥ�bǲ��>�K������O��9;I{AoLB���z,A.�^����C��[~o��T�&�ާ)�������!��J�`o	U+^'���k��o���qidtr<%:���d�.�EΈ��5gV��Ʉ���r�]���NZ���+�f~J��&����3���d��2!?\��}�8��j�q�?h���Z&���:�mT�F*ߞ A��A���R�.�A��>Ok:���4L�'�௅���)�h��'��+O�+�Mw�J�UZ��D ���k�{ӷC��ۧ�<�	�1f��D�A^[8"�Q�[�#�&���n�Vp���_������*�o�]w�!��38����~�:W򈤵����gfQ/H�c��E�ʑb�[M�2F�h���=m�'�k|`�Y*��=�Ywn��o��l��̓y"��Y��>(W{4�h���QE�d�������x����;n�8�!�;�*_y�l����Ze�*�;_þ4t�����_�zC6-#�#�>��B�-Xғ1J]�U�F�i����O�E���ׄ�<�J�y*���-2XT|���i��D����bL4�^"FÑ/	�YQ����
��i]����9�B�Z˕O>��i�� ����>tm�	��η=o�[N~eo0'�����,��,ZW-�V�$��%ZM�~��I�^�����˸ǌx�6���mO��G.�f�����LU�_�!�@��H϶Z/D�Z�F�r_~������}/���N��ɣu debW�V���L�k<=Z(��7��xn��T��/�bA��xa��7e5�6$X���s
*(�RI`W�B��\����w�H��rp���e�ds# ���x	�1gHC/�`g�i<�p��Yh����ϕ�2��_��E�|�S�։�8�	M7Y���Ӯ�{p�s���2u�ܖ*?�$R��}�aؼ��vI��L k"H�@W�3�Q���H��XMu���G�s�D��G�8����g�	Kx�6t��/rHP�('\����D���]�m���ٓ
��6V�mI��ݺ��d��a>&�$���,�̜6��L�����=�IBL�ט^W�wі��m�����"�[�?��گ���q�3o0�Q���lh�H�)�h~QĞ�pc���*���C�����$�QT�>�B����"��#8L�"'��b�Zai\D��s��_���;Ԡm9��(�y��K���T� ���`��V�=�E"���� dM8O���<�����|ZCӰ��I_��Ɔ\��"d.�9v����:�
����fTz��N�Z!ۮci/��}�ߐ��΃t���_���7�H������y�����J��]���K���E&-�C;��L7����2g؋g�~���~Ӹ��&J��p�ۅ���^�$�z����.C�0���X��4�)L���c�G����6�c��y��{��K�S���*	�\�m* �-�Ƕ���Dǵ�|.��5�GlJ��:&�3���t>ysp2$1�9�(�����v(5�k�1��x�b��E�u|M�ݕ����"^��8�e�|^����A���>5�W�$�p����=�X���X�����cw��}��=q7��~:Ķ��\���'jS~��l;�W���	��w���k�0Б%��soU��E�;���Ԯϱ
i� Eh��# R�ۼ\,'��4|
��ș�ZΛ��7���N�41q���l#u ��MW3n�����Y�����Gt�s�\~��b�Ό��b�$�%9E�������R#���Tk�N�2�˩M��dt�BFcEc���]�ЄYqSw�It|��G^�s�Y�m��z��,��~5l��+I�SP��7�3�x���OW mTc���ʚw�&�5}�WÒ5�bˍ��=�g��">�$G	cѦ�R_XA���.�ֽ6 �jt�{�ifX���	����Q�I�#���n�;�����Z,�P���+M��E���h+�m�*�3�;������6|�G��VԑŅ�<ȗ��;�g.��̍�7?�E���rDa=�O�c.qM]�DLE%��XY}?��H�LR���&aI%���la?l�c����Ez���
 ��=@�������G�T�y��N�ʄ"L�<Si��[��g���0�l�i>Orj"���@v:t���Q�����f1�r�b4�� =��Ec)���aj��1]u�_L�p@��`n�����y7ˈ��&I�\��j-t��h�����Q�:�L-��/���0�	m8�_U�u���l�2��E�1��v��D�Vl�sR^�K,ⷩ�A������(���Z��bc縳����Y���;_��� ���Ɣu�����~w|���i����$��FDS��5/�&AY ��m����0aֆQٙ�A.q�Z;���Io�K%+��.���:�_�t��þ������ﴻgԬ�<��(�5��~�6��u՘R�$
qi�4��Y��u��n�
�5���g�5��z+�����]� ��2(�y�Hd���Ș!_�{4~�R}�!�a_2�;-�Y�S��8YSp�F����C:@�c�����		��Ȧ�]mƢ�{{�J*I��\��K�O�q�=��+��e~���;��/iˉnt���%8ű~�w��f�cÕ�a�D���:DV���2�)�;�S@���b&��J'tY���N���̢1ߍ�d�W;��֎������	)E>��@��tbuA�_v��l��O/���^T܋D�{���@��;�V��|�q2"�XŅF�������j�_6��/(+�>l��S�_N)+!�M'��N�ߓZ�M�ܝ:��-im�5���gmx O�>��.��U�I�7�ˊ��q�������zڿ�!�G��'�b-�}
�K�D�G[o7��P�]{�kf8M�ٱʟ���#��B��e�q�n�х��u	(�:��}yE��ݸБ� �ŵ)4��]�7UR��q��_�G�z�d\�?��B=�}�$�l��"�r0s@4��Ԅ������HU".�L�/M��������ʨ7���8͜h�t��)���_����T���v�����HWq�7z+I��1J�o�����'7��F����ʥgO�"Oh#�A[cg��w�I�]A��ȘnϲP���T�Vy~ts�R<M������|�kTJ�_b'%��9�^n��	�~��#�!�)r-�h�\��z� "��v/7�'��Jr�?,�{��-zdP��¯����dXz� s��K����hF�h�`�ja#�T����ǽ�ӞM��$_�ƹf���ؗX�h���4>E$%a.r��}҇��*L��D���m�5��Q�Eߢ1v���D�mo�Ġ�b�u/�9Pp����	ђi�%���AM_�~��r�kQt����+���|CޖTxg&�������J�T?@c���+L��OjH� S�ʁ!U�Yo���S��)��OXo~}�����᮴�]w����|��D�#9�s�b���?1�nOcz���dӺZ���/(��G	�֖d�a�e|/s�� *|���3'챵Ԝ�f�~�ƍ/AwK�������H�nE_�A��.��@��3��̸�i����vkS��Ob���5��CfҮ�P�:�;0\��>��pJUN<R���t�ǧ29��	���C.y0�c	P��p�܋�t����R&G;H�������j�}N����5)E+6�Y�&h� g�ˑO��4����G��E���5��;��	%mS-�I^�c�w䇪.���t$�.	e%�M�Q&KM�q�'v��H� ���H�:;7W�E��rk�XÖU�)�^u��nC���_�;�������ƷJ�cU@�	�|�lۯ�'�4'����N�6�sG�Y�N\Ͼ�3���c�cc����|���=�:w��T�SE��1P�L�߰���vqb��,`l"ݖ�D��j�C��	_]7��]�9^[�
�IR��W]w8o������Q�o�W'��)�㣏����u�"[���
J)1���2QY	h���YB�����`&Mf˼�o�%�6�4��a�;2�?"��ھ�4yi�U+�J�8M�nG����&/�����%ȩ\o����U�2�/n�E�C�,jV�ڠ��E��B�w��p��\�_�nv��ӧ8�s�J��R�#� -�<X�W��^/S��*"n��n6洓�~�w�̷�Y7�D ��lc��?��7��&�􀳖Q�X�)�N�(VY���%�sQ��zYCMeq��h��4����>m�>�ID�Ӵ��/#S� ��kԷ���6Af����9���j�	F����0�T�YfcԬ/U���w"m9^�/To�E���
9�a.{�Y���mP�m����!�o�Z�vG��ث���Y3}�}Ы���#٭�`ö+bH�����,km�/�٪%J�23ڽ�.��ϩ&���Z�����	�����H���u_���`��,�L4W�����P���y�x��(z��9��A,du��乛L�x�T��0��#�
��LZOr�1��|}P�b�ˣ�ط�%�W�0���TD9Ł �.��{���������u��Ї�3��DX�$�4k�6��|,�׬�,f!�X`�g(��P���[Y쏹�a�2����jM�fu�D�·Uѿ��OB�/lK�/���5���\`C8
��P����?ˣ
��v�K���gƛ�����̌BV��]m�]mk�CsW��zM�Wn�*��'��5�r6Z�5����mߞe�Q����Rb��G�7wF2޶?o)�ҳ�"�{*�:�䧦hޭ�����0���a[�&E�~�r3u��,VDS���_�=�*D/�^6�����ĮoEQ����,���핞F&`�%��j�9?�'Nh��U��Go�bY����~t<��?��}�֧�;ś��������~,�^E���h`�|"��wj}=j6�.~mL���P�,a�M�o�$E��Ԧ������Q*e{>�-�&Vo�B4�b|�3>��e�0�	���^�������~��l�#�|���-������ؐp�3]8t7�[i��xB��]ť��9%��m?�M<gy�-v]�ޙΗ�1���-��j����(�����`��TG]���I7'-�:��/9Tq�L��K
%���K<E~�� 﨟�Y���9}T�d�@t��+gl�7�k ��`�\���v��]ǹ��9[Q���u�<X,�rҊ���՛B�N���y��e�a�7j�m�9��翬�l�q�}�F��u��r�ꙵH��9�Qlإ�ΥE�aM�M�.x紞3�ӓg3������,,y	�Z������y���Ϗ������`�N�lQ�����yq��Z��v�\^.��������6��jr�U3y-n��˗�3xK��l���+����c�1d�]���k�q��1&�=B���f������,)�8[����RJ��1��F�0��Z�u�G�끛�c�|�E���ȩ��f9�k�a<�v��,9���"���@N�:��B�?(�m����E���Tc@璩pտ	2����0c��LԢZ�(�jQ7��t��1`�Y�K34˳V��DaZ)Ǌ>�)~I���� k�D��x�kJ0I7&0�F̣Ƿ�ER��\9�A�T_����t�_���3�8b�HU���mƹ�(
u�y~�w�q�d��	r>[��ep:B�u�Cv�(/5f��-;s��zJ��s�<ℝ�|�A��.o�G��J'~���|�������؊��N��c����F�ab�X��p#�)z����EB��"-�i����e	x-�F���>^E�57GNj��qa���̇L*�|RF!+���HQ��rŶ���oأ(lf��9��Ĉ)�?�X@�0`���|��\A���sI�=��x|�!zV�5Y6W�?�Sl%���e�ݯ��0J������
X�
���MǛ�DV���4��!Gg9!���<��μ ��M^��3�nL6��֍r�ܚ�ڢ��V���s�������Ϡ?���f�=�v5��1�@Yp������zk���ד��/fF�T6����'E�v?`��E.@���=Y[��n�_��7WJ0?:�*��ZoG��C�8`�۱<19U��:"�`D�D�b?�;�&[�M�9���_gM��m��{�}�L�>���|�_X�IB�{���qf�
���jk<���kci�����{��]ko^BWsfh?��ǡ�-�.���V$��_��W�7O�?wx��`��(���ȋ���_.6���v.���q��G��[P�眕8�L�l�?��r��t4�L�|δ��m2铐�[@���i�L����K��ݸ)c��^d��\���?�Q�v"�뙖�z^��hǲ=�2,�F�ط:�kK�.�0��\4�fQB���P\RZ���)�nH���TUg��I-�
p��{�B�v���X}*Ÿu������y�@//G��D��o-�]x�x�T_��㖺��r�`���y���yFSg�4uT�r���z��,�F_}��߃c��.���ܯ�+H΀���k!9��[�Y�f�TA��|�=�����ÊRdƩX�!u����7�V�-�I�\eZe�BO��<����H��hO�֊�<ڿ�K�
c�+5�2�B����ǈ�E�ȕ�<:�m�������u��8���%z	����d�k,���pam}o�G�eL�kI���ફG�&l�'���3V^Ͽm�+V�����v�PY��O9f��7\#������@Ԛ�ԧ�#?�.�<��v/�o�x+�{��9]���a�U����/\�23y$xX���+�'�C����;�h�7�D�_:N�ؤ�q����p,.`P 2/>'R�@������l5��%��R�r���5'����E��eG����&��pP��^�e��V��5J�l{[�m�6�VW��ϡ���Ʈ�d�H��Y(U0V���^���$�ٵ&e����&ȗ!A`,I|�O�ΏJ�S�b�C5r<��qcݷ��&�M��[�YC��{�3�H�1ع��/�䇹
Z�1NnS`�\�w�nC�ʙ� e�]�c�C��p�\�C��@*ߥ�U�9���RlB��'��Iu��4q�͠���^C�x��RIZ��b�B�����q!	ֲ�քi���� /
;ɗG; �2�K���C*wq��B��2���9m;0uRsH<��pRVB��6�x�e#����EnL���w2T3�\����<���8tn��VFZ��QG��;��N�G����5/Y����1%�a��ƒ,aNk�q���أ����4:����ߖ������s��߇p5�v�;�G��*m3���D�i�y+K����vu���=vc#f�� ��������k�q�΂LJ�:`܏J����C-z<7-�,�ձ�B�N���"�җA#�&={9:�����{�kMk�V�� �e@��[����oS�ç��hv]�p�f��D�R�0h�UR�vЌ<i�v��؟�ˀZ�#���2o�h7�{�����N�+�i�m����2i f�&<f��:ޥY|4z�L#y�M�V0��@�<�X�o��.3`/!���j�rf�����ɠ���1w�H�L=m��>��|h��}�4n%I/ �OJ{
';+�ZT���@>R�XC�8NR�<E�b�
��SV�dA8�*���n��r�x�:ex����WwO_�+�2�
������w?~UV�Y���d�P���K�����]��ȸ&�2�/�i��^ϕ�v�Ձ�+�z�̽ց�g�%�R�O������F��Azg[��� bG�x��z�x�Bn3��1�4�"AQ�<9�/$���r��g��O)�W��&�"�h ���O��J9��||(���`�ٸ���������{>jL�V����7�G3��_�}ZI�r��;:F&'>�'D��N�bm8p�^ϣj��H�#�j	Q̱;0K�c��L�.�p:�LYޖ�CiO�U��������#�f��n����' R�SnW��	M0vt!,��@s�́+b<�ڕ�ާm��_SV����e��N�C���*_;���w�tM��c���I ��F]t�����bS�oeQx1e��c����ګ��kW�������H�������iF�'Ku��ݴ�~b��UF�q�}+���U�	u�������u2l:�ޛÙ����,�8�7P�ߓ��������c�g���xUKkV����jk�ޣ�����V{�M��ZU�w�{b�رS� "B?��y����<�|�����''��Հ�L�Y����l��M�a���k�^�����o�fl���W����bF0値az3�t	ظ+��x.�3�u'��d,I��~'�L_͑S�u����;�Oh%P�+�r� 
��x�Z}��@+@ �� �B*���������n�KP|v�����s#Y��S2��uRS�A`�f�K�s[Y����U�F������� ���c���� ���9��%XW�hU� �͹bǮ��'�n�����=ӌ�j����8����C&G�>���T��g9Ѝ����I���!�<�-����(�\�j���C�5E#f���w�C�C c`~�ۃ���0��8�AB�u�m������W@?"x'?�b�׫r5Ki�cr=r/�쓈Hj\Nw�Z0�u�z�L`t��9 �u�<����k�1<�/�lJmB�H��]\L`�?�_�����3�90ֺ��Yҭ ���ӓT�c6�t8�O�eTM8�������c��LWsP��cI�y�}�J"]F�&��3�����A��0c�NaP�`�b�����m�M�����
�!�J������x�#�rs	O~�l�/�� c�so�a�:���-Î��f�*~��fff�+�un?(�Q*��4@O����q�m�� �%7�ް�b�%���K3C�$�~���Μ������&�(��	M��#Moz{�Y;z�^�M�O�|����s�Twn�Hj��]I��c��3�d��"�LMH�GE�F�Iz�(l'*�|:�+bbB=9d1�r�҃��L�`�"�#�W�O��X�0x���h��q-u�x��OJ[J���p+Ώ3+��1h)�bW�0c���$�����i9țgq~2�si���!7z�+z9
o�_be.�+>ѓ�+@F��� �1�p���K�/�2��� �x���y�<��!n�m�̳��v�]�s8�������.F��f����5���dG>2�#�ՙ����^=a��#m�0"I6?�$5х۫8��\��3�XmTHG�y�(yd����B��9r�P^ѝ��'zf뽑�k�iʍx*����(�|�f{39�����@�o�H?�U[��<3<==-�K����G���0f���?0�!��m?lsp3��L�|��J�w��/��.G䢷���9�#lh>��?|ٔD���zO��@��BU�k����B�zgJ�\��vO���$�\'D7�tdZ97�e`
���W�����>��P��]M�*���G��c���$_�9
b��ę�밍[�g� e8�4�8���O����
=�q-B�@ ���95������E���zU�sac踞�[��~�T���[S�q���T���a���a�	��Y�C�}[_�
�c�c�@��ʸ��z�����O\ൔ�*�]�ũ��i}�b`�d�&M�ؒt�W ԉ�?�M��(�͵r��ߦ/p�ど���H6�g�g*|��p����t�O�~'vM����9��l,L,����h=�;�kߕ����*��`gN�>Ya����Zz��xS'}�f�k���BÓ��%�'�m9]����z�LRyl��<�z��I�����n���q�����H�~�E��E��Ս�v��/䳊��_O�3� >t>��H-���0�� ��Z7��<�@�l��[n6��2��K��}%����Y��[�mv	��l;y7	�S����&�K���y��O]�����[=(.?gt�&��CO�.��>W茂\�(�V�����,��H���&$mj3�Q��>wj^�t���x��,X_�֙�̄c,��n�Iɗ�I�z~'�vEL �G.!�������6%gnC�2o������GX�&&n��\6+&����]jF�>�~n�3� V��o6�X%@��d(��vy�mTo-�i�-4���%|�赑�4�8߈��X]��ڊ������"]��Y|a���l,�c��aÇ�y�a�\���~�����f�и@��'M~x��\	��^�w�n��F��1i,��2Gׇ1�@�S>���#�`�����&�#������囨�\�O+`#�pol�H��c��S�\��A ���m]�:�Q�YZ���a_'�	��5�.3sgݶ���g�v�o��Kj����f�R���O1h�U�i��قe�@�W���t�H[��2A��*��:�Ù��q�{�����ÒT�V�|�2X7����>�\t�龕�W.�Q1����]Ԧc�].�	`X�w�Ѭ��+TBrkp�h��7	L�F.]�:�26�.�)!�>�^P����u}2�=���Eƣ�{AD�_>��0��L;*���!�Q�Y����wL?��/S\��]l��}W�YC�ԃ]��%?��A�=���I����4mF�| �	��C� �N�Xr����L�'o��Y��n�V�����j��N�b�CNG�����D��$���C'��F�F
��O'J��E�
d����gv�WZ_�:
�;	�� �	�Ӥ�����MJj�(��ǈLC�#l�U6o�뵲���@��l4� �:�x1�^p�=�\x\�^��^@9
3�+
��^���S�}���$��oɪ5�{CY|\;��/Mך9^/�C3<��>����E��	�l���$]�Y��jL �RD��&��vߠE�*e��NM��ib��;`�������Sss�<_b+�h��G��c���������B�d�7֑��Fyj.���S�ܣO�1��w(xrSf爏c<��B�cBC�R�r&�q�'b���^���4�Tb0����o�4�N0��_��l��t.z �08��[�w�B��Ĳ���헰^�(ڗ����^��U��rTЯ��EFo$Xy�?�~P.e��:�kr>�Ǵ�Ȩ��m1y���S��i����E�$Zs_�Fs:E�U�t��dn�Û�}��\����,X
�;�����"e�eT�WM��%X��܊�� 
��;d�D�^����X�Ǉ����[�{��j�jxh��g3��
T��Y0#�t]�g�	��?�V�^��ˤ�!^)r���p&/�}k��.�yr$7D7��k!�,݇���qػ��N�=@�����V1����C�m�X�>�oMk����
���(��gV���{$Ǌ�A�^�#q�6�]8+�jJ�z�A.���M��͜�7w(������]|ÿT�&_�:�Q��d��š�r��xxlp��5ؒW~�~���������byL"k`����*B4�F�Cj90;�k����+1�o^�ƌ�kte�L�.Q�Υ�6��Ont�A�����(.@N������P)��%�O���-�Sm8�qxO�j|W	��~� 6�*�=1t��7Sv�֖u������+@�>�Y�<���7�|	Ϲc3�U��y��*laR�*���e˺ Z�}�ZJ�J�>?%�~�����/imߢ�D����I�ȜYޱ��ה�HJ����Ӂ�#���w�K�V_عR�	_��p��#�.t6�t��*������� �X�9�:���A}]*��j�@^T��h��$��sN��Rǁ���U��[���wfp%�#+D`�����Qt�z���l.�#���J��{A[4� �'u��(7�ƈ���_�ʋφ�<s1[�3�ק^��Ǝ�aר���q���Ih��i#�Q�����y0�=�1uo�s��h>�&����I�b��bF	g���Ľ|�DGZ�y(E�u�g��ؒ5�bm�cf�RnOhc��WQ&ᓼ�Q.��Xu�,�a�/���UT��Ѩ��B�k�apܛ�0�7�;-��UmA;؈d���������6�/&��Po׽�?����	�R����L�
O+��v��{y1���ӱɼw�%�:���/�1&���k��Ȅ�fVkN3cx��ʑ���e�0=�\/��g(|ɕ��mڢp���|oki>a2P<~�̀�N6$蓕�s�Z�s���(-��хb�H!�q+�t!����v�ٔKT��h�=�L������r������H�m�Y�o����O��@�[�*� �	)�
,Ydۧ7`c`N<#`HW[|v1u���o� >M~ی�t��ZM����|V�W��!ޒ/�T&���We�>�%=�?��Fҷ�Ѩ�7�r�:YI��}y(������jsۼP�5?D�:�HB��yq`] *Y_�sdK�'���Y:���T��SZ���ǎu	�l�#F ���RQ"���!�O)��.��w���*6͹�(x[A�V��u$�E�U]p&�J!����{%�f�1D�ߡ��^����,N��dl��{���_���z�^��z��.ul��-��^�v��2spɨL��{�ʐs��=���@��y�p��p4c9'�:�5H��Jx�S��|����Pg+�oy�̕�Y��
���AwsVsI�����4j�	;��¾�sJI�a63��ĭr��4޿`n��Y0Y���[:�Ss��j�n�h��]�_��a�LC��u6`�e�FN�����WrӘɪ�R����ߩ�m��O��U��L��[�U��f�`�e/�Q�C/���4�Ʉ]��ָ"�����VӇs/_�-[bA��w�����t��F�.��-49k���X�[����2�������;���ў������ّ�	�Y�/c���h���%;����e��r��y�?�?��Z���Dw�^h��V�.uc;�U��3j":�2��sS��Ԉ"���s*�I�bn�9�����Bjz�#l�)�Ns�)����j���|,iŽל�����ԍ1�����֡i��%��no�'�a�@>�2^���Z�0���{���*d����FS���3��R{��"'�uO�y�Ɓ���`z�0�})��8bƷ��%���9P��ķ|�Sb��&��<��x�R����e{���C��@�vT�%Ij�=�³�QR�Z�>{�?�NA�.Z#�䘁Ƽ�ko�"�;��у��MGޡ�K�.�k)cb�uƔ���U�m�&�6s���x���Wu�}����(�ae��OMξT�� ��5�W��q{:v��[�	�0"+0����s��A���KH/3@�d��1�
ҧ|g�h����VEi�Ds�M\�K�f�!	�~��?����U_by��IYȡ[I�Y���P��%������#�@y�MFl�bq��Z����)Ȗη��w�./��qf�t������q�ʼ��j?�:�Ո�ӊ����h]ۋ��C�,�������7����R��V,�菘��*�4:#מ��u3~�����LÛ.�,��~���0�P!���؜U�`	��(��v���wA5ݒr���e��*��,���m&�����~�t�߱œ��ɴz蜼Y~m…�#�������ն��y|��q9�+�,�3]�z�@'�q��"��?)?)����'����2=�	��n�g�0�6�C~���S�o� d�y�sS-�aoA�'��oY��(�6
���0�2��o}P�=:��CJ��u��\R�4�e��hy��2��0|JA�(պ�b;�.d^�,'^�ï�ԤC��k��xh����u�X���L�F�8�5�W� �E���d�vO�n#]�����h}?�JqYH@~3Y�ލ0*q��硢&����ǵ����N�Z q���ɧ�j�Pw�OF��n�Y�ߠ�%H=��?���]h���4l����ϸ�G�a�zon�V�#d�)nw�΋�n/�-������1���ي�<9(]w%��1�K5�u�9Ԟ���PߚU�����f��b˾�����㖄g��iL��g��?�-m1��5B@۹D<X�o��BY�;�Q�ߴdω��D���D�8�}��4������h5^�Nnc�����0NÁ��<�r�S�8=xL 'e@�F����*ne:�J}�Ѷa�����6�̔�=u��A�	�qv��Fb,���m�\�GV��`<?X(�+qd���Fԙ~� �쐇�o,��٤�iy�JG���j�i��Š�`��*Ens[��H!�?�kab5y�-���v���-+�1���Z�|�i"� �A�#���� A�z����m?���j��B����J�fL��6���x�>�n�����l����-rnhtu>(���9��yŽ�m�)/x�C�y���p�L����a�hN/i��G��指M���!�=Vq:��+��X�Ǔ�lᖏ�¤�2W�1�����+��_J�r�sLW��O�w���}r���.ik��#1^����/S^R�.�
B�+~�ݒ���3�뛌��jC����#^�a)F �i��S!��T8�}V�G��"���G�T���>)�4������3�'>�T�q�X���E�W["R���D+{�Tmפ]K�U=��d8�;o0�,��F<��mtJ����Go�����m��$�C����f���#{�,\��ݤ���_�b��b6+]5����Ql����s�BZ��>��'��r&�|2nR|����yU'�:���ѷ׶o�i/���D���`�X�d���n�c[���(����?��^k�S�`�+�V�;Ƴ��М�%�"�ߗc!ƥ� ֠�=�FqD�}��_�)r���?H�9~�L?�d� E�VkޫL}Y�X��{��3<x���Ђ�z�Q�SW(�A�$�<�u$��;[�J��\\���C�^n�F1*ᰯ�Ĵ N��_�iS��Rz��)�|#f�����iq���9�6Y�������W��ιkt�T�]F�s�����G�Y� ͱm��Iض���n?���h�A4�z��"��@,��-N������f�����9#�����W��٢����v�K|�Ț~'�B��%QI~ OA��<7zV"����9�Q(���H@���*�)��i�D�V�=�s��%�C><�@::meom��~�}$(�z��u_��IBxmN�n<@9a��c�/�*\*;�G7&+�S����M0;��#vw:��\�$֎)�E��U��U1�����t m�#�>��+�u�e'{���M��~�7��W>�%"�j��דR� r�U.v<��cW4��->u��A��:���g��Y�W������@
u)�l?]��^�yp���"�F@�@6##�2-��7^Y���/e��4jh#ٔl\��#�����[p<���Y���Q���S����lqLPٺ�ESȷmt���qJ���R�0I�cQjԝ�N_�����Bێ]��;N��ܗ��]�R�$���lmS�59�9�M;&�d\�2]:�8K�߲�����i�a#�3�x�Eƿ\��m�lu�����Ic��l���H%�`ː�=u9j�o3?(��{���|�u��&D�bI���2�<G �����.u��GD.�$#��h.���/8G'�}|�)O����}ق�ѺA��Uv�p����s>��x�e�XUd��׫�)��˱+=��^��>8���:��;�������Sao�y�˃f�Uu��'��Ҟ��A�Y�D� �ES3�����^
�ב�ZZ$�	8�>_uo ��9�-%�}ؑ&���ϛ8��y�pUe �^2�F.���x������~G�w5'nL�?�/M�*� ��X��ݰEm�������:>�
��j
�+ۅ�(Y�Do���}��sw)�og�V��:�千�@��2SQE��y�?�
u�I�)\}we�������ot� s+ᘫڱ9ĕv�¼u�i-�����(K���Ty���[��a2��:D���]ԛ���)ձ�b��e�7o��
O��N?$�]9<s��\����Ɋ�<[f���J�R��>�Q{r��� 6�~<#�S��o�T���sx�[3UI-H}If�v����usg{t����⤽�WnW�����<��#so�-�㦛Xz��F�� ��a��t��Mu�6����yi����sZ'�՟T��=���ю�_�~w� ݥ��^����/�'����x5�V%��ڱYzzU�Y��ݨ(n�Y�ZM*T���׭��|Y6�w7�\�/о��{*=�
��Wk�"�����
|����WN����̧/Si��o�B'��PHDAM�k�{�]w�(.�[ w�a��&�s�*73�{,$	��ĪY�� ��d�]�:��
͕1�r�>��9H�!��-ɍ8����\�:0��DXSҒ�Q����M=�=�Ab~Z,"4�KO�P�(tgn�D�KC���.�X���Xj�/�z�W����[ݐ��?��t�L��rO���
�1��jn J4#L��K)�cJ\��v?�6��GxB�R�V�'{?!�|k<�Qg���9��@ɞ-�/H��W@o:}Ģ|
��:��(*+�I�di�r`g�N�5df֌�	��I2m�k�ڤo����'y"����1�a1DV���=�O�}:�k��������D��gK�`�\�v��+��v�5�zK��=tau��T[ɃM?�9r��8�@9fz�T�k�7���_U��c蛧�lX���?���8�g�2�E��X���R
R>i����6�}n���Z�f}R"m` ��5���1��������skq��T�Tz�lt����"#��_�ج[��+��_,W�)��~j��D���G�do���6Wo��]˚emlln/z�6t�B	lC�Gi�I�kL͞�<�l�3�+��2y�Z��x����5�Z��a����b<��4~��o��[*�,����rȔu��O��ɱ�~�Cos�-_���;��wΟH��ϒ��p�w鿾����m�'�c]g��7�Q��0�s�Wt6�|Y������ݜ�ᢑs����?�2�dZ7��t���W8�]�~~�W�X��ۓ�y_Bɩ�(� s}��WwAF�o�0��;0 �UF�2��2W��~��h�r�<��� d��<��k����$�z�F��R�^�S��� 
�ZLhٮҏpd?��W.t>�u]s�JcQ���.�]��ݨ#�eB"�-��*�K����V簐=��o���g�)іl�Rv2��_��ː�9O���=�UX�e;�Z� Ț_V\S���%_V�	Y�bk��_��k}�펶�f�,;��ӎ��g%�����+��rr�x����G�kl9.?b*��-�)���5aM�GX��6�fujTw�v�j��9Jb�YPEz9ѓut�B����!�j����\.��g3.Pd6K惔�v�M�r/��}�Q��`z��A��v���<�L��T���Îg����5��y�]��A�'tt�) ��.(ȑ�A�RX7���~�%����[�_W���������1R��Q����vk�ONY�D�K�.�N�U@�����&�{ ��!����R�)���%
��F�j�?�����];,$�����!7Ws�Yl��ĥO%	Wo)$A�z�����}�
.�ƺ��9��g�j��Ag�=Zn�Y_,.�Y�k��&�H�6���b[L5n�7~�2 ������f�`�DĞn>g[�J'��M��`*ff��T�+T�-����n�Ǜ�ݸҰ^�7�U�m��\�Tݿ�ݓ�Y3}�1����&�ɫ�ޡ�4��%��7Ÿ�R��hj)"��G�Hq�*��Of���}񘓌���I�?Uw��G^�9Z�iW<���u� ��&Ul��ަ	����5�iUYQ�4Y�,�����?p��E����>)4���&ON��֞��*���y��uM�"���l^�Gm�a�:F�R�b�nE�}V�Q�q��HC�z���1���"�<Y�Ť3��3��8H�~Д9�L3��!6������2�k�.~`#��6��,�C�Թ��p3��7���C'4n�D��ޗ��1��e�	��-C�����4@>~s�c�|�,��M8.3о; 
� ��$�:ZHT[m��~�������D��s��:��>����"��{�*+���z�kp�`hP������Ёp�4��r���=���_ڣ�\��dk�+�!?�q�Fwq\Uv�~O0���g�u�6b�����L2W� �;V�r�x�"m+<nQe�|3A�cۀ�m�[��M0!��8�z�����]��.�An�� }iDɤ��L�m����ۭ�>�bu�����d�wßzd�WR�����FzvQ�H'��m� �R��$�zg\������7�c�$Ga�7��cn��u�|d��DD�2�;'@�"�i�Ƙ%�cɑ9ǎI��J�C����9��x������$h����6���S+�c�#��[�P��fGB"�"��Gv1�ے����5���<s�yN���S�$�c1��;{��ʎ<�^�����`������ݤbL �7�g�)Z��Q����`
�B��^v<�E^br��/�ei�M�ika�;�пҗF������)�G݌�kCQ�k�d"��������./�:���Ͽx���B+b��W���a/����¬�]��خ�{D�y@��I�}\��Og<�$$�{iCF�=�G�*�Z���;{��46Ica�NJ|>���Al.NV���a��M�}��T�;/	�:�gmq�~��(F�'�C
�!���;$�`�-
�i������w�%�4Q���ŏ�ng�ο/�Ή�)f5B�8of�1jHJP���1f�9Ϟ�1��0��(Y��7%�%*�-���iG&Rs�g?����5�L��ͻq�˧�6���Wj�Y"f��/��B/����I�J�2�b�����x(DR0XE��}�F9����^��$S�D� ��h��T��Ld���(x���Q58����Iv���iRM�s��֡�uk�F�=���4�����*
�����d�x�mz̒Q�CԮ�)n����VĬX��U�'��^���iE��;�d��af�7�ZŹ�{Z��F��dSvW��e"!�\Ŝ��[M��-{�;� ��Q����{ۻ���=���5�7|�¼�Bs�;����k͇�d$K
8-s�8�J�mR�l���b�q*�W<�O��=?��cx&M�>�ӖE�Q��UCl�'J�2�\x��o�9���.L��p�2����B1���p�]3�'l���A�C}H7o���lݝm_nBب�&SMݯ00��*��:�s�`Λ�}�&�֠�����&�l>6p[7p#G��j���*k�-J�mvYI˽(���qf c��9�l�L5�0�<�^N-����^�&����Y����m���s������9Kчn����ԃ>j�y����?�%�� ���{�uT=g	9a�yK����Q�m�����c���ܺ�����ʘ��C;&��w!���^����f���oB��O�0;�eͯ�'�t��Z�E��������Z�\��������@I"a*��Vz0���3h�u�������L��Z �Jp[��'W�k��[��Uo�A�c�x����35��JӚ?r�%|]����ʹl7w�;�7�����^��6�&��%k�U'|%6��R;��H��8�����a��%G6�7G��a��q��ַ�D�����ހ�����,/�U^|޳r�9��w%�� ���5z2�z§k�\[$���R?.������q��^�tR����x�b�%�tj���v��9[��)��R82+���^rU�o%���x$ �Qa��\�����X=vc�ʬ����V����.���ﴺ�vK*��=�XhO�I�o<��9�����nx���Y}��fnq)<�֬
�N����of����ֈ��x(��y��ԫ;�
����|�e-��&$%��x���>�ͦ*iʳ�Uo��O
ގ��v��Ļ����#Yb�;��TF��6y�������2���l��%�o@SW����%��	�|j�Z"�%)2��4���'�n��>��ʷ��m/�����b:r�կT���?���#���Y.�}y��(�cq���X��]����V/����-�6띺�� ����rګ�Wt��H���fʓHT/|��དƮx�u���K���a{8���kw|��L��Hs����J�����=��V��Bj&!�U�"�����`�G%�4C;F��2X���j{o�7@���7�D���VV%Qg���PP���lA��Na0�a�*��&Eb������1�̔.1mK`⻥�}�JI��%�/l�߿4��tvv��O�K��xe�YF(�4#�۝kk{-1$�9��-�W�3{�+��q�.jɏA&IY�#�j���°���VÉ_zE�l��@	�i�e�wJ��j�Y9#v%�M��QV�W\D3,Tx Wf�6�������㠿���V	�b1�nM~z�������C��F��jt�	N-d��J��£�ڏ�a#��+��h>�v���nR�"���!V����]h5��l�R������_���^W�͓>ޞ��Wuͥ>����9m����k���3
��O�&!D���=��׻!m����Y��n� y���w���Z�$�x^��C�����j�ջ7����Cg�9L�8VN<[e_f �)~�O?�Cu�P�@)$�@v��q�̦u�i�����bT~��E)����+U�.��;�A~ٿ'mS�,���{?���ΦG���F�R}�tT�l�+TIad�qϓ �&���W#G��jf8u�=$	��QO�OQ�������7����`�[V�����不:�|�^t���iW50F3QIvHZB��Θ�j���^�%�Z��edI�v��D���$r�D,�@\�q�U��m=�����$�D�o������osh��F��u����(9���b�Q���b���!I`x8��R�+��7#����>O�8<YH��Vq����`�[qpKT2���R}���Y~��{>����]�ZR^C��ylmV�n��-�jt�53��Ӭ�0�J�#c|&$�������/�X�����'����|֖�n���ߐL'�p.�DW_D�bhh���V�Q����t�I�K�5����"=�%&MIaW�Ĕpi����	�~���� Us���/cG�b�i�4��/h/�	�]�Rд�#�� ��o_ �
��q��m�8?֓A45��>S�,N��)^��At�� J���ɡ��Ag��֯|cA���{/�������t<���|���Ib��j[\�VP}#-@�IBRJO��Ƭj��􇊿�a�x.D����Z ��5	u/A��t���l��[ɦ�\_mO�RJjv�T2Я��x���ͧ+2���xR�����ӆ���kG7Ė��`�@ ܄O�&L?�Ȓ�n϶���j6뵤� �_˶�_��gX?)d%k.u��$��Ծf�_���]�'|��;���J� � J3�7FQ�����<� �:�}���HԷ���@
6��|�bΦj�4].J|�:��=�.�铴y�%�s ^�
���@#(���Y219&�8�Q�/���Ʃ����y,^�/�S:�o�t��k�����2�h&�Z{��)ڣ�&
�u�|GLn��Y�����^��>�&���sS
�;�3puiqL/e|]EvC�`E�'� 8��[v~� �[�P'�5�gK�(��y�����95���pS��	�M � '-�'��|��G�D�p6�:M�����0V�b^]�*�/0F�l�����X���~%p�I���-oG|)��V��N��J^l�8 ��G�K��C��	 ��������1��QMa��t2�5 k⫞�{�t"�7�!�a��"�d�.;SR�����	�4׮��!V��A{����4�ً��y&������'��z��U��,�o��:�PHxl�z]��Dl�9�[��fr���������=�G�b3&2�&�)Q$$2�G�=ҷ4 �r��G&�������b�c|l�4�w�z������vi���N읆3`x<"+�1���3]mm6k�'|U$-���yg��C��"F�~�������<��_�B󴾱O�ATP�y���V��{�׵T^Q�WּǍ�LQ��ˑh1�`_Y�hn���O�_>k�ɶ��{��<��+d��g�̥�~�z���R�/ֳ�z���:��G���6�(d���J��*����R�8���L�|N9c��(���*�i��w�*���}�&n�i���k�4Ã�eg��O����l�����:���'�}r���N$��@��{\�/_���	�,�Z��c<Cm��ƥ��0H��m2�w�;B"�(u����w�P���f+7���I�nƙյMO��<f�Պ9���̂��n6�Ȭ9t��j��J�9H]J�8�� ��nBC]v.�!]9f��~����>Lҟ�$`��{�\eS-D�G��˶���xTc�8"�]�!�	�`�ޙ�4T���um�Qa�p2�����I;�L�űW�8�X]�v���\׌��z�;�|V�h�<m����J�i�ç2ό��X��%f�/��l7�������%"[�w�<���������T���-j�8d�.n��ӉeGΣ��ˋ7��������Y�{���"��:�����H��.���~��E��hgХ�@y|ܓ1j㊹��� ���Uwce�>�7cW��ϗҕ�jF`��n���>�䂪�M�ɬ?��̭Z<e6O'ビT������]���Y?1w�\v���j:�cg ����Z{I㼱+U�K�y�|9nS6뭉��b�0�_$��ay)Q� ����N7���ͳ��܎��%��|Mi&���fZ���=�ɽ����(��ö����e������	�ts�p��$�}3@Fw��>v�T�R�hY��>�1^�@Vrc��6V�3y���qԋ6����i}<�}֘�W5i���!���b����:5=�y;3zw�,s��L�K�hS���.9�{���\��U�'M�R�����A���G�OP�vR�����W���|��?{�A�f�We����W���\^�~߃�m��06��_ ������iV>��j���;3jW�3��ޒ%��zk���'9d�Q��XR����C��&W��B/���B��|8B�����KG_j�'l����ͻN\p�m8����V�����5����[�����Q�̢&���陮�p�}s+|��Yi��^���I��T�

JfO�*4�v���<�� �Ŷo������л������{QYU����`1k /sc��p�VX]�{�We�F�_�('�O��s��vF#�ȹ.����
\�T�i��垟�Hz��3����#�nۍQ�D��	���}�I"��vv/��o�g�K��6���i��$�Òf��f��:O�� �,��R��uށ���y<^��v�@��"~ƿ��%���C��t����L�*#��}�� ��[0�z����3},)L��_��F��5@m�-lW��1"�E;�_�H���uPK� �K��8]��U��� a�Yi%[�:��z���^%�$ڎ;x�S����w�y��uJL��l�O��)ƞ�L,Oj���c7�Ze)~q`H�޹�)>����e�G��7뾜�a��\�S}]�4*)�x��0�^�����4u0�D-l��W煼(�y�5����a�����*@"x�&��P�+���<gg�H�٬�O�WY�ͷɕ�������V�����d2>�β
�p�9IR�^����� I�i�'Dw5�P�P%4У�[)�2�}�:��'�%~�׀fOm���]*��'��Ӆ��S�Y5s���#�X.��R������=v%�͟�2�e�vQ'��{�
�Yq��-�_�C��qNGW�\��f(�3b�/��������s��B;���?�P6;��V��V�c�׫<�+Y/��δ	)�!8->IR�c� �e���D�T�� Խ]oX��/��a�t��:�J�j�p�6������nN ����e&(�g'? [�8g��w��B��R�r�4�)4��W�m
�1~���f����U���?M�ɔ}���N�RU���}����4�H�)���������:+ŏ�����ծ��Q<�Mv����8,��B���r�)B{}���������9Z����^eU�����Y�M�g��������ᗱכ2��b���oX��Q�S�X�A���}�������aT��ď�p��
�
��N�/�x��6��48'$ܫ�Q<4��B�0t�tg9�-`�ځK� ;�W?;�2^��"��GdF�f��B�I��J���T�*+}���1�Q>���H�t�,%�� Hww-!Jw,%�� ݝ��)��twו��Ͻ��9�<s�}ϙڳꔶ�[>���V�<j]tJ4�>����4��w=�%0z��;�B�Sd�5h�|e�sd�������U���gh���pVkCn{��2~�|<��,�Te-��$9�b��gXa�"CVW�����*���:f�$n�S�FI��+�3O1M�ڂi��4|�ƅ'�ur>(k B4��9�qP�;_�48)��Sxt�[�9-�T
/�����W%�M1�������[@�Rױ�C���L��S4�[�w��Ѧ�& �}��!0ԴbYM�k�9���}��^�,��7�_%�]��"�"�q�^�����9�S+)u��d�����o�޺�h�vm�G� �㫿E�~����	�K��o\��B��'����L1�� ��o��{o�(ހ�;Hm�!~�&bd�٧��`�׻���t��v�i��W6��H��(1����yn�xd�mK�=~���uk�X1.�S���I���E^�Q��㐖^6xW�8T�v�qq��\��u�C�����n@{Ϋ/pw���X�vg�'q W҆g��0T���3������ٞ2�MR����#��)�N�O=�C,z��Gl6���g":�;�x1�������]ܼ���pk'�]�|�.��\�w��
���FFF;�G'�Oڢ����=#�XI�ׅ�j5���j�mx�j�fDT%Z9Q~�(���Y�����g�`0��p�Atm%���x�y�u���I��ʟ�򶵿���d/���'3���V�����y$�?8ͅ4��[�A���V��9ZE��6S-��1���`t[*�9x�\zqp��{��d}��bʣ?�Q�R^�B*B뺕�1t�B�`�ޗfI}���o�X]֠m�v�����	�8�\��M!���^�\��u�",�J~�E3�Uiԋ�+mkQ~�^�<��_���� �/�۟�J�35�|��e�\�9�:�����hne�=��(|BBd�%��`\��H�s�ؤ'�̧.��M��k@�V��f�A9ǴC�]xY���'RL�i�mM3 ���tt�˯��F��L|4%c�=�����Y�ͪ���~/Bi���&?�]�Z�]!g��El��6	-�Nf~�w{��������,�@">mO�^����.md�B��N� � �r�X�QS#`(����.�|��	$��=t,�e�p�#��j� E�}g���Blx��y�3����׽�h�������(��sd}(��L@u���T"����O��_��̌�}��#��5���Gmb��"ћ�մ�Ӵ%`4�d�d����G1���JQ=��d�=֠����x�,`��_H����>tߡ�c*�|+vF<�)pR	{y
~u$*2�q�Pp��!_����#ݪ2)�H���ڏ��)�D�)�	q�|h�uBK�Ss/�z�pRH.�C�F����B%uM�F��U�x�]��K���`9dJj�Bk,W�¦�����oz�/�8c�-/�暋g��5!�a���pb��q�?�yW˱���(�M�!�>c�����Y�S�udܨ��1���;�~W���Vٲ�
�벥��e�B��%F CLE"S�ZT!t��D� �r ��zHg�9h�B�z�`�,�<2��Ģ�����8��b��0�~2�L�B�����Ot�me�e�+-%v��r�jkP�iA�eNa��������HO�ɖ��]W?i��/��������d�~�l/�j��y%|̜yR������+�gyM(�'xP��w���>oZ\^�.��,��If1�KE6n�q.�iS����̫D���/����x����<}e�߻Rp��8����$I	�����O��	�����3Xӗ��k0��6t�6�+U?_M�����%CmOO���*�|�7t���|�5Bh�e�ɩP�H� -��eJR}}��L��;@.l��1(����yS��e\��<�c7���A`j��E���!lPF�ԩr��;<������,�dI�r�4�٣�N�=)�7�[x�.p�o���x3��'�^���{zэʭ���PU��\����2�s�� �35�;c
����FF×��̼B�]vs/�O���o�81��a�x�w,8��D�w����gc0�����'~/�
�!�]��r��P��j,'<���X>��=vs������+���(^˝ �^��|KY`"j�I轰�C��w�Q�=�^�@��U/�lSR7�+�t{+���5]S���&p��Y[����I"�s���/�?ye�<��[��ӽ�$��FM�6�	�\��)���`7(R���D-���8Xrm��X�A�2�&�u�ז��&�Ğ���\���%�������g���"ed��v�P����^.}��Ʀ�.�
���_��gƟ�Ov7���ޮn=�a+\��%� mm�9A�0��0�U��c㒂�6v�h('�����)/���E)N�_ڱ�"���.�� ��"l�9�wb������ JQw�����2���o�R��,/y�T-+�Nd�'��R��;�Hwi�����>�2Ƥ��7�dA?R�9Y�(ħ� �n���-~��}
���nz�|b�!��B�~�4	�r8g.��Z �*��!�����/�I�N��#��.���hۀ�s��x�C� �mԇ�y{�	7�M'c�˂���7%�%E�a�N�	c�zΞhx}:�B����\�SY(��k2��{|߀7(L�7�d�,�r���W������y$��˂��`���o\|x��]f#���d�zٓ|O.Ѡ�p�_�˨~A)��]t){���c>�d� M'��X坂���#�C��V�oL��b8���8�"��g�I���b�!�'�;=۶]�	S����w�&h��Β+���U�X�����Qǔ�g:s_H�|��<���i�1����p�g��#��<��Af�$"��5/%�=k.� 3�2z?Jj�X���M	-�R&�r��LԺ)]
E>_��_A?DiOtM��nSR��u�q��@���Ss�4�&���x/�y���|I4���W��1S�GB@�W�`%�����M�H!��wY�|fQE[���ͅ!7�'�w��򋣋�[|�xNy8U�3�K���;m�����A�A��\^�T��N�e�>T-'m=h���MG�$U�@���Oƒ&���._��P$5}WC"�t���#�������J`��FlX��Ө�`���}	��(��� 8��;�.���1^�o��ʡ���ts��u[^���׉Gx�*b�ЎƩj&gq�\d����DBaz��#w��u�/��׭01Gտޮ�4�m��}���AG�g-)Bǲ6�HY�nh�He��r��+�~���Q�9��DQ�z0�O�s���2%����cY��P��_iZ9��5��䉮��[Z��3xQ� �dٍ��}D��5!�M6�P-'�/~&����N;�2��� v&>wk�-�~��b\|'M�������&MVYQN��(�)r�3�>:B�5�,O�M��o�pX�xOZ C�4�x(�Y�$�o�7Vh�[�G,tw�c���t��5[�s�B��7�h ���<I?4/uٕ�-���Ŧ�ك8�%�M,J��זJ/��B�T>��@��R��:-yI�E�<�x\#�!5ܚ$|/ �)�����6S��>w� ~w��}�SǠ<��R`�^�Z!�=�y_��:�z���ǔO:P�Y�F{�-ֆr��7Y�a��<�]bQ�KĖ�_�� 3k��\��
r[+}�����Q����{Ze	���#��)�e�?�2�/Q���k���F�%2�L����GU�m�e���`�q��R�e,��.^��&���4���t�������}������ (?f�V�g|o��d�{�2�Lvr�mp%�^���O{E_.>�)@a��ј���w���0�߂���Ͳu!� yf%���%�8&�G�?���~{2ͽ@�"��D��UC�0e9T�$��nf�V�u�~ �$&a� Ι����;}���')i�?��~B�ʹYT� ���L��v�\4��'0�!7��8љy�f{�aN���>����5{Nk�Q���1�P��Z%��FM|��;�F��p)մ^=����=5]Lkg�NY��r���P���<�]��P�q]����h�%Dh�:#�5�P���"0���A�/t�DMp٬|$E��\$��k-�jx���2dh�ΰr
�ȶM�*�iwR`���#TךX�����u�욙M@���j��vұ�W�&XNT�Kݵ����. � �0i��R^�2���d�?Ѫ3Y��-b.�B��F7tI��v/fMC�ݹ��������Y�A9���u�v�-�?�W�J�P�����l1:�$�75
e�o�~a��O�V�ϓd����Ͻ;+�&�;Ikԩ�:�%$k5R�L�I��b��;0+�bحd��~|�4��`��� �zԲ�g]"D�!�`��yp��4i�E��y�$'�Ir�;p:���=��$h���M�D�5D�گ�(JL*�I��SԚό&T�pP�v��WbNvPP�B͇|u::rƁ+����X0c^�d��W"�'��F�	���?�d6�P��"�u4���d���E�,@���j���%�&N�tp��oP��}���u��:�5��!2��"�+m>��2\����~�X�	l&w�{��m�1@�u����Bg�+�cLҸKT�x�;	���sDo�����r&�lP��Q����3�>�sR���3"�J��)���;f�=�B;LXD���^����)p!���g�Rj_��֝L
�e���g�,�%VzS7,A���z5�k�`|�����/Q\����I���%��HX�Q�BV����;v����{��]�)��?���0��*��~��x�7Іm�u����{3��G82J��C�_,�ֱ-�AZ'=�KR�U#�B_g��gJ0����E�ꚇ��aU(�^���o�]*I�@E��9�&p��1Θ�ꉫ��1�I�o����ќ	" ��0���ߙ$�-}' ��:��>dF�����<p�� \�N�U4���N����;��u���V2p�Q�u� }�n=�5��)-��ƺ���sN��� l�����E�T0w��^s�Q���l����%9Z�ݎ����%u؅�1�'\&q��8���|���Wf;�F�$���fG֬�i��߬����������:@Q��{�&}��~�w���b��X�8j������'��4M��,s^�FB�tg.וZ��r�;'e���H��,}��4�w�x��L��*�a�Ŗ��ܛo�M�]�JxC���
�k�����+�H>�@�b~t��#h%�yL��A�ʒ��	��_����Y�<�j��N��_� ���^!Q:�6���z��E�h�af�]��B*1!�{�n�xZo3�m_X����O��d��=^;���+e0��K[c-<���E���F�=P�Z<o߭�~C��1j�`<�
����b�&�nb��w�Ø����J��Z]�C7j�����Njhd�����7N7����$y���.;��ۮ��Vō��A��.�Q�=��G��	��[5���~���e)�-�\�g:=�k0�{c�v|o��wj�r��(J���
L߸�N���GK� �����R5($Ug�� �(��f�c����3��X�L5��mm�6]k~�6q؋`��rT���?�٣Ǘ��k���NCONni�D��/�rK���lKa�*M�l
2О�bi.�k�d�b�{{�#�Ծ�B��
��4��P�O(!�$�z���_B�5g���ϲ���N�%���F�üA_Yu�ct�tD�s�_=�:9�2:�`��￡�4�{hFL���$s	C|{�^Lgm�����N�G�]�U-�~:�5��u||���)��_�\"�w��faW���C����7�4�:'�_pf��%�AK�B��	��;y��cc��e����GU�%���Z��[�W�l}�Ė%��#�.���y/6ӈ��
��4��t�v��X�_���nc6Eӽp#���Ip��֞\��lƷ����Mw�H�
�@�F�w���M�s �T���O�5q�GS����Mf�MB���|GГ]�;,��W������$]���Lz$�@��JG�H����
�o��?
F8~!�s9E��D���#�R�%�a6�\	�$�.��U^�S�����(���% ܈�4*�<�pj�=/؃HD��_�r?>��Y2�1��7���o8���X�;�/f	z������ëx�gr�����!��ݯ�N΃8���5]�?s�ł��=����F���B�9h�g��I��Į,�"�ʐ���*6ª(��r߿��!�6�y��D� j��G���C�Q�q�56ݦ2��;����~����m!�?받��t'R]���Eq�G_�[�6�b�'3;��wv��ʎg�h�Yc�N��q��&3ݮ�V��{B���-D�W W<���Ig3�y�����H|Ww��wW� c�T��5Q��M`4��b���G�e�������$�1�z�PN_�*�s|CEVsL3wP��ϳq�3���u�`����
q�z̭��qx�Çm�@$ �i�t=�-�����r��BW��wQ��"B��	�xZ���|v]tL�~��=�rҳ��u����ݬ26@�Z���A��w'�cB��f&k8Ͽ_n��J�0�Zh9�9#�c:2��_��gOlN��~X�!o;ᇸ�OCv͓���3p�Gi���R�/f���`��,�d2�=��k�[���/v����x�)P�Mx��AB�b��p�9��j�����ş��Q�*�q5�(��]�_'��gF���c��<�v�>l�w߀.Q� ��B�Aw�/�״���?��~N:�w�|�;��à_*}�z���}��T$J���J�L*�\}�z-~��o�:��	�!�Q��.��$�~�	���K��*�ՇG{K�B&�j	@R�5��o��~�-��q|�q��C����k���}PL]̆<�d��̂@)!��Z�Q5F�/qQ!D�5�+C =�X�n�����o��;����Q��9�I��� iī�
!J�̢ts�M ɕ<�J�giR�㎒��S��(��f���h����>�.$��|�:��\Lr�MA��;Ŵd<�]�R�]v:��xjC�`
&���5k�4��.�y
�r��-nYզ��+$f��$"^8^��#�i^�b\ w D�Ùsrn�#uU�n�Exc���P���D��xpyy9 K�Ӭts��ApS{�+�NW,,gj3���*���m`�BXl#��CTZ��ް\z`�Y����`�4�#�A1����+|ñ��Y�����-�?�H״34���|��������8x&8�	���_�aXz�kg��҂b����P6N\fC`y��m��7�c�We?P����C��CU:�MêW��f��g4\Јfy�[d��̍G�E^��&�_e^n��x�`���2g�o4�̫�)������1jS�sQ��p��K��.��a��F��>�̤��o0��r*��C:�=M��p�	��b��O��V��W{��\������N�mJ�-#�.[�zF�8��Kl!���?����Z�f>�]���v�3gv��{#�Uh�+����c�?�ň�1*o:M��.H����Y��uF(�V��-%��W�K�%˛����{�y�<���6mU-��8
�5|��R�����c6y�N ���LƎ�Fn�p������]��L2��,��6��	�upcEjk�����G��n�`�i]�(�^��~w���W��E�;k9+�h�+IT�b��G�zLȗx���� �&�.=���
�+�c�5�;�pEJ���T+N�����r�����E)orL:��ر����.c���H�7�/��5��\�%c�)���&�d���L޿�B@��A���#�^��u���r*<0H�iW�l�������6#2��(S>�j[���0�Fyn�ە���S�],>���ZN�,A*��0y���Lk`��+r���*���h�&���Y��b��j64��_��.�C�@L���$�r6ueD����-J<��m�a��-[�EJc��b�bo�+R9g;~�ͤp�k�q4�R�[��um�>�ǡ���AX��������y��N�V[�i��$���1�+�����u�S$J<���~!$�J�̋�E��<A��K�4`(�p��8��;������v�[�#Sӂ���Y�"Y���݊�q�~K{��_��]]��G�b�5K�lvS��{{����'����N�i�r;.PZ�<�n��M�#����-�v�W�a� ���Q��3Y@6��D���`�r�ۻQ�E�m�h��U2��9w�c��n��f�l�'�d��y,#m�B��t��NN���
�F���vf���b4dx�k~�?+�*ޣ[�#�XW�@�Ĉ�qDG�y��o��ģ�_���7���!e�8I>���]$,��kU�<K�遶��-��Q�2JA% 6�\��ZE/��e��������"�AG�<�+j��O���M�.���rב���$�����Fڝ�*'�d|��+���p���)O���z���ڒUɅ1v����'U�ve$=��<e���,��
b�;%e�Q ��$f;:Y����x�6�Ut�nn��q��P�1X����[^O��)��PIVi��G5*̽7��s��q)�h���HTI��]_7�q!��_�i�v�<I���d�0�{�b9Fi&�<�=���C'�nU�ޔ
�#�S�j�?;o����@FT'�#泞���1%��߸8��s�6�<�֨X��s��a�&�Ʀ?ߴ!�x��J���Xe����=�Z�����x������ k��Z��Ԑ�s�z��&�a	R(���:�~� �WY5�)�Eʇ�����rm�ȓ��L_u�Ǟ�G?3�,��$���~�n�Mt1ϫO��:5��*
�5�o��2|��y�P@B�����q�|8����tK�櫫m(-I�m��
����\fJ�1|�3O��7)��坅���1�@F���8*XͯןĩL3�œ��uǷ�a��G|9�*9�ENaկ�3��ڨ����-?�sI�NV[�c��t_.�_$��.?0�i��H�]�+�qE�5�c�a��e�a!Ä�EX��5I�����mZ�f#6ժ��q�/NET�xs��Xw����?l�8+����yK����D�h]�MM-�/N��QM��&��SI��-�v�낼�����ë��[n���>wԎ���/.�3~vD�5a��&�/i8RnCЈ�Gu�����xHj�6��=c�o:x��qw}}��4q��k@fڕv��k�(�\��E�?{L�nh�eo0�3�R>���jY��hDL����J;�zK_��H�(KY3�L��zcS�PU{ �Àvy��t�i�����<������`V���� L�/�J�9Yn\^(_N% Q���E�1�הKM��dM�H�5�Y��ɋ7p��x�b�b�4��0\��67�І׈D��U��^\���.^������ݱ��������o������oh��@{�.��9���/aA
�ƶ�I��:%�Il�ge���4A�|)���G�_>:zA1�A��N/%����Kz�N$P&�|�SQJ�ix�X�K2��_'�Y��j�!]�����L�c�T�)�(tߞ20ՋBk��P��ܩI��l����HڔLʃ���ZZ���b������[��4ԘU�� O�t�Py���s��K�'y���X���T�x"x�Δ��ّ	��&��B���Ć_[���FY�`��a�#������ڕiJ	�/�v���aO[#�v�qM�����ѵ1�UKH��d��А���tө9\���{�d��T��N�O�Xq���{#�įp��r�������/�>q�w�Q�\��j6v�ܨ��]UF�H�=�'��T��!�Soe�E��H�pW .�z\���,�2�xKh��-��~�nK>'���c3B-�τ�ީ�@�M����ݡ���Z{l%�� ���<?���SO*��銰]E�%�򋲠��Ѓ�:��O��E�vđ�Y�E��,I��>f�|�#���=���`1����$@�)`�F��E����߅>k����b���)���z�%�ĥ[�ZX�CF3���ȗ$�g"/ܗn�Q�R,�����E�\�Q��i������b���vKn5�(��2������ĴP��ծЫn�C�2Yڋ]�b�^��,�L�#	(̞+���8V�b6�ᯉ����!��'��	�͂�zb۟8-jJa0�\��50�H�N]�]D����������4_���N�e}���~`�6Cv��^,ƙ��ͤqa�f�$�eʺ)���W���.ؗ�7�W�o�����j���SO3��6���-LDr���Y{(�2�`ήi��TK,7꾴�s���2�9o�p�V�~V;lF�A�A0�yR,�"7tn�y��⊅6`�Cx�76-�R�Ȏ��}ĭ�j \�l���]�3]���Ķٯ�����q7�.�m�O����W��!\mޢ���v��Ժ&l�lM��?��7�m��?)C�;>��6�,"�&�1{�m�/�{���ԙ������h���/�#h�a��7Z�s��~U�aK�7꼢����H�C������y ��Ṹ��M���m�$ +�-��j��j����q�X2�z���_*������}a=��
_b4��ۨE�6��>���G�����G�se���9U~�FҴ���m_�5��H^�3��J����$�0�q�~Ghm}'V�cH�~gk٬@�g��x���X�����I��r�%ӷ-��'H��O]ґ��g�y��g���~5�e��Z�L�ms�b�H��:tԃktA����7v�+��G�[�n��m�x[[ÿmS����!��|��/�*^G�Wy�=�f�T[�4u����1e�d���:Ovw?��j�� ����;u����Mœ��\ʋx�����h�kݺne��G|���3w�;Bғb�4��7)�[���ݡ;�ڹ֋���wp��]HƁ�t�M��54�-^�/���_��:l�8�b�G���O?S����.4�c��h}�w#�.�|��ᐶў��_��v|���ޗx�G�DK�_�rgd����T�	��A��2���#g^��H���+�Qw�d� ?�Y��S��uЗXAG�-�����R���$�/�M�w�� gm�+=���q�^.d���f��waC޸�U=�:��3��Y�|Ķ�_�qb�G I#@�vsN=�#k�b��lB���ur���&���1� ^ʣ���k8��4��~�<p�u��߱��k��O�R�HB��>�}��ZP��^ߙ�J������,N#��?����.�g��yx�&�$�с���.?�(+}G_jDq7�~��'���$�z��ğa\�l�:������n�o�I?�S�d~�)�+؄ܽ�8U����C%��F����8jsM��7�✌hݯ�|�в{����i�o�ה�ɨMw8�+��Gy��~P�Ju�����̂�nȷ�v��)�^�ڢ4pT�{�GH_��ߢw�/w�5�)"԰�Oym�)���yX�u���̵�es��H���/@��h̅�˻�̻LƟ��uu�aV����M�L��'7v�[z�ͺ����!Q�9��Z<<�(�M�T�^�~��8dR�q���!˃5֨�;Ճ�i�&���}4�`�_��N�ђ2�*%F/�'%���K�i�~_�=�ͩ�]��-K4�Xْc�v�wB$�7&H��?�N}�?�Ues�(�w&~0�� �� ��O��tj�)��ac��&,��;�b;�YE��8���uC���G;Ҟ2���
���'�dF��Ծ����O?���B�A����0����ŽÜ��$ĩ��g[�xL��[wl����s�ӽӳ_c[�)��oo��3���HU^�k46=WY뮧'V�Iy�c�[�����yq�OZ|��m3�3�ZM�9��@*|C����=�V���p����/��~���#�=mŜ��+��Ͻ�s���QI���kRh�i�&��#���^~�f&���Ab�o��V2�GUh�H��'U����?��������[b����z�J��$D�����1�{��������(2�v����oD������AO�χ�������V��	V�y_��[Ƅn��#��^�	��s���u]��n�ڸ/x�/�q���?�(���4�f�uѲ�a�����03�����U珖:�!�;[�۲-���������?U!*IYSꮆ��S�c��/��C"�q�m�_L�2��JT�=�p6�c}����O��Z=k�4)-[0B0����>	�fa�8�3���l`v��jOZ/����l7PX<z<���_��?y7>����>ε]�)�ïI؈6x��p����N�w�>����q���ġ�GƭY�����E�V��O2��4�T��'�'��9���z����t2����m\�y�{�r�0�u���4m|�yo�X֤����9�����?+/���?�iON�ՖS�ȯ�`�w�÷*K#*���4g۝�o%�*���ڂ�:�~=O2�܏������T��8��Ժ��WQ��򀈨7�]^]!M������M�ؕ 8�yh/ J��/I���i]�zlb�-`�+�O���`����[��\�?T��bү�0u�sۆ��$כ��f|�RJ����6��^��r��937���h�^���rY3@�^x����w������xX=l��tó�n�2��p�O{&i!�X�O���쉆)���cB�i���,��&�(X'��F]�ᚨ���Y��B5}1b��7$��n�{g�.�DKհR��?xc9U��
x7�ڧ���*ȩf�����X�D՟ti�g���>/��1Ոt���y@v�0-t
{�i�(��Ћm��CSy��F��| ���ρe�Y�#֙��v�aO�R����%��zP��Hj����P������/@����П:���)�����+Zo�*�M�(-^�L�e(��7�S��-�_oұ,��55S��3��0��ܼ���M8j����N��*�5�Q����H���ǿ=l��%��v��g���"��ǣ o���Z}���GAf��'�\K�`����8�W�q=�욕E,�3�_�T=���NfZ$3j���i��z0���T�Y�pb�%8�%����2Ꮁ�it�f��<�&$t�m��U�Q@�3!�E,of>i=7��h֊ih�S�RxМ��Y�����Z��n��BD����Hi]Iǒ������c�1��QA��!�П�� M���7������R��2�/��_�l�$s6M&�O�1u,�|����|�暥��Q�D���남Qa�޹�0��11w0G�+R�Y�f���6���ᗞ���[r7�J%IN�7��gaǣ0�!��
��K�O���:gbk����P-b��H�x���c�,��q����mBA]�^D�׎�t��w��"�v���d�ϳ��Rz�F����s�o��״	��?�����مJn��5���<�/��.L� )�Ҳ^%�P+f
�^���G{]
�2\�d��<��^x�:>t���M��кD1iMB���:��UC�Sr��oS�:*���U�If�p(0CLy;ܪn��|J#�vԘ[Zv���E[���PT���/�G8x��!5�E7�q�(���\�:�Mgp������ᷟ�s4��;�
�����^��;6t8�؏���w�j_8��`���๐!�>���q�V��x��Q>��u�0��L/.ӊ�%��&����o��Ga��Ay_F�����!��Jn�5܈e�=���/J�cy"���,,����R��q>�B��e���bg�v�An��x���W�mS�DZ�}�0�^I?9
y��hX�O�Niz[7�57$��1�z/���`N�b�[������K�J���6ZN�]\1��!��@��?n���[6.�����"cn�ς�KE�v6V�G��E
l1�7t<�*��=Ng>�W- ���}0�(�oe��I\F�,3�дN�G�"���+*�ɥ>� Be~$��sf,۹@�����;����GS+{���+l��$�<�Q�I���ա���9��/;�i���q]!;���U-��%lZoJ�`M��E��灴^�����6Ϯ#�������v�$Q�4��ZS��j���H����)�Ȱ�s
��i������@�؊i|[�Ѷ�I���������H=薺����w����g�����Uێ�!W����w4R(�x���01��1�S���7P�q���Z�	�i�H�m�-x�o��"Q�
��Z�6���C�/�k��շ^��O�ຘa(�Bri��.}����BD 'w�M�m�_V�;��w�0���������W�I�-b�1#v��<Rz\ִ��J��eUβ����9n�����v2Y�7�-�1�keҾUC���wK��^��~Q�Тe��'?
��˃?//�u��Vha̒�!�q[��Jz��6�]��Pr$_X�����48l|�(����
�E$�>��0��k
��1��ֵA�\���g��Q�S�5pS�����͎�������NA�C7�SG�]v���TH֒�`�|�%�,���4�\���O�A,��4�}�M�q_W�o�w�k��#�
w�����Ts�tXͮa�߆�X)�n��r�xXٞ<����jg�<��{�Qۯ�U셾��������<D��B�B�jYU��`�k��w?��;�U�{�b��vǤhג�
��0����_H�3�SA�[@��JH�)����e�>U�:��)f\���/�"�mF�46`8�T>���^Wt��\�H��N6CV<Xf�j��x��a����5D!��|���*�)Ks��	yC]C�Zr|�P#��n:�x�6��q���*�UEZYϽ��-������j͊BD�-<�2�!�p�ꦞ�m'��1Z�q�L��W�㯉Cow���-�^��au��M��xeR]�;�{��N�r7�u��#����_�>�V�p�^�X>`D��,\�\4g+5�cmg��*K�$�}@*��W��R��q	}}M��u`gi��&&#��~s�r�+{��G���(�T�������y�u'��?�a-M�Q����TT�.��.e;�cx���Y���ՅEX�`�H�}���� /�U�\SP��3�sV�n-���X�ɢ�UU����P�����|��:������}����죷r��_s��7~8a�>��K�+~��	�X����z3�zRQ�QSeu�V�X�k�#V�U)������j�|�����o	�S4N�~�Ί�#aO��(I������9�;yZ��6���$�t��d΋�_�N-fA�T���=���X-Z�&�[�2�H�ot�Sa� 8Փ9 �>�����_��_ ~Y�Ƹ>�Jդ�JO�Y&��>�����QOM������f��;�L>�h�w�iS-��&N�Ḭ�JK�U��x�Μl:�y�D�:Y��e[G!f�	���ǈ�):""b����d g��עy�b����s�MxS����}󈗉�	-�<b�]�SO��c��3j�-�P�z�;��������c-�Sp�&�j�c�������
H�5X���>A�.zfq4!qA����7<AEY
������<f([���J{I�o�;�����r�9Z0*U��a}�� O"�"j\���ĉ��4n͛M�'��F^� �����}�$ø��K����:��"�~�U��}��������|�0*�wW\�.��/�']��c�׷@t�M�~���[�,��a��T�TB�,K��q�Q5�)�ox6����mJ�v��2#&�_�����1��PuJ\���*�"�SE�&���塡[�����,��9�s�
ʙ_�mz�����M�h��Z���֗l��M��@���k�s�&��xT�u��@Wo�9�9�#����6+f��K�G/cZ��ew��լf�e���.Bl+���f��d;�C�g��
����_��$"|r�Z�h&͙�n��0�t?�i�8r�]��
ࢿ�,�x͉�'�ZkuA�ΐ�6����W^�`�0���)��G���f��W���p�gi_HWg,t�"�?���8��\90h��Z�����2j�k��/�r7N�"D���a	��̡�3�S����3�_8;�$$����%2��2�yݫOvh���#ص�U�)�Ò�L�cRd��ʼ!�ūy������Q�*�KI�1Es%}@b�X�C>0'؎���a�-��
��a$�=��	����,@pܝ�%x����`�%@`������>����TM�:gw��^{��G�����,Rk�0C��狍!��aXi���V/k���EA� ������g�1j�L�fB����&s4?l��ٱ.G�D����l#XE�[��Wy��y4�Ž� �&Žc���ٰ��TW@�*K2$�s�������!N�=�����ӪhnԵ)�O�~�w�����T�Wr|��ښ���3a�ǾV���yPE�Â����ݱ�:�,�d�� �I�m,�W�xК�֢�"�6	�Jr�K"����"�Ȣcla�m5�%��`^�,�>��ۧ�@�w:A���MY���<��2�PXAJ���.�_�э}�_ӌz�G���Cr'� ��64�ɓ��9�7��������2D��D��y;��Z�_��኿��i@Oh�5,���"����mh��WJ�(�x�|;�������#����@f{k���_	�]�wd>ԇ���,�Cd������C�k������ ��~7K�?Af ���������T61P#������b5���	���P�5#��g,S�OQ�]���%"Up�/� RB"��װ�{�Km�
����W���4E���+
d�-��~r_�;��!P���%��,�`i��@��_��������&�A��+��e6HiO����w,^2c�Rs[F�F�f�tF��u�E��P���R�*��EqY��V�ց�'�O�Y��6&?�bO���z;�CV2����`����&�4P�0XR�"}�	�`�3�Ǿ2?��7���������TA��if��'�O�(a�����K���������EnY݅;��~�C���F��#�2j��F�R*���N�~�@v]��/ٯdL����h�׽������ֹl���9�!�-6H����߄O3�t�?:�y��pLg��")]�V�mL�@"����{(�h"�7i�2�����I^=0e*�w��W��j�Ɨ�v�/6i�t����N��d�	��`�?5=���D�<���)_�xS��k�sy��m��ϐ�($"I=�L����m��aW8`(�q�o�l�N	��${�,Y[D�������qW�L���0oRJCUx�	�E��N/6��:�E�{�Fq�0��ۍ^�^����˟ȇ�7�Ƿ3^�|Ħ�/��8�ɍ1�z��#�g�k ��`'�܉��؆-�	8|�RE��],�nr�QLW�;t�?�͕
�䛼���`!�|��J�bH��0��%�~܊ �L
��1-�TTЀmH ��*�q� �d�}l}�}��v3�?���������\g�]�����$��c��S��> 	?���V����Rt�骴^��X����'(��pg��Ȟoi[4���d��$���b�A�<��JN�/m2��m��n�]<I��/��}P1"����\���P�RVl�͸~�iP8Y���Q���R���U���Dw���{�%!u�`�a�P���!&`9�( ��0+˂���]�n�{#�Kk��X(%�q:��1�HVY�8ex�qe�G[ʩ���8
�]�j�:𐑋��T*��B��h��#�1�,4�l� �ӿ~�߼�ȳf=k�)�h�q��OR����;�`+q�H+|""N3�����̾1{ikU������5���oj�����\|_�a�T�\����6��պ-!mA�q,�Bf#׊�:3~���� [TT>U/D?��Ǒ�G��q�R�*��o%wǨ��J�%�yP#ʂ�ݵ�w96Ocd�J�� ��тU�׷ˣXT(k�ZH�
>	e���hEvZƏs��2qjw����ɠ�1h���V;�F��g����e����K��,�+����<I�,���C�Yf�+������^ӕ� �����rY��f%�ZCJ�@])�vҀ��	GǚQW'%ƥ!�*�a�.v��է��ۏ�nJ������h��_��Hw�~�0���;PE�7�T�0e�VB�z�1L�=��Ԡ������J�*5��z:WK86>�+��`vp��> ����+L!�V��5#�.�=��la�/<�2WǳFnx�p،��*��;��G��t��gS�T9�X��]�!�E:K�u��Z�_.ɹ��=z]ft�����%�0�R�}U1q�"r�����Y�`�Yf�jmr�=݄���%UGp2�'u����{>��e�Z��&1�,�Lt�&�� &-��x�_��h�3��KW=���)�)'����s�+��>�<bL�3�ڭ�s����6d���-������Iu'Msr�+�]:Ն6�N�vk�s�w�f>����p^g���c��l��e7ѧ?��aG�yJ�<.%Úx�VDVϻ�n�g9��(e�냈=�9��e�l�$C�okĬ�d��ogtE"!d�����nI�N��������i�PJ��L�tu����l��]���>dպ��zHL#�,�a�W�.�L�͇�kD@�_R���!�(`��U���O�K�"!;�u���0�f�#�>�G:����$�3�A �q�����xC,�s����O硸�;�ś4ÆcU���`@:�c�B���	��|�=ͱ�!w�*�A��?��.��{Ǣ��8�;��u"��w9N�IV\��~�[3�����a�?��}5b���`� �`6�lm���w��z�H�Y�O�t,�U!Xy���y�]�Knaqt�d�-����|�"z���A��&cwՅv``���`:�>s�&�6�h��>�Js�1�����#��0syꉂ��9w~%����a��M�")+�
�Gr�o''@�Hp�&��T��A�溡��N�#K�if���MBK���T6�����^�Xl!�6ق6�+4'Q_��6}j�ܡ�Dԙ�/a����ԫ�{�M���)�ĥeo��ܤ���;���B�\��O���<˦�.�G+�rjBԬ�g�����|��U�*ԭ� ��a�ح��f��Є�0�3��C�&�eK��Gh.��]`%�̕�)>�]�ܤoDC0TT��;�I�22�>�L3ph��G�v]4��'�c;ڪ��4{��Xq���+n�Bx�pk�9�*�f{����`���	~x��	��Eį�}ȂF��
Wĥ�R��WS�88��8�m��ëiNzK��"�%#>���K��d���Ξ������wQ���64�M�jn����˕N���+�cX�rI����"�f�D�� ƛs�3��Ȑ���_+n3����?������� �k���.φg�>���g�l �g�P���_��O�X^E�ɠ(.?��)1�����/�苂b��S��g<��s�wy�x�%�~���c������;a|U�}R����x�*��u�H<��U�"G���k�2nMĿD\ɻ�Q��:?���2BQ�?�VT���UBAO�%�m�x����V���||��v���<���jg���r7� �&7!��_7�sN_�<�|Ω�����"j��6�PR�`,ذ��������{���"\PT �:�%�C��F"E�M��������FG��W��w�.�c;�U%��yA7"�F��"��t%tv�)���eޫ]1��4���~�5|��g9�M����ٳ��gU��,�k����)��h�J�gMy���xi^��-��c|7o��bxG%�G���P�_�S�b������ k�[��H��w��p^H��G[�7$��L+R��S�0>rs2�� �\� �\f���]�T�u!eW�0�H�UN8�+l�染rq�~�I����g����ʼ�JrO�	35=
�1bO���j�7�^EF~�[��ҋ����Sh�|m�S�xܒ����FA���^7�d��:��=#�����,tC�wxJYH\g��:<�e�0�ĝ����IO��AH[嶧Kz���ߙ�KQ́~랞�C|�DM�v{0��D�w������e@O�q���F�)�0�iY�����#�	�O��-|�8��#�Ͻ֞��}�c�����;'Hn��^.�x*�T�}�b΢�8���ʈ,��5��J?�����[2���ו��DS�t����gJ	QI��6덞��+<�<�[��N0͞�ڵܤ�q_ ��H���̇Ƈ����^��]uw�m����HwЄ�6T���s�� oQhNѕ�e�?�b$��AQۏ2E�MI���e�u�\p�$D��X:�Ɍ�z�T�h��vk�����{c��'�B�#s��_E�/������w")�XW���G0���w3�2k���m��a�`�Us}~���t�dj-ʭv��˄�R���ܾ�+�N�jb�@��k�]YK�&,�XO,�.�R�Ŵ��ڀ�励-E�u�_�<TH�t��8_��#�,��Q�v"^Ge�=�OWM�ɧb�/�H��������
z�����5S��%'���`�,+`nz�6��2�0��vd��p��͋{�7<L�����c�H']�s<5\��sakb�?a�:h�§�xF�om��]ǭ�0��sн�'ς���0讝Ey�����> g���6�4@i;�!�������X�6!rf:h��UnZK����,M����LO�q�ٓ�х����0�Y�g'5m��ϒ��T�,Pjp���	������'�hg/��1&�SB�Y&��X�] �����(��}mc����_�0�O�����
"�T�Q��dG�cs*X2*��~��[_��o-I��5�G���ďB��.�!H��SklB� U���"��z����~��q���U��JyE>���`H0�ۭ��j�f��컳.�:�Q�<<3=�}�H���I���PS]�\�]!�mp��3�%)·�`�~��e�-���(��w�=�kBY7���mw���U�zSE-�{kL�'62 ���G��Ӻ�sV����Ƽ>���{�n4��O���BF�t'#vsfgq��Gg�,m��������.��E��j�t�Xr������>����{�:9t��^�ϙ�����VQXx_�.��"�N��n
p�3⻸U&�x�\GC���vxT�%��م��ȱ����rSY0 c�?^�~�󮔍^Z�r�;(�a��ij��HI!˥�R��(PRL[��{�2h�&���4�����,��:rC����`3Kl��1���3y]���(A�]����\I�'�-z��7��g��/����@�`V�@�aT.��!ܕ�`��ǖ�c�����R9]��BrC��u�n�ک�=��|�����s�t ���;V��ր�j~~�� ����,0+�, �1��R��H�����Awk�Ly��YKzg0���ן*���i�.%�n:a"]�zT�V$2EW5��虿G�l��qל����>��U��r�Ò��v��cU�Zi�%��Wx�҇R{|��'pҚ3�y:9�L��zm��nU���綶���)�[�n��	@�-�ܾ���/� DhЂ�}	�r&�Q�PW&_ހ���k�Qbg���G����ٔ�n����aʪ�;HQP�!�o��J@e�0�設���S��\�&^�e�������6���{�l�jAJ-���G�t����U�eaw����2B���'��~O����S��oB+?�:��<�Q�IHuzd�H��V��
Sl1I]9ؤy��@���p�H��y�����;th�sR�5S��_[0�ص�fJ>�Z%jG�Vm��5`k�z��8�_P��7����B-�d��C%���L�����伧¿�s��~���~	���Lt�;�tC�������qe�[�m@��&�nlH�e5)�cr�����)qu����w+���'Z�v�Zd_)�%��a�M�2��N{M\oA�?�ODf��Ф�b��屎^�d�nٓuر��X���'�����"0�z�U'��"���ذ�us�8
	�+T.���9����Ѫ@��F]�o%vo3����˳��$3��ut�e���철g5ڴhl�$�9���m�|$l���MA݉ѣ�h�H{���N[;J����&G���ܞ�A�i}��C3��[�>d��VX G�Um�_lI�,
��&����������<h� ��,q���#\��&U�Jrҕ���0�����8y���*��WT�*
�DEw�2gr+��x��H-�yYGP'_�J.ǕJ��Ҙ�Wp=ѻ�ܲGbk>�ۼ�ͭ|?
��hQ'C��k�?�C?ʂs$��H]���Z��Uu��;v �0��{��.�Jz``ʏ����4��i���J[���s&�:g����� �4�}��Z�t%��0o>AMC�d̻�٫����zL��v/�1�5 �C���;r�F� �/��k]��=n�e�����X��?�>J���P�N���amH�9'�ʆ�y�!�Z�KX̶�HGy�4��Ӯ[�9E�ʯA��	��)�{Z��������VnBe ��	��*ˑ�灶�n�r��d7��`�aV�gt�3XW�⿍6s��3R�ʁ{'¤��9��!z��&�ß� ui�����p,1�Y�F�T����.��IG�4N2Uv�4A�ƈ���h �jOk��=���T�T��
��kfgQf��l�O�/�(�.�˷5(��Ĉ�����[e��Z����NR(�bd�=�K+�f��O�G
����7y��� 
�xL��w�܌�I$G�g{����
��+��8~0H��{�x�Lr�drW�Q���,`Bl���(�h���ު��	ךM)s�>��D�ul�om-L�$��D��^D��tߡ�Lubzφ�V��~?�*��_+	f\=KtR>ʼ�QI���x��+�rJ�dR�֐�yF����I��Ym�<莢�����rɾ��ʻ����4���x��`��l�٫���~)�r��r@%�>�ծ��'К"cw��Wm�	���8��]�&Wp";VC�9V~�} E��2�yK�:�����_�����������^jv�P��o�i3����d��k���݄�ٴ�{��rE�I>�[��O��@���]�J�;�+�)�NKz��5�?qL	��ʟ�lȑ���>���2T5�FZ��?��R4z���R򖸑Z��5ˑ�>��2�� q.}}�f�����C���(u��Q��9�ޝ5�^.Uk_o�L�s�h���7)����ƈ��$���I��w
9,�ٕ�YD!$੔-2��]�nz�Ю��;+v�ڐ�o�s|��PNT�m>$�U�'�/���U,V��͢�'r&鎉��L�RU�U_ݔ��ռ�vB�HY:��9H�\�Z��4"~��f1�Ġ���b��J��Bp{���rلU�|N\�lC�g?���K���+�V������
e�9fX�l���S�l]r��k���R��(��B��]n|8PH ��;�E��}�s�v��a�Y%�|aE��I�X��Χ���{MO��C"����y����|�����ͥ'V�ŷ��(��y��ѣM���KYl��k%��S��$��B��c�kI�x�@���8;��l���������ʡcl`4ˢ��4c�ͼY��h%34����[d�i%s��t-Df�)D�u���f��'�52)����\<E��U���󻎅�(�G���+//�@�k�H�9rgX��S�N�4�|R�lٞ��������˴�H*5q��mrͬ�	�lk����0>��w(i�/����p�ӱ��� �F�T����wN½7˛�;OM��z;���d���a�����~w�|��n2����M�_�����������6Bu+�k�����d�Nku��ό��e�n�������������O�� ��SB���MFk�J��v�G5χ���́�>_��5k/�y �0C	G���Y;QߚJ=W���q+X%ƨ�lQ����.�HA��w̡�3��% �^k%�W�F:���Q����A�E֤��p��D=�?ך����O��'f}��v:�����)'��í��92ӊX�]L�z7�����5�X�W�`�W������인J/^r/�Nu[O�[��L�  }�W�Ch��e�F@��\�GԠ��P�O���B�0쌢p��tY�0�u�usZ�d6grxc��1$����{��B���?o� Qg����A{�ڼ��r:%p*�>���B���+תؾ~���^o����0w(Svk���1�1��ӑ����W�L��7�� X!�/3X����X��Jt=,���@���e�Gbbv��I�J��E)�ɽ? UH�*,��T^*i��������̉����(�)2����C�����$ )!�|z�1�7���P^9��OT��X�T�v��:Q�)��Z2������W�S�������@F��,i���?��"?9�}�9��h�B�-����f(Ú�Z�W?�����M�����f���:�3���*�H��e��	���[P�ߑ�b�Hy��uL����
��>��b�~~�G7i'�S!,ʄ(^����9e�'��G^Q"S������H8�BS���GL�C���Ɯʽ:��s4�9�Q�ƨ�Mg����~�,�q����)�.�fX��bz�GN������*]���+�jE)�WT|�;�h��=�\CO�s;yƗ�γ�)W&:�e �x�$��vm��T��B����ki-ߪ-~���$*�Ѱtc�C�L�I�#���a�w`�e��M»fr���6^>
?���g����MF4,��_�!���:YM&����4�`Iu�a�KȢ{�0D�skC����̀�ӯ�=���lߋ�]"C����<���o��n��`c����xұ#A�0]���h�|��*��r��3A�A�S�uA(;�3�o׵�]_Jw<3(U���!�_###�6���4�0�����E��D|���Rz�	m������* ��
�-��y�wI����4���~���6)�x�]T�zW�c��O�����ߟt����!|�z�zzD�&Zc��D<:�)�H�� �or��ޏZ�t?/'#��K��5������w�r���Xֈ?O�
,��+���h���C��?�W67#T�3�`���i5��z3����L�a��U �n8g����eQ�[��e<���I���m�š�>��J�	 ^w�ʯ�S��S��Q ��x�Hi}��}�EB���l9�;LS�:K��o &�צ}����b����H��I���o?~*C>z��yH�0�G��qyYpdɟĜ���s��Ov�;�E��_�ܽ�)'���N��*5ۜ}ӦkD�������.�J�7|.7t�^���3���V{t�������eT�{ڄк�v*�q@nW���?t\y��a.��U�����d+��|B�ɞCj�<�n���M� ���Ȏ��A�.��"2��*tjҸld==[��ly�ܬ����v9���]�F��y���Y~�>�x'tHX�i���+��ט:4���
��nm�������S��Ke��i �~:�&���{���'yl�U�O�<N��[��������}Ijr(Ijc��Z��/��O 6���fX^����}�g���t� `h�C��s��$Q���Dr���N�Ľ߃=R���%Z�~�f�1�jj�r��Z�iT�'f+�ު�2R���Κ
 }4^/	�ls�w���^�������c�>gC�e��k�wa�װ��;C�4�v�a'��W+y��VK�X�|�we�T�x� =�P����&f���X��6�F���!*���6�l�~�S�j�-nZ`�`ç��fe�I�.|�8���sս�b�r���|�b��۽Hf�r9�N���;�9�)W�Yn#$G������dk+h��Z}�����c�2Y�z?+��"�}�)�̈T;�s�~QQ$BYvۙFq؉�P}�CA��3�l�����%fpƨ�jIZb#��6C�-�a���R`.y��%ڃ���]��F�_W��X ���u�9ci��c&�J�[d�$�\�PF$AD�Cٟ�T��k�il!Wvg�J1=[�����М�5�a7n���i�W�+�Q1�Nh>�������G��9��l��0��Z��!�H�@�C�/�ߡ7���V����Z>�؋�aK.L\��$���d�<���*P�c7/@o��9�AI��ZÛ��Q\�G)Jy��Ht�p��I�*O����[��H�d��M���1D�P3�����208�S��k5rJ\��x���G��#YU�٘��1��m7�<���{�l��|��Z�m�j�.�{t���	0,�R�M����_�Mb�9�;��\����;��	a��>��Red?i��7�E�^�'+��M�2j@{B� �
��A���Q��C��K�>����3%Y���4��c0�6����]<����VZW
��9#];�[<��ݪ��%�	s*q͚l�G,�c�����y>�{X�����c���_+�]�ðE���$�����@�>�[���`D	����
��YB��4�c���o��1��u��q-=)����.v�,���3��G. �wg�1�4���~�'��W���9#D�r-`���6�2Ry�r�J#�o@��{Ţrg���5�O���3��z�b2��X}[�p�yBy>xͨjiֈ���gr��b*�fN����q�}�-�)ǺR*4�!�ll�)E	ɼ<18�� M0waa����$_�y�@��z7R�����`��"h��|N�a�^�C\N�G쀀ʄ��̔������u�3�fVY���L�W�a�&��<iRϪw��!D�ֹ�m)L/�]��b��קf��lY��4s�~]x,�H:��)w���9˦-e'�?T���Gs��q�?��gq�gL��ܵ	PQ&�n�#��~�B�Ó�b�2J�r����e��f��#�6b��~2@���9���|< AH�q�P��+4�.7�������Ƅ�s��R�?h#��<}z��g ��&���<4��I�R0�㭷�s�.x�,�1:�;5ϧ����}	�K��;n�.l_G�/��S�b�l��!��~͇��B=3��(ˁ��C�Zc��wV��j�nD��Z�2^���ͳ�tqW��d��E_%`��^��E�����_�Ϛs���sh)yW�]�"	ޟm�w�cL�kM~�`�σE�;
kfh_zѩ.��-^`"l=���}K0��n���,����\ܴ��f+�����2�XF���W�`}&�N(�#�Kѐ�-W{�}����M���	��2<��c��*��kU��}ǻ|,�<�3Iy�ohͱdJyT�LA;@����|�O�E3!p���:�0�#p�;��,ј��O�N��HS?Q��RWO4.�*�/��^p7NJ"$��-��$�t?��:�k���z��]���an'��(�`H�0���ϼrK���s�z)[�����~�vb���5��ݥ��o6#D'�#'j�G�y�}��~�u[H'	���9�c�ӊQ(�����L �V�Pa-#�����jU5=����������[l��Ք~����V8!9�/+�B���,鎅SE��]�xz���S�<H��E=�S3�c�-�9�"H:h��>G�1x�+�-��Z���*�2��������+�W
�pL���,Mo����T��9����1����\ؑ$ZG���oO��.�yVJ�7C��$����z���WD�jC汛��)F������:���u,��QX����IOb3�L��]����8lB�d2��K���d��>�
�[������c���9��d�J���-t�Rb.Q1L8��~��(��{{E>7ӌe��a"Ղ����9�\!��3���~{�y�.�l��m���,'�"��M����?,Z��<4�d�.��#�� @��N1��b������nB�J�m�)��Y��ڊ����hѤ�km���2���� ������56��-f���;q�\鼋�E�]2f����b>����Z�/��$�6~���?��|���ui;"vy�ɥiێח[��D~����x&�%��T)�. I�D	�*�<.�ET��?r6|L�&������C5.���x�o���7�d0��'����k/�q�p���N���w���`��5�0�h��;��z�!	�_ArרOʼb��߼��,*�K;�|l�(1�2nAAV��q���\&��~8���>�v�91�k͈փ�Fz�r�}��¼�wr�tTi.�$���X`�Fj�O�v�r��S5x���1�������Ԥ����\v�*����QUѪ��EJ�mI"ç�����~E[NE��Q�&�>�y��023�&�jt���*H�#�~�3X��ru��"brU絟�"_8�-J��&�����{;��{۫��1�X�|�]��=�X~Q�K�g�V��,�8����_u_m��eX]]������������
߲�u�0%��GK'�O|Y��V�)�RC�Ї�Hc�&��{�O5HW��2i�
'@?�Ϋ��ّ�o,�@F�Øl&��o�҆�vq�����s�!�I��k��aO���c����ϼ�*s��/v+WY�� }c\c�W:Z��,�هW/�[�mO�K�a�{��
PAn��%W�����>���sOK�Ig0�Ӂ�W��Ο������0�C���K=F�"t�=�%4^��'+��5�;!y|:B�]�Ȉ���~�ɇ5=�ݏ����bb�V�Q�Mf����T����Y�	�V�I)F��4z(-��<&~���#Y��b�q��I*��p��ٯ՛w�:ێEb�T��f����͵'"9����þ���]��Ӝ�,�n#��H��$ȗن�vv���`���"����&1�~��.o%�(9�Z9��uv%��ҩ3F���=�}��`�(>�������8-i�V�9E��.�>�3�ȿ*���>u���]��d�}�c�.|��wL@���������`i�IӢ�7o6݆�����0d%≸�!>�-]Oww������ހ���/���/�#�-�V,����t��AZ�/��RqC�t|�7?|��0`@�d�hD��?���d���|H�!䃈!.���a��<�~1�k"��A:f�N����J�4|���&�X��.K׶���JQ��ABe����%���+F��ێ��:��C09�T\�s��m��VV���̶��CB\?�2���ϥw�go���(��.=�$�".>�%�ؽ�f ){��N�s�.WM"2K���Ez��&R��s�8W�nB`8�8�i��VG�v�.�)��K��w���Ǯ��.�<}���ƣ?.s�]�/���U�R���I&��dJ�eL�����F%�50���We�y,�L��`j�S���#%��\�f	?����N^J�u���t�g����˳�@aC�M~�W����tJ	����jw�~�8�r�����]!	2B�)Y���N��M��	&��%�j��o=�u��ִ�So������]�;�ʙ�	��=��6�q�a<+[ۅ�Dl���W��
**�(((G(�˨loIz{N�&Ұ3�:�P�{��g��,Z��/��hKJ翓�8G�:��d�Գܮ�1���Cvke����F,��:�+�T��m2ۚ��3ٚ~��$2�)��(T'���:}�v��ٺ�S�]h����������)�P?�'���g�Ek�N��XTT���)�Vakx����J��ی �# +��n7�Vg���I��ñ ��e2)��B١g�<jAq-��ĸ�x���h�m�]m��B��}l�HF`4�<�D�0η$�=��I�`+�#�L��@4�t4���f<S7�|�,x�{1���K�"�s��GOL�,^���O���|�A��1`YǸ��s_��668
�<��������-P�W@M��e/G�H#�W+�K
H�<Lّr|�
�z�8�X���Ԕw~�!�H�	�^= (E�C��H�d�����q���<$�Ή�D�ƈ~��ȓ,�[�³r����	�-�r#���dt�q?I�?��\+�I''8gd�-< +�!��7��r�垆ag�H��x.+����6^�x1se'AҸ�}���pӸ�i��̭�/�믫������q�X��4,��j7V�Ν��KR�;#�U!�|q�O����Σ�LLR����q�x'�x�&�����58����%Kd]P�]��Hkg� M�K�S*u��S����^Q=[=���v?�G0}�Z���:mu�"Z��e�}I���P�.Ǳ�]�G�kM�a�Q�ٲ=%���=����@"�eA�r�Z���B��Mr�����xd��J{th׳���I3c���!������)�f���m�#\��7��=���W<��R�8aL`hӨ0��Z�lw�쭒�S]�p��p���gK]D5���f�%�����ڑz����;+����[�MB��܏������0Yw	�
��"���`�ٶ궙���S�oY�[�HU�Ӌ�N��W�
�Ŕ�P�y5q&�[���̭��k1
�9`�����Dqi�>��#~إX�i��K�@�J�E�~z1B��QF�>"<Q�}�B��f���^b�y�#�3��S�o~����浊+'�G�N�-P�J>�
�iǹh3@�m]Co����ˎ�;'Q���2~�� �q��y�J�����NTk7��[��~�0��d�)I�6<��_�'�@o��K�Gə�P�hM�eG��JϰgՅ��"s�rj�wo��孶N��L�B���h׊}ފ��cRY�۷����Z���t�sڥS�u���*�/����rv����o2m�S�m�r5�4t	nu�	G�|`�[��������?��:# �:�C���l%]#�*��_nƙO��Q�(�h��ԖŽΈ`Z{�Q����G�Qݭ�R���卍�I'[��4�'�\ؽ��f�"�w���А0�l�on~݂)�^�J&�n��N�/ޢ��in��*s�9>ɶ�H��s���C,�3�q����1�e�g�$�Ӂ�"3��C�MU�&L�u�4�2�����������S���/1v�Ki�U��+�QKlj�%$ĀMe\aBնR���+���b�^��ڞ.�v�q�N����B��e������m� �  ������w��<�����R/���'K�Yx,őY(\��&�����שm|��q���R%8��X[a���X2K���˧��!����6�d,��¡^��i�i��d�$h���U�w��-��AWiL���u]�[�kMC������Ű�3����iO-�Yk^���Dܲ]��Ŝ��S?���S۳��*��;m"Ͽ^�(�G`�ө���v��ϥ�YXc�=�#pG̉.,Ҽ�fT�QX�mƑ�H���Jx��Ug�:�)8a��U��v.��&n	e�uI�u^و
�!1q2�@8�;�Q�Ol��l�e���j]�a$) m�R����PɌ�K���J{�q��Dk��1�ulz���C@�&�}
�����%I-ޥ����,]�a�� ,��VH��+�s���d��+i�����M�ȶ:P�`�	�T#���6«�R�r-�,8��j#�S�I� ���q���]����+�����98��?�*���"	�im�p�r|��v�B��~���I1�B��ӿe�l�F��A�\q.�M�s�M��z�JSÐ;bʠ��}%��Y<͎5b�Sv�W����j�<�&��22v~�vj�aVj���fټ�(�����ʐys4��?�Z�Yki�%gK:�(��3�|���׫����A3R�_oV4ޠ�.^M��gC��oMvK�E�a�ɀ\}GW;��v�}��jhp4z矽�pm�&�-� �������TWN�9i�MÓ=j+��]�m���	q���|0���I��M6��O E�N�C� �1�yD4�g��X���?��Hr2O�[$�*����A��'����7I.��.�#E&��	�k,���n�G�?<=�a�3�s�����y�		�낱����J����$zm���U]���eɕ�,T�Ay��VI���T���}���Hx���R�͂G�w�0r� �����O�ı-�T3�H�t�9�<,�]�Go8��	W����2�i�RE1�3A(! ��ͣ�]�0�����@t{���h���8�BJ�j�
H����#�i������#���ߖ0�j�@)k�r�)�L���V;q���3��h~9VƄ�L�������'1���\�͎�( F�L�Z�s
�`�{��u���I^�_v��\��_�r�hD����Y��d���n?ՙ	M�����i�/��F�5�a@�Δ���N�����oX%���'�/3���s������Z����iA�8�Z��ݪ�?bsF?C�\z?v�V��R��U�z�CIzVp�Ҷ?7��x7����4�?�h����T����.:�h�E���:ˇ��*L��k����u�qQv[��A�kHA�KB�nɡ�;��nQBB��[@�BJ�������?�3��g�}�:�WbF���H�;�U�6j|,j$��K3�j�G�/�����U?M��`F,O3[xz������X�T�5H_s;<Yϱ����<���^�^:�X�[���qt]��GK�@ʞ�D���5�&ʱm���a����z�����k����I��d���!���0;��R�A?�1�ȖG"_�w�Wa���jyu[���n�J��E���1@��v��m=a�k��E5����R����gA��wBV[�3�����rth����v��I#eqS��2�-T:���@��F�@��<؀ȞXHz �M���wg�G�	����m��#j���_W����'�s4�$1|a�M��ɿy4o�/O,�6�uN���V��?o�!�Y������k�l���G��dJ
�ŧJ^x �59�����*&�L�K�9����7	?��{��>DE�����R{%H�}��	���u�-�!�Ⲩ߻m9��=�%v�Z6�O�e���%���u�\z���<��"�����\$ں��j�'��-o����D,�(��k�iG�E�si�+V~ �F<�n��iX0;��A��y,bX�%�ڏ�#�
fD9A\�
�D{����O"n|�� #�Ec�+J�FO(�_�B[�բ��w�SP~c�9g���sJ�ܪ��?AD�W��<MWi�)!��	בή� Y�]n�u��֪ʕ=?����9�ߴN}8w��H����Q�^�U�?���?%��?2j�#Q�Y��o������$��-�ymR�iǇ�$�sL�Zhg=n�8k=E���aQ��C��d�x��0��ꄊ��r1P\���o}f�_��i�	:I��9����憀��Dy����#������\�37�}�.�B>��&�.�aK$��@�߼V.�$v�T2��!jk����I���\M��JIGN���#��g)�m�si�d��/�n{�#6��)%� T�s	E��[�LգX:�UG�ˮ�73-GT�6�c�c�g塀���힠�M;�W}�.�H�áT�7��m��#0}y��t�5��/���s���d��2����5vƨ#����S�6ǚ'*��W���T�$�uՔ}�s������>���1��s�o��Wl?뤅1��9i��������ve��=`�"��� ����p��Uƛ�	qD�8 ��N���l�5�l��뿺,�g�(�`��;6ʡ��C3�_gv�[�v�����3���n�C��!=�y�H,D�����7'`m��rSJ��A����|*�}�M�,Z���������n8^1k�m31Y�iET�|�R��G��T�11�n�5���ܪI�{ =U�XNl{��#w�v���f��L9�+�v�g��)ˎd��&��B����u�A��d���fR'<02^�wG�}\�$@m�u��Df���yS�����X�Ĳl�ڵX����}#p?�X�q8[M���N�{�U����?���nߨ@�El��c$ڈ�r�#��8*~��P5��*.�&�a����Uφ�a��Fb�\5���
�f{�ߡ[ٔ�Q2W��?����y���x��l�<�ir�m�.Y���2u�>r�͓[@۶�8��7�-���u����m������iM�<y�\��/vNJ8�?�Ƴ��z,���$�0����U�Ԫ�>��d�{<m�����Ã��]b�+L҅ԡ����s���x������:��:��pBA�RR	v\/�4���6����To����Vq�if^��=y�ϑ{ͯ��N��{���5�%�;�A��u`amB#�߮�T8�|�u�rX�U8�*^���i����'e#vH���@�b���O�Ǥd�����^�u�Si
��?�7��W�xi/��9e^��1��#�x�- ��鼰`���
.�	_t�$����7�>��w�����P���(�O ���{�VӁ|�(��UA���x��:v��K���P��-0aʬn�lɫJ�2�8�y����k^��YH�\�:I+c�O��7�ث���\��Y֊�ݨ�἖��Uȕ^!Bg�|]����x	@O2��Kg��J(�|'���˃����.V|W�(���T�f4��a�!�i���W���Ϸb5�n������,�!
�yhN:���w�x9G�'e���61�*��S��9����o�RK@�{�s�&��0%�]�6��"����=]@.����mV��w���q�y�2;^�v�K���ʋN7��� �A��k	^f����`�#� a��b8P�EE
[�E�r�.m3PDXy.�2���R=���8�.a;ӧ_��Ew�'ߺ�.���6�Wy����矼��(g�TN�����Ez�М���u�����s����uc�;C0��G�6��X�x��� ϴ����g�B��)��]'���5��/]��d���MQ�*� -���3������j-.�(��`e�9�~T���~�غ:Q5��%0�ؚ(8�ٜ�Rw��y_��c�m����tb�kR3>�yC�Z�ݣLa�>��T�2�5D�Vk,��D�u���W>
���R8�ʙwt �aY�U��@&
�,[Q�1j[��o\�|�J�]o�=���p�"Q=.K��G�#�%��m��oW4��2�v��JP�۫�Bz���'㛢����H�,��嶳�?I�����\f?�2i�����s��Ȣt�ૼT�u�E��9�[=����~L�+S���m�-�_�}Λ�̠��a�ٍ�C޲�٩�fMj�x��}���*�GP5��i�.�3Ҟ3�W{)������<=�^�98)��8����ݶ�*�O�c��v	˻Q�y v��[�4V�w<��	Nrl �fN�rՔ�n��R�]������q���\��r�*�i}�}	��%�4�|'2v� �O\�_}l���R���7�Oڳ!v��w�&O����=M4�E��̣�rW�g,��+��F{lӅ�+3n�<ko�/�Da�V=�O3���@���	#V����7v-�:���*ŏx�R�c�Y|��6A�}D�HKR �ON�+��L�'IG9�?{(x�J7|pYퟷ�|e>g�O�|��d�;8����[4}ْ#�[�c5�ĹɈ�q�|��^�V_���,A���8�+�gKXz����9F��Q���[�Y���X_=��'���f ������s��������jt�S��Ti�Z�*t�L�k�glo��t�+�ӌ~1��ĺs,�3�;G�rD^˗�QS�!��'��k>��P������?&])��[̚�F���s��
Ь��n���Y%�sk��f|��!��r��	�����)��@��]�W��^'�a�Q�,u�ћ�j�C��n�0C��B%��H�"�܆u˲�b[�B ���m��jyǪ9�ܝ�k����3t��*�ڻ���:M��~�cd��y�f�K���*-;c���_)�@�)��9`�~�X
I6bWe��^�>K���Y�ʛ��T����)̘��|QD�����S�S�.���(�:�X2U��Y�c�uKzh'�MVրۇ��K�vs9�{�����N,MϜ;���}q�bw�r��L�����j��b�udsР���;���
�ƾ��+��	����AߏYn�`����p�𾨄V� ]����G�E��65���Vc�,c����o�����T���G7��O�B5B/l-�����֛}��%�EEr��AQ'�x����ߔ���Y\\�`����饵�?}-u���t�Y�E�	���9��Dn��2�x����J�0�4��^�e��������S��
�^̗�`Oz�����Zѻ �,������C�9��s����L���R���1��1��g��t����(㔦�;�3�$�������)6�q���Y3��*��N2%�`̐hu'�l��&��Bu0���\��F;�Tc�3�ʠ������CM�+o���B��x��4D�!���	%u�O2�cY�\;f�a�Ҽ�����_���i�;���9�����w�2�,�(��{zÞ�W�~����C�[�R"�SJ6�^Y��1���{%��w���F�:���)b:��k�2��\����dV\�G��y<��_�fsu�?�k*���	��'�c��Br�v��Ƈ����A@��~�I%�C �@*SG�����x��f?�-<*���u�S����ס�Ɔ�r�1�ei���BXi�5#H�'hx	���)�&2��QP��GK��?�y�:��n�fFN�&5�Њ��x���h�wm��o�Ve�eY(py�ڱچ}�+_���P��F�eK�	����A�/����ʂ��'K
c�� �&�S�OR�`��M�+q[�F��������f���.E�� ^�i@�$j�c��)h���CT�-������d������yL��ͲqD���2���#����ﺾ�v��N���P]w�Y�*&	�H%���@),A_a���k0r.i��v~#>���?�t�@2���wYG�4�&�7:X:���a|C�&c��q��4��\�rg�GK����ejJUa ��S�~�l�m�"�&)	�򗹮�9�?�%Z�٫�ݸ]�����]@z�g�z��`�b�wgq�G��9Jof���O�Ҿo���o*cch�D���4h� ^�'�<�`	$p��y��Ү�?��/qO�кW샇Mo�7�D�b昹�}��Y[W��	I�9G�Z�M�'f�ӭ$��Ǔ3����v��j�"?-�|D����M�6�m�e� q��)��ъ�Gs�#-�]�R���sa_.��_z���z[����YD��e��L/ի�r�11�f����!�;�T)]QG']��#��z�o���kbVгT6��`dLeoܾ����]TT�	�4�	>�Ln��1j���#N���%i�[��ldI���3ޖ?Ν������6j.�����ޮ,Zv���q�2�s���@\���4�i�X��'�-��t�҂O�Y��!A��x�B�`��FZi�>���Rվ���C�T��
��V�L��ږ�+���C�����	-�VV�#B��_�I�,���OA�eoK~;�,:Ru���9�����}3�d��\�8� ��V�{�yA;N�Ԫ;o?�j��?Gˬ���8ϜJY�8q{Ѧ�ྛ��~������>CE��l�B�Jtn�n���Ư���ޑa��б�w�ܢ�Gn�ۂ��Ai��lݱ�m	v|p�e��=R��AY��}���i̺�vop��� Q��J>;Gj�R��nU�,n�b�����v�� ��q*�um�w����BN�-��)c�vl;o��A���܋ �Q���ϵ�
�u+D]Zib�Sn�pd��v����#�T��;{��MYU��]��]q�
׋<�������>C�UF��j�T�{_L<L	���Ů�K���ڗ/e)W^���u�-EM��?�Z_y&&���W�럆�>�z��5�~�s���u1#�}:�7u$uٶv�y3��93�yh�Ԋ/Y������Wl��w���?8�O�Dq��_����9xJ�z{�ځ�_�F'��`�=>�|�LJ0��Y)�"W!-m(�������ͪ����$���cX[�//�Ok)�{+>�{M�����b(�	޺8Wc�ױ�Sa�$��r ��r5�e���k�/����m�G����aSpD�X�\lNN�����-�'-{T���;���-(	�+5��b�(�iCf����'���Ǻ�+ 9u� %�V��e��*���dB����VC���p�cl;�}B�"�`���3�/��f�l�-&�\��G�y[�گ����v/��+��%!&����<5K>��� <�_;�|��л�O���x؇��Ii��-�T��ee��$#hظ?�%;�"��	���q
�K����?jU�����yWP;���V@}�z=�_^a{��z��X4�"�GO���c-��7.7�կ�O�[O����z�{	�=��Mi�`rʢMoF����my�a��_B�a��D�x��o�rA������%yp������@*؏������K�������Mea݈����N�$9�S:��d���Q��i�ZSUX�����߸Ww�z24��(Sz _.鋻t��y�ތ�=�tݦ���:݈r�[j�){�+\����0� z��wp�� Gyj�S�%���a���L�h��ƈ�j�3p.(o�z�����5��ß��~Ǒ!��S*~U�?�+ZIB�\��ĺ8�+�,P����y�VLf�#R�Z�"�L��ȷ�]A>O']l���+}x�ǎl�鈆�blJ�p3�2��� �5g�V4+dXt�{kȷ�VEҨY�4^d�8�U"^K�J�\�p-���ͨ�'ʇ���VsW�f�n���7��ם�Nb��o�Pq�Vܩ2�H1�~@�aa��C�@��zW=��J�n���礯�(��['c՚f�4n�#VZ�EC�Y��h(4�iH4�hl�O;�����9�:^4aW��X]�"�"��zugh�	��OI��mB�����8"�4  +�O�L�d���=o\���@О���>��H_���Sh֒�Z�񌏝�7)�W����*B��1k����;����[���������	=�ԍHT��)���l�+��X>bU.�����Xj��q;����A�Ա����7Ib�YI���^���.�
h(�*AV�Y��S��qO��4u~ff8�^8=�ܫ�RS����F���G��~c��Y?��ƍ��?t�$�HJ���lɽ�UϮ�w�`o<�χ �N�LCc���T��w�3�͇�D����� �'f%b
� c^mޜ��p�ZM z@���\���c��Wk�f�x�H+WwIzWJ�D��3U9(�=RݝȖ��t]��$�'����߮Q\m���ԠF���	����˵�MZ�#���@&���C�LN^�6��spay��hw[�ĥ����\~�-�u\¢N�?|��L�QSŸ��c�f�����캨��ۏK=Mع*���x�����\��+�T����/w|���oU9��>7l�g'����3���&�� �Gσ߶*�Atz�����!���<�5�ߕD�O w�4���Yn�:�D�[���:YA��Z<������6��V�g�a�\�$|�Rl��B+�o�Z�1���W]
�ӹ�U���vclN8�5:�އ�r���ʦ�.�+�:x=�:rq��� �>��A���s�~u�������;'܁ط7r�Y��=s0�F�	� !��{w_:�d=�!Th�AYvZ#�3�)<����$�g�E�UQ�|^�F�	���X��P��J�����(k��}���������Q6�<�=Օ��Q�s�S�^�����&�Ou������q�g��$<�~G^��S�5�)����0���}W�~���C�&	���
w�N�k,��j����I� ���!r���S2�5�9"�
�����!�¦�Z�61���� (�B�F��,`[���%�$ ݙD���������؟��1���v�g㈓[��F�BG�lQ�m9�*O��������z���f��{pwG�O��Dx/��R���"�n��~\;D��1�7ܙ���^�۳Op:˾:��b̥�20�9��TU����aI�?�,Œ���<����o��� ���PA/���vċ߯���e�5�
�C����ߓ��r���8��B�}�f׉+�V��V�<�ۺk�8��.ͫ+�e��%����I�G��Alw
�_�]���<�K�3C	[��e��{������;�j�^��q�4������q-�VN:��j��1��k6�q#�%�|T�li���J;:>�� �]�/;��t��(:y#�����`QO�ǲ�oi��R�9r�x Ҳc����g��g{�\R(0�Kr�~Z�'����/mE/�`���pWc��4�t�\Ow�O�V2�!��6�Z8~ A��֕/�5�	$�h�7'f��x�^,!鳼厞!��A���l�����<^<͡���9�<�C �v��6�
��ņ�0������R$e���,���{��t�v�#����Yn�)!�qW��j6Z�{��k�$g�)d�����=�3�c�Q7*,0z	|���OU�tli������ێ�bH1G������F�����$;Q�?b«?Ѷܝ�)���kP�kn<xE�1d��'��,����Q��>��� ���/{7�0\�;�Z�8��M�6τ�fm/���\�"�W$�����lRq�-�9�̐�$�tqU`��y�聺�W^Z�|�����R;>���U}���%c��/E.}l)�O��,�T�}�q
-iJ�z�(�U9}\䷩V� �a�����tW�W}�����P<I]̺"٠��߇�)�9���7�G��7R(���>Z0��xM==��{IN�a�H�i4��.���E�Z#�|]���!�dDSC��o8?���y֡k�25�.F>����H���+̔�f�Ub�9^�r�aoԧ�t��;���~������y��V��"���~l8^�N�.�(�@������X}�)�v�42�����,B�wp�h1*3�>m�?e��LXx��ʂV��ZՅɴ�\^���|b9��Id%| ㌣"s���&a��`�@��+�#�b�dc�����T�I��E{�:��$�a�]��E�$j���4_�iaI�m`�JI���b:0'�b`}^�_x	��{hzaU�!rk�;�b���T)Qu���z�:��x�t^�p��K}���;��g1Ƒ�á�X�n�i��a�F�ޠ�8�ٓ�S�N%�7�S�!�S�u��)�|�` ���P�_���N{G��P1h=����O��h�r>����O�6�G���fS�O�����m=�a4�j��(%}���<�1D�O��������<�*xߏu�X�a+���q�nY3���Np'����-_�*��:�����"��޲U��Ӛ��]�L�%\O�ɼ��ܔ�Djj��n�g���V	A���čh��W�$.�������t7~�f<�NC[s�N����t������ղc�vPeB���z�ӛ����NN�gCM��y�F���"CU\X���2��CSR��|�!Cdi����o,���ݹe�G��cҌ�(CW6@������S&�N�l3�(�,[n�v�E���)'u�Oln���
G��K=%�e���d���Ǻ��T�&-��@�}�< ���A�l��f6��elzb��m�fq=��Z�����\�ܥ��n�=�~T�>��^��]�����}c����4�!H-��S��Y�]�����鬓�����ӄ�b$�l'{�Z���_��]�҉�L�~{P�9�m�
��tƄc8p���E4��LT��;�-Z7:�T���x�wc��B}n�a`�V�h`��ʰ�p���K�D���c�ѳ)�,+�����(�}풃	c�$��2@�Ggg�j�4@�	�8�ā�L>��=�����_cc������`*�e������aE��
��R���e�n�[c^�R�H���G1�b{�%�k���8:�Ōff���m:
` ���K��iz����N�b�2���m���^��N�����E���.�UMw�R	��T����+��j�N��FD~��2��\�c�'�߿.��f߇�D��!�ך�ٗ�[bMﺵ�S�����A8�!7}�I�	w6�׊���v��ay!�&#�H�����G���V��ϚF�e��p��z��zm��fu6F�ɽ��k�	�%�f���<�P ��#���'�;[[X(�{b�@�ъn�,�kf�
 ��
� ��3&v���ц
��\�gU������c��ڥ�,�I�[�'^�����q�sL�-�Y�녎�'�$�*q�D�< ��J��7*��3�R�I�X�o�b�V��]�JO�n<��h���~a��0A|�kb�:��ג��5��i�x'�<��f�ȝ��G������ ������e�^�&���3���?�B�����5 �x�<Y���WA+c�'��/)���"C�w�\	6�dʣ�j�c�U�MgJ/�J��[�K�4(�����T�f��tżR q9�����N�_ruT&�o\Ԟ8����g�q�9�+k���2L״jF&��2Jt�[��o���%���Smj��l,pAm�~I��8�h�ܖdW.�j	K�	F�!� V��nT�4;�������o��1{�Y�I�f����;JP��سR��"�ȓv���hff��$��l�m��NnL38}2�7�4t1�Vn�ww�N��P-�����hܦ�(�]8�V���b/����O�y�F{��NՅ	���KP�|�t��eM@�@u���n�o��qk`q���P�i��t�޾��Lf��2tyvC�~���o"�酅�������0�,���N	�U�V/H������㥠��.�b�k���[����ȡ_���.4=���_�qd\�[��CG��5(0r#G�#�X�b��$�x8#4�tSӹ`�l�y�ө-"[)`j�r�p�C��:����vϮd10>v�O��Z�'!V�>�aj�-�llv"}7��
��hj�:�hG-������Px��8ޟdl�۔��dcEo��[�d�UM���RJ�$��n9I9���}����l���yS{l�7�����7���^�'j��>"W��P �e!���2���:s2cp�UT')��2�B�j�-������'�d�rhQFfW��$��W+l%���Ol>7zM�n�/ϛ!Q��LFh��7�"b��"��m��@l�H���
rA;���kw��4��}x�Ҙ��.S�L�:"�F&)�^ږl1�Ix��Ϥ�c��T��>5�юt�ȧ���9��S-���m�(��$y��`,>���Iw=���QH_'c0�7��h�e�į[�(Tqhw*s�1�2��~���E9MȹZP['!I�-�`!=Zf�0�?ԡ(�v�q�)�t|���,ȵM$�HR}��n��%��S��"L�uc�6�y��%Ͱ5��rHam��w?�"ĺ&�]2����u�AH��ɦ*�}[�p�<�������W��]��A�:��.y0lk�0�t�Xtm�_*e*,E�t��X�%����R6��QBI�7��{ߡ$(�6�P~v�ő�Åx�kEV.�JZ(�[*!B$e�k�X��7�3�����d��;7�)���7�꧈m+�$%��Aۊ�"e~�	����bJV���ָ�5��E��ϕi�����j���2������Q�O��v�C%JV$3kw�VQ�X櫵|����6	q[�@|�My���e�qzp3{���7�9U;�
����::�=W^����L�9tbN��H��Xu[�(�Lo�oч��j��E�w�
�
�0�cqkǱ�6�x�	�L>$~��.ŏe����j$C}�	Am��S�'V�*��N̡7��?M�n)�����>_�(��ﻡ&Z��&�Q��@+�9Z��I���^�y�顭���sf��>���dd��s��6�pd
�o�*��9��±]ݷ�_���4U2o��������{Sm�����{Y-����^7k/4�ǥ����#�p�����n���x���b"ymbV��������f~6im�;i�j�8�/iSR�3��g^���\b��)	t�b��G9�Ծ$�E�c9����[��hv�w�;�N5�5.�v0�l��ȹ�I�T�hf�-�R0�D:�诎J��
Rɠ��۞^�Ψ�~=���^89��s+++�-�܎o,��N!�4}�b�G�!"ѿ�T��`WZ�X�:����)�>(up�v��^��Wj�c�]]]��5.���6�؛4�遇Y%."ps�s��k1<��W��b4�/��n�'��Ԇ��C��H�'��V�mUF�J �ĦS�;_����U6�Z}�Va��ܳY-�P	E��7ה��/���~�c�٬�8�~!�~��DP�g8�:My��\o����	ƪ�3�ӻ��cb-c'v���0��%��o�<+�U���C�=fI��c_:�o��W,숛�W�Q��-.��9���o4A������w�ED�=<�E���|p�!�RoJ��-˶5�q���r�S���}��������h�<Yi)U{�v��4��Ŝ�Os�J��:�^�(x�tb^׼�2r#&:���$�&����֐U醮-QV2�S��Ȁ�y�N�ܙVh�n���6tc�!ĔMhK�w5��T1��F�u��%Ħ\��a� ;��z4
�͢IƬ���I�P�)(���d$B|ˈش�9�V�$�X1�q�@{�#�'uК Xs�sPO�����v#��R)g"�Tv�*Qjw�e �g�;|y�k��yԴ�Ք`l��4�1�@���^��_��4�)}�j�qe�t�o��r�8�N.wy,���:��
�K�~�b��*߯�sa� �F��̌�����+!��P�R�N}�����&8n������+k�2_�&����ӥ�xw���дy����KL��2�EK����WLtD�F	�܅E���l�b�Nt[d,mpy������,�]E�Vt4�T�	Vwdr�;��EdY���ߔY��nJ�;k�`EK� �W�:�#�ve:��b����-x��C�6�;�)l�N3Z1SN�~�n�(��iٌ[�0�^\�>)E3�HSfi���za^	g�K���ߌg��KRђ-���'P;����� F`wp��(�X��T��H`��=](���ʔ��΁.YPW�Gfu��Ύ4������:���C~Y�-��Q��b<^��m�z8Vk���P���4�-u�V�m0�*�_��д�;��5�<�-�p�Q8�X��ru:N��p�k�KiP���&��X&�9ƣ�,�Yo����nb]!Ŷ�I�wR�a9(���7�
r�]d���u�r�Խs�F�����AT�!qe�t��2ce}�6�0+����4Ժ�N୺�I0a�%�����;�r7�:��)��]$���6��V�6 ��Q8��>/��}����w��NO�§�~�y�8�#B�L�����c+2����o��m.�g��2OV���tWR-v��p��4�	�,�ל=��s��z��݄>	��ޖv�j)n���0&K�C�
�ʞ�7F��o�������m��O�퍯{I��¢Gw�h96`�2)usv�L���?t%��\��1d&�S�����6CC��}Ϗ�~m2��������D�E_/���|��� ��?Et��샌<7�Ev�׵Cz����VO�YcS)���	-����N�c����/�1���c	bm�/�;e-�*S�b�=r��Zp�"M��!�G�]v- 4G�"�Rס~�I>%J�<��,��=6È�$#i?Woy�vI�NR饫��([���{�q&+^������})h���Y�?��\@m�����I���ޑ4��-s�/:_��dV�B�x	�
�v)`�|o"������~���xYD��~��]"\B!��Q�ͺ�i�l���tM㪻>O%&��q;sl�oh�">��ӥ$LE]�x�����4�E�W���tp?^t���a����U����x��U�����u�5gŅPƄE��c_�����Du��l�zq7lU0���a��h@��6~��˫oY�`��"<�L'Qs��֥��#�h�J��|$��爡b����T�'��Y�����i_�su\$}�f��lr�vS�0,NBũ��Ѥ�U�E����	�v�f��I�>�Z��L����_m�vF����(W���a8�<�sl}��
���)ʱ��'h�	P4�'
���\9��\�3���v<�ܭ��`�����H����!�M]�@���95G\���k�q��0_	.�A��pՀ۟���4��̩�Q (�y�ˀY�"����İ���&�'%[���ʻ���D&y�&I'o={F˞�z�iNeN@7:��Լ6�}�@ry
�G@�f��4~�d><=���U�_p >��z�9�!��f�Ie�d?9���f*��ڗ������_f����W�p�(���X�H�	����XL"v9�i��O���sy��N��	���i�I�F�o
D�[-խXg>��{~�8a��l�A��IO���;��]��W	u�f�t�-<=8�R�o�nQ�S$��^�7���TJ���m�g�K�c᧎%d?�#��j�ĝ���������N�������؍��ҭ���s�+�Wl���^6N�*Y�I��?�����]�(�X�B���9�|�{��Yh���� t>��ĕ���W��wxo\8
�:S���!���o6�����FS�̷3�˂����>�gC��=7�+p��m�1�pt]��c"���a�"�BH�NSK�3={�γ�H����xY3��#�&��hD��Q-W��)�VJ��4bߚ�� DZ��646Fhg���L�aI�<S�P��`��^���<�D���O��j���g7��:z�z?� B.@sN��N	���ѭ�sN���=�����/�4+�!�P��f\'���"[� �������;��iM�?nZm���z��VSg��V�9�-y��M��L��6�_�<�<v�5�ʷ5+�B��d�>	��۞U~n-Q����[@5�.'E���v�$�k+@�FK�#���~2�)2l�.\q��q�SB�"�Ԉ�(�r�˥<�h�?dxJ4hI���s遏P�Ҽ����KaK@oWks��!kK�}||z^}Rκ^�U�~չ=���F_�#j	�k&,K��m[�w��V��|S��������j�܄[��U]M�s*|fy��zz�'s����20la�$��@D�%����jy��Ja�i��%.��2��s�)���W��j %u��Q7U	&(�oZk����oU����;h%��(A$�e���������7�R���-4�z�Vt7�2߲X��,8�X��Q�U�f�a�x܈��$�Ⱥ;ۺ���~N��_d��|�.��ѼȰ]L�RH�u�� ���[���G�iB7�����	�,��M�|N���B��lu�:Z�4N�\5��x02f���#��i�*�D������G/�������:(��6x���L
ۊ�����b�Ր�9��� �ͱ�����H����('U+
�')��!S�k���6����я����Z�C��觛� �n�S�~��I�Q�4/6����#}j+�?Ic�0�I2���%D�qt�I4Y"�mp��P>��Ó5����!0���UI9N�LB/�1׍D�Z��ֲ�U�%G�Y�9�IS�WU�D?9(+�L���~��rA�A>O̜i�Y�g��D��ҍ�"�~Y�s ��b�l׻����/"L��-z��j7T��D�~���œ:�����l2�ZR��?�b�(�}��c�w�ǌ�?���Ɂ�-��Eb�ɷ/���<~j7>��p!�����t4��H��k�E
}�F����B�K5��p�����ʄ��u}�ۼM�5)���b�}�[7.v������^��I0��5T_5F,k	SC1i���$�����8&�a>�ޙ��"t������+�QIⲒwm~~>��nA�z��L�w�bo�ЯoU�7��Vה؏p��%�IN�E�)�����N����%p�}@���`�"�B�K�
蓦�Q��V�z���p�����"���=-��eP���kd�O&ɥU�\-��ڥZ���H��&��M��p֎N���~�$ϩ��1���G�~k[��	K}�����C�jmyw��
�ęqn*v�Q!4x[��y����[����XB����cA���E<c֦~B�.�r����¯C���*!ğ�T�xr�(A����c�t�-�M�E�֋��Ƕ]X ڲ��u�r�3����fuS%�IV���9��x3�Ho��=Bt�`�m�r^u[���t��N)�,��h�ӹ�L~z,�Zg&�	�.��x�t���U���f��"wuE3^�<*hB�F�.�>C�r.�|��Yn���Gf9갳�$-q�H�-��U��Bp�`?g�<�v#�--R ��0����Dl�n51u�k@$�^wKD&bd�|~��ݺ"��A���26���+	��������&�@�հ�������z���Y�l�MH�/��4�m�|��� ��6,���ʓ�7�8Ǡ�DU<l�+���юa��zF�O���.	-'+��X%`D�TD��)9N���6�F��xSH}��۞�>���L:M�9݂�py)깬I#E�x���x7;���Y�3>�|^����a3� �w����?d�*C��^���#��x�(�9
�(7�*}(����Ej�M�?>|o��Ļ���{E�2�|���V�7�����>(W�?��2.�'Z��t��)�)"ҽt�����%�ݵ��.Hw�R�q�������r�s�<g�3�̌N6�"$� �A2�cL9�c�|�^���������=�^�=x�$>������G�ƥ(��[��%Jh$�CLKL..FC啽���zD=r���v�̀�~*�q�sƈ0L����e0�еٴd�{C��d���R���Y�L�I���?ԩ+�ǯ��` %e����O��\��@�֍*%7\]�l-=��-�l.������ V`�J�;�q�v����v,���+4��Ca� &� 	w��J[v]$���Q�����U�w@U����a.=h�	g|	d J��<\����w�tO@��Z�-s.b.�����"E�3�'��g�+��	���jt��C"I5z���}�~Bak���]���T�x�OQ���������2T\���r´�s����t�8Q>�?�H�E�ר^�[mI�����>C��r$e��C">@��2��j2$�k�Kr	��������~��j���|WB)F��:�� ����� @�K�4� �A`�ϴW�b���*u���(�^��������2O�a���+ڬ��Da^O��\Z7��j� 5�ȸ!x4����o���V�7��ͫ^
3A)��DG��>S߭�C�L_�2�v߆x��۷7�(Y}u��ٌXwe�7n�zڞR����s9m$�ǈ��-"�O�D�b�"T��y�	Q�2#�X�Z �Ԟ}@]�08gjsD0��)�S6�,��x+��X�~�5K��*P��c	�/�|+���=B�M������#��*����ź��*�=�{�k��U���j�8��z J���+2��v;�����#�ø
n	b4	��eN?�U3$�Na�H�i���q�Ő�_7/�k�,�G��ǵ��"�*V�k��p���窆ՃH\��bCw�FO͊���i�R���En�	��K4I��h�o@��;�U�1����G�q��OH�t������1P1�
�Ǖ"Q���Uv���Iփ�C
��]Q��v3"�@���X�x�+����Z���n�� �.$����8 #��m�t��k3rq�"� grƹ�kcJ/�X�i��os	oG�Wj�-(:���̂��
�{<�\��,�e�����o�������%<�����A��'�����q��g�u��Sh��nuLk��G��X#���!k?�@[%̙��1����4�K�A�ן����B�� �'fec	!WE���H-�8	H0U²UI�uL�����/�$
4"6+M�a��0�'ądc�~�0hO� Fx��H53�G�G���Y ��R��u��r�̻e��h�x@�N�3��K�K��S+Ga)9,(<��ݟ��ANMt�H\]?�$����*����C�A���Uj���
��v\�5K7���6�2��Iy�.�+��!�Rnz?���"z,K��\�+�WbwJ$�#g'�����)��AV/b�� ���v���+�I��'̕s�g�3Dƶ�D%vM��MO��r�N�W�(�z%���\�I����F˘=�:T�aZ��}}~�θ�'���ݚ��KJ%e���}��I��}��a�a�=�"j���ɵ���oｩ��6�ҹ̗2�c蹓d�.eH��(���u��9g�g#|l�D~�gl�D ��8��;Vg>�h��4���"����E��zM��}[|�F�����*c��:8��5�0������?�R�{�&v�L��yU9��89hǝ�g?O�<7�SÃ&�!ق1t��	��x?,g����R�DT��1�+�}X�����nbJ|���7�?.��<��{�\U�r�������+�e����@����I�<v�x�/|1}0Ƿ 2�e����i��G�+lT�I$Z r47�����HEC�s��C�y�»"� *雈<�' IcW�'���ލ���9C����Їo���-��#�gk�S������Q�4&�>ϫbw��ƽ�:�
�V�
jZ�]���I��K���;xG��62y4���m�[���o[T4䥠�RF�$:�]L�1�w4l~�p�J1�*K���t�*����G1�/����P���V.Ed��T�J��!Ϧ��z�i��$E���$ߣWc�ԝ�eD�91��0^�b��u�{.6D'f,.>��
�2cLX~X�&���*��~,�d��Z!��Qű�D��l���(T�ߟ�[Wug��ԛ��"����*G����n�`�A��.�N�C\|l(&+���_Ŕ���q:����t���k��a=��u»��㜩���9@��I%��LH��D=���%���4��Ո2�o�6y.����� |9S���9��a�&��z�)��v5#�f�I^z? w�=�>�)ƹ����<?������R�F���I�:z{&y]�ƚ�(oު������A}�_���e�����F����ܯ�.���]}?�o� <~'	���E��x�bjq�H�Ϊ���}�`��&*-��+hI��]`�,�WKX�>���?�qB�\��v�=D9ﻼ@�����0���{	�Ǌ���$r�}�)�b!��8���8�~�O���9�o�-����q.^[�"�������o���U�e�bio	"����&����NP!�9����f��V`,3�Ou%{��� ����
*�(�=��8)I�=��Z�a>U�E	����i�ud�Dl��0�
"��pJ�#��Ļx�Z����;���[?�)`{� )�����	&�|*��2˦|�p3e=i�1��4ȘʼU�����	�
>UZ"s_v�g�y����i��k��>\v�c��ت��ݧ��R��#v��H;�G	��q �Bg�߸��U�=r'���$]��U�m*D���~7�\��oF-�����n7����z]���PP'Ñ�*ۊ>#��d�|`p��7!7(���/ݼ��x��-�>�۽(����˫����6cQ��$fV&�&bY8D��b��P��։����O	;�F�s�tF�.�*�'����U�u�.�I-g���B��.�3��������*5s&jD��JI/S�qC'���]��'uTD>8�T�Ay��k�9�=WՊ@֯B���V_�|���VFB;��=����\�l�Я�z�M�S���[���Џ#Y�2��-�Bs�ߏ%ֵ�F�wֳ�}�]sc�5k�*�x\/XDN����+���9<���W~�_q_;��3����UDYV����
5X..�Hd��F��H�R��3�>l9z�v�~���[�ao.B]:/�L~4�"�DPP�b[�VGs3w?���O7U���ȉ�ؔ{`b��������&h�1��I�DJ�v��99��ܓr���2��������=Nb���Gڙ�NϜ��i1w;9�ܷ�}ec��|C�d��mךf�_�e&���;%�y�\������SS.s�#g���Ό�,I�����=�t`��~��2ظ�~�]j�	}L�����ź�^��Fh����n��_xD���\֎.	��|�^uRN�<,-hc1��B�s�?(�^nuYZ��O�shՏ���<�,�K�)�����C��'	��&"8N��e��X��>�L��[��@��L����쩴��M:������$�Sp�LgU�I!�젅&~nմl���V�i�J��!J������g��R��=U�%��˹��{��O��R��zڮ�റ���~�"H9��/,�7��"pF�kr>T~qI�ehfTL��J6/���W8�2<�d(�9ţ�kV�CA��t��a�pc��_�2-���d�`tſ�d�-R�?����U���D�p�Ĩp���b�j�xU��Q���4/�ެ�G�.��9�9*��;�[�2ͪ_&��#���>�����$M8N��@�ꥱ�����\�t��_������ � q'�ۘT9����@܍����Ϛj�ښ��O�/}�ԐG��hpi�-�E)r�i�4';qT,����.����x2"V��ycV���Q����Q�mS��9<	@Zi�/ѕ�V���mo/��GK�
0WL��S�}g\3}�3)D���A��!f!o�qq�����P�
��c��~Y!4�.��b(QH1�+LB���$���'�� "��x��j�W߳s��zO��̌���o.���Jc'���5}����KϔD[�;�Y����\����|��)$kN���N�����Ї����C��v�ԗ���^W�V��pĞ1UwАa<V��Đ1��%Z����V	�����R��	头{y.� ߄�"����J���z�,�{{�UO��6yR��s�܎��TSrf�	��Q�t����B���п[���8���/����p��1<(�!I�G3��濠p�5W���ϰkb�=2��\�M��a-L�<CG]����(��?-�) +l���Yr'�+k�,�
?��I��_M�L)k��6>��<]$M*e�vX��Ͽ8��؀�F}):�6�3 ,�%G�Z���=0U��2��F	��4���AţS�S�����_v-b��tpVD��O�]w�,��7+sM�H���Z2='��3`*��m�h�kQ��%��6��}@��
/i�.�V@����Ѐk��7���`eW�� �S��=�}Ic�8�8o-_'>S��_��J^K(,*����oC���	����$�j����u�XvO/ uxxP���g�a�;�M��';�ܠP�Pe꠫e�Mb
_�rt��񳹷̽f��}t<o�ϥy�/u�U��z4���~>�lj=�ͨK����C�]\�����<��z�O�h-�4806I_�����}ʹ��*a�ztɩ�V�̦k�1�76�0<'���g�|�~��xJ�XA�y������.��ڞ�[��� �l]����MN�Ͱ�����Num�Xƹs��X��7k�>0z���W�rml�Sw_����5��^Y�c���Ԓ�(8� ,5|�b� B:�������>�B2*
�:��-]���'�LwZo����:+,��=�Ń��tL;WAL���M�g*���2�c0ϱ�����:e�E�>n/^�>&�%p��T�<��Y'!BM��UK��Fԭekۧ��~�{���,I�/@h�C[!-����O�fX̋wE��|�����t6���F_���c��X@�NU�-@�p@J	��$�v=<POV`�Ɩ�6k7@`�7 ""���s����~���6S�z�
o!�ɋ���L�19�T+�(�Ԕ���`����:(u\�zɘz��eg<�=�S��qJ�2��Yc�o#���Bkd�`��'vP�3'(x9���	
�Y�<�Q[ו�O�ā�ż���g�����`�R���4��������hX1���[�l�����.�`�Q8��֡���E�݁���P��Ub�g�<bw	���~�� �E�sA��g���*�=�$����s]������#�g=<���\0d)R]~�ZnJrH��f	h�nr����8��U����FH�B�󅆊p�	���J�s�0xo@������g��[+VR�|L���'����rg}�S�&�\�Rr-�Ug�T��k{EçZ^*bz{�>��xZ~�x��i�����k��>�`R���q3<ptP��ٯg��Xs�sP�d��K{*^�Rz�^u���
r��(Õ����呚�Go�'$��r�|�������p�d#G���5ù�^*�{,�Έ�o��Z�B���flHQ+wj/p�����70��Djf��8)E��qE���s��W��UMU�?x���B"�D��A��x��P��<���a����-���4�6���>'�s?�(����-u��di���/����`@��왷����s+�3|b��� �����d��a��{,~]�@g<�f.�H�b(���+v���
��?7L2wx�:�T��4���`��� h�è%�|��sE��Vޓ����������L:�N�Pl��5�����!|s��=֯���E#�a�IQ��]�f�Ԃ�mld|ʙ�����1X+�؁S�4�?���o���B�TX�޶�E�3�،�x�A���oh��_��=�?g#���!_,��L�E��:�s �
�'a�R#���3��8*���l���r��=س߉\�`K,KU��j�i� �Z
��]n���tGycRn�G`ڦ�W���$�S<D.���F��o�#����W6�p�=~�l;���B�����2�d_n�!!����b"(C^���\�]�l;7�CN�ZNk��\��Ww�@�Na���`,��ϖ՟��=�k��911�Պ�/ψah� P�K_�CM�&���7�%�wݲZE��p���]���Y���w�18���rw���KSۀS+�qY0���He��l�HB���x�}���qzgnU�򧞎�G���p��D�%���\.v ���,�u^��!�X�}V�D���ǮWc,�,�t�*D����O"��_���?��M ����8~�/����]5j)��m�*go���U�CW�a,moiU	�N��HoBx���P��?���ŃQ���zT��ɠG�����Ԕq�`n�����%a������#�N9b:���'�O)�_�f�sQa�g:hn�D�
h*ʍ�bq|��O�H�m��������t�ϩ��r}��{&6k�.,9���	�fF9��fhɌ�*��t=���
�n+�i_�������fy����/�E�*�KW�Qq�.{�J���"�7~Zۥ?�-���O����R1�w��+չX�EV%2��3s���E�Q��P���!��zq{i���_Q�s��{��O��j��.'�k@f����v�3��,�����]*$ED����Ԍ_�4��%׆�@D�"�K������=��6(2��ӍB�ka<�;喪�>�a��[��eZÆ�>�󹞓Qw���kf�鎵�&<��V�%����Y	�O�|�����w�)���g���#����"�~2�q�E�/�~�+��K��d�C��Se�#�Ћ�}yx��ng��Jɨ��J��HX����<b���4�O�ճ����0��}�]ny�ݬF�UՑ6}u���5�r6���_��_�jwqv�|��pj������'�X�
��EJ�ԈYJ��	���'8�l|C�[�:0`}}�@/����^;d�=O���,�u3���OqO���
�i3�;zÛ�:��\�o;�f��G��3���%]�2��P��=�����=��|�{n�i�!���HԈ#+�n�vA�bv���'�vp�����ys�����r$��Y����wWˡR��\G�hae�E�d�	�I'p��M�]��1��_�;�m�qE^��74�}O8���.ώGd�d��@;t�1��T5�k���t!"\m�WhO�>j&ĳ�;�\���l֤�T��[6��\f����a��z�C�,)VY����	|q����im��o��i����n���x����hK����J��8jf����y�U{Ã�E����<���#���	�eoT~Ԯ]gg������te0�iU` ��XK>K����p�s��+������5��(���lIfg=?��vkqw��7�����b�1V%���
?�m���u��D�x��q��'9�Wi�5��!�����W�KlTYSŴ$��0X�� ���"0�tߏi������5���14!_�-������A�^[11^�i�W$���x��%��ь�sj����k��� �M��GU�g���_T�5���ص����1Bfs?������"�=�n9{f�NX>�� ��n&��b��1��<0�/ȏ����వ�1|��\�t竡Ԩ����	өl]b�Y���2�p��Be�LYy�D�3j+����A��\<�2~�����mk�l+\l�[�Y�|G#��3��i�Z��� ��w�Ȧ�F�',(xa���~����_͉"{=��r�D��!性r�*B�}�\��,,����^=C��ڏ��	*�du��a��2���8oI#�f~�	��
��y+�$�\��hR�J�f�ϯ��a&[�u��l��%��JL���t7{h0<$�r�8.hV�U�Ɏ^�O0���;�&���#�(}ht겉b��U�&�����?�"�ۑ�Q�nm��O�	�<pU��t�A��ѭ�tv>����i�E����n��\�z����}��xG�b�����ӌ(=�^�Q<hU��MD\�cr���2a�)���QMD�;�
e�����e��K�o����1�H�(z�4�nYo����)>��-��d�Dك��r</4�����,�V6	ZS�꨹}��Nq{�_%t�ݬ��ͷf�܇fnJ��(����}�o���qL�\�g%�|��f�o�����Q(i���-�j�U�Qq{߆��Y�n03��P��ViɎ+*��pP��z�fL
k�W����%v����1���92�Y{��-�%����G��Y�H����0R-Gck뻩�T�4M见m�D����$�9��������`�S��Ђћ�%y��)�`Ȗ�\`�jJD�).r<������q�o��[�I�(�@��<����Z��(�,=ȕ��M�r�P����
V�X�}|o��m��C4����?�J��W�$o�d�]!v~�6^މ.]��Tt�������=��ܫ��[6E�cխ?��_r�g�D����0͊K���H��3m��͜7%i��ȕ�480��w^����Pdu�mƩ�(��	�Ud箸R�j��s�g��Y	���փ8F#��3�t���x��_0�CBӻ�%6@ �	�l��x��� �@^bM��̆����I���jd*<��>��d#���r��[�w�<��T1�j�Roߋ��G/�U�$t E�ط��(?��"sbߪ+�=����ӌ���k��;�r�ow&(������!�g8('#���bmE	{Z?���e���t��o�S3� ���H,CLp� W���˩�*9�O$����?�p�˟fx}`���,&W}o�h��*��W?t�
���hi�*���/��7#3Z�J�+��b�?8��G�h�v��k�[F�s��m=�o���b�һ�/���e���R�Lm���7d�hM�z������-�/�P��Ld�w}��S9ˀ����8��x\:ԹMU����Y�w������z~���򬕙?C��)٬��>�$3���N���#ژ��9�O����֫�A��Z.��"(IQ���6$g�f�7�o�ait2a��ǉ%꼞ٲ��M��u֋�w~:�Wi��UΤӞ^�ݮ�d�z��)�au�'VA3�4��
�m<`���Q��v��{�8F����V8��5�+'0]�7�a�}�B9�O�5&u<d3�5�̷{[�]a�;H]z��mԃ>�,3�~�q���#3ʬݖt�L���֦z�x�����?s?�0g��c9����s$��Q��+���7KC�� ?�_�Y�j"w	8Y�w�B�J:ٿ��V��r�c�0������ܪ����ڼ�FWщ�K;�R���1e���'�Q����˻�x
@h��5�,Y�`������BR���E1���4�S=3���� BC�#���C.k(Ξ���"Es�/ј�5��)Ή�/���W���,xK��_�g%'�]���l�$(�����/`�Ë��f�����D�A�h���Jd�E�6�\�τq%g�h,kz?ΞM';��ƾ������:_��9O��G�ٛ���co)��#7��fC�����,��J` ��JI"�_���O6ʔ���zО_�'�\b1i �o�����&h�ZWaM[��Qç}���Q�l��X��0�Q.u���0��aGT(�C�b��`��%Y���+kvDm^O�9�YD�:�ֆKe`6�a����ӐuB�Xʓ���Y���(}/�W�����e�&Y���X�>�SE)I&��Ɉ+���Q�L+��HN��ף�rY�(���`[1��&i)�V�5���'��h�^��(c(�������+����8(.0����K?��X�)n�!��*¸/��T�����K`l+O��H�|n*.�u�U9�O+0���PB�	��Я�Px�Q�@U_�	Zű���t�h>\��y�T��En</����"�2�?�[2��=�4�}믯�}�G^pD�ゴ��	���^H�ы%�h%���\�p�d4�Gq�����0s*x�eIc�p�*/���1��|~6����=�pԾcҳH�*d��f@��H���C8��s�CU���F|��,�+N'�?$�9��^b�xK;�H��1���	wǧ5������w]-JvX�Օ������Ww�xf��)�Q#��O�!����!�b �q�闙��"��9��l��̑ue]~����L	���ncc��A���I���N>	�yM��:����~����;<-��Yfᒐ ��ھA(.ĳ3��GS2,��s�{4��K�F<�ZB��������AqL����F��;~c�V�����(@����g���V�*w�ϫ����Ֆ�p�[����n�C�s*�Uc<�H�o�_��9���9�&�iC��O��g$�8��_��v@L�L"5x��� ?��5���W.��A���<O��;-5�}��D�U@��������<0���q�	�nJ�c�l��y �]v��_��Xˮ�<F��A�WLv^��2TtD�Q�_H��h�韫�q�����D�5j[@ܴ��Gt�Aq�
Ì���4.�<�ڨ�j]t��X08��~�t:>��{�I����ߨ�y`��u��n��9������mF��QH�R]0��N��T|�⿪SG�ۓ���jΒo+��#���َLM\,XR̦G���V�`�]�l������~���.��< :�}8;��MC�*�t����%_�����o���dM$���׿TBC$8�_H{�4�d����N��p�ucX��D�.P��$��8����<��]z�$h+dS��RJ�p%�.��/���=/��F��d4k��6p[%+�aC�q��o%ݷ����K�$x�i\̵$�%IF&�c�s����(�.#�+fp���	�ߢq��D_�i���Cyy���o��i:�$	�7�.��ݼZ��1 �˙���n���&�$'�C'Pr/ۍ
�2���iU�b���{J��
�%�|��y%l��j�/��pX��z�8b�<D�	�S�"{���x0��r	C�^��U���ܖ��I�^.�憤e4Vg���]�h�M�$RL���H"�sX۷�;>� �µ�})� ���Y�����m�'�"s�����T�N�D��k�P�罫"E*l��I1�R���N(hC�^�k�ɾ��S���7slB^��G��z3Q��iB#���a*51L���Q�cR��?�c�$I� Q��""���o�f&a�KQ$b�F�S�	�f��vƇ,s�K���wr���bgc&���[�-;��E�^�f������ލ�5F;̡7���Qx�³;��!u��?�ѣ�\�k��?Ɇi���s�����%ȳ���ܹ�Ey��߁H�a:��#�Ş���PI�f�r�Iy�'�|ad@܌D������ʳ#W�`W�l6��R��j�kӲ�v����D��tJݘr� $�m� �V�z �kp\��8� .�l�O�o���;4�"�-�U���E3��y��jeL���n}�΍ap^�}�Q� �T*S��v�`�<�#baZK�8?��w�y��j� �$�ڠX%,�L�[,_mMO0��p�[W$����x%��������Wd=@$�v{��0��խ�AX1��j�H7���. C���K*y�RyW�P1��e����� UGPqj2�C�' �=��aÚ֮1�h^�1�H�2z�߬���5��d^���2N����FX~2�&`Օ��c-��ʒ�O�AV�K����#�W��}%��ܓ����p[�D�s��Ա���AN2����׉���]J٢��V8��2�	'��G�w��ߋʹywV��+�l�B�~���m�Ň���}�p��p�bۢ�*ÿI|��qTr�R9I�1������(�ʢ�H�� '��L��{-��!F	��xxx�;�%���ϭ"�����,E C�wƋ�w!�.a�m�����M��p���Q�c��?��F�9Ă�5���	��*4��!����ˢ�C��~��IF65��Ѯ����R��F�zÚl�xE����+��O�xҭf�?�l�ߕf����� ���^ο��m6�3�]Y��Y0!&0p���
��m�	.Q�RW�O��o_�������Ɣ*V���\@���@�`�o���c�r�V,���HL���&�m�1�����,�|G6CF�h|7'�5J��~2�dN�	q�!���f!����|~��j��Q��.�[%�����˜����;j� 9ڪ^m �U�d:(s�0��'�A�o�N�?3�qjZ+��V,2Yػ�^�W5J�I%�����b8�=�R�X��A���sd�6)���cI�$��[
i�c�(�.�=-p�����\�gi����<�W��<�S���TN���|� ��<��M�]�m�~��s:�ֱ��ȘБMyf���x*R�(�Q�Y����K{N+>AY-^8*`�+�8�HC�&۾�7u:�ERK�*��>�t�XS`K'M"��V�8�5�U�"�A�c"=�Ѡ�4�I�k�c�Vsi��NZ��y��R�ᇛ��B)l?��ę����r��}�T��c���g��IT��q�FRR����8��?���n�y֓���)��v*"ֱ�]!O�����T�c�j�މ��&�xԉ�>�]��>9���bC<�� ��H��~ȇ���(�_�~�F���,��ԩis� �,|�Ł"��8�۫��Y�!?Xq��dY9�{K��7U�Ʀ�s��w]��P'���C��?����"\к.LA����d�>��ڲ�eI+�>"C)�'���욬@��l:Fu�ph�\�oT�C�ǘ�F����%��ԡ���MX�=��L�n�d���m~&f�t��L�8�-'�C��I)��|��KB/���Ҷ1���)C�f�)Ig�Ka�����H�e���VF�R����^k�mG�.��WF{��q#��F0�x(9���9վ㩻�����<�aR(s՝�����G��8Bd͜��z��j*۲~EV�����+/~�a9�^X���jr�BI<�$��^�&"�P%���g�v���f�E�J�Q�5��!�&{#l�,J�]w���{���b���������I���LQ~7�R��������A��8�cvcֻ�it�5�r aDՁx���l�>+X�Y�d՘�Ϫ����fp�	���Z-z/�� 	�7���{�AJ��]r��h�<?s�9[/ӧ-�rᏉ����P�A��� 
.�PK�k��-"pWj4�rm�qz
�|���L*_�N؛��YA��K��F6k:�:N˃Q!�_v"��lx�(��O��F%��Z3}�~=1Z�H�#����b��6��n�	�X]�-�n����d�i�P1[�qv�����n����ͬ���w��k<�8�n-�@��g�Hē��٫N ����w\���r.>�K�	o4nsA W��$$��ye��NtUS���ؿ�߱��������d�^�I��a��!z:"M 	(4틬ͻ�Y��@���|W�;T�4��jV�^J�pcd���%�H伤�z�Հ�@�g|�(�Գ��z5�ɦh����y�����GLIiNI�Y3�j�1��{S%h�3��ޛy4��U`�N�U�C��B+k��c��	��p�qP���_���h����=���>�]�$^x�o�ɒ�Gn�dk0 m��a�yд��$2\�U�����;0�p����/��`4��Mz4������.V�� ��f���	α����i���C�G��ǹ��5p:]`;:�#��aw�����/S�r7�h1����}o�%����v1�a�~�-���K��G^�޲J�=��ެ^���Č��i�Jy�	�#).J����|UD|d.����]j�Rl2�FŊ�4��- �}pM7���~��xu�h5�D��#���ۮ}���s?���W��j����A��^bN�X��b�����S�H��2Ѳ����`W7
 ��r��w!�6���o����� #���x^�n^�}9��!#RzD�fڕ�b��xB���J-R�)ي%Q��2$~Q��]�A�37?�A�ل@�3s�3�Qu��5����
0=wy�j�'(�&H\�'rwH{mE2~.�֎���!q��+Pܫ�wq���b?�:G-�^�d�����|ڂѓ{��a�W�h'�U��$������ue`���k;���L�-f�e��'Cc�B������G#Q	X�>����~�Z����b�нiDd�}���*߯H���;BB�� o�;B=�IBs��%��+k��Z���w���>�\ʑ��M�&�b��:M���}��h-B�,h�Լ����-k+O㢷�O5;j1��#���tJY�d~���,Y�,�c��A��Ha ������>2��pa�ȬԾ��C�&5�}��ZF�UG���-�7���ju��<*�^�v��u��7�Zm�r&H=�Pb�=K�X�I܊Ն�z�@������ջ��� r��-\���@��]��
\��3$���dl����j,Y�o�P�_�%JaX�l~�����-:B���O"Ξ<=Oj��;Տz$��� ��V	�I6��TS�݌)���K�G�%_K^I�!�������y<�1�p��-�$��Ά�Tw�Zx�����#0b*Ce!�0AX�0g�j"i�!�W]m�h��O�C/�����LUWe�`��&P��$l9�!�ٞ����f��+�G�P���ٞ%�K�&�:2����ئ�O"O�����}�8��>lҥQ���G('{isLi���/A
ƾ�Jy�ϧ������m)�8j��W�ڻں)��\L���߅P�-�h��\x��f�f��eZ 2��Ki��,�]����&]3���?4�D?�6���[���%�Z4�-"�ʾ�[�*f�k �RY�{�����i�5��:ہ��'D�䅲3Bf���,�.��aўs�G��YU[��� ^|gO�p�re��yl��"P���
��Ȧ�px���~G�1w�4N��BW1!���^tZ�����7%���D>Q�����逘���5B��U/�E��¿�۶m�4f����!_��@�<�ؘ�b6^��wd��ב��|�@m�c���~�œq� �﹎�糠����*���P��xeCx|s+��ڄƽZ����LYDD�~���*��߃�����'T�g�݂��K$ �ebk�7r��#a��s������_)���C�ԋ�jH������/���Ь"�DG����1}l�~=	�'tY�sj5ҟ�q���6-1�B�sF�<��њ1�b.M�!T��2cm(Mu(�E�8�����hD$��S�ٺ���B�2:��-�t�2V���J�p���Em�Gݟ�ך�7�w/��s��1���o6*�~9�ѡ��S=|��{�6Q�!%D(��v��a�3œ�-���}z?��J�����%�h1.P���q�C��Ԃ#ٲQ���d��eH)YZ�|PL�D��oV� ����Z��Yp|9��_u��.��'c���Оغ��Y�������kyS�E��k�V���A����T?U��ԟ��On�J*1�)�
~?T��$~O�	��Y�tY���,��VG�.��d�����~��/�[L�+�_���9��ɼ��m��Jɽ���αܐ��$�L��`of�5�k7őA��p��H#r�f�1�����s�v�<jj�M���4^t}�y2'��^�
$�uw�7<Đ�պ���:'~���X���*t����iғ%d�r�,�(�c{!��������x^��.=��)�o �M ��V��	$����-��%ů�	R�U���l7!m,���1�%{�29�n��� 
1��n.��Px��P�%�W���k�L�NS�l��ZJ�;U�b}�]V�ׅ�Ѱw88�6R����}n����N������DN���B1Y4s���+<eT�VuTngS!��8��S���+���n�4�����ƈ��\���l-�����A�g�	6�9{浄�D{Z�����EH��K�J��A�ޕ[�>�p;<��w["���J)$7O-'��~2#W���\1���g卓ړ���h�[���-�;�l�aM����!m�:�^�A,�����Jp � H@��n�B�uX�D�z�5_�у�0�S`$sy�:;���b,v&�@>*�Xw`�#�a���)���ղ���U���ŋ�h�\h��F��`9-Z�Ⱥ�R�̂E+i��Vv�1SE*�(roP�w��bA�s1����3���g���dĔ/z����=�����l�N�~�KO��xF��;@�q�ӯ�F�6r�`��23[�GV�r��9�3���f;=��,߬N��m8˿��E�(�45��BO沾��e�JZ\*_f-o�Vv��,Y�L�l�C�E1]od�M�Ȯ�̂���@�0�{q4.���|Tx�4f��m�]蹗��������������#*ꤣw*P8�Ut4{hLc�n8�Rk���ޚ���gblx�8L�VTQ�9�=�o7��L�z@dpΫ�4P�0ҹ<�)�BtH�BD�L���f6�o�z��s&E�����q.m<�d�<��eG��	�-�l�;����	��l�# C��w]���B��9�=o-\��&��!�8qN��4;�y�B��N�m��0=r8;I3�IiT�,q�@F��u��H#��r,[)aT�UȎ���t�5��|)%c��#�p�ۯ���2:5���Z���)E�!*�0�[g�\g�EW���v-� �<�ˣ��м�W�듦�ĩEm��R�U�9��m$��������MYE��pL�5�����z!�{�u��t��k�.�-eZٹIY�eLZ�4�/�s�K�R(:��ZO�\~&��`km�L������f9EeT�X��LZL�
�0NC���,;C."�h͜����ʛSi�%Ʌ�&�e:�I	��}���4j� �t���\�\���k��	�w�������g1����a�1���rG����UE��Ƿ�ׁ�*zT���vt�9R\)�v��@Xl�Dj�xW���I�O��0{�J}��o���s��ہ��Ut�-�9t�����ΧDzf�R���$��(�,.h�"P�m�s�d9)�8sԪ�ә���Z�RE�r�u������P�e[�rrl�  �y^�{�ǰ��h��<�\z�RX�[����YD���ף�b%a8�؝h����6�L86~1�w-㘲	-&&Jcz~⌳�� V�aR&j���Gut�u�М����G�) ���{�r�<e�Vj��)밑�F<d��K��U�|�L�l�Þ�B�FWu���[DL�C���m>e�-h}�,�5T�}���i�1#h��F������n���z���8�1aƦ��Q:�P�Yt	���]���֭�**uQt8H#6H���t�7��!.�=��f4��l�2$DE�/�,!���@ey�4��U�+�e�������� ��k"	mI��=s_�r�Mi���Dy��m�0~l���k���C>�h)���{|_6?Q��˖���)����.ޗ�3����Υ���E��GM˰�X,��~�J��M�������ت9w�������w����Q�����b��P�#n��{�n�^v�[N�·��9.`�Iϣ�hU��%R\87�KiUk�.��=*5{�w\s:���;
���06�41l��D���`N}OtC�c����轅����h��{��!CGw�~~ٗh��ǐ׺�l�=�t*򝙼fs����k#��ƆEa����^~)9vH�`0}�����<�Z���o/�:+G���-v*b��91� ;�X�h�cC]C�3;�A�f���&}0s1��gh��֒��$��d0]p�i�-,*zp�1�~�̀�8C��e��N��J�Z!Q�G���-�-t����Z���&���?~w!�8z0�q2�d�ݙTZt7���덞"nW�dJ?������g7�.�<[����&t���6N�_ v8�qo&;��O��r���K�#q�s)��pyL_��n�?��������ѐ�)2uΔ1|@w؁���pH��St���j+����o�_x�����qޭ��J�F;*�����_�y�n�ڇ�6�r�5Z�	������E���I/������T1� s����Ш�3��_v��]� �f��Tt�E��YZؘ�?�3��N_Ы���_qm=j��&vvء�7h�@�+v�b?	^�v�"}i��&v�1���~�f%c����ΣA�,t_eǶX�p�+��E%-KUTj}�\���,������`�K���=,��������x՗i�����7��G��&p����4�#؛�|`�J�.��v�/���_~})5��V��G�*�+�<�p�!g�di�DaH;�vְ֢���l������w+M�3��y��4�Τ.7t��Q&���{�B���C`P�r^��1�y@�bӡ��
�]�s�/=�o�q(���l����6�N&Y&���9���(EgAcG�+lW�Q0���o��K�GxWKr�b]$�����9O־{�4��!��̌���O�<�h��}����Fa�9�4�@�m�@�?^J�����*zM��8�~�a"
m�[T,!�=�Xb�6L1���W�ZB)g8iz��<���l�����H������+�Т�Ki�]wA�,����0����;b,_���	���)6���H�]��ؓ�xn�2����Ɵ�E�ޜ�:��'��Aƌ�p��X=�0v�fg#`=�7�cOO�_��	��ޗ8\�q�H�6ۄo��%C����}t=����$�a�T�xp'���;mI/����2�P�T��z�Y4x@J8�,i�G#Z�E����d��b��}���Z��q��t�?^Nxo���@�{~2m��@�x����,����Mg3�����"�u��2N��y ����P}}D[�E��5�O��V@EϞ;���O8�����䋼9�YG�<�*㑹):M�Ɍ�b/�������K�<͛�${�rĻN�qS�c?���:+<3�m�������b�LStLW�E>e�����3;�Cj~��1��@��+��#�3o8����b!�&�e��aҲ�t�ew�kSf�������~j<��4`�`jm]Ei�9�n�!6�"v�,]�5#���Ɣ�!�?o1f8�2A�3��z8��}i��G�ج@ib�/�� 7*�S�9��i��<
X;L{ -X�J�^~����>�\{�E�����������(6����u�<$,��| F�e�40��:���	���yG�[a��ْG�Q��W!Z�0FL����-�̱�&����.��4s�*�۷%��wfӿ�;�?pwr��l�9�B�l�#1*�}�lQ�b�2x\+
hĈaԚ+����@r�n������=�wa�,S,G�RHC�=Χc.���/�B�L;f?�9e���e�c\�$^�b�b�@Ť�k��e���?x6"g��X2\�IS�9G�f�.Q��Q��'�L����ל'j7����~���I��a����G7A�%��8�خ�&����g��?�C�*��9����M/��lA���ˎK��H��1}?J�����_��&�����HUL+:d��):��Ȍ|����{.�[�i*�+Iˤ�xVC��(�(�F�e��S��7v����8B���ͫ��f�%�1)�-��	]Gk�t�ee\��dk>�x�>������w���[�C�eG��|ˊ���3�B &����X��}i:}����X�В��]\��Y�(�θ�d�ev�M���A>5R$�Q.U��6 �-Щ_�G����;��9��Y�'s���= �}��H35��)���Y!���g_��<���r�C�ި��!�8uΊ���u�L�Fn*`w�s�ؙ)9.��ak�j�N!�uV�3֐6�h ���ӝ�f��\D�g�S|��1i��cH'�a'C�zu�4��w�Z[y��&N�M-M���v[Q�i��ʻE��4���^���@2u�}w����-�g����'TuŚAg'��Т��E��r֋z��:j��8�8�B��<96@�b`ѓ/�M��i�D3����h��,��x0i�AQ�9��{�`m�z~3;�E:��}�'�''R(ځ���+�$+�Q�j���c�>v����w�t��#a�D�2w�}��ߞx�e��rb����G�7HÇ����Ʀf.[�b��ޥ�@��s�G�O�E�?pWz��I"_Pt��o�s$m��P�C�<�"CGWtγ cl��+>�Qi�iXnc/L����S���c7sR"J�
���(�{`o���6�}����M72cG��B�m�(:I���Q���kh�I���tӍhΜE�`Ys�@EW9��=h�v��9�ie(Լ��"J�#qi��a�y]_y{:�����CgƼ崪��v�=;L-�E.:��Mg��f��_d�,_)�X�"����mz��wJgR(��~�(�f��"�3�D:+��锸h�֧(�z���;�� ��n��<������<�����Q*eЖ�7�g��(�*��`���b.eL?��4���M��k�Ԭ5�O��I���`�Ie2�c�.;�p����KL;��H�-9��ޗ�7�RX�^{k&��lc��1�	�Ե =�5�B�lv���#/d;�)��͘.gޟ��tEW�{���c���gyA%;������+��(���*~ؐD���S����|����sw���M�d�bCP]ӻe�;i�¥��f���9�fcK�e�Ub=M��(��Y�C�Q$/�Ȉm����JG)�
���#	2C�D�W�`��bm�
|���`�x�ٲ�rϿ9����sdg��)�`Z�(��a�ǠPϐ�5���ToL#G�aU�[�'����.���{��[YƲ�Jk,S��C�yj1�~臢r��ޠ���56�+�gp��<2�^zu"577�����-��K:j�x���8�00>�k�=v޼t�b5C��i���YsL3K��@���+�b�d*1� �&��syz�����ޯx'�o���ֻb�G�O��P&�l�r��L����g���d��{�!��&�'���D/��Q�X���DZ@!/A��6�)�<Z���y��E�W5�o�7L�^��Z�����{����'��vdl�E]s؀/ո�%�FL	lW��9��.�:'%��0J���b������o��� $��?�m4]
��或qҲ�92��֬mQ!�чs�@%h��Q��̜���5��c6�ZA����W -m	cJBJǎO�9��s�a��C�{;9�B�s���F�F����Gb.}4�{�)� ���)�S4���{�2�_���om��(�tp��-�\�Xw-�ذu����2L��4eR}�����g�$'Q�<(_�r����d:���&=�)d'��¨@^�S�j �,Г/Ϥ��;����kg�.;lIC�fXU�d7��<u.W�"نN���A�uj�=�nCϼ�~rE��M��?\�i��2�n�i~�FP���o�T�ä�}���N"���hw#'%��@5ۉz1��I����G���y�#���?��.0�֛/�4g|`�.�-���+v��FK"��Ȯ��{������^��Ea��H��#G���d�&o`'�I�:6п.M�F�L�4Z\�����7>ȿ�?N�����34m�v��b|}}��bAt���i¸ET�����m���h���qW(X[L�;�aa&�6�^bu���ԐBDl���ј9k9��ǅ������描д��d;u<v,2d8Y�ِ�K}�1ϸia�6���X+`�m6�tڡ������3��4,L�D�fyʘ��4�����ϲ~�NЏ�6����b�s���"�(K�)��b�?г$
<�N4��g�P p�~�et� =�ȶ2b���h�T��%#�:˺��Cn1�Z��7f�·�Ƌ��#��̹��/�[��'��4'�-�2Ѝ��U\�y��K[�B��Ci�bC�D�p�\��dia0�乁�2��9r�:\?L�q��]�{*~�kG�x��7RS��g�`Zl:�.S��Qar�x����o}QU�(�����ɶv$8���"ݦ���zcPʱ����)���������k�N-���(v�c�r�=š/ʶ8֨>3���|t56��Ƌ�+j�?����.�[��3�G�A�7��y�I��S�7]u�?��[�ϗ��.�쬨��/��1�?�a��o�(��c�
�?=��J��
��ȃ��1���)�,����ٴ�����QO�MKѹ�L�lh1�lXX�L��o�^�Cf'G*:����'R�귮��^��XdŘ'38�hyK�(Ӿ��a�y��z���ň��������M��ݱ!�ٴ-�pHm�d�ܥB�@~�ӋoL��zfK��ӿ�n�`6�"N�V?鵂
�'�:��16Gc�|)��e�����Z�B�j��`��$zA�6�t�������
}�I�ׇ_��@kwL)��@7E[8T;�a�ΰ��L&Rc�4j�:�-��b2����pvBo�N�S�yk]�5��|����	�˳����Yyt�3��i��Ȫ�䴀�S�.ՐS�.�o�@�r8��.Y���qb�΃�@�@]%&������6a�}�(��h�7~r�,�o�!��HEgQ�x���S4u���K�!?�.YC'�r̸������=J��W�F�fi�b}�晟#=v)�M��%2*zq���(��y�[�{�t�K��EV�^BϽ�6���~b:�ePT�������#���g?8M8�ZE�?������,;�I��q,--M�?!e�u��B�\LϾ2�*��K��s�����(��ʪ�l9N2����i�V��>��KE-���?8�b��`��L8��TZ4D�%<��:��I���)�飏��s��?��^��"v�1?�9!��P1v�9LK�BS��8/��׎�4S���Ґ1�7W~�S�'/�r^l�� �T�0
(�j(��,Q\ L'��|}U�R�3v���%oE}Ȼ���]Ay�=�5��亇no
��,�."��"[��.[�]�7�X3�3`;��Ͽ:O�J�	�i�ݷ�e��!�a�^�b*�y�u�,�b'<"�a OU�S!��]ϑ�� /�ŋ�1}p��ec��0C)+�,Z5	�"n2�f�)�u���R%+�~�";�1MQ.�Q��誛���V��\y�?��4�[�U��[�S��-�
GåA���A)�f���e�m�����|s9��\V�S
�O�wq�F��鉪��0u���2$C��"y��	[淮�͒�֓��1v3�E���=���ʟ��6�Y�8����l1�*p�)Nz�)�F�z�l[��䤴ª��+���kv��]B9�=GK�;<��c\�,c�;����Z�$R�x��8�-�C��;�Di.Я��	��Tt�f��S]&�BK@N�XG�.�iK�n��ӈ�02h�si����_Vh����j�L�V�'�m"�ڄ�]�X��|�ޥ_*j���ޒ��NZ��Y'�v���x�:}�����wX_�V�Xx}�,
�,9�b��e����Cn;�Cv�]:x��K�T�(�t�~�X:�[�����)��D	�2)���,=��GU�-��_D�O�G��)?]ጛ�A;��!*'��"�D�xt�Wt�_^v2�Q#����655�by��Dtz?E�� v ��wE_��p��Bs`�E{���ٷ��*@[7��eJӓ/~�Ȓe+&��*�
.��� ¢��Q�3`����	(�b�f������*}�Z��y�I\h�P}�jjA��H���S
����豧�#�NUr�=O�Ӷ���ٱJz��+N��kN=�>�=h;�N�_*j]3��S�B���Ɖ����%��S��Z�XWL����z��������B��]~v����G1�3����e��<���ШA�Cu���TW� ���U��ф��Æ�e����z.�a��"�ѧ^e=	(���Nf�0ty�|1E\	˰y�C߼���U�t��'H[�ٔ�&��#x�N��y!'��8KŢON�J�^$����Ql;�ٳ�������p�U�v�|�Y0w�ۗ���S���eEF����&Mus�2;����4|6��ˤc�؏�1�HT|L!3fS�b-�FR39��Q�D��ޥs��S:k�b�����/�t!|��T�1O&���
��2�u.9>��Jv�Ҵ� ��KE���cJg-J�DE�'���7Ywع�#WT\i��OH�ߛK.��JKΥwߟAk���%�u�"��D���n�ȏ,��9�Ը�Zc�!)2�f��u�M!����>�G0?� �<;��'L���k׏��1�Y���H#������)��<�R��C#4h����Cŧ8`�h��g�'#^E�Q=&�x{�,qJtS'��4ݣ�W���8�F��s��k:�D�"�I��sY>]�I��w�����'�yQs�w#J�{��7�xf�#3d��Ǳ_�)�I���`#F�5н_L�����b�ۤK��"m?f0g.��mPǶQ�_"{i -�g��y�\�ڪ<�3���D�ż�\�I��!GE1�� UL�ا����a � 1P|0R��C���":��j�W�DϽ�i0qʇb�k2�7J������ȡW;^[�A�����s�mX����1��Q>'eND:ˉf����N~T�Lyo��zJ����(�8dW< J�M�;h7< ]��B�"D�n>��y��"� Ei1ݨ�kz(z>��Չ�"�G��P��'KO��(�Fv髯�;����Fэ()����ϗ�3k~�0�
6g�n䑙aC��bt��i*u�ӄ��Z��)�N�O�u"˥�m�����~��B:�HGi`�,��_����Vb�2m�XU`'�f�Ӡ`�8j���;]�M1;\���^��E�q�{�+��%gوʋ�
��A
Q�|j�$*x1=��V7O��>��I�*��©��\B�!Сc>�Gi���y�n��>h�3&놔Y�� +[\z�E�s5s�#��@End�e�Xȶ�aO�|�	�/�i�gܹ�+�6���;�,�H"[�KX���zX6��/�i:����3s9�u��eނƗo��'��Yɯ݉r�{�ez��|�y�0�S���{e�G�eD�k��<"��@����B���)��5�(ǩ���9O��xn�̘���;�������6����8F�x���B�%i��S*���w�a�!x��7�rN.Z�В�<(���ĩ3Xz�9|�B�#��OZ>�	�m�f��S�o�`:m2| �uC�%b����ʊ���ή��%���p�|�/�*�+��v~�`�v	�bR�1r�N\F+�� %n��<v[��q[g�Hl�)���7zF�C�׭�f6�|4��
���f������e�T>\��� ʒ�=��Z�j³���b!�Z9�8�ـ�0rEW@���e��]$Sj��\4��������&{�C�d(B��58� F4����[�<�;�N�{E��Yj0f*q00Z��ȣ�Tt�Z�!��
[�0X0�{�L$�/X�A��"5�ձ��4}΢�����y"�@�+����k8��i!�4T�#�fؑLz�ű�& kT����CSޯ�F6���^�z����F�k�X��d &��q�Ѡꦬ�T��n��؎���5��
T?���W~aW�X�0��e�����2ؖ�]jjY:��Ƨ�������蒾,����Q�x�>43o����.k���hjV�hYQt�p�0~�s�gDa����L�qD��,��$E��ug쪀k�bL=b�t�H �t�aH�����q,^�8�l'M��T�p�A�
3LI�4��46�xߐA���D��'�;$#�L����c^ә:jmm�l��^����M��<�շ>"�qD^��CV��;�|����E֗�ا�~�n�w�	9�~@6PA��匈�����h��o���F� �r^���M��c�q8m8O����u��$,��O?��=�b�A�M=�yJDE����(�Fly,�\��T�u������xiӔ���i>
�����!�#޻4����}�A��,%?l�+���4
y��{�OE�3��mv��u���X�)���}v�ߵ���e��z6|6�V�0��H`0�\�1yviK��)vV�j�S2q!�b�e;z�2��"8������~��v6�h��Ft�H��Kc�\gg�B���0������ȗ~U�,Z�B�BA|.w�d>��O��aL��F�6E�3f�p�'�a
p�Q}���)��І��V�����xs
*��oؔʤ�.�-.g��|[�ܱ0���Z��B��/|vg:�]��b2l�Z�f�����H�XW�l�J�m�i]E��\c+�gƳ�����ǋ�������A�#��,�����ʄ7L'lT��.c��h��dw�4i�e����Gi��.g�*�髧H��UM��2x �\���d���j0ʇ�g�h�膎9��#�$( �F^D��V�����x���C|a!���w �2�#v�cӢ�K��K�.�)����8>�;��Ð��Z`�ȡ�-��pO��	�
�eƥ9s$�k�|�Y�-�_$;��N�Yw��v�9]�ko���/j�f�9�����������"?l,	�K��)�D�6z>��.SO��`ի����������NE����%ђ�w��k���[�01`�D��"Mq��!V�A��%��a$���$�ۢ^�^�bˤPT����<]|�Q���!5�o5r0ivș �Ӆ+��N�f�4mn���KW��8q�#3Nq:D�!���	�5,�7���Q��jg�k���D�"Y�T�~����fX�<�b�f/hI~PC�����l=a�YL�d�aܡ<C8���)t5�q����v�1:y�Kċ��aǢTbӠo6��-\U{�͇���u����;G~n ;��N;�z�і#��~Q[�&�z�`���/P���B�TbF���)r8Oɲ�� �,_z-���a8MN�X�sZ�� ��5���=O����fYUw�0��j��<���83ּ KgS�z"�����������u�n��ʴ�ɲb��7N)�ܔ�!�]��N��� *4 ֨�onɉ﵄��m����u6����
R_�HF��3Q�q�УB���o���)�^dz }�.��4��ꧾ.�����u�ŉm�b�9⭭9�/@�� k�|��$>V{1H &?�.>�|��e�g�4�ö[&�e�t]ڬ��{aK�[�Z"���,[T�"�対�������A,3u���Yr,[���ȬE�]%e9�	Oَ誎B��Zx{@�]{nMf3�F��爐��+�V�\����X��\^��4��4��'T��5#c\A�,Hy���j/�����"��l����IÌ1�9j�x�������zH�#�I���+_Pq%^8Q�������eN��k�k:'��>����d�:z��C�S�E�O�1%ܲ���`����z�w�;�JE��>��{�0��xq춴4���Fj���|?�t�I�VtB
Ծ�� ׏�)�i@Ʀ��~�5��+��c�l������p40��p=O��J2�4D�Q��LbB�HG���X˖�Z"
�8�NP�Nb\=�/٬�AR+H]H�M�.U���c)����%���y	Ht'�L���PH�M?9�FOQX��r:$� =�nX�J;������z�ߞ�7��K"��G9�}K+�0������k�u4'��u6�rE��4�R*K�*:�ibz]�+��؁��O[�"�6a�Ͽw�(j����4�ړ����#+ց^V�6��E]I���g�(kۯ�>��-?�	U�|������^<�/�sm�q=^��laHf\{5�N�P��ǎ��7���Y�I��M�NEo��g���+�{���b�jF��Y�D�DZ�x�*����@���F��T9�z��J��햃��Y3
��q���2+@�<��-�'��h��/%� �Kт՞Y��x��N��	 ?�FUc M�k��.�Xjq�K-�^U�c���H���϶]{�Oey��Od� �ì���x�o�}��p����:
���(����'���|+�R�����7i��'y��d���P�x߃�Ss�y��ǃ8�v��R����gR*#�2�j(dC1�ȱu*�����Ԕo&3͎h�������نN9z�ҏ����V.�a(!�N�`#)N>G����84]h˝,PnHJ��m*E�������=)2���f��1L~�����!I�0]���6��N$"�G���1򡡢7��x�8N���C�XCti�s�i�2�ځ(�~��t�>;Q1(��D:[�	�,��R:R�sr�9�|�?�e6/ʰ�e�#^�y��_��O�JO+��i�h��C�w�0J��9�I!HW���NT��?&�Rz��V���Ӂ{oQ�e���1ǆPҒ'Z�8+�Kߥ!�tB��Z�4厸4�������Jcs�߹|��~�3�+�ˇ�Ԟ#�gƼ�x~� �+Х0��Q9�5Ck.��<T��I����mȈ�m��$�/l�`��T�3��Ƕ�����8i 7�X.�11h�!_/��₝����5�����ڛ&�P�x��2ki�ѻ|y�cfeB=�#6�D�M��J?�.Gi�A���Z'F���υ[$�:���1�Nf�9���i�O�;�X�j���;g�
�4�l~� r�\�h�C�Y�E�Q��;j�!�X���D+��KLy�ڌ(��FӬ��J�PT;�/�6&yo���i��x��l,�-��^��5�0#�9�y�VyaqO��0Q��r�;c��wR+L_\d-�)D+8��d'+OzO��x����,t���e��6�^����Ov�<�"���N��� �,���3g�VW/[n6�.��!�&v��l�����\���(k]B����z�7"�lm�m�]�����ၩ��Y���q�k���r�+�E���yf�»�8j�� Na|���34I$ktd�1`��Xlk�Qt�ʻ^����O������7m�-ofg�3i=�w���C�R�4����gϲޱ�&-�a)� �&��xۜy�K�PT;��3$yB�l.Zl4C=B�'�;�6[n.��#7ۘ��4;XIF���%�p̡?����Ϭ9�E���MT����#���ź4z�&|tm0Æ!/`�ӄ���k-FZy��$�G�})��ՋN7��D1,P���y�
^۔M�)d������RnIM}�������ʋ�0�������H���l������cR]s����C�i�^׮�Ƌ\Nw�:;�1�Z@}z���Vm]��U#�N�Ci�SJ#I^�5zӁ�s-���j���|J���GA����>���a�Ѭ�K�)��y؉�Q	�	��[i�1�8����P���R;�|���z.�8ʜ�DO�n����.R�x�0�����5���=�do>Ȅ�y*�����a�&�Jg8���CLJQ�^�6��!�I�O"F��U�9�=����s��Ŕ�U ǞJ�MT�T̻Tg����Q!������y���J�*��W��b��U7��hX�	���+�F�	K������=�͊��m�s,̋��)�����_�Y����HI��O:Im|bT���}wߦ*�`Ml��P2u�yeW��\��sX�!�B��1`#��[,�,_�B�eS%N���	�,I+�@#?vy:h��J��n�L�ǖI^d˧,���@gR�C�W�1�²M�N@W������DL! }�Sm;f��^���"[��y�P0
��Ӌ���-�V5W_8������Xij�=rk�Ҳ��<EA�RY�u�b��(ې���_��7� *��Wș�7c���,9ҭ\��E�$�Q�a�'im���p��gL���BާL&K��S�ʥdi>����NQ
,O�"g vP�@А/�͘Mź����5vS�l�!E��i�i�k,�F0,��'�,-^��ZaE���A��?�D�˲�^4��v��y�����4��"߀��|�;8`h��c�V4������-d�ia�`�l	��H���r^[�}vے�%��f��c6F)'CͭMT�͒$�Z`�G�9�4�8O	B�
ޚ�� o�禯� ���"�Q�إ���´9�M�
�b�e�|8s���X�*�^��j��c�#^��ya�7���Vʌ�Ri5Y�B
���I~��<�fS�'���r��b6 B6t(9�E���7]�fx5���wf�c����A��"�(YG;l5��H|�n��w�v�DB�+����%Ƌ�W
�%�壩U���J�pq����BA`\'zG �#6%Ψe��P-��q��c���(���H��:�X|<9q)j��VO8�1睉(�.W��|�����[n"*u�$�;�!�����t�k������YwB�'S�ή�$�)qߍgQ�t�]��D���ʹ��9��9��ȋ�\�0'^~��1.|/�1Y}��ܸ�e�{o|���=�Z\������:�d�n��eR���G>��O���je
.�}�օt�/�;�'��$"A���8��s6�ӡ�n-��f���֛�q�g�s�%�S�%5�g�^�NUJ����~��I��ís�Z�4h�J��(f�a�:�=6,M[mV��m�5�5Xmy�h�.���i�+fG����.�JQ@_^}��G�E��C&�~�L����Y���{mCi��Y1s�A���#�����qC�<���RJ�`3����ɰҔ�0M�E��<Kg��WW�F%�S�߁OZx~lϿ��[��%�k�kEr���Q�x�|x����'^~m�Ė��U��ǲ��0zT��.�N�p�,5�\(rـP�	E���^SH������U�O���L��D+�t��Y~�
-�׮�������:�Pr.�Ƈ��i��y�!i�%Zƣ��7��;E�0a�4�XWX-��S�%b#:q85<	���5��<x/���V:�=�-���D�ȏ����6dߞ��jq-��S/NNfrY�y�t��L�gȇ����=�0�S����^��﵈a-���e���g�����"2m�>�U=�@��l~�:���F:��!9N@Ma#9l�ǉ+#֍�_�2i�
��
S�C����}_������;К,b�)�ȱ2�V��浢K���,�<�B��`TFl^�!�@Y2R6�~HC�0����U��xaD��il(!b��(�:� Z��NE�B&�h�cXު�PB;��{oAN�����ɆQ�����M�Q [˰�h��E�rSQK,k�(2��:r�p���
�
M*�y2��h�2<��wK���u<ѭ���'����΄��m9�pQ�q�x1�)��9	榨�,̳}�"�e�u}�L��h@`��0�"{��h߽�;�셽ǎ�⸅
1�����q���ee���kE�9?)�����q�To��|�!^ �6:qv`"L�/t��ԫ ^��.�9_�0:�Ҝ�Q*lZT��������%oAQ!(G����I�~��:M�b�`�ir�f�`谣��Y"v����5��@7��\�r�_�n��~�y2ف��ّ��;�]��Zz1"��OYdF&}���K��.` �����.��a�	��h��S)N�";�l(-\����*�k���a�[sY.r��ى@ �Xgyis2�u�]pvJ���AU�\���;� 
<���#*�Pq��#�K]��c*�^z�-N�ꭔP����a��,�/�0��l�S�y�?�m�q5��/~n��uƿy��l��b��rDe�i���F)�Z��BJ�������ۮ�it�5���L�D��+L�sO��������l��\!��p��n�GW>U�Qa(G���������Þ����!1x��S�,~�B�4rE��&2Ȥ�~rV�W��^�J.�^���R�I�E*eS���CkF��#���!{�����3z������
.�*-�b��U1el�Bͣ?ލ8'�Z�����2��d�l�����b�;���:���kU�*��wk�عn����c!Z�9=4V"���E�Cw���)�a5����t����:�Xg���ꜿ�����<t��՗��މ��g'<%z��ވE����r4*�E2ɦ���~����7��ڨnۧ�����"���5;�[lv��l��/�)k�_���8VGDIWs�V ��?|��3ǽ$�[\ׅ%$�����R�AJ����b�!�����f�n�n���>����9k�u־�#�9�y϶����*�o��i��]i����&�e����g��DJ����냧%�۟w���Wv;#��,f��|���=�ȁ� �s~��jR��t^Zь(�o�1]��̰nK�=S���o�iLؿ�~,��Up��#z��`rd3�[ǚ�����X���y'�ųx$�-���soq��Ƞ(�C���z|-�n5�Pv#��6}��Y���M�縖������ϵ?���˄H��d���݅�z!�|�$[��^>d����~�*��ZĴU������=��gUۗhce�ǁ^�G�w]Z��@��5�_JEؑ���s<�,F�7Ԍ���Z��ĳ���ٽ��gZ���bq>���5M���T���j,��8��Mz.(�P�#��.�C=��`���*�Oy�.%�'y��/b@c\X�0����&I��ƔC�c|�]��\�����P_ϝGGa_@�.x����Hz�lQ�����)�,�s�hHC�y�����^�rX�ލa҇�S�B�|"�"����d�8��%���E�������	U�Wz���ty��ٵJ�����`��������o�e��5CX���1SG,ѻ;��-Y�O���.b��Gc*ZPk#�|� ��n��@:��ƫ�;����$_ �)Ƒ�¢�E%�b�4���֥9�ڗH$�(3�k#�wf�W6����W�����cJ����"�%����7/(����B1���+�܅9dc��݃�\-�f�$:w���I߬X��ԤU�j�E�;LK}�3vf@3/�:%P,��/#�� ���8��|Wn��p�+b�,��Wt�l�f�B%�Bg����3�P�K�n9NFag��q#�|��ir�z�@�]0��'�s�Ώ�I߭��9�?)��EQd�O�@G�y�Z��9O�U�ڤY�үşBq��hUzЧ7A~�a��}$��&�J�<��Bo���	Xg{�V��
��QX�`�y��*G*^���v��B�,_>W��>B�s^�}���+���Ol&��G~����G��_o0�fW!!C���7�������{9��8��=�
�Q���Q]=m�n<���Zಎ��.�c�N�Z	�O���\�'e�������󼁏�_�<����v&�]��꭮����8�Y���#E�5qOU�w޶�1g���j�k�#' �����Q������	2gf}��� PW�ڣ������&���O����]�7\�r#�W�Iĥ%@U�r�6�(v:I&���&V�Q ~�����y����X쫴=�E�����#����S{e:�:=X��4ܤ]rj{�X#�D�O6^yP9
���.��y�{
��LIŘ׷��U�,���W3���T�ͯ6�d��Y�bH��|����ä�SR�� ��[6&�C^(E�"�����ˬ6���&ry��<�+�Y2�T|�D|pd�<���t��Zb�;�ͅ�ׅ�r*�"R�I��'��yآ������NT�~~l0��9�h~�&V�\����5g�����)U�]m��X�|���Z)C��3��|UU�tN��������Nw�¾/��_�\J������)ibB�@�S����}�\���c��R^�Z����l��|�	ZF�hsUU?�G�R>n��Z��ba�,;�;%�����pbK��u�,AA�����!H@��zI�ɀi�4�ϖ��{"��A;�ڲ��!X�R�k-?�4�x?���0���k#�x���s;�����%Q'��r�S𷷤ʝ�{T�y���?�b��͉��N�A�ͱJ�ǌ(g�=����~Gh{x�2�kئC(&]mA=U��QO��vB�6���1b��J���|�"�l���c�o��w��Kc޽<wT\����3�.����pe炯8�Vl#}�&wW9�fX���!�Q���u����7�}�Ij�SǢV�α�G3[̧׮'* N��<�5iS����Tg]��~�������}h�\5��ͣ��ug����M�)T��Q��ly�S�ib��I��%�ՎF�E��-n�<���˙�Ԣ=���i�S��/W�M\0.n�I��
�n�7){)�$�_$��e�N6�GHt��K,g+lk�f�$�z�V��	���m��+����1}��L?��r������rj^ʣ��BPn�XX�v�B�OX�1^��A)�j�%��	5��ͻ%mU.8п�H>��xzO��0��)���3)h�D���nR_�QE�!�]�+$|�q|+�.�b�x29��m�^�~g���
�������}�����Ow#��@?N~�a��%H���&G�@�=�)����Uʩ�g h�8��kO�2���ʉє]��K~p/�![��F��?�&'��������\�jK0��j�b*t��������Z��ZAǕ޼�+��¢��Ґ��	������#3��?8����fAl��XN��B�s>Ҩ+/�����L�S�ݢ��*Bc��s4jk"�h#tZ���~��eF�	ZJ�=m/b�L���
AR�=�񡿱Vm���;�♁��󋱹����g
JcB�@p�/������gTI:I����gTY��>�V��1��#x�N�8�����:+X:������I��q7'Ϲ���.�RƇ��5d�0	U1*�<�.��3R�ܪRG�{�N�B;�٭tۑj�0^�'��5�F��^oIr��O>�:����Z�����9[�N�h���l�*jZ����QB�i(����vE��r��ws��@�%A�&?�F�� ns㗁�.�ސֺ�¾���j��C+R���Z��
r��l�ƬC�P�v�������i�������C�'���Y��L<��W���퇋�԰���'z���	�m�;��7�הF娟�&��z~�r-z�wt[�J�
�̉���r���g�(�9����<����2�)<���&�/��Ο���'�F�n��g����F�J�&��9e�*[�_*�" 
i�nu<������ޮ�Gֲ�D�G
���$�]I�"v5��r�k�t�
�ЛO �n�$2gݜ�9U��2�:�c�'���}NWt̂�%Ue�&H
U4�U�}[Z�[Ϋ%�pq��/C�y����1�g&q���qK��݂ ܤ�+/��ŋe��"*����n���nO�I�f�Ac#�W�� �/��H�KnW5Y�uf�}aJw�ſ��.�Z�Pekl]�mF�c����u������&MCU�D�B}�^��~��b�F�S ѽr�F��Ʌ	Mקs=��������H���o�8s�~*r��r�r�-�HՍ�>�"���z�6�A���6��r�����ˊ�:5���y"�d�-z�#ErB�'�q���'K-����? 9O�sѶ�NY��za�O���֣44�Ǧ<������ʩ����Z����{�ޚ�2��[�f�L��(nTti�렷�}��]<����f��"ޒ�i�������0Id¬w`ύ���ԞR�[�4�#���p~������MO�{t}u��� �Ҙoп��n����L��:��͇�J��~�!�	z�'S��F?��j��$,2��:gj@�Gb�X���cs�[L�� ��vn�2�Y(��L�/�Z{��20�T��x6U@�;�GP��[�����ZX�[��#A�&t�f^2�f��>h�.����5�5p�y�	�J(��k	o��m<���jy�ٮc�e�°[�+�n��0p���1��/A��ē|W���s-	��Um��I�L�j����(�g���S翼�Q���D���gb{-�)��x%���l_�l�Xl0�{I����׉V�'t֡o�����.����z:��$�%w�����E=6$c���ζ�G^��3*b�协&�Sy�J��*1C1�h�C������N�5{0�I4�I��:��+$��'����=C\_�r��$ČY����3�xr��t�����mW��Z�:H�#'�R��s+M��L�ú��S�Qy$�b�8��i-:L���^�鱇��Q��NfW�3RC�V��|���ޞ`�,߅*�7��'�2� ��6�F� 7w��_�ſ<�P���yhޱ��BK> V���9�\�����aT���w�ڮ�^(X����������4��MA��n�	�i�8����� ���L�g�������솙�s��8+7B'h���r���;=�����x��Z���W��
mk�7����Z��5�2#@ū}�ʴq�F�G�m�T��z�/�YF͸,FϺ�ч����m	F����(>�HQQwʜ��(,��E�֬�8>k��h�=O�n��z5YMΫ�[���-K�nU?����P~��ﺍ���	�w}*��x�Yf�0�|Ғ&�H�>`"Ŗ�D�5��b0q��i�㶿b�U��4�F�������^)m�km��/��m���z�"{e�4�b�nf�w��eR�O��?�*��x�p"��&h?���q%63%$���@�%)��#e��k�8��r2�����Ҡ�!�"�ŵ���G�%��?|���^��o[���ezZt6����_nD�_�5���+r���e�mZ����2���p�Y�3-_T�I���w�L���1��W����O\�O�F��kْ� )�{=��#�.e�����^����^�;�n�!���K�9.�`����gc
��}&a�\\�TI��e2��۳���i���m4� �;C�Ė�FEа��[*�?�V ���ۡa�K.�wE֘�|H�a�X3�m�b��9߻��s��`iIy�J�?c�9"ض��(x��醹�;��"��8�=DsM
ˍ;ʆ��� �T���#5*�%�hxVT*.3[����f�]�yM�b*ڣ<�(%%�Wa����"�C��M�����;�������D�y^iW�-��GAHV��X.ᴒ8CH�������p^?�I��d�=N'��p�2��྇�$�/�1N�.g�Q�4Dy�����Kjzf�I3��@�,c�"���S#K �W����J-���$0���i/ǃ��I�Z! r���<�ʆ�[�#�ÚL5��jF���𵥛��'Ѧ&�46�ŭ��u�[<�e����d?�tr)3
+f`�O3с��x�20n�i��l*�x�q�4%�_�紧��߄��]ݾ�9�4�'ؔGw	���hzߡ*�b8D������t�g�Z,�2��R��	���A���3�To�s)�-��-�|+	G�p}F��_}����:�����R�F'ť<	w������c�A�(�v�s��BS��mlQE�^��}�wi�Hh��~���<�WF)�v3�i�tL���R��IV9)Y���U�h�CO?�:EtQ^Su�����1� l��b�����W*�L*�PMڠ9��]��0<U���lR�b5_�w"�0,}��q~�׎|y�ކ!6P�@��JQiȋ��x+?_S�nf�<AC�bhC9s-��ȚA�ny��#j�nPZ����@U�w�e��
�}�1�'+C@��*� :JY�B�A/R�;���Zm�nx���1��%#�A��#A����A*uQ#/9���_�D�|c~ش#|7��g�m�.�-B4�Nٚ�E
ǃ@�FA����U�>\��� q��eBR��]|�5�1]��G�����eN��.������ż��@���f�bj9�D�E!��_���xO3��_��^?�aW���J�HP/�6C��:��_�qP�c6��_L��k��i��S�3/�9� ����3
C�i[N�g�����4+p��Y�+���i�v ���d�k%������aN��7S���Ѧ��#  �W�oH���Oi"�w���h҈�K���BJk�������ua=�)�0^ɍz�DBT�46:,��	���H{+����/�T��$���8��X
�JrC)rW:�/�� WrI� �l�o�m��{~��&)i��8-����(ulÊoK�|i�$=8�p�^3�]f/���.n��^�;vaW��%~?R	��$�~}��C�M�����U���'��E�(�^�!�"?��1��Y��	Bl7��f�rqg����ͤ��n�ʍ��;1鸘o��b�����E��͒�=�m ��bמC���h�[��w.U�s��QZz���}~�U���qmvFى��ᣭ�r�Y�E���R�Pī�!ɺ��Ě���(Lty#X��C�0�Z�µ�o����Sn�޳|т�|y����'[����*��L&=�j5��˪�ϔk�G��"XO(ge�Lv�3�uɚ�6�w�2=K�Rmc��p��G�Rت�8�l2����iuw52{���a\�=W �Il������\f��w |_܊��TX�i)��* �r%l�q���4�9�j��:+�hz���;(�0�sS����%�M�ʔ��'.q<�I��b����1ۧ�q2��i�2$����;����{��+��Zq�&�S����qUv��������ˏ�����S�5��S��0a�?j�w_��tۢƳ�����D�2z����@��Y�6<37H��p
�q��y҆���F��ߎ�q��o��f6�N���� �ً��k�۬;�͐儝�E�]"�܎a����<�6l�#��q����F'g|燳9�N1��P[
P�7�|J�w�]�Del� �]R�_���3j�*1��f��/���+f�;��M�#�_��n����i�+ϖ��&�_O�O�?TPpnK���@��'��B�HJ?�O2KA����e+������y�U�Gy8��W�p��t���5�K�"�>}�:��U#[���x��~*n�>�0�Xk׿��nA�a��ID���/�<���/$�2ڗ#��EyZ�.��lq͛�J9sI?�\���S �l�xW�w	^��c�b�q�L���X�Cr��C%��%m�~�M1!&��Z�u%�Y�����F��Wu���,����jw����Ʊ�'!��g�6Y9���-Ix��)�Gj��u�V����ۻ�XB��%yT�F�J�HI�j�j���S���bQ�B0�:����U��$�[��l.�8k@J�(��ӾN���	
�4
^壓�<�{��������db�L�XOY���9��k�L^��RX �W	"�RW�b��{i�\�k�Mǐ�0(*)�~�Au�O��碝�q�j Y\�v3Uݵ?�g����e�o�����F�%���<w���J����J%[��F�����.~�KEf?�w�^�7,B?���3e�~\��_r������=�1 4I'����������tx�e�����@�ɬ�x����� ��9�����,�I��p�g���`KR�~W�L�U�S�7��,Ɣe��#
�8�Z�tX�+V��(��Ү����U�V�M�~��/jw�L8�5G%�����"�:W�G�T�@-;`5�W��T_�c!�����$���?��[i���8
��.o$�6�������u&�KrЃ�d��:,BH��	P���Qo$��*!�����BHc�5��IvC������D@�y>��)�0
_j��^p��l�ddBO������#kk�K^� m�c���I�*W�[*�%5��pLv���U=U�\w�|��&2�on|�F�x��fy�N����%$����Թ��H%����9W��C���xꖶ�I�@x��-+�ռ��V�3`Q�LL;���=�� ����+a��A�s���}�Mq2�����xt�4�kD0q Մ�m��*yC�%}R������_Q�at�_�.3Hߌ�0��܇!n�=ɭ�Rb��E�0���.�Qʺs!b�	k��3zݕ���in�H?3�lg�E_��"���M����}��=��sx��k��k��7C]�M�d�
�OZ3�a�
0K�#�=�Ʌ��(�[�; ��_LCު<��"<��afgoPB�����p/�ԅSM���^Z��=�1�g!�7��1�T�5��>'�_9�EӃ��L�����o�7�S	��Wd�O9z�����?Bq:7���t�R�\%����`���ƕ#�-F�����k��!\�Pi_f�q/*��w�@�f��>�?#֒�e�.�f��a�#FR�����&�l��h��:�p)��_�6�O�^�r) ��B�Pb����Z*c�Q�K� ~�&��Vv�Di���)�@�����dm��7^3u��qPQ�"��-SxI����/J4konޛ�ز�B޿	�nΨ�KGO���hЅ({wB���z`��b�b��1�2a�ZU���%7?X�Ö0��5{{w&+�)њ�Ǭ9BX�2�
�l��#̡�](R��]#���[0B�q�&W�N1wy*~�
�Q��rR� �3�۝���RVbq�Q.բ�����b|F$L��ؘ2V���S�^g6�Z�K�h��M��)	g��!B�QL%G4���~[Zx�N���A����Q�YX�IȜ��;�J�R��:��:6��3�,��b�qd�Q��̇�~��z�q�Ȍ���[r1B��
���&S�[�&S�'F��>@��M:.�B��B����*"�6���S̿t81KB�JP�}i�6`W;��.���F�����"QHxxoD|����59��7'��q��� �u�Fk)�c~vq!�m�M�M'y���z�-�B:�%�ӽ�|�+&�%�z΅��--<m���I+���Y�nwg��&��7	���~���Ɏ��Mq����.����{a<Y�ԚWO�!�3Dڌ;�<H_Og��F�E-���r���2��%w�Ԥ�^�+z=d�M~'<`�B�Jʥ��1�P�j]���
<�@e?��U�1H(j���:G�ݪ$'�	�z��~_���m�EI,Rr �h�^V�U�7������SwK:z��=iwI��=�*��*K���ݿ���O�g]=��6�`ZVs�5t�����9��"�>����ò�[
޵֏^̨q�?��[d��I�y�|�愗|Ng0PP.�|��@�|����w����m;�@1r%�Eo�p��;��@r��}V>pf��ك;r��b���֡2���!�<C�)��q�Y����l7Qi��A~>���c��`B�C缄��.��u��u7�ծ�(N�"r���D�g�}���qr^
n1���W��"�r{����=�<ڏ�d������$��T������Z�Ԍ�{����� �@���t���$l)������cЫN�f�¥f�U�[��E{�<sh�&��!��1r����"|�d������������k�+���U���X�YH��s����+�Q��{��38�hȲe$���mg�_�C�
W�L]_��!J,���s��/f�d���{������/UE���U��V��nԄ(E������Pl����y�o�����aKw�[���������F���+���52lZ��o��u�tn���T�b֦�e�T��oI±<����Yn�I�P�}l��-	bZud!���H���b��$t�o���ۋ��(&s��'����q�W����c�Is��t S�d+\�!iJg��`:���w&E���*S$�AM�B%пѩJN��m��}��"hZQ�jH'T�7�P5�5�ܷ*�6 ����/��� Gb;���j�� qI8m���(s9ܯ\�j@��[{y�+�(�ܱF����"l�܊�+2qݹ���i�g�_��},��3�pQyU#o &~e;�I���9�ѭ�- A�W:>��>�K���8���7��XC"I�m��d�\]Ć0c��Jt��J�u�;pJ�W����V���pm���L����V������`�9}׵Yv����� ӦOJ��mUш�Dao/�^�AJϵ}0��p�	�H_����)�mvk�fI �ȑ���|B��H��C�l��O������%�֬U����VX�b��[]�t�����$���D�_�L֋�H/�0��:�5��YΆv�p3�K��Vn��d�{�_�Xv��d>�7�"�\��f7��4�����#�s�İ{�%�h�鶂���d����]����|"s���=�#�P����+�<&�f���-��Ķ���\����T8�}��k�M4L-[%��B�L5�~̽0����<�+,��:�!����"5����YS��f�%�ulf�f��]{`6��i1�_=߰�C��6!�<��W*����Ib��~���<�7���0G���3w���H����Fj�q�9C�OF�J�G���S��E6#鈞����Dnc�D��M�rݜPh���o/�-gY�F�c�p��ۖ'\>d{�;���`
U�m�4x�0lea
2�J��5aYg��]�^ןۮ���|�o�4t��@�t.?3��\$k���9G�W�\[��<�d����k�����\ � {��&8I�L��9�·?��5�YO{��S�!�a��=]�o^�)������?��(Ro�8���d��0��O�.cT1��C��(�p�������[h�V��R�ɇ2��z&�v;W��ޓ-�/��C�z?�"7(1eV
��c�/9��*I�,���=��&0/�!b���*^�e����~�-�/P�Zܑ���f����"t;�*� �^K����] `H�T.-sK��vFHb:��>C�;���ިL�>�[�*۰Q*D�����#�6B��v����Ǥ�3��jnKb�����+�p��R �L��uѓӓtf�>*�#k��y���k��!����e,�2ȸ2+i�g)�@�(��"1\�y5�ֈ��/���	ރ쁈���\";hOV�(+��K��+�Aw�l�����:/�J:j�䇚�.��g���+"���=�H���D��>�H�t<J�z�l2��qr�q������K���5����fW���N]�cke�'�]L�9�6Jߍ��]�z-�r�1�c��u�3���N���I���H��vXӆ��A�*[4Ro��s�(�{*�ӂK>�~�6�E� �<>ȊJl�R�?�\7_��O7ϴe� ��\�n�u��ɾ6"LTKH�&�n�=�2���6��+`����r��)��;x�s@���^�\�f�%H�)��>}�gV����j���3�.�$��m��"��FsT�m���8��Q,?qt)�&��f����	hc���Wv��
P�:p�p�6f�|Pe3����X��b�Z���p`��l�)g�����&L�MZx�����h�/л&�k}E@T��|��M�o���Z���H��n�vJ,���3�0q'j-	����O]k0��~�Cݦ;ݹS���Hȟ(��>ͺ�ʄL*hU4��� �Y�r`�79�A�ӝNA����S^������<?�O-� z:Vn���o��Ã������d��p|U�a�rw�8�Zԟ)�DA�(���55֦��/6��n��ة��O��Ut�����������έ��{���8ɿ�98�FZ[V[��²��(Զ��pn~��;'C]'�R��Vހ|Nq{�(r�k�5 ��wY?�Z�o�.	�	��U<k�I�F3��u��I��@~$ʒ�
��pk����`�r���4��'�ƎMX�^o={���P�R��L�ն�/;����5��dko,�>gE �m����UC�ן�u+��ZI)�T�6�~I\�o�s����"���ZYĹB+���܉挧�ƭ�����\K��Xޔ��!�?��MV���G�|���u��ٱ}E�äc�s�P����Q�.��Г�
��������E�hO�{Lpl��"z�j 7��	 ������N$�~�$p�_��ƒu���ȡ���
\[W.X�xq؄W�Z��%�����Yi�Z)�D=k8	�z'"l_�i�u��U�$&	>nǼ�|ϟ�q���z��� �T�rפ8�W�5���>��x	�>�E�4����N��`͟[U|�
i�χ꜐$��5
 S��bk�!��J	��I�譸2R�߇�r>q����'7`��q�F<�}�1g�_x�q	��X|!��[��&FC=�{��� �+�UE��.�>_e]́��;����^z��ۜռ��·^����9E���3Fz��A��x�s�n6�=�w#�5F�e��I;7S7� ��e	U�Y^{��7���`��>��箆Y?�5�e��'��D��(��y����1x/�%��J|�=\V�"�^J��m�.���I
��х*�{8��J5�R���0���W/E+���#�H��̸��e&-�ڶT�ǣ���ѤS�q�Ns!G��)r+efW�1�:aS�CÀQ�n~��,�%x_^9�ui�~�ItNG��*~����'����ؓ���.\+��'��s���!��w����(�^h.�ʽ/�3#���f�?�P��f�qU����|�pX#<o+�gc����3�:�u���}�b��O+��w&p_���DG��*�g�n�
�l��
䚶���~���vl:A����GI�R��J_��l)[3�m�2A�i�S���/$�,����Ez�Ys���D��G�p���b��1���=����U�[?Y Tm��Kޞ_��R�����N{�U =T�Z)�Ɛu+&��K�l	@�������*Y���+E�x��5���ǚ����"�����L�����	k�}��p�΅}�����2%�0z ޖ��(�^�l<�ߏ��ї/禣�	Mk�O�ؗ>CS�_6D}����5o�`*�bb���z�^��}��=޿X(��S8��*T��e[��n�d�/خ���3�)����0S��NcID������F�a��a�E���w�|� B�bZ1J�\eDh��u��-�kD������$�W+/�\ͮ)�S��yZ>�`��<jZmr����+0��1�s���5(b���o��������^y_F�uʑ�US��I.��Jl�/��hI�}Fg��8Π���6:H��v`�PƝ�$	�j��b� %XI{���$��T9ʪ��W1� �RFT�
êu�yt��6�I��2���Oq�qM���tJ��.5�F	}���J/F6�`o���tgԋ^.�˽C=$��g���.����~��F��Mo�ꇶZ��/a��3�䈢ЂoN��=<5cĆ?�GR��o��11�+&��Ky%Z�S�`��X��̌�麚�M4��!���[�.Ϛ��rGT���e�	�Z�:�L�/���;�>z'�۲X<�(V����w�D���'��:�A׍h��J���}:^g�Hj����	ɍ�Q���Ҵ����������P8�x��6����z� ���� �GT��5�tޠ3�`m�n����؞
1X��49ˁ��I?3��m�M�mq�S�nİdI� ͚��?��GM���=r)���Iw�V��?�@��?݈A)����i���1�����Q�?���vb��������d-i��}��&JcK�}��"�,u���}yZ�O֟q�/�V��E���z�/8�sv|8},���VL��J��m�W� [��	u���J��$���ݤ��\/U.�ߦ�☗O��/Y&��n��~
��.S������Գ$Tl`�>)1;�m��1_�H2ه����1/V�i�xd�щ/��J�[i�N]��<~?��9�n��GM�������������p_�?/�m�����T�3-(��ڻ�����}wOI���v�~�F��tYVd�jf3�� .37�.״�I�����9�n�b���	������EW��X��}�d�O��@sSM�+�SD�2���<���t>f�K�}_`M�Z*��\��/27�(��4X��@-A�;��Chu�ק��h� G������K��e$��'sXAa�b�oĥ�����W�GY�!)�h^�ڻ^+m�N��0�����
���Y� �e�L5�u�~�p�&PZF����g�;b1΂ADo?��(u�!�4�(b�uǛ��,�P6=C�-ns�W=	a��6���atr�w]���'���Y���*��zh��B�2�7�Y aF�N��tC��Y�mZ��2�I������x7X�"���8��׺�S���U���-��:��su����.���JDf� )d>�Vk(�Y�W���zb������U�V��!�~�-x.��y��� @&�5��Z���kc��1�ïr¼A�h��m=lg�*������ 7�a~�~�.F�͞�N'��ˋp�ܹ
�ft��d�}W�;l�^/�����9:G�q�ܟ|�����`z��O�����_�Ӵ��a��S�8��~�i����g��F����'ܢ�F�������5ﰙ���TC#~��-B9�i�C�g�n2HI��ڐ�yK��w3JKuLA:�yMY#�Lſ3z�T��{�>��-T�0߉c�P�G���X��$CA���~������\[ɫ�����8ʓz���,�|.Q�f�k�*��39jM��X�yR
�[e�6�����5ґ���:ù�D4��5�Q7���%ue7���IB����j#H<^��B�sd��t�u�D�/��"�Ro�E;Q�Nfl%�քn�wQI��19���j�D��[6S�=F�at��2EQy�O��4���M�Ǉ�M���BW9EHM�gm[�/T~�i��N�jI� A�p-T��X�Zk�1�6�p��/U#�^8�#�����ڛ���O8�S!_��b���(x�Y�a\��&����k�e=�1*��Nq�!����'��Lǘ�,���曲#+�^*~��F+��f0��/�sm�2G��{e��(�\j4���[�pFĐo��S�Y~S�w[��KFG��7��j���˹\��e����:!=�a?��I�u�:� ����������rh���)>���&�n8s=B��.֊BP��mi����)n^�ds��7Qq��g�]@�� �P��-=I	���=����4i��@�����X�_�4�5���sR�}�i����K��)H�n�T+�?��O_'DֱS�lZ���BY�
��ɫ@�[X���Ljܳ������v����J�IU�D4x8( <��s�'����ԍ]k���c�,��b�[ݳ$��g������f����#a'1�����hC���渵�������	ܕ�F-5Yb�Q�-���q�t�����'�Y�C?C�nlDq�:��ņ;�PDӊ��}��9�c�O�v�� s��d;�� ?s�?_j�";��O�|S\�Y+���9\"K"=����:�&��Jsv�`����Tr�uY� Ϥ<��ڛ{�$��Uk�Hx�㊮������#��	 �^`)Mx$�������"rE����nmo="6��L=��gy�Ϳ=U����������Yk(���c��ִ��X�c�kʆ��
�)��Q��x��W��6,�,���5/��P�Tҏ.��i�L�5��C�i�.]�Z%�<;`0�\���׈9+�n{���|�zhs�,m�ҮZ�O{�1k��ȇ59�G\�uEBa|����N��j%�u/���l7p��2�: ��x�j����;˫�j��	���:z�qVY(����azL��ʑ�ocOMS��צK`w�{Q�i��O�m<��C�s��R���"�Ǚa�*2L6ETU�Q7������b�T4 !����*o�����e�֛1�̩�/���f�����/^��6���_&��_P���5�r4b+5i���ԫ����K��R��� ��ZT_>Y�q�}���2#���a����������h>�������m�|,���c����Wd����9�~X�c!��&�Η������CmW�������H��J�@Tf����q��va��Z��;�9\���p��A�y|V�#(+􂸪&.�Q�� �5��2�y�;%z�gԗ7�������?.C�_��Į˾��*H�ጟD̽�	J(�y>�92�L��-]C�6�Cn|
��|wt	�/�0k��z�ɞG�=R���!�G�x�]LT~�$�(V�Kv/��kD�k1H���}���(�ڏ�O,�/���Ґc�Bh~�Z�Od�9n�_��xB���n<������;�	��c��|�~��.�;��Q�'}1C�3�I�����AT�k@�*0ƶ�6����5�Z!�y¢�{��n���P�b��~��F �88Y��n�7�'�7D=�䠸���B����6v�3L�g�u��J�Y�M���xzˀ���i�-��]����V�Hq���ݭX��N�Bp����n��~�����Z3kfN�I"h��rc}̣z��B�1?�����AF�6��
����W��Si``�ġ&�-��v̢8�$����M�?�w�p�����\�M��dZ0�/.�nc��g�j���a好���o���N��)��j�e֯�].�w8L�7)>cx�,��������<~���tn�ʮ�Mun��e��Yl��q,U�/��'���I�]ׅϿ\3�
H}��X�L����_�$�E�]po�̐1��8���x�S��i�5<O��R��WWz�@9�C���7ߚ۾A�#�+�f�t?A�X�H�i�'h�X��Y��`@2p�?#�0W5���������XS�z;<��ᾑ7(!�t��^`�˒vD��̝vh��Cıi�ln�=O !Yēr)/U��)�������aҜ����@�Ô.���&1	��o
��j���d�Ͼ��A�'��1&
�I��9Hx�l�>���n-8��l���VD��P�f�h�� ��%���*���{��szLi�X'NO���� h`	F���NB/�Y�Q�ZCXXА�.T���w7��Z���5���P�|k�b��>$2�-�+uf�β ��N)��H���1V��D�#mq֚��O���1�jKٻC}t�� �{�K�D]L��	���>��,X���E>��'f�~f5�u��M�5��LV�%:�&htnl���JBxiND�m�\Q>������k��@�,H��h��v#*M���{��-o��2�o�2	���m��l25����s���*Ĳ鱄�9��/zg���G���-b�]]c�Y>x��V����g6�ð�&�iDx������I���x��"���EQ0{�q_��=<�2A����,�K�{��=�/4��b�;�dMh,~��n���Su	��A�X1μ�$|�dW(��w�I`WOY�ɗ�{0���n��fa���p�y��@���װ� !x��;��$�^���AW��w2��۳�Z�W�Y�S-gspE�4)$�k���Z��O���P/K䮡]P"A��_�J��/����[�:�W����S,�g�U���9��b�����#� � ���$wG����'2Fy#�d77�s���v���כg���x1V%�"���v��1�푒��0 <��d�Y��oH�~T����g$᯻㭑O_	c&��[l'*DڎAC2A,��o%}b�w����k77�Ҧ9��(�i3�*]'A���y�~���9jȗj�X�ԕ�?a�Q�,�9޳?���}zN�2I�v�Z{��<�\g���l5��*��)�	�Q��;�z=ј���9&�޾V��_������`�=�q��G�+�=��:[�i��å�&�w�k��p�SP���`�jQ��`���#�w���:־d�,o��?hζ°�1+fNWx�t!����̒f�n͗%�[�Q?�@7&nh�@��C�w���ݝ��o����:��-i����+
�ф�_����ҊLVP�Z�i��)
�awݩvs���V��뚹[uZ�F�M��dN찁���Y�����){�tn�� VF$i�M&5�mM\���Y�!���8��0�U�M�\�3�bF��5_Ur���������T�(��4�^�}ޟ3�e+��Ҕr��Ɨ"�4����@"�1[C����$�I�{��,ɷ�୻�(U.��-Ŵ����zH��H��R��B2b4)K旅�䔤�ڣ��ߣ�]3'0�5���7�}J|w0^����+��5?���O�h]��4��_J8K����GI �YE���u����f8"s��s�E�h�c���j�u�Y�Iw�u�.�%�e�sR�2�������ݸ�1��y�"�)QE
!��剧�~����f^�&�w��H���ix�_��ON�I�mg�_#�8.G�I'�$��Ő��K3N���n��y��Lɷ�K~~[j�4x4X�`p'��"�H%�Ys��U���G�C�x��ůhלV���Qބ(V]�����,L� ���V��?7kt�/ﷂ��fS<]��	����'��8"�ai[�S��~�W��؄�ݕS�J`.}6�r���{�K��$��@��ܲg ��C�u~�ǡ������]��T��6��p+'i�[ׂȝ)�;��:#�N�6�_���ʆ�����jb7*|��f��ǍGD�}}��������g�ZH�h5�Kæ*����M���!�u��\T�=
v?�Lr����T��@_5p���n�@Rnح� ��� �����������9�޻6��P�&��+Sm�Q\+%$��b#������ �IBys�X���?�0)~��3��i])2���]/ �F[�],��'�D�ĕ���`�"�T2fd�����r�Ԗ��� ʋon�V��IS�k;�Z%�!_ώ���V���r�Д#T��O��nă���<��4��0�I�%7+6�9p og�3!��XyD!2���5�	���3s_y��|��	�� kiu�e'�V�ם�i�.`v�h�8盅~�e��u\��o��P݅��e��>�r�/�'������ �����������EŞ�Vm�G8A�fL����Z��Ut�c:O��1*ӪN\�qa'ܙ\�"

�� �UH��EH�.�h��y�:�����^������g!+J�Lh~��Ũ!afO0��Z[ꍰY�1�Hx�+�/)(�b�[k�!]w��}Ꭹ�H}_9�����IJ��E�{r�.�uW J�?)��e)�%�R��V�A�J^����o��u��`ib�ïFyauv��;�`�gOp[OHG�1^ocjY=La>.D�g��
����7��'�(U&t	�y��S�D�.��:�e��Fq�`�
��d?�ׂ3����S:�A���g�檖��1*�l���g�.�к�Rܢ%X�_����W����(� C�����������m��1�x\O�U�Mqe��ˎ��k8�.T�kQ��F
y�*9	�v��; 3p�h68%����E>&4�(?jL9�!Ұ]���皱�5����Ŋ�q��&�r�ӱv�N��>%�d��Y�����Y{�m�LC��4���i��8Z5%����?��TMՉ�eC�z�BO��v�z�b+��6կ���"!O��~S��C^q�������,���(��W��I|���Oc�G�0�F��t%�d��W����V���4鶟���7�)�G�!Br��UJ�}`l��V�RV���A����<.�[f��Ӂ�Zjx��"��Y���	�ifA}I�6z���,ۭ��N�Б�hw�?G�@�}�:m���u0F��kȑ���qx1[9��(����3qUʂ�:8۟C�,���Fl��r���n�W��=�P'�1n�߁����w?ٚ(��K)���)�1ZjeG�aT���bd�Baa}P�B��c-�1�N��b@�)������Ȧ��;��7x�8&e�a�5�2�#�{�2�+y�}�xv�g��9�Z��QxMiM
/TԵ�X	���M�o�B��u�Q���#{�.ط�=M_�t��Һ}���k�3""��h��a?��o�����Z7����L�f
V6\�ӝ��Y�J���!vA1nsЃ�e1vkЍ�?
��|�@���f���@@�1I_!�a���{э3�'��1rV��k����3�N��&����c9%��@�z���_�P;���:��bG�ԜյZ�rCm7y��������u�� �~tr�:~"%�Ѻ�"ߓ�*����F_h��eE{~�c��L��8���	����	��3!LD,��E�]o���+�z���u	"I�K��Xo��9��P"o��B�g$mȴ�.5��X
��2�wS�o���:�ѲX��Z�V���ӌ���4X�M�������߆�I�1���!�<���	Nc:qi�*�e>|'��/�;{�]��W�����6�[��{�3@���[�dFp���^
��+a�)\sPY�vS;�퍱�X
%�(X:);��k�1l(�i�<8Jׂ;z�xr.�|���=^��bQG7��5\�C���J2p���z\�|Z��Ռ��(�m�G�����}���[t��S����D��|��y��C��e�3�PX�jq�ɨA�c�-9���p,e*�-����,5��,�ۚ{�,r�9?��$j�&�(_9f�~�R��3�g�t"�;���q8�"�B�\wBH�%��%���+�U�v���ϥs�1�kx���{g��a��$�U�}P:|�j޺�=��(�h���O�1���b��	�����f�{O$��7ir.���Rݏ.a��O��C��L���͂�OPK��kd�]��;Ě�|�/�/p�m1�%�;-���w��{cl�R��;��N�(�S)��Ӌf��o�A廼�Ftx0�Ɯt4�Nh%RǼ�U���2�U���=�To4�1��N�5��jI#Ҋ���I^rBq�s*�{4����&Uh�`�1�2-�&����/�gm��"RR�V��5o�&����{��| � '�ú*��J�e{Ƕr�cK�9.��5RD.+���$�۸�J��\O�w���,/1q��59+1��z�bsV:��>B�v`i~�rv�����y���XZ���z�UR�P M��oIZ1a�Q��1G�Gkը8���JWL$6A�����wm����z���=0>)�J��C�W��1<���>.��i �!Z����y��m)�}1��O�2�e�vX2Ɍ.u(,�_!�ŝo/���$���u������>�dHh�)/�ȑsw�b��H�����5u~~�X+e�)a����+tp�r���bl>.����hC��\�7�=�~n(��O������¯�'m���������y��]A�jX���+,mj0�xڲBN�S��,@�	J��
X(٨.�T
G/�K�6��Q�ţ�"�S�p#����������#
�0a�vdI�UԻ��M�DZ�����:o��\�Vy��G�Xf�K���lu}nD�V��t�����w����F��v!���Dr�sz:����a3�w���d,.��P�g���R����ש����M��5�r���-@j@ϱ��8��j�g�m�6����dq�)X����b�f��M9/X�|zv$9�a�n�%���ҧG��iIu���ޔA���k�g���×��q�ޠ�Z�j����6N�§��;�O�rF����!b���1|�(n��T��K�������s&%󙮃��X�G֎�-�����{ 9�iB6�j��T����u�W�O<��� �B�=��Z�C��T=��%1������`���0Įh���ж��QЬʩ�)PYL�b��?G��������@Q^ġh
#�H�������[C�~#!��[���V���a�'�%i&��r������k-�*��M%N���tv���Ho�Y�ժN�c�ߗ~b:��#�8��A3�`s��tb5}S>$�R�۴���D����,[[p�ƀu��[|:	^F�69�
;J��d��U��jt$��5�x?�Q�U�����|��d�� a���\����Ƥ\���]�2�`8Fo;�g?*��9����="�]��_P���TP ~/�r��:0�{SJ�S<U����Eg��#0X�"�����ˈ{��.�Ǣ�应#r�jɯ�:D�7,��h[��Xl�K�K��l��:Y��Z{��~�g��S|/�	�hK����qQ8�*�U�N���rw���g>J�Tjvxu��"���.|�~M �6���f0j9�Z����|efklS�����]�ˊO��S=S�Gxd}\~�r�i�gF`�N� ?��U���Љ���<��߭@d&����ق�1�4h|Q�q?v��ˤ�
s@�$9����ކ7B����|t��4��A�K�#��SL�ϋ� �H))�w�N)DՒɸI���m�8'}��)�jP�ϱ�T��Y�7�є������H�^r���gdu��
&��p�o��h�QϜEה������`�f	)��i>�����BN��B��/��㻡D#���'�ÇI�zq\s�X���j��R}���3/�]� �.u�K�1S-��E8ґdx�g3����~����Q�s���ss���q�޺(��v�*�V/`<��ռ}{���mǵ(WZ`��^"F�9�2��+������2t�|#�CQ����/�$�v�a�|��3���j�/&������yC?,� v��|���j�	�K�
����gOK ҕ�4��,�r�Q|t���Q:A�������v�@U`gAIX~�C��C�GwUD�7�K�^���-j�������R{�UDƙס&K����[K)��$P�5K�r����B�D��z��YԵ�m"�0�`��ET�!���G���w����/c���jn_�ۜ4��xc2�d�-�о��j��k��GJ_��ee��o��EF��H���TB�䩕�T��L�8Y�I�6m������E��UJש��A��Fi�>�=��7�U޸6`=F�!��aR�O+��=k��XC��O	��J�Ru�A����vXƂ�(C����_�����<�ٞ�c̵*�h���f(Q�F�� P�y�����X:��\����k=��LM�3_�)F(��meʋi��G��㖠+g��#�n��vn�*�����Gf�:�'ް�TKz��޿n�mX�E�l�f
��z�k�����Ѡ��Q�Omh��MB�\�;��8Ȇ�U�����%^%���w�2_����;I����"��%�sY/�P;����X3���F�u�yc�"��~`�m=�c����~&������\,V�#�TV��2!�� 嗣���&�fB�d�σ����ќ����cdȰ ���oJn���H�HV|�DyP6Ӝ�lPg�d���8��������a�R5}!�6߁����nϛ�tg�Ҭ�W�����wh�P�7*ħ�e���������q�o���Ÿ����N}J��금�eK��M�,�V��S�\q���U�#&	&C��@�����
���m㊜7���^i,X�YR�	*v��z�87A�Ix�}6�כ�'Id�L�Ě�h�O�&io����Ԇ��3{~���-�&���)�@���'��xN��|ߢ*dT�5d*GRAU�J���	�$��M ��u�:�'���4H
��z'�xvY*���M��m������~���ԋj����o+��o��d�s��:�c?B5	k�	b�k��W�a�$J��|�<�F���c�|��)����}���`�?���q�_��w�j�M��� _CL@�~ ����}�Xt^�.ɰ0P�Ϛ��$���_T`��|E朅|���q6�u��s��-a�nƋ]�**t湤S{��@)�{�G�5?�B1��mPC�E��t 
�QU$��i�-?*t�o�Y', �O�_;�Q��3�M�+ X��i�26rI�q�v-Yp���`S��2���WC�s�����Z0�����N����v(aD�G�b��Z~��y��}�懱���� �b�*��D-~������H��G��Ǵ�"��{�3ls� Dӑ��� ��2��$�]UQ����v�w�Z"�%@��7�'�"z�t^<���䲙*�ܤ&��T%��n����9L��O	���+VL-LR>5o[���Jm�16������JJ�i�� 0�nh����|��n�R�(V�/��=���]Ů:���n�Ry��q��I�ǜe��A�B��F�a���P��$�di���S���4�߳�̶'�?�ީt�!��)b�?dt�5y�P�m�)
K[�QE��(��@��a��Z:����z�ww3ZE�Xܥ�Q^���՛��V#�c��w{�3q���	�<�v�UBB�+�]c��M�ɷ�Bĵ����S%�t��m\�H������XQ��bt�`�k�" =�%j��
]�2g�}ß�`�'���]U=��S�40�#��
�*j5$\�m�6�R�
�o�K(pN����K�W�-��ۉ�N���w���eAQ�G�Yp6m��:�c?/�LGr�a6`~�Ӗ�吸����<=�A���"�;+o82
�	�2�C��j�UJ�g�g6���K�H�JJ��҄��U\b�f���j���p-�����_K����
yܹ���5���VY;��"���O�>[jEQ�"Τ-��ㅡ�e�&�*,uj!y^�M2Z=��?���\vL�i���-��3���������_b����M1�o�x�<��kQ����pl�͔H�k���h܌o��-\nȯ}$4�w�r��Z�7��>9��#'glr@o����H�Ʒ�aǿ`��yl�� q�?�p=����_���li�Ϩ��bN��m���1�Oc/?[{I��vOoiԄ�-��OԜ3'�p�Xb��P0T��(���}��&">�C�D�R���U�/GY�n�	�V
�N-喝����K�ˑ��e�ȳ���i��X<ce��� ���]�Or��l<�� �o����!�M�Tb��4������,�����TY�����B"p�⚄$�1<d��[S�x�;�c�SJ�G���Q�z���8�r\�����Xf�0�2�x�H�zC_�.3�T�d/��o
i�u��e��a2g�IY�oت��	��c%#�;�t�Cuq�hCA�&ZH4�h�x
<QW^��P��,T$
G]̈�=�$8�
���O��r�P���H �wN��uU�X�-l/���������EC�Z��R �lc�r���?��|?pFU�B(���ް�����Uo�	x�^��~M/p��݄yV�%������(�+}�9�8zk�W~���-B�d���M.�"�4��:^.#<Z��/}2�	@a�o��E����ȳ
͎'�x}p�P���(��C=	�'ƾL�������L�^rBs�]��3����܏_Ӑ�t���z���@ۖ�=w%'�(�.�����sR7p+��%�0�l�&En�Q/����R��q��M3C�޲�z/�ًXd��0&�LD{*�T�E$�Z���EdNn��u���-�"�G/�� ��B��$?�؟��aI�p��	�tko�MK�4���bi�k�a�&uY�u��8\hv��a�`��@ȝ�ס̾�.����|l6���Ǌ5�9�3��B���G�Ƴ�����|�j�cg��g]��MI�>f�s���(��8�P���h&��#{����'��6i�ӏ�v j Q�ר��@7�*L�����ӝ���Nr����pD��L=�B7�3q�ԨǠ�	��NY���"���īIu���D�&��l"~)EAi�ݦ��ɨ@a����;�&c�X�6�����ϭ={o�Ǐ����.+ �.#J��{��lob�C�IB���ZIfvEĞ��f�={�L�{��;�ʠ�n�ˊ	}̺�=.��ߨ��Q��m����)�j�Vn��띖H���g�o�j�!�Ao��7�fH$��OK�b��Pi_pb�D�ȢIO�MT>�\.�Se�W~���^d��-Q�fua�����'��{m&'d��ը�%`�pk�F��#��/.&�t(i�&��⧔yDȗN�R�������*����\ƛ;�qA�W���+�ۇ�3����c�����)��p�癏�H̀�M��^�Nl8e�o�ڏ�=���k�Z��3NY��v[2�Q%,�<�0I] �[ ���.����v�e���6�"�xp��>!�T@����+n(�jɐl��`ȴ㏯����u<("@�:�_T��K1Lѕ�֕Q�π��n{�u[D&�Y��!�`�J�2wY<���fx�h�mGkl�qV��R�g"Ԧ��K.���`�D�ɭ@��PC�_é �mԜ�Ν-]pV5J��b�g��<���Ӯ�/d>����?�x3�-W��7�M�T���g�o��:˯��ڍgmOE"��u�;�~qFX&�������w6'�y���v����U���2b�"�& k�?��GT�� |�\�2,�oaT̎�y(�̂��xߗ'�F�9�{��0��Ȼ���F&�{�"u?ŧ%vp�f��S�M3D�Ǩf���� ��k��6j�,�˯��m*��lN�(���2�*��n��7<�Hq���Â�i��5l��d��Zٶ=V�!QD���g��[�>��u�w'��T"z��w��W�a3��b@� ��OBR.Wb:�X� �|��Ԃ�1�5q��}5H����RV��4�T�&_��km����װ�Ŀ��/���^��ގ�F^+>��]��H�g��`>PС�;@�F2%�1 i&.V����~�!����@�-���� �X#�Ӹ!���o1?���6�$t�e���
�Y����˝�d5_���Z��ƾ;��5AY"�#m$-T<*����(y��h8m�WO������:x��Y�$���7�w4�QY��F���Qk]�4�a�-���X���}gi�H3/�mO��~qvu_�Iy2B�E�[������{�r�" �S���cQel�\5}�
�C�������#���=�����D$�Av��H�ZE��/	h��dڅ-[0P�a�u�r�gٯ��:y�}#=�vۈy��@vg�Ti�����p��D8ZV�qs����23V7��c	���\+x4K�:�A�����P[�t�+�-��^��=�# 8�ơw׈�lI_Mv��i�߃pl��4��5�L�O$�U���#���5�F0{$*2,DC����!u?f���zu�͠��)�D]j��K՛�C��m.ػ����p��mo�d�G�n&��@Q}��Hu���.K8�Q1:Q3���Je'�c��X��g����S�:���J��߄�aJ�h�2�**b��~a��#���M�K]�M�����i��?�é)�y�����א/�뻝dP�F�X�Lpe�^��2����9�z���avD'���o�����L�(k*x�,,���uC14ؠB4���I��&���:t��}7��"���X��7�6��7r�Qt�9tL�p����n�?��ԩ^��+���}�� @]�gNI[ɷ�?�3^v�1O�9�-c�i��Ѓ��_,Ce,�6lWp�E0A��	��'��*�b�E�<�� �ێ��(��(��-$d?�{}}m4Pc�8h}��q�M�$��n� z���=����J�V�݅*k:�$X�����Ǡ�Ǡ��Z�X6�R���{0��� Dg�+X��㹛q����
2�a��1�!��kb�������9(9���+[nwzay4)��Q�:=(���4��=�nXzt9d`A`�wX��y�xXػ}�����Ml�����խ6���P��s0�y�����da���4u�&��3{"d	��<ZE�S\��\��oJ�V�S���x�Pۭ�f�r�O���x�دj.�O��x�`�l2Ըx��2��
.���XmUjT�f����
��'��i,�{����R�X�&G�߬(t�!��~Ӝ���x�Mj~�ߒ���!M�◓k��M�.9�(��A��ιf�eMq�g*���lmejJ��0����>�<�J���S0'Ts�o���<=�d»��yl0�*����5��^KE�B�z�>��z<����&7cW��a����Y�ٰ�a�ben*����G��D矫��d%D����z`kп���>��}�͊@���l�R^�+����o�P�˸���c��r�3F�MX|3�͈�SZ�u��G��"���N�*�C!����9i�QI����2Z4�r쩝\��fU�`�\�-A�]��]���������K���o\��%)6���:93 �F�AȚǽ��y�&��Z!K�Գ~�t^���a��w>ƝO_љ���ت�m�/6�a��2�|��C��15t��ݜ����=��[$�at馇�tw��m�#�j):�s��{�:f��nd��ĥ��#�$C��_�B�˛���<.�t���N���\�h�\�,�y��?J�w���'PI�21������C��9W #���1��k�t��ܧQ�͑?�4t����*�hM���zkN�OR����y\7���"�����Ё.N����4�@ �f�8�9�vw�н�尾�ǵ^�8��=)�KpܟK���&ik��9��� ��2{[�����Q�N)��>?�xU{kS|6*���X�mW��$XIC�n�H�t��an7��=��TR�(� Cb��G�BꚂ����L+�klF��nA;5�D4\Z�V���P���Ȑ4�qRV�;[6���p�:���J4�2�A���k�fZ��P�Q�����ZZf��z���9:/*i�	c��tP5g�ܮ�SV�����q]'�!1��s��Z�;��!s�OC�M1d��{��â�&4֍zm$[�<	cT��l�"X<�׿n�2p���w��Ե.	��$�O���\vl���{L9���k�^U0�nY͡�����P;�;��ӟ�|��O*�c�Ũ��0��$�$��ǱY����E칀��j�]"1��O:� �{��T:�R0�ªޠ�8i�����k�$>���O�g�B���(���iL�i��g���]M� �����g��vA ӽ��^�v���↊�z�X�����&EZ�0�$;���%�<%��dutL��ca�h��qh{��ob�C�z���@G���.���~�{���k�b���I�m
�#���iX3I�� \��j�iKf%0N؎�>_ ��aC`�W�4�Wj6�uI��-�����&��J2�=ƈ1��T!5�t����Ϙ��Ӹ0tp�7���7ŎL��chʋ�T�J/x7���A:�a��FbK(��<�� /�J�˖a�nH��}s��#C�<���;S���mi\F�b+u{n���G��M���y��lm�����#1̠�G��红�뽟i��R�;�^��XK1.^�L��g��k\�M8AN�㸲{��|��{�nRf��>F��n���V�w����D����Y�k:P� P��u�q�\^�;�L�ͤ�n��%vD!�~�6���6���z��їؙi��Y�A�����C�v������[R���D�e����7�	�c��P��y��m��\hO��E�L-(�{}5���-"��Qt�!����}�u����(H8�,��� �N����1%G0�d�,q�C��lϢ�h���2@�@�cF�!�������A^���"�����L1�����2"duL(g�����ɝ�\��g�!�Z~g�����b�	�����<��)
]��+.4r�`R/��?5��q=�{ZS&�1L������������ud6p�L-_���2%��4�L�N
R���HC'���?ރ"���#����Z���B�]鶷�⦮yA��7�!�χ �v�)(�+�ں�}nV�k)O�|N;�oƹN���;})7@
�����)�:5e�TK��L3��K�b�Ci�υ	�m(g����U���D�Q����H{��ė$��4L� ���}��K�|3��|<Y�^*6�"��P�1P�3���t;[�r����x�+���]�2��,ı�����"�D�J%B�l��V��f��;D�|����D$��ޏ���I
�%�@��b�|qp��O���G�y�s���c��l��<s�~�A��v".�سY4�/KzA���
��ߚ�ڲ!�Q��}m��}F4"�M�����ia?��T�Tt�c�Q-	��H��6�'���Jf$A�z�L�{����d�ft:�Kev�`c�~��N����2&�<z�u�K]�6�(��2
 8���R�{�&���BU��t�{((ȴB�;T`��]f'v��EHK�����H���]�8;ϙ�v-5�RJ��,9����7j��WM^�W�Ӊ�',ǔ-��e��] m5����m�?;�t�A��,㙴�#��>�5�pH�ߢ;�P��yL{�$QĿ���0&\X�fs�{�SH�a�'T�E�-����i��ݶ�WKsz+�;)��� =q��[� ?/�V��K��Y�Htb�z"�ZQ_��FJ��lB�9$.32ʀ�+����u�w^��Me����U��2���4�[���Z�j�[/�y��>B�'$"BX��,D�@�����{��NQR�����c.W�YZ�ߑ%/�&s/��ϊ8oy?aj��v�������D5q�ۖ)R�g����Jf��j��Ly�g�EɉI�Ӊ���ހs��4~GSܚ�*�MTZ�U>4O����#�ї��OLm|����Yz|�\�m�mmE"��|�x�e��3�lR���]1 ��p.�юpc$~��k�W�e�������f��~'���uyq��m�*ΘHı��_l�-���q.�w�򿺍���B�����o��'�N:J�5-b������f����^�82������R?H���#=�}0�Cm�����sfC�����ѫ�=˂*����J������,�=*Y�FpLH��̽��U�Z�r���nNC}E�6��BK��1/���e����zwj���wa�9JƳ"����h� i4�r�j2 K��A,�㻄�;�m.�C����&�YG�_��T�_�������D��l����PRS�ĝC�O�?�+v&�����>�:ųQ)z�k����-�b
=d����z���iU����n�8o''y��K���e��ϭh_��+�A���-`^�8*�_��ezs�E>�ښ��L|��.������ٜ���G]3�s�\x�e���f֕Mv�[����q�Oy��Q`���Z.b��v��8�1����(ؾ�f?z4��F��w�I����钹��������}*�6a?T�Еo�h�9`�o�\���/:k��Z3qYd`PE���x�H�P���W��G��l�YY��A�:����2,�Cc�ur"� Y����#�S�ɖ��z�[���v��۷k���R�~SP��|��8i5��Q���5��˥6-�ǸJ��bh��G��BO8�?�����Ds�!qw��m�S����u�Se�bo��R�9�K�w ٳ�;(sE6�C�N$��y��-SJ�׀��&��d�2�f����Ta����.�B��WPJ�������p)�Ս��#�_ yL>���xچz��K��\�ˉ+"w�@��u�#��~�l�;��`��>i���A���1�ע=���<�o� �у���ęx�֮��p�O������Lg^�tޭ��Arݎ������<�;�qk�#�i:�
���|toO��̤��av`?�t���RϝH�m���}�6�e�zX|Cf�f���+��@lh#%���F٧֓ߘ���%p�χ�}M�W�!��ɷ���φ� ,4-D@�(���NL���uQ�l���Qo��͒tL�q`��D�g��:bm�&�U��U��p+�$��
��	��$�7.��uv�&�܁B�|\1\y�`	\�?�Aŀ݇{��9V/�q�����R���WZQ��I����܁�����]�,�l)����_",E�S�T~���Dl��̍(��F��$�WHz�ݩ�/�t�"�β��f+d�cSU�S���i̝U���Y�S�]�4�ekOK(���.YA=
:w�?��v�0�?����a�_$��0>�D�s����u׮�KF�E�:�D����\��l��w����Bt�w�ҥ#?6e���@77(�*���$� ��'u��B��)u��l7amg�5�*�C�3��࣎��������c����oq�y�7?[i�o{�@������+�4f�7��'I6����:��HJ�[Y���\C[�F����[��UQ5���u�:)�+��6���Q�~������)�H��D���Y�: ��E���Ȑ��]!�SD��m���Y��e�uū\������d#gd�y?���9k�R9ʡ��W�%�G\>}��DY�o]��մ[Ũz87gn���{�򰈦~�y���[E��^�Ew������5��LsB
6k����WT����@x/�!I͡�]��9l��m�%X�Y4� ��������3���H�s�F%�J�/�B
� 2 T̻���8*)��ok(�y��:��l�d	F�0�6
�����R��OȔ8	=D=�RN��^�'C��L|p֨ ��om�y/Y�r4O�����@Q����(>�-	�-喎�p��^��0��W��S��"�6�^(�עAj��ݚR�)��2��b|JT�c�U�MD؞�M��ղ�^u�����ì����a��mD��4oA���R۵���.2{х��"Ru�K`�7�be&=	��<��2^v��G&4x��
+��lKq�d��Y$�u1��ЫC2�ȳRȮ��ܟ�����Լ��-� �8�����lh��(( H�"� 5*A:>�H	R�J｣����ނ��!t�#%��;!� ��$�z��}���|;�ff�5k�5g�f�@h|�����|��[�2�d��K�d�#o�7ת���̹
΀?;��3��/O��n6\����xI��p˶���������J���z���j�?�}��Gj��Ճ赋˟��I�"��_�'Tm+����m֥|7K�<��S	����wS��nx�[��x4�}�m��܂�2<_�
��u��ffE�H��!W%��k/I�z�k��J%.�m�%ʟq[��H>p��E���g��G2ۿ^����o~��a�ῐ���?�M �<D�e:���<���5L-���Du�{:���u��w��+s~���Z�.'L�K��0d�j�� ��7�l��� �Kfs�NN4hu=�t�^[ݜ%�f�.|ё�/X ��I;�9�r�+���U�9�,�N���S�ߠ&N���B��hV䨾$^�&�K����V��j�\�
G��}�Qj�[����Ȋ?)��wKd}�S\~��Y3:��5��a�;;77�C���p9�D�-�o�4gTBr�\�Xj��NГ�%f!V{��i��r��s����Σ"�*VjE�J�f�iK�N����޹�uY Dw�Q{$�|�x�gӠ�5jmPx��4�H��M�-+��
%C,xk���l���=��޾V
���Tr�2�H�G�6/�9^�rF��jJF8����ֳ���O^���ޑjK�@��LƵ�~y���S�[�t|Uk�"����ֽߧ��n���3L,�Y ���B�0�0�-|(���Fd)��	 �?˩Q�!u�IB.�`�?���)�ov��A����=�����]�[_QW廭����BN�YF������h����D檉�l���l�:�~���ו�d����\ZE�~�"��kYd���RA3e�DU���d�ef�J��6�L����������ZL����x���\�D�o�`�4��s>�6�4Y=d��1�D�c���sg�Ds�`Jo���=:� P�H-OZ#̺&]2`TүZ�^��H�X$y����@aED�������-�@�5Zb�d"Z"����3�%о �HcM�R�z=݁�\i���
�)�4WM�Pm�,�]#E�</�x6�����R�g�������x�lL����U�5Ʋ�l{M�W��E�iS��ʄl�T�@t
Q�d�F��ի���)
���~�.͘$���e� �)��,)B����X�^�R�O���g��r8��r����%W
�̺-I��E�I� ��=ΎF�^Sw���f
�_"I�C��GҲ�t-Y"�I{�i˔K#��y���n����<�e�q�U�8y�(Y����7�SJW�5��y�;�$����+\��$�T<k!k�7�v�j����c{�<�ͱi�?�������v�-yMaG8_Z�a���I%�vX�1�m��5��UwL�h[���G0��,�@F_�;���@�RN����5̶l�6���z��H5�6��͈�D�ה�W��E
�8]�w�b;��-���(�Q�ՇX�E��Q+�U�WFް#��A|��z�[������S#JZ�����b	s��A�������6'���,Rz'< %�G�H�p�;�8j����{�P�{At
D��*Η�T��d0k�=�
ˋ"	̀&E��8���}�<{�q��h���L1���p_�0�ܙ�.a�@�s����5蹋J/��,���`^% �A�j�>�I�!���a�:3��LحN����)�{X���7:�i`�Z�<e�g���$�<T2���.=p�>������q���B%hG̐����
�&\Mb�O9o�Ȯz���y�"�WxƙP��������gk��(�cE�Y�&��C�˃�Z0��DA�1x��_�D�k@�ǎ+'�D��AG$�u�(�p�W~>��U_tX�����yw$�S!�M6ؔN����A¡�(��F���	��I=h���am��؈Қ��X�g��9����a���X�&��f���+�8E0���K?�G���; �Wc��Ri�@��j���c�ϩ�_N������")��dBf���!k-�ٍud;;��)��[���ǵ�7]���J��m����=1�C��������Ҩ1�wr!���-��W������Ȏ�/��n�T�%�\pᅦK������'JsۿW66�*0�~[.�i��"���ދiG��4X�)��]�c���̧Zl��d���@5��&��w���e�.O���/�j�7�9�Mdh�?��<BP�#><����Y����ܵa�mʔ�6*&l�"�J/�St�v�B��� �t�T��n�ݑ�����IL�����S7�4���U��)���F��m�#��֬��=ʖ��8�箤�����T�c[�2�!Ԣ�sL�9!�gA5��@���GA���r2,b���}랰ST'S������@*��iu�^1W�!�8'��%�+j�
�x�a���"�ݕb2U/�IX>{>�{I�p�Zݖ3Y�Rի*���-��6 �Τ>��o�5Z�^�x����t��L�Q誄j�$O�x�"�-�2e��!��1Vi:��Sn�̤Vz��oF�bc�ئX�8��x.; ���N�(����6��~5^>MI}�NZX٫A`Έ�ң�D�Ÿ?k����7�܇3�B��z8w��-1�T���E�c�;NO7�{���#�u��,Q&&�_��7�	K�E<�%��b��}�z�{	ߎ���л�aC��k9�?��<�?��Od�7S�v&L�X:��+[ܬv�4��c@�3�>����5�����K�+���*eJ��I_̔~�AZ�W��
�XJJ�!���X�e'�''�K��Z�C�ŉ��^�p='��ջ������M~H�ŭ�,n��^���'Y��}�Ӝ׵a����M�]1&|!9ƞ@����o�q��~XY�N��Z�u刍�Ό	�Ẅ�$7A�sZ�J��@T[�[w��A]õ��.m��5���'��nc�-��-����<�ƍBם�L���rc/Gq�̧Z�M���쮝a�!�_#���fk�oE�~m��ǎ�M؅����8�U�$���B�Y�l|ME�8�`�H;�y�)ܑ�\]Z����o1+���1���EQ�m����0\ɪ�L��$�������\�$�[X@���K�a��m{nF��AEk��z��˄����{|MM�bm�0������_�P�����Mm:��Պl�.�p�&@�O���hE������ݣGDף���7S�_��G7���sx�Y�_k��с��! :~_�9k̥�N&��cT~��A�T/"GtY���1c���Q&��u��.Q,�	��rD�ڻ�T�����^�������4t?��R)7!�@��$�I!Y�{X�6&ݵH��ݓ�}^��d����JSCMQ�<��"���Z�e�wSM�C�V�j1�4���ҩ�fa ��0hD��԰����/R�*�><5�h�S�ƺ-��Ox{��o�ڂڋ�͢�Y��P�gA��`��q��R��vʷ����m9 ��؉���	j�2n�)��s����:���T�i����.��i}��3�D]0!z�Oi�=𖧰�l�1���k0|Y����؃� ���֋�ߨ>	&��dR˭&��}�~st��w%F[�9����l����u�-v���9�����O��oYCKj��YՏ|^�����z���ޓ�͛��`;�����&�_�cM�(Qh��c�����|5�_�e@@�4�)Z�6��Ƕ��/NhR� �O^��'��܋��+ڶWj������so�ZQ�k+*>�.~V)%k��	](�X�i#��<	��-��ɱˣ�A��:q9��6�-)�����<��v*�y�J>��~sk����&_V�(�5�D�0>�i�S/[!��o��k�*��1D��BZ\�U���k��J.v9�����L
�h �j�*����M�Юնfa��H
W]O��=�P�[؀g�)ָ5I)��=�:���H�*���*%��Ū|�㱱�ݬ�7�|�F]'����ՆO�ls/�˩��Cr@d�̸���Sp�%���๚@C��a����yy"V���K15 �on�X�F!�Ǥ�Sg�h�R��.�l�ø�W^�ksAz�E��+�aJ�qmAL��Υ���G�Z��R�PW���W`mN��Vmo�pã}��%�3kh0
��m؁�r�ӄ���L>ǵ��6&����ݠ[���x�xn�Δ C�y�U2�)%V�񁆌���%��E�2yVQ���I�i�d�^m�l�	� ߉fOd�<��@�j �o����{���"2&����	�t�*�P�ܻR�m��6C���8��DK��l�]1ͭշ�$��fV�l�R��ψY��7����p����F �����_B C� %�ֱH&�8X�+�SJ=7~��FLe߆���y��Xc�Q�hp2�A�|@�SH n��q�g��f�.�~�����'���I.i��gx�^�o�j��5��R=N*��}�Gf��G*�KV��Ѹ��a�D����E�o�!Cd������ý 3q�2��}n��6n`Z��B�W6i�񡛨s��l�M����b�?�`
:�/�;X�C"�^9]W��̈�)^:����/�Np��;�s��N�5����
)�������Y��xy�x�)��5PwK���+��Պ5�%��{���-��z��#�7���߀X��|�c^�Ģ0�C;��K<�R��ڝ����r�p{�"X�|SP�'�ug�Ŀ'A�u��IUI?��}��H�E�u��xfoK�O��E	�H�MҀdG�xu���*���ԣ��Aqc_��
E�?�j?j�����@� `K�c
��*p��W�μĲ�z�>�$8�d���y�r5��`=����Z�5XA�zZ]�F�y�͊����P��ђ)h'�y�i0k��I'&�U�F䄾�� �/�(%">��V#&��W���c�o�����_�]+5rc,+��F��+�Wu�kn���t�K*S\#�7x���3V�`Q�O����-USj.)�AO�t q�͗S����.g�G�i�c��y޹�M�y'4�HZC�{�i�˒T_4��Y��~g3�r�a\i@��u3l��*���s�%/�?a?>�$M	�uLq��"�[ IDs��W�x�Q+�����<d���E7����{�����;X�'|G�c<gN��./Z2v��As�qcᾞ�c�R�<:^��/%���Y��]=[��<g���ѕ�U�����M��= ��(�F�E� �p��[G�����}��IukW�K�$��W�e�������7Ҏe�pĤ���Ճ�������?��+=�*�]+g�)!$�xv^
����
�������n�H��Tmr�K�]~�%��{2�� s:r�+&.�
a�ɣ�F�
}}P�����J���+�Z�pN��n�c��*�~8�xj�O)�{��ǟ �Ub~LFHWB�2���i����6�:S{e�!Co��t��\��^�X��+Xb$lk�>8���k��m��FM�(T@ڡ ��E�ɍL"s�~T���e����m�ig��������-�=dÁ��XL�<4W5=z��ZO�Ƙ��!��%Ţ1U��r�N��qz��6��������t�`����{go{����IGWM���`�t����p�%T_B�����t��3:���xx�w_�v+�G�
����8�_���e��$py��~��=Dx*��/Y��k�mң]x�AC�;�$�꘧���2|�톨#���;i���!�ߡ졒oǭK��El0�� l�<�ȴ�}����������O{H�x��*A:_��b��?���A��S�����:�8.!&��ƽZb�d1
����E�Y�>Ŵ�&��6��l�{�e���W�U� ���,��ל��AM�_Ѻ��o�8oi�&�6H2�V��$���f�Y��o��9���m�u�u�hl��$��Kq5�����	m~�{y��5��cr�Z菖���oB�3�a�xJ�}�����L3L�Ę[������\�H|���G����|���[_)�v�fw����f��!h�A�n)X�9������&Y�B�x�@����
e����3\ɮA�g���	�����J�=
(�I��C������w%y�We/��PK   (}OX5r��W
 zX
 /   images/cccdd3b5-475e-4e4b-8694-ce23b104edc1.png|�P\O����kp���ww]�.Y�Mp��� ���<�������[���N����_�Lw��9�Td1PIP  ����  2 ���p*:!^(.r��  �_(����3�'o-/�@�3A �� �?�_��_�g� �����?F �����Z��������b�Gܿ�< �	����)�)%/��i�;��w�0PU���������������#���������o������aN�����.�#������쯩�^�a/�ZOY�J��L������Z���J���ZPC�ݿ�?3���=<\�ٽ��ټ�ٜ�l�9�9�ع�X��`u�u�0�aur��G����[�ٺx�:;Q�57�p��y���5�<����ǒ�����s@��$�l���ak���K�L�?8῔	������m�x���D��������"���nRΎ���	˿��-��&���X����6��_M�uA�����_.�v���f�o������\����A���z�����Pu��sT����߼�����
�����&�*���&�(�Q�K ��"/-��u�a��F�����jq����u�ŗ��S����!!a�����ɂ���zi t�V�s.y���t+�h3��ㆺK ��s�ѻ�oぁ��`ď��y��z5�ggg�̱� ���8�oFSk�۴,�~������Uy�v��qNNO7NN0u*^m�{N�):�[!wS���y3�����?��	[t���)[���DH���I�ۣhB�R�[r���s�U�Q����C�܎��E�DbA7��|||WYs���kMg��>ʇr���3!��}��������,���R�s�K`��.���e��ht�����mV�Y��Эo`����}�����h�����޵��3� ����^O^{�Ɉ�L��g[�4�cݴ�@�Ss�]O~8����gYVv�g�j���*�f�Ɠ3o�����c���ƪ���?��1�}t��K�P.ˏ8=�ݕl1��ǻ�;�ڐ>`��]�.w�NX�-����6W�w�~�����'<�昻.�D,{�/W�*)L�.�2�������kw?��=�*�&�p��Z��mVR��`�J���{�$�!���A>�X�2�F�Ӧ�\b4k*� 7xҫm?O�q�� ��>�l�ʛY�'�_�z],��8LMB��!TgfR�q�%9OxF�%�C��Q�F�ݼ�,��T��0T5b(�@ޣ�����6|�<�k���yzt�"n+rBSPnN-f��8O_��8�/J�Q�5B��C�����U6������
"���l�+i�І�!���R�l5���5:!w��� 2h�a"��-#�(w�r�@@����/)z] ��5hГ�c����o���ۤ���a�ۜ�T�Q;a.�P�ll���RJ��4�ق���틩�C�լ������h��N�+��ϛ�[<߮�ŉ 4��w��"�p<�8�~�E�/� ��q��6D�G�9"̠��N	3���7��&��	/c1$��	A��_�*��N�*EgA���^�H�=�oи��Q�!O�B���C�;<^ 
/x�$�����X{�!�=�8�郙���Ӕ�U�,A���ǛS�$ִ�Y�i��+au����v��JM�2;��z�\LT��3N�W�먏�i�FUs�Qz��"`~x�.B��py��*k�1d��_D<{'\@���Xr^{FoiA�H�ӟu�!�i"Z��Wḋ��ӥ�t;jG�|ɁԨ���a~?�\(��D���gw��jy�(�{�Q� ���G�יE��������8�կq%8v,��h��ף������^���@�/���Ƒ~�~���o@s5�PT~PX�؇��V[��`H8���SP��3�6�Sl��_��T]z��*�ց&ޓ�����
��ҺS 0�j?y4z�-B4����eI�q��MK|I U���Ⱥ��"�%�Y:��p,f���2�˔L"��d�~8�y����Kv�{7@(�ū�>;��������U��'��\��q ��My'��nT�D�i����b��^"�*3�� :G�T��k7�\�ČU(�:u=�!���Y�<�c���z�V<8څ\�2W�(���:J�mOpe����9�Yb��I$�d S?ù}�C�c� 	FV����6%%"�F��Y��'�����!/�r_��Ю~����[��:g�9#��R�%6w&��5����h@r�ySM=��Ʃ�LWl��6X��2��^��l2��(��f>N���z����|.2IU�N1r������;����r�s������q��I!ka.�d�kV*��0^�����W�v�.��!�u7OO������	����,d
�)A��i4�����Zњ����u�^vD?�Vʂ�_h��fb��#�8�8j��c(G�<>K���:Ӵ�Y��'�)�'-^G�X����%�6 /�	�{!�+3�$�:/S!83�
���M��:/c�$=I�j*xmgns/�ڍ�ܵg�;�d*�>��r���A���.���$��zM��tT�R�Пؚ�������:&��ϋ�C�O�]s�O[p(��U�H�B?�ߩA��ω�뾵�C�GS4�v�|\��t�W+�6g�J3�>p�g��B,�r�Z����B�Ƅ= �����{T���%�2cL T T�iC$ ��|���Q���8�C�$E:�����)C��r���������]��� ��������tr���o�(�%�|NgGt��e���90a�ׯL1��dD�9�t�_�>Y�5'ܷ��`�Hi���՟߳w>J�ՃJ���bX+�眉�\��YM���4^�Zj��R>�(������4��_7�6��7,�Y�W����t��Dl�����'���r�G��$�w��2݇A�v��7\�v]��P7`�tMc�׃.Ԗ_���yd�T����:�}���?�֪�x/���ǟn|��Ce5;rUt蚫�n�5ٛRu��W���d<�JP^�^�Vh\±��/:8i��:�t(�lpj�-~l�aa��N䟸TEw���5���dZ�|��i8�q���[ҭ6*$`qf��1cv:�Tg}�=��;P�="��0-�,7�u��3��{D&`挸�\3�-�^k�Bܓ(�ξ�W��p�Fr�	�WWn���H�P�'��f_w��|�^�ԫ<}�ť�l����Ou���XG#\/�kU��%�V|ġ�ub��T�>���9u/f�,;�R��ℳ�|�l��VI3s	�l&dT��'���յ�0�8-�I�=��D�k�[Vz��M�3�]IOu,��|���2"ç����]�}���S9i�D��p��#�!��H`�����AU�n�9�V�^-r7�hF���v��[Oj+����������X���+o�Л�"�Y�0���T�����@@��I9��Qe�?���5`��[�"��J��3^3
j��]s�]'AhB�x�C�
g�4�|�®)Y^��tH4�
 ],���M"$�B7"4��r�wid���1�T����v0�
zt÷��䐡o;�Iz�P����e���ԛ�CZ�F���� � ��^����5���C�����T�:J����g��H��� ��頧�W��ѾZ��Ş�ޅ)�a#����1�1li�7)���d]��{�(771�O{/�Di��@�5�^���O����}�h�*mN�Û�?��N��lM'��ג��#7�LL>B�?ki�I|�f(��5�Viؙ�][�h�.�BI��h����'�tu��F��vH����G�pQ�:	�X �����cp&�en��͙'f	�_��z�<~��;^�,�٪I����c�zM`_�~U��L5>�7C��Yj���u�6��M�++�me�;��t䋬�D��6�6"�$J�V{\l��	�~�0y��/�����g��.�1E���)
	$i�kJ���x��P��?�K�#�G k|	�B=%��	kXXP<W�5.���E�iuuՒ~h��XE��}�$����7R�� eL�7�8Ӊ j����w����f����T��1����2���x1��x��Y��/(}�E����K] ų�T�c��W���1�0M�8\+Hs���a��m��C��G���'�$j�+�;�.F���D��b����cP�ұ���������.�.�V?�+�EZR�|"�J��/�uѨ���ʍcKX2az���8L�U�/r��]׏��1���Ox�Sۨf��Cl
�w�a-��!:�kH�1�l�ˡn��sq���Q�[[�)�k�߿�[Q�(:d6��{;�)�Z��}�Ԝ���Y%��-7���J7vY�u�:l��Z��t�ޣ����Nf���6��� =�n�GkIFH�m�}���qd%ަ���g��:�;����<��G�[�ɻ�����hfe�(�U���r1�q2�+mi}n����߲��!��:LBD.ۂ!�L�̾+�n<��,Fc�����M*�0�(e����ʪdOl����{�Wz[�ޞ�?[s��Y�5�P3��oj�ҵ�j��X���w���_�ë�����?~��s�x0|�Ԅ�M���P,�Zr~ɘ����b�E�j�O^��{��cQ)k��8	n�g��!N��E�����I����ֶ#�B�I'���;-{27ɭ����pЗ��ao�B�'�p�ؾ�e����v�v��)\MbFs��&��U8:z��b遦K^��%�Y�ڜ6��_����C����h1���u���x&��� ah�����D9�^#/�">і�a��>��+�^^���Ѯ;pnBhh��A��Kw�Z�
�#:L�{a�r����TH6��QN=�E����Y���x.��b�eLT�X|ʃ3�͵��޴Fh)i^@�}o߁rὢ���>5����qwh���n�7=�z8�2�'W�qO�wH 5����+`i�Λ��9wfS�8���E�ډ%a,Qf�)������]�T���;���7�I/������K�d�Fs�{�������e#�	]R.� �R<���w��Ԟ��]E���po�p�ͽ�����	!v�'�D埖^Q�x�8��dÝ�VM��g g�L����L�`���O7͌br_2��Ų�=�V�C��z� �����h��p=�Ƃ}�C�D�h��P�� L�z���zF�JDR�Uyݖ�b��:|CM��q���W���O���^m�KR�At�s����0���򍯋@a�&x`�
_>��j������ ����)�wgUm�xEu|\j���z�r�LN�����O�� �kr�O�^�L�	ΈS���R�Ɵ_�޿S�{�V��	�ŰC��ܧ �r�dd@7�c�(fW3{=:��P$Zk�v�t�m�zΙ�]K�h����oo �̥�����;Ř��_W��Ωj��G��>�<��v/�乮�z�����a<
��E$����9-0@�yMoK�'�6'0U=�v	�D3����p:�7����պ���G
�1��9�<
��p�'�{���s�>,:�6���NM���j�%w��!�����ȧu���9���1��{��#9�_�������,��f��^�a���j;�vY��)��2�,�����K�;�2ϧ�ٕk#{�0d��dQe.�@�ho�6:�����;sE�TUʩ�Ǒi_�`��c��#Vb=�@a3H=v��<M9�yn���7����\A�TUImX�f6딴L¾�VH�D���iN�h�b�;���+�w��>�AS�$o��[�_���r���̑��� ���v[><v
9�K=�1��~2�(�~w*�W�����(6���TO;� F��Z�ۣ���W/�+�n�E��L 0�]W~<-Yy�A{_��;m���Se������E���W4�W�EB���P5����z#��,�]�Rk��֯���d*�� �!C:�!����\3�����C-�藥��eC��ި��ù�>D��%�&<B��%k���;��?�z�0���JƘ��,�E̴4q��~�æ{X0�/+燐�:���̰�4!�Av�A�1�?�H2�cx�M��^�w�vlT�6U�b,�=��+ܖ��wD[&��&Ѡ9%6���Gom)p��+�ߪ��R*A�K���,�[9y���ӱ���3S˟������� ��f�Ft����{���Cb1b�e����3u�I�v"�s"�����n�b���of֮~�l�K�rz�e���RAv�c�r���ƣ�	h��T22������+F	�#�C���
����*^7(հ���/�4d����Y�s����M5\�+/��&��"�}�~�D�/YH?��FGP'�0�t��ت`$��om�!:�^�Hr���쪉���=�SVZP��P�����jv���N�yv1v����N4kn+<����?;��:l���K,����3(��]#������T_���t�|�|�2PW��y~݀����^�������I^�hR%��6��o�4 ����&R1,о@����n-d���Rk/��2͝���+��M��.����r�$e�Y�z�V���Fw�/.�x81�@n<��Oz�M�H�̓�B����=5X�Cj��1���&�o �"xS�`��Ի���'�+��h��n��O��JM7S���U�<��&A{��t4�jܺ9u��ĽS]��XZ�s9�tq
M��)y�rm��k��f�6
��?9�QRR�;�,���y���s�����rx��Q2|&���K��A�nD���è��'�4�E?Kr6������f�O�z��}���!�:��ދ�Y��)�O�Jt��ch���E���{��������v�U���K2˂���<G{��
\�$�Sfbz��ʹO���.;��[)��8�?a�l�ݶ�C��$����B���c�.|axftF}���'����b��k��tݑӔ1h�9S�r��'��" s�����)E�~<W�Vd������7�引���U�i#*�t$�k|�vx�\5]�ǲ��٥��Q�GIN�.��g_弱��B� �1�"�,iDq?���g񋫔��ͭ��n�]8���\�w���P����G��ǌ�x(�\�y܅K�v��R(���:j�K>sd8YD8����$?���;��P2��<�YW�z�R�=��eF�MD\��[pZ�������m�3׫�q��fe�Ɗ忾�x��W#j� ���_�������'K��ޅ)�z�w��i��/� R�xk����_;��`՛s�@�~j���$������L4�;c�[���z���S-�k�	����'��e�oЌ�=�t�1Ar�}%V��禓���%7�P�)�ߵ[�tQ�GQ��04zk���V�;W��l�=���W n�G`��9�3�	��UYZ�y�0��)"8)*�ȭ��@ߪ�HX�ӄ��G!I*R%�,�NVdR�TJ�}���Sp��ntډ���)�J͒�֣}>�_�j�eg|Y����l��.�g�4��ь�2���k��+q'��6&���K?�6�=F~��D�ĳ���>txuijq��Y#|2i@7c�/�^mA�����}�x�#���a�U3z(��W��ETm�+/ҷ�l$�r�s��x�z~��h;�F?i|� �k���W*K����:}�۝?��o���V~�2�G�D�	�7S+fR��.�<L�0�_����Y%�j�}�h7x�~ж��:���d��4x�o2q����<�#�
֙"�p�?�3l�Zc���3����\dF�D_q�W���\	y�T��s�b�lC������M�8$3S
�E�ҷ�= �.jN�&��秲A?~q�%�`5;�Z�lr��������u��`R��#^��
� sv1חn�P\�d��XM���������%��W��5���9����ۖ�+շe�����-h6�Ns{��u
�'�˳1=�~V27���A��$P��ES�+�E��瘅X����%���A���\2��!�����|����y_�iy;���c��ӭ�qd�#5x���U�v���J ��Z�'���;mY:���A+B�JQ��(��&A�X���m�S)��V�D�ˍl0oe�q��]Ns%Z��\R8b�˼�:�@��*�'D����$�巑���M�� ���ӗ�5��\4]����w9�������xo�jk'�s����Y���nCD��e���D�a�JY���"�Q�aN,k�%�1����կ�"���@j�35�mU��f/xߊ�"/^a ��6��g����u��hW�B�p@1R}�w7���G�^�_j{�O
h�i��j�o�7л�7�"�2�@]3��u�.S�#[zj�;�wխ��uq���Y��K2�ڭW��hBf8���`��큐m|�l�c�k)O�O�d�ŅB��Kh�p�֞"D6���w@n��@6���L��y{��]�_���w�?�����Ϊ�*����jտ��e�B���.]�y�����:8�M/���C!����YaU�|#ߝLY����� ������=8o��0:�����;���2?3�Z�`@Q����X����N;���N|̷�^��!­ue��7˛:S�t����T�l�xQ���\�G2R����L�^o��{]4������Ht�:��Z���vB��R*��F�5q�.���ɽ�a���um���#�%X�������]s�w��m�Rݻ,2�r����6�b��y�1݅�xr�$`�M�9�&�48���,�~=�}hkK�h��x> �l釉9���~�
͖�)Z+����l]��zml�2R�d�>�k*3-"?_K�������X�f���0c<���t��.���?����Z^@l<'��y�<V���u]xn��H�l7ae�,�:���H,��o�E�З#��,128�xy�'�Yqi*���:�3�^�Z���m����*���ÞX��@¥(i�ꯖu�]%�����>It��'�*`X�ޒ��\��)L9fK%UW�������d�"�y|$�f�kie��f�by�7�j�kN�q�����G	s�w�a��'��5�1�F/^I�H{�_�Z�7�a�xݩ�c�9h|4��@b�� �g��,��[�V��De�螶4�r���c������etL���9�*g��"�?� ���u�L��΃���-(�OΈ)�%?2KQE��	%`�cP�����"�]��¼�;-+��I�yQSz��fT�%̎���m���}x��b��%,^���HR�K��T۔�Uo��Gܖ����l5�O��_��E���]
�0ԣʹLNVvsu�;
r��MRu"�)��"Q�Uo;l�ײ��\��U�!CL��}�s��8Է��x�I|E��͐"�c�I�YI=V��wB2I�Ôba��h��C�@#���y$a��q
�S���5�� ��z0U�cOe�P�!�+jؼ�p�)V3�?�4�i݋A�h�����'�J��T���$��?}a�I�\���ج#&��?��&G�uڗ�R����O�q�Ix9�Q�&6)Ö�D�K-��� .p]��rw�SϬe��]�� �^�^]'�K>��s>�#��bGoƻ$v�[�_L����I�E��ǄXa��{D�]����S/v��B�C��i��X���m���^�&,Xj�kK��>0�+,��%��6�>�,�`���(���	=�|�^�����K�$lB!��xc�=Y��y�Zw//�B��P'�^��)n�5� ���H��:�,��g�Xs�ș��B�A�o��[���p\����������$V1N]���O�rԊj5>lc9��]�'m��p��Sl#�-�I 9Vc������dqa�Z䦐6QFc��3G��;˃5���������X����R3a��T����/�ՙ�a���n� ^-E}d�Ud#4"�(��<$�E܆��J%C#��"���#K��Ş�K��W�7�n�R\W8Ə��*Ek.�>��h.^�H�Bg{��>�t�9���� q�AoI��ړ�'�g���(1:Ğ�:o�:����U�[Fw7:�jG���2~�Lk���RS���-)8������������	�g��w?��x@Æ��]fɖ��N�Ԍ�����f�	վ[�Ś����Cv���~ﵩ%�U�TU=2�|$��[��a>&�H_;��Nuq,Py�W����t����X����z������ů�B����~���G���̒C�)�쥲l���Yq�������`E	h�������6�cy�jjd��GL������rGX�ƫ�u�MQ�)�>������|� ?Q(s����3"D䉄�F"c/V�� I�ZUe��QS}���Ӻ!LR$�W��q�ҳZ�K��Յ��IbޝC��������^�G<���l3��1%?~,�(��<Rr1����N-��I!���K�������*�_�W5�o���.o���T�里��_���V�&%���f��g�9�O�{�e��^�B{���d�gUꏳ���	����E:�A5���2���v&ߒ�P��Y�k���6���4�5U>��F�~��e�I�Z#!Z���ͻ�L���?:n��b�&j�	�!��ن߄�6W��2���`�8R�,1�`"����X��IY	���Z�K�?TeB��0V�E���V,�K�;ݍ?��4�%U�r�Z�i�E��:��۵�uY@|��aA�^��%)I��Pn�)
�~9�i]`��X��/�
j�59�-�h���O�	���=�iU؍�TǦ5���a��� z>p������ñ�3����MwR�(ի�]��(� Y
���MmN,91�'w.�q�\�_����I!�0�"'R�mI��r�4�4j ����2c���)mQ�s�*�
m�݋@'-���*�nts(*g����-���'EbM=�����Yl�G�+�2�9��v�w�nl��oF���9m�.!��M��y�f��\K^<F���P$��JWߦ�%tX�=5�ح���f!�8t�9��N�r���d�;F��>n���{��10'�0	$W?�M�(������xo��()(aѩ5y�;��*�﹖+-C�j~��x�4�?]r����/^-�%;���Nt�����3i�9����_���c������jQ;��û���C}�1��ވC�͕w�FӾ�[C��gY8�O4��6�/�d�ݎ#[��A1S�����۴T2ט��T���ݴֵp�oTM5����9��0F]��)��bi贈C�=���gt{��F�9Ṋ�����V���n�~�1�Ђ���b!����\@j�}���|t����Z�9i� ��a���Ǉ�\[�"���:=�!�z����Z��K�����@f�)�o�f���>"�w�y��I.<I-���p?)w�'�wP㾭)W*M���+��������WQDL����C���t��4q��
/�D��E-�0�ʅ2)J~��1�i6=�$�{-��9)�ЛD|����#���qN`xnt��۱�c��B��H���>\`4:s1m�x������q,�_�U�֪�.����1�wZp�{�"DF�*r�k�����Y�1�dwx�����͌a���]S��7���/A�g���U?X��̛��"�cC� j��\�,.���F�~�>��X�?~1��o��u$j��λY,W�<��)�G�Z��L�D]o�C���n/ǘ�B��
?�V=�Hy2�.4�Y)Sw��L�ٻ�ߚԄl�9�孏Z�l�H`�E۰�����J��M���7�i�1n�o�F�n���ﭔ�׼AC�F�
��
<�9�40r$:fO�-�&���xߎl���=��Y�q�qM��S�Kz0,�K�I_maɂ9}�����p�I/2���Y�y>m�\���Ɛ���əG�Bf���Y�F��WO	,�s.�cۆA9{����)���?���G���/�T��b(�"�Xry��?��#�u@(�e���/��,!��hر9�͈wI�&��@���`�'���垈�G��u�z�3��U1�귆?�j%7��5\�u�m�]O �v4�IErKf5{N���b')7�Ӽ��;� w���(��%�,D�4sq�=�]���~�Z�)�����X�����C�o>,��>,��ڝ���
��u���I�j�Ga762���R�S�}��l��������|��[_�74MXG-F�ܱg*MC���>	�^�d�������(�bc���[Gl2��^" �v�E����S�q�%B����nޢY@�|�z��y��$���~b�->[�
V�����d(�!7��񛖼���v���]]���<x�'�i���5k�Z�F��,ʅrm1z����0L�J߶Z<D�2��3�/�쬮���Ez�]��blU���!���xdF����O{�ȝ��Ik�ϝR�v�<��:':>���}��e�u��ւF;8�nm�P�M�v�߽��b�3���L>��)��I�Kj���B�o�s���ː��p*�2$���ɲ�?1$l��<X�;X�x3�&m�-��ޯq�,��/��,�-8.>:|O+�"�>�%9:5c^��X��c�p<��W��gp��J�������}��렓�<�W�2l΂�V��1�_Th���o��C�zɾ*ݕK{��i�R�	_����ln�65��V7Ü�vិa�����Ȏ�(���[�Q��,�Y/��W����Y7�]�<���,�ͽ[n�����6�b]sYG�w�r=K˹��|xQ��9�0or~����m�D�e/����-L
��ZD�Ǐ�<~ب������!j?����9Z���32�I\۬|s��^k6�E*�^q�$
�
m���5�i˴�FbW~��/�`�ֲ�
��~�R�B���(�!W���
�$߮�J���:�	�)hz,����n�vȺ=�}�'*(`��c]f3����B���ys���� ��80oN�[���B�}X �xA/�b�3O�-Y�7Y�,��:��\�|ۖ/K��׽w�����(�.c�g�S0�\m|���{��ϊ�^�Z�
.E������Y�w=$�`���#8��$�:��";��h���������q� �O�(�����B٠Tl�AhY�ý$"6���x�%�4�_Z(N�\��:�Zҩ��%��U�d=n!�e�E��������/W3�F����ѷBﶘ`s�z�����]d��u};d	&������y_��ۨb�0�[�d�it$����R�1s��)A���Ǵ2�F��F�Ead3���bj�2�-���=��\(�y�ɤ�P�ϥ�Pjn����=?(�t'f�¸s(��se���<�h_Y=bs�S�8� ��ѫ|�mp�C�:��=
��0N�&���\#8�!<�z ���r��+���ΡNo*�����5�ޛ�Y6�ߪ���!�z+��;��+'{� ��7L5IJ��]��'���QH�;�*mi�Qf惡,�%G��s$xɌFu�������A�ڀ�|�����OoD�ͮ�e1ی�ԥ_�\��~�P"�������H�z�!�7ծ��X�A����Rn?b��Nmvz|�q�o4<��G��2�H�7�y���gX�u��[+��<%L�ŹvuH?��WMTӂ|Qk����e�U5M)�~�<�ϒ�BHc��)`�����B�D�l]��@.���Q)1�u�lw#aI�vo��-n���R�+�{�J��4|�|l��$�<)3�uӚ��B�5��	c�j�� ��u�%�Q�]�zy��G��W�=_X�S��ե����Vd��.�iI)N���/%n˲"5��c�Ʈ��/M�-�_\|���A�V����A)~��.�7��Z5��IE���p뷷���۟�z6����a�TswP2�]����EpE�+�;�/�8;݀��e�ɦ���Ξ��������V��>���KRrǙ
r鹁GE�
G�[*�|;���2hAbc�d���*i��g�0�9\����iM�\���7bY*�J�¶av$_����N���_���C�ե >���D�ɱiQ�BS�i�#%L����^A������ᑐ!YC�>^���&]#�|g�X5c����#���F�<%^n\/6�er��y��ٷ!7CB� 3U�$\.��\Rpv�y��E�l�ؑ�цc�B��a�Al��-Ҭ6�F��r��iY�[14]o�m`jxK߆�ݑ �x�*_
65������O�Hwۉ�qތ�c�䭾m�+m�K�X�o��,69�"�L]�6��u���4����ˮ�KE�.h=W	���4��@<r�fL߀q���(��_�ġ���q��Q�2t�"����},΍�[�p���J�kD]�b�/F�i����`�)��
��@�r�x��֥	��[�h�O�C�E7Q���;5a�:����� g,+���W��N�8�`��x��^��-B�L�����r. �;����)M��ч�Io(�n(Ӊ��:�su�P��J@{��3� ���&<��n�Q���u$��[�.6����䨏@_�4������U?�}�l��
�$ժ��e�yXo6�'<8�%6+cr�X�o�vk֪�Q\)�u�ɐ�m�Q����c�Iy{�Iܛ6��+�Zݳ�	S䨎֎��3ow�13^<�2�oh�O���d~�\e|�[4���I$�Z�rI��lv�_~]�,�B�d;5�<�����|*o���'�d�!�" ��,��~nSy�]a��ϫg&�dU1�+�����JY��p����h��� />�~kL��a��P;=�@2,��޴�+S��(�o��,L�y9���u3Ε���Su�zI�d�j.��}��4�Q&6�m����,4zy��<y�*ł�q�W��\�X�� �,�
��w�բ���p�MdWI�ʬ�)��?B�md�����?��D�)��ۂ�ͷW�2�h�P�63�$u���ۨ0~+��.�����	�k&��D�#�@)r��Χm|^6���E�E҃Ly�-�T��'��i��G��Ȧ�� }$ r�e�����0u�����R܎��2�S�3[�L�3�eȩ%Ŏd瑗E�洟��:���im��ˤ9��6�'u��.i:���	1WuDMQ�wJ<R�#l�D��෢�i[�� ]Q��ռ��vɅE��bGuࡵ5,;7�/��A�H-/����w�H�wǪg�b�����N�!�
?�0��w��ݯnY'�&�"t��G��dG�{���ɥgWRM���C���P�$��9F�Bj��]͙�[���@���*�p��s��.�$���#b�_K�`3���:Kf �`����>`��6}.
6�c�c�!��Q��z�1�m�X�'4�?�g��������0�N�ߞ��_�:Kl�������?��qUU�b�D�z*{���с*[q�wo�B��/(�&�[���������W��B���P�'`"��~�9���kB�QL��:p斶7�V�s�q��}y�O�pj��{�o�QKS2)�� ��FjMKI�P�$�r���6�V�O�ko��_��֓�Y��A���+��0�ԥ\&�
���~s�Yb�#&ȿ/\����|���Ŗ
w��+R� ��²�G|���]
e6�,
<�F�d��Z�F��2��9��"�?�������4l.J�đ�\���g�|��֎
X�J8գ���^���"Up�x�W�Ri�4��]z��[@
���G߱N�=f����C Kn�<���g�O��/W �x�ۧy��k{�+����{DL���'�F����� ޷e]s]LA�.ȷ��&U�g�:X�����nrץ�����k�U�{����w�e΅���6��p��Zi�갗����z����^dG�0' d�5�H��0�gg��E����=��=�Y�=�)�RpU�;G]�ş�}לlt�)e�HP%��V���G4V��,c�0�X��ew����������0mh �d��4�/��0C��Q�<t�)�n��ʊS�(��|�����7��CDh8��nI6�r��>���ݺ H	�u�����U������:[��ӄ�w����TF�K��t���&�BuNMN������Jؒ�Bt0���ceM�멗d��]E	J�A#Ro?o7a�uO��~�6W05$�м��pu���ج�Fo>������6G�3p�߶�f�����\�t�㲲�+2�+�%�f����h{�b0W^���"��N�a�o�'�6��{��%yX(}�8q�AO��-�LP�:r�ʥ�2RA� "@ݿ��'�6H�a�����'x��~�������wo�����ͫ �؆LA4�6k�c t�'5`C+�ޕ�45�T�mWpw�@+��?ï�} �3|��% �GX�1S�(��a�Ni�ݗڂ�m,r�Ƶj�+UG��`6�	xYc~��JK�4��ڳq�S ���0P�2d�j��,�/���y��+(��"�wZcd��tzg�:^N���$��	�Ջ�W�����i5���{xx|"[��z#*a�����GP�!���ic�~���|�Oz=!�Q�bHu�a\�8�*C��h(�]�|	�泏%����Z����X�5-�ijء �|�\�J�,M�xj���+��(��0T�m���7T1��h���kX<=�2�ܵjj��/e��0��g��JX�5�L�͓��2G.]�46W)�Hr�rӑ}i�m+9`�5m� ����J3d~d�|�����HH���봛���%���u�]+�T֚��HRaz�*N�^; ���- ko%��ܞܑ�F�圣a>ڊͶ�s���i�� Ƕ�<���}����	�����^�m�c�B�`�٘ƚz;٪:���v~�
޿G��~��=���>}�
_���	0[m�����x���9�"�45���S�B��3�D��& ����Ûߜ��^�c�XvǄ��t2H�)m�� ��f�x�.4��m�Q�< t�I�%��*-�z�7�2�|k;�����W�0�W1-M����p��5���{��?�1�~�������?X%��V�M�����>�=L�BrR��P�?��!�c��0�\[��k	��Q3�{c`���P|���2Wez%�[c��%���a*�4G-�����p�>_�C�nA��U���~��\���z�BH��nm<jm�y����rq����v-�0�zqW�����܄�v�ԛ:��݃ހ0g�ȉΙ�U��H���f��P�ΐ�i���⣼�uL�j�3��
�$�A ��m�"ceʗ�!�g��y/���>�������E�����A�ZD�:��c��Z*qg�p����"��j���2�_C�z
@����w��������3� lI�%�����L&�G������Z@U���=|��~��7����_~�� ؗ�p�
�C�v
�pŀ��g������b�I�5h�nG�HZ�M���`/_]Y�]��7���I�N� }"��؉K5$���T�!76g���
2�w�g����9�A�G������o��w�6r4n��n;.M�P� ~���R}&abk��g�
��5{xM��T�@�84�3�N�1�/�՗�PkL�! �d��~�ҋ���O���-�?E����0�d=k�Ŕ�^.n�z��nO��IK�Y����UB+`{%q���NA�i;a�x��$��u#�i^�tфfKZf��q|�ν0L-8Q�yY�f@��k��w�..��u�,�&y�y�PY�cd��Z�6Y��{���N�w�7��Iow�3��-�<�lHo��2T�WA�S/
�y/��J!�n�i�w�4�ī8_;�3�� ��O��}���\���G��W�3�z��젙aS%���6�M�vw�ک���x
~z\�]׿��/�ga�> ���'_O� �P���� 0D�sh3_�Ԑ�0P��㨱�I�<���$�:!��Cv5Q��ӧtm1�kF+g c}^��R#{6�n�3��"åg��mn=�����-�V"+;t�����{��Ћ�3�c�ܳ��VTA�����/���~��̑M >�����������_���R2U`�y��	B��؆�m��A'������,�oĶXdtԾ��W�˰��;Cj�oj6ES@����g�aF���k�o_�����>�N�Ԯ�i�T7W�?ލ���9W�^�nH�.�[�������x��fM��@��g�F.rv|��0���9	��g ����g��:Q���Z�gA/��+�=N�I}�&��� �� ���T%����MG`�~J��$�N���|Ҿ���#�!'~㘱J;�3m䀉y��S�ʋ{e�T�|9�"��D�����8��d.���^�A<�SbO��h��݄f[h�I���_`���`������k����khॆJ%t�j'd�cB�ww�d���_����Ͽ�/�~�란�y�쬛-n�Ŏ��6םz v�~l��I�+ѥ.��@d̘���j��C��g-���d�ؕ��j��V\���x�`E�>�?���w�s�۬gi�tU��ά�(Km�� �>ch�p>���V�&߭�ݛ<�v�;&�����#�����;���#�^]�r>���ف��i��+K=�l��\�H���4lŹ��m�Ԡ:Ǜl�1LS¾j���s1��>�cJ~��W{f��֦c?��0Q&�o��J;:{�r�G?���aj9*(;SI'
`��ӂ2G5�@AB�[��bo�"kK�.zvK�����^�z�
�֊�Xw��6e���Xr��ڰ*j� M���hq�ݑ�{ɳ��RY��W�"FR�U�1���h��H��f &9S}>�/�V�ju�xb�7|Vm�\���_`�LV�Kj��ަ�a�����̞�AT��]V�r`���#�L�:�c�\���H�	&q��R�Ė"�ڊG��H�l��H8 `�������/�X�o��+��o_�:I�F�,b)S�Y��c�#�������ߓ�ן� ���	������S ^�+�=�
t��m�.�����X��D���<�m��[�]Θ�46@F���㢺�)5��X�\���4d�o��E�Ҍ{39B�#	��"V�������9j#-s2^��*����t �N�Q$zڙ����ވF�\�<���!��A&�ƥ��� �q���n {��kh^����Z-<>>+vs}��X��r�A��56 áB��B��?}L�ؽ��T�߱�/�.�/�ynpuh�䫦2<6L����x�� {>�T�a'����5v�$3Gjf�����͌��jС*9�r�n�y�OO�zz�q�~>���#�S"�`ǻ��4@���PF̗�^$�P��؊� S9]�� !KՅq��HO� ��_���b�SoX�Śb cu�/q}�2Xk��.��d`��SiÁ~v	�|�OBK�|��S��zJ����nL>�� .�۞�<6�dj%u�D�ET�X�y#.@� �A&u���\����<`�5����߃|����������ܼ��-��* ��vbd�>����+��/h��~}�>1V��n�x\Cka�h�v�3G���n����	^[F�Ml@ѣz��w� 0{�%`��`7����5�IZ7l��س̚�t�D���{�"0�%��$t���+����������]u� L�;���Ewd��-�X����&�p}uV��qu�_om{Az�6:��H�Ǟtl���P\z/.�*P�0��:�:��0E�t�4�T�C�ƀL�9��1-b�T 0\��C�MaO��R�k���N^�{�'���U���a@� 	��pF��#�⹴I�|O*�0O�Wz�G�y�!��ս\^+�G�m�ڶ�7�p�(�C�B?�D�`��7�����7���v��o�,P���mzB
U�9��Ԭx�$�U�L.����,��܍Pjk6vO�XAmdLټRf�W��>��� �X��7�]ew�Sw�oc'��a�\*����~[H���AS���U �O����Oo�b��_����B�n������	===��/_�ݻw���A������l�xL�w����{���^ςڱ�u��m�#�yc�G-� �Rxu[����L��۬M�:�X�L��O�8f�r5ab�,�y��T�7�,��QՈ3N�R8�mC��~�=�a�G��ղiY�& �:�@W�xT����r;6,Tǭt�x���ȉ&���� �qW�H�E��/�.��z2���u]e��(���NNg	T��s���/K�B��ae�q���[�G&0O�*��`KY��z_t�of�Ź��UY����N���ck����2�����³�6, �n�G
�c�-*Q:!!�������+<v�m���_P����/����C���F�h����x��	�@�r��e��0���R����3*T3NX�ι��>Ԇ+�G�LI��(��!���< =����Y�Sl�b9Z�w]�O�C+ZENQW��w���䈦��U &�����(��]�VӰ;�F�X���p��A�|�ќU�3D�k2���[��Y���
����N�Y�o���|V	�T��0��_�ޑ���޽�w�?�����5<mZ����̍.�v�Ac�+\OD�<a2��$��+���
@Y,��dc��et�cj�c��J�D��e�����'�7t�NK�2���ܣ~R����<��=$���'�7':�r�u�51O ��6_�������~���Y`^c5@�{��i`D�)А9M6\T�W<j���p}u	�9Of��h����]�G��Ȍ)�Ƶ]ێ"�,�ɱ$t��y����>�3SX���9M��ä��[��(��o
[�*þ6��8���	yPF@�/sm�m�EnY���X���!��ph���@U�
�ɹv��Y�W���fml�'����ϖ!�' ]�{�e��X0�����®..���/�~�W�^ӎʧ�kx���ٻO��~��c �;�d�AA������?sH�@��|���=���9�}�N�4?7ʂ9Yt3�5�����|7V����?���I��j����
�>�"�,X�M�Q�8g�sѸZ_bk�6�H+�Dc�*0��0��]��ĝ��E��7N�5J���6y���3r��L�f���;a����~2�����N���\�,L���YW�F�_|}����~��=|���l�6��й���ΠYp�BT�[<��� �����B���#��r"�h���^��3Kj8]-���9�̙gufd��DPf�X.5�L���_@�s�D�S:�E2�v�wF\y���OY���tf�4>F`��tw�z�磀�e[dĴ��6��m�z��<Y/u0�ŕ�.$�&.G�G֧�����OM��:���z�����|ɅH�t���v&y��QF_��t����
�R�b�'K�7g�J6����^��)��P���uf����e���V�Wj�g�NKK1Fy��v~�ͬ��se_�{'���6~F~��6����&bw�5��2>�*�ɖ�iD1��o��P{/A�����������-\��\`����.�r9���+x��K�1��� L_�˯�?������l�[H��;Q?z�
Nw�"K�<"�I��d{.�l��E����l��~�6I.ʁټ�cut.������̨������adGGNm1�w�8���F�H�&1zM�i�8���+X�e����5_b٩mo����%xtq�en�D�\�P�UB��f&�[3�6t����� �cZ\��KN��d"nFۮVth�/��' 6{�
���L~�M�8^����:XE�����������#�!2��!�3�r��;)�ƒ����M��$��pAX���L@ �=O�]��}'1�5�@��`&����f٢�#,��@G�m�N��h+ub�����'���v��)�u0H��H���,uu=:���f��'�AYC��I�TS��
w��*i�����V��@m�B�A�`(G�X�z��ŋ��۟���+x��Op{u	w_��fu�f����i,2��}�8���1��TW}�����a�t��D���P�c��8�@̔|=sjPQ�<$�}T�ә�;�R��sf'Vg�քM&y���<�+dAJ����@�
��������>l���{(��d�����a�ˌ�'9�6�;Y�6l\�~�B~�8���s9�ps�^��y���t6�jղCV������|Y@Ъ�4�-Q�Ҵ/�Z-:qA��2u���*%�g3��o/�͛����=��[��Œ}v�6�HH�䵀|;R�9̲p_N6V.��Qumʘ5ed��)y���>˽&�ԋ���v%'�Y���D�0>H$�]���O4z�����C��u�ۀp��o�>ëW/���k�q����yv�U��[p������}�_��q�a����4����V�9#R;��	ڌ��r$k<m/@�{����v��t�c�)�~MW�fJ�0S&%>��՝ ��k:r���KY���e �a�p���>C ��A�x���8�tm|��׸p�mف)n�%w�ĳ�wY�ķ}����.t
�����P'='[� ����<�6aJ��߆��`>f����� n�����EG/cg�#��y/^�^������-���/���]�h/�抽X8xw{�w���'o�o�8�<<�����a
/��\���U���((��� ���_i�FT�L
���{��Ta��)��1B�֩T~c��}�~,p�����!�o���i
�u��K��/I ;s��bY�����:�[��h�EU�]$��!g��{���_�1ݫ~MI�kYP��&Kd��/`�N~����1f�S��p��Yo��q��v��5j<����2���h�����/�~u��\��A �Eu��\<飑S��1H�U$)�L��4VA b�� ̉�O�@Σ䇪{eZ<�\p,��'�?�`� ƺX���-��ܶ4/c�H�E�H��;Ӧ^n��/E����8�]�HSD�	�v׵�&G��z�3���]��_{$�w���^�Iq�7�&�ȱ��y�<ɜ|}�ə���$�ض�?Fb��ǯ�:�?��Ǹ��r��]��z�>��ۻ�~!�C �m�l\��ݎ�y6�E��X��
�S��7�:JG&���&����r �!����јk�XR��u�	eS���K�Ʉb��<\U  Y� [4�x�
�l��:T������D0�\�zBԃ�u�{�i1k0a V#M�>Y�I �T�0Z�|4��1 �j[����|�YQ����w���w��ݖ��ʃ�RGm�x���p�}}{	��[���: �?�Ώ�2�&m7OD�?=��׊������h��g4��'���kW�J)�O��C_���a?��}L��`_~��W_�S�4�l�N��	%��|�G'��;�H�.�O��>�.�2����	%�5�~O�h,�Pf�C^�QO���pk(��[�t,���b�6:s?�L �B�VB���=Ђ�b1�:��<:<\,.��2�g?�&�pO��/�	�$�����UՋQ��>��	���N�%�Z.�)`څI5O�h���0'� ��n��x���\p`Fщh�n`qy�AA�fb�v�ލK �u�z�%�]��t!�6ί7���\i}�X�ZE�J��P���ű�8�<M'p
|�K�fԶۙ��:��L���w�wd����/�gl;w��@�RQ-���x�Z��'öWx`�����_�}�O_�~�^����h� A���4/�T�D��1�{m��st׊��\�gi7�U[��L I;��:���h��ڸ�!�L��ҁ#�sd������������3���
uxV?�y/_����a��`u� x6<2>Kl�5�����Vd�.�Z�t-�1n�UƌU�h\ �l؂��AXxe��n�d�>N �G_��r�]�3R�b�6���U��62��uQ�jǟ������������P0\u^�U#������ܡ��\CZ�wg�^����I�o �BVl�@LKϦZ#0��5�|f��Y�4�ʰ �LӷL�|�T*�1��tj�*���9�(��7�۫{��4�ֿ�.K��?=>;����T�/��������Ӱ�	�I���Ga((i�@tފ,�2��������K���?�]�r�2 �9���%�ݟ���������	Pi��y5̟;:~���Ͼ5��L�F�D�	|{6D�i'%�����&7�pu�$����>��~���Q<��W�p�^���z�;X�9�?��7���nv���Y@���	,����w�U��uZn���"`$g3[�<R��K����H]����fxϘN59ao^v�&���xɖ�KY�5� O�����&T�0�].���|�c�7��x���� OFv� �����g���1_O�zܸ ��3-������R+KQcD	٪12���8�L���}F+���?.����@.�a���z��F}@";�$�GF��:��;��o�Y�W���#�Ce_]\���u��� ��s0�w��{��03^������Hgk@ю#Q�F�2��A��E@��0��|=�Wd���"��0�..f���C�A�$j�xĘ� ���^�T��qG��޼�?�����?���Đ�\�<��R�s�"�=�d����:��l��/U��6u��>6�
q)бA����>�k��+Y�S��l\% ����7:,��`}�<<������I
��Sɧ����Y��]�i� �+v��H�U�5�02���!�fB�.���Im�F���m6t
.�_����[X���_��.�� �3�S�x������j)+��կ&*�S4�/��z�88& �������<<>����>Ѷ�,ȯ��]�c(�e�6�4�81�wE~)���\�����.�ZzN��n�����H[E0Բ��6m�SR�=hS�
S�U�	(,�Ue��X��F��������a�r�y ֛��&��}͡?�Ǉǀf� S����׻{���+|�|�:ʜ�촨&C7�с�̤��]`C8�$#�X�N�O�I\�d�q��OP��ںT�H��2`���i'����qsVE����0I�
�l�v���lp5���}k�����va����-o_��Y =O��+��_���� ����h�$��_���*L��7@���C|WαM����|��ϰy|�HX�����7W�����1 B�����<a��8T�nB��d��������-����5���-��`�ܙ��d���	p��8`m㔩��N\X��>���ݑxd�|�C�8x��5�"	��i���)·R���c�������=�ԡ���!雨;{�޷<��?���K��3#i���X����"��Jp`���_=��\�6G8o�B�A�=>�ӂn�\�0�Ϛ�(���~)�a��-��!�A����sSXX������+r����F�s��W�K@3�,�rE�m���t����ku.2Uw�+�Q�,�2��4��ٱ��/Bޗ2W��ڠc�5� /������F��Xź�9�e�f;�fF�\|a�vmz��x1����H�8������?�*��D���cS�m\�����(����:�|�r��P0��=��y'��nM�]h��_���}� �5�//��b�s�%�u��t�rGtٚ�p��}R������B�);�c�u�]���H��"`���A� ����FA�IC �_�ʓI�(D=�+`�h衠�g%O��Ϳ^���4'(�u��i6���������2��j 1�[�"���b�J�ˎ/R�e�x�`���~�F ˝�=��<|��߿�O��u~@���� �E�,npE�6�ìC��Z+T>&�#x^Z��ؾ��n�%����~��_�%�|qC�j6�Mz����࠶�� ���QuNh�-{�W�A+2�?�gq��c�/��/*(T Vw'�vZ�c*��
��a�	%��c�l8�J���ZZ���1vo(V��ڳ/oC�_q}���m�	=R~l\iR��H^��ް��<�u�vn'�8�t�����d�c:�cȤ9� �b>�bP&��}���#�?�m��S�!�J-_N��l��r0q棧��:\�e`"�U��]�l�ء�%���V��&('�~%0��D��,�tAm�*�����Jv�ِgR���1@NkA2��e�W�֋���3G��	?��u��b "S�z��nb�V7jt�|�u;���1Ǔ0�;�|0���;��܅rl����'��z	�7/Cԗٜ:���������h{j�d[d-�@�P��Y嵘�J:B9�e���(&{�6�t�����4����M�Ҏ{3���_!*m�2�Ýl{��:UD��i�/���'r��� �F��"ӄ �t��X��!�Y��� d�!���\]�,��&ܲ�Y-�J��2�1׺�4}FgZ��{k��+|�� �>�joon�A��-�7� 
�!�Mhǝx��ҩq��F�hЏ6_��o�s�����W����':�qN_�8�Q��r!������"vZ���Huƪꔭ 0�ܡ�:,��'	��|<� �o�u\���S���E��j�mھvO�䥼������g���!�|����t΀=�~ӿ��g�����`å����鳹�œC�����LHZ0��kޡ�����>j��Wt��a���	�6��4�����׌K`ٴ��;gsqW4�1EO��Κ�H�bp���<��x�{b`
	x�ؖ��pFm.v��������1dȄ�N~�,�޼�*_��h�[���iW!�Qv��T׵�'ؠ�x�BƇ��LT�,�
��g�����%Z�F�2��~X��J�'?�Mʧʤs`�.b{�9��m a;2�A;�Y�" �ZC�̺�{_>{�Y�y��4�������ghZs>�.d���vA@� t������U��1|�'�-2���s� $�]"Q���,� �)����F�=�ޥ#�e�b X�*�XB�J厐|��<5��]qL8�zh�<�ԙ��\���g[���2���j�ػ6:>e�#{cNe5+A��ȼ��f�s�D%����G{z|"@�~z�N�\\���&�h�9�/�r���i�U �k�SAn-�_�ۿ8A����������o���4!aGG ���V�;��a�bh��e� ̊ڳ-"N�zX.v�rR>9�8y���së>���pJF�0�Fij������PJ��>������	� kC�35t����'�o�}�a���\���Ǹv�v=�G�ߐx�?�7�w�BD[��}��4����4jg�ʤݎ�f���V+O���Y��$j��U��a��3$i�Z���i��j �-��9mO/s�Ϟ�B���;�̑�$U�)l���	�;�f���lݒ,@��*44��y�
�no�uR���DR��LvQ$��ܥn��Q�K2ݳLb�6t��n�W�m�������.D-�\�b\����ݱ:3aN�8�f�8�#Ɲx7�~DSEp(�&� C���9Ո��^����D��7�-�`�~�w�C���qhV�����|���O�C=���f���74�:�+z��5��'*`�0��SH����P�À�=�@@�`%�Hm�?�J�ƝԶz5FcIa-�A؈��9�E}6�b��v�T��y��"W #F�N@�'��w�.)�T�����?<_
�,>?[B�%����gfd��c��40餩��F�ual��^m ����F��#�� �%P4#���/ޱq����G��Q5go�<$�/ܘzFZK�] �!��?���?�@;D�{� о�/4RM+^>�۝����`TL��s���9����m8�;B�S;�j�(|����W>�Z�{zR�������:�>0P2e���٨�Pkf���)��@L` �K����♹�'�g���H�N�c�t�e- ��鹻��-��ɏ��9	˄���-ϩ���o�����Wbh^�xA �����V�tr�L�Z{:70��ZQ�4�e�X?g���+��\qF\���7*�}�cW<o�A�g'��5�Bp����(F?e�{����^��#\ݼ ^
M�Щ(ʭ�֓�H2����HKͰ�����?2]� �|m�@PPXX�o٭�������3s�0^|�޼�8y˰hB�@v�2HF@��+�~4�/:�4F��c����܇��>� �+�A.����"\r1`&tH�*V��6�ΆT���<���{�y4 [��G��Ƶ���+X����;�X�(?�0�xf��HC�Î�-�CNW���mjT^J8qN��A�o���*��U����%��]@C�w:�>�+��e���^(���⑳Rt� ł]l ������@�"�th��/<���#S�d_���exa^������gV5����S���.�l �v#X;����wG2-�ݱQc�ZT�zsB�J'E0�>q^�z�_�`���Mrӡ@�����K'Z=rʹt*=�Զ��$[/�gٸ�����Ah�F��ҥT�PQ��cs����>a���Xz�Ʈ��[_�䷏Q��c-�ӪBs5�T�s({�q��~�r�k#ة[K��� ��!T��bF��Ϳ��93w��\��sI�F��Q� L���Y��8���,�w�F�%v�#�BS��cr2�6�LP�5��h�L��B�t����j�(GAJX�!���Qn7�V��]Y����^�"��w\��5��5� �;�wS��bަR��L��ML�HZ2��$?Pݸ��kѠ٤�����'�4>���k.��FG��'��|���$�W������K��)0�sx�,��\.ft�&�Ɍ�gG����ē��x�^�]�}�(��kwkxz| =�n`� % �e� ��"h�(�B���p:��N�1>dZ� �8l�gu(�G
 �Z$�,��J:uT �l���ֈ��	` ��'|�L@�ex��3���x�h����*,�4��\B���1B��Ry愒�p��5�޼dZZ;h����;��QNO+x�h+:y�^<�{�+�AFq�#�ڛ���f��"�yyuV2[x�}���n`{�H�g7�t~Ն<�o��ky����VO3>f��� W��no �� �ʌ���bɫGd�f<��A>�z�����j ��#�<b�����>	�Q�ݜWR�"x��1Pn�ק۬�)�����s�LC��M��S幌f5�Ư��<$-�V���Θu�72�|���?y��ӣ�vm��״�zb��ls�6�K�-��3�:&� �d&�@2�&�����5싳{���z~Wf�MFtbO��m�n��61���}B�4"[�j��ޠ���E�T��Ǭm�l�������Ǟ�[��(Q�E�Er-��z���';/rZ�"u���-�>��stt>O^��"�Ş��b��>�;0�k@|~	TmS�K������6��a{>m��ѩ4-�#��&.(/3:#�%��i�}	��^#���7�Y�wɒ
��g�=�$G�l1s !SWU�Q;�w�����o��<��Y���%R���k�݁@�̬��;*3#���p�~��ZS�Y���T'H�M^��X�\�
�/c��)HZ��IEVGB�����������V+�ǂ��J��ťt�U+�E���*���*)���(�Q����̀�?Xic���0eq2� L�
}��e��~�:�y�4nd�[�,��i��M�D[.���K�v$�q�k��SLf�<uD��ʧ�~S��e($��US�^ � �
+�����<�f��Ю-׫Z�j^�b�gP¿b=J;�S�!\�8��nK�#�OsN��fS��i[��2��p��=�k�5]7��X�W�"��{�ݤ]��ZF�����v��ʐ��5����{���S�p�ܣ�l��O�~ߍw������������AӉ��r�:����۹��I2-F�įd���b#\�z�DƒP�\nN܇����\ww6���h�NX�-/��l#�ò�t��e�:�[[���ԓ�q�.��2&i��'��0�[�*��)�� H�Ǳ��ھ�dB�c�r�M�jIasL����}�O�Z��8T";�To����+�x!�?�Ѓ��������%�*v�N��ɹ�L���$QUvO�бLT��?�[+ �m�L�ܛ ��o+v��.Ƣ�z�ُ;U*X/܍\E�H`� ���F�߄��@�b��)�Li�q�%qE>���ֶ9����lF{O��g�0�\f�7ף�� �&��^��9eiP��� ��{�u��5��n����0�PH�l0~��j,^I��nW�q*��E���L�:�[�}Z��=�e�j�q�6R|���y\�3>�i"�uƀ9�����^�k��j_1M�������z�؍ 	"a����M���F�u���Mh��{p�8�R�fĮ�/|�)e6Z�J�oٌ8V�o߾��"ĂA����O��p˃��k	������Ug���6�f�l��-�3�f5���i}��m�k��w
��[?~�9n�_r;�`�}`�Ê���{�Ex;��� gn�3�?ĮH⯝9A���Ȣ۹��F)���hd�Z�j�ūe��z~�������d��D�*�/؝F[k8٨ό�c	�qZ���ה.�1Ko �v V����x�O�UaInI��?�Y^]h��߰Z;C��L����R�kG�.43GYu���ɑ��]ڈ��K�
u-�j�wN.>�ǟtM'%]̧tqyA7ח�~L�
�E���ؕ�G՚ׇȪ��j��sq��=@R���`��$��G��Lk��(U����aJ�1�"�'���ƵG���ܬJ��@��#�p�:�m!�l�Ѳ��.����f��l޴�ct��0f#�tgd��gʴ���5-)�S �)ł�K�UpR�U�Z��V��pP�=�� ����tK�``G:�k
�խd����a���.ŷ�l_��V�Tv}N0]�hv��~��MB�'�%&�?*x�`E�*���Y��I�V��{&G1x�\�u� �=�8ǔ�i>~�:�����\@1z$�H4 ���Y1+bX�γ�U� �L&����fo�?�D�\������ppy��oz�v(F��~�����0E9�9d�1=�/�e��������{/���>�簃ǎ{lK�Q�}��q���r�Ϲw�5𾁋CF��kv��.S�ƕZ8��� �BC#"�Ni�1��,
%fqD`�`,��/&\jm����Xl��m396�Z��17]��4c�|���?���/�i�X2:$OK����U1sN��RH�jT�lO�]����F{d?�j�/��,�fͱ�P���p ^���UC���`�/f\�U[�x��M� ���X���˜��^�L�+��W�d��	|�H�O"`	�Ir�VI+
g�
���p4����k?>��.�S�=�`	'Ъ����m�l���z�F�f=��h�~F��r��Cƴh"�ϚbJ�z�s3����׸zT����i-~)��c��+Ѳ�S;�5�����_]�����Z�2P�����.OiPe�`���֩��Z���\�i���5Z�N�f��܄֞�SU��d�Z�fD+�Z��C׉H`��!��.{ �˗��W{v�z.6+�O�f�Ť�f��b~yI#�SV�v#�z����0Р5����Sd��+���s6��l�Xt��ȏ?�,��l�Z}p�1j��.8�}�p>öļ��xV�	Lӡc� 襌M��q�c�u��%�=�����;�X��Tiʔ��1���Ϊ��pM9��Mm��#YJ>�WfXU>�� K[�V���g^B*0���%�F�"'�\T�	ΌQK���͇�Ļ򱪊AۨF�c�Z�[�u6�ַ��e�z}c��0�[�Yo�?����h'����+j<�C���}��9x���BR��mu�!uaRS������:�mp��� c����V����ӑ���9�{sM_}��� �fv;r�=d��`��Vr�`�q��e@�@v"6|��*�&�����

�(���ֹ_�|#�DŌf�����~��c�Q����6ٍ
'�E����.)U�3m6���"�o#� ^,�ߪ�&6�^�F�*��\p�:~r��F^r_�Ȫ0c�l���S�@OY2 qj[-� ��ͦ�L�M��n%8r���2y�ep6N(�b�g��Ht�2� @�Z�PP,�����Lz�"�Vq?����l�$;����6��y(]�\��u�Z�ӕ�	�6���[�{�9U�W�0�
G�+n���KV�Ǹ�}�|q��ZD۾kZ<�YA�|�{�6Y�x��EPZ�l����EA�}�c�>���Wj�ks;������6 r*�q�|����`��uN{���9�s�x}n��{��0�6�ӹ�����fG�7�����3��*��݊���~-�e�؟}���F�9
���ߎ�K�M�bܵ��gm��5�;#	�繨��h�K��l �ƃ���s�5DW7���ǖX�z�)�d��]�A��[�~��x�dio9g�!����b�3��jP�X�,V������|_f9�ݲ@%�޼^dI��S��-W�d*��݆��Z�j����ftw=�7���Ż7��W_���5�C�8e�y�vK�J���*�{��k5>͠F&�'_�t)ml��b��̞��K�P� �4��.m�#AU�1M�]zyLꈮ.oXt�`ƺ��OJ�e�X��_l���E���H�+�d���-+:8|�h(t�,[������T�Bi%w���@��Ɍ�-���!�<nV"�a���D�JuK�:=�a���#� P��w>}����Gz|\��Ӓ��XmiɊ��d* `>wͭ9�Ȝ��m�p�	E�8�	��qf�H��֤r�)��l"hlye�O�����Ґ�i�,M�=*6e�.>�(��<�4����� �;���[�	�����?�m�H��Լd�G]5�����|�DWml��R�7�i�l��Ui,Z� z��E|��=�7��ꞵ�Ky��q!�E����=�����^��!�Ω۹���}�C��A�>�Ծ���\7�P����T۩m�w�S����=���FF�MJ ����K:Fv�����]7羶��1�1k]���P�l;�0+6�i�>��MX�y����j�Y��~rAh�r6�2{_���a~z��~.�ͻ���4 ��?����)�cQ��+�(��M!3�mk��6�h�+Xhmo��Mﹳ�@�{^ߏez����8>�V�w� 	�y�њ�X&�w(�1�mR{ϒA�����<7J-ǖ٭��%JĚSM�� � ��E������￦o�zK7�s������+����'��K~Ul�����&����F���8z�,`�E����CÞ0/�����yѦ�	�ͱ�##�H5?K~!�m:��/��:�:`�}���M�f�@� �,W k�{9���7���W���-�0P��͆kj©�-��X�L	/�����6%��t�[����"UP1�(H܎� ��d��ެ�j�
�1:a�U �>]��' ��'�xO�?|���%=�6�\K���i)������ٿf-�����O1�s��ZӬ*��U�-�2)>CZ��\�i�S��R�i(H������!�kb�,59?��A]�&��+�e����^`A� ���c�=v38ŉ�(122/K6��3b��E!'Xh�>��3<��S4�������D���sc��mǾ�\�a��>���`�wI�S�S����צ�>A�N��apOi�K�}m��Rd���n���]@u$�ǐ������u���׽��8��	���,<��*��8]�9�E� Tўp��M�`K>R����U��Ĵ�G�(R]����>�lb����p�6�e�0E�,{[��	��t�ۃlVFL�Ү^�u�N��Fw��"��Y�ϗܔ��X����*8�qS53�`�Fx�'�����7o�_�} �<`�Y�Gu�F���m��q���S&L=0��Ţ}�U҉��B0x!�2��2��X�s٪���gOψ$ I��H�	膔���5���;?��&\��-�H�ߐ�g,� l���9�������t��+��oظ^\A|l%� �)_,*.x�:L�g��T�$�Wn�F]
S��
�-�G5�%���e�Q���8��;��I���"Po���Jٰ���'z���V��p� �Zs��(]!�q�T"d���7�;�q@X�@��PS��#�!�,S|����)���Y�櫗���c$0��X2&* �yI����uQ�e�(�3Ɖ���p휙�T	����ዣ�ꀩO�ד��� � ���������BW2�@�ִ^�8VL ��x�]�Pi"�嶴�����ݎ�! {h�c���ɿ�R���v�ع+�Z�@X�c�N�[����J�~z���9�t�����;@]�<t��6}�M܊�͍.N�9�4@�IK��c�?ǓQ�2�0aH�ȏ�g��8��#U�6"�	�a��<�_��� ����h	U�"�$�ޠ<P\�-vq��������"z�қ	L��=��ŽO�/?d���fF�� �L-��J�&Cu0`-�	��a@X+�_�������%���_ӿ��+��7_����dC�Ⱥ/�X{`f����c���D���r(&wTL��yc�e9�ܐ.�}�!���I�A	�S��x/Y�R/�dO]U��%��6�8�e�|I��WtU�9.m�7��B�؁C�J�Я�s�_4� ��� �ް�)��" ����I!���a �}�~)�#ʳ��Y�$	�7M��DҁtX��gV�K\b��=%@�KTwT;9��e0��y8����ꊞ+� ����>�| #��EP�$`����!]w[q�.��W9_�� �_ZZ�â=��SrR6�0W@WH�NO��=є}���S��.�<�ic&o��� (N\qm�f�zd=���]���t`�pz����6�lVK��&��'��_k;�.$.Md�h�ӕ�m��c�O���� ����?����@�����>wv�vl;�����7t�S��g3��̟�s���t����������ͭi�Z��*wa�>�����r:Y
�%�.cX���Eb�ew[�-A��8��>г�ϳ�?b�d t�no(��i��F~��2��������ݎ�49J�$�QÑ��Dߝ_�^�e@__����}����������^�h.hF&dB�$�R0մ6���IX�I�2�I� 0������y!��T5H�f�\�3Q�C<_��� 0�~���@��Y9.��q��πpz�����G�rDf�+�8V�-Îwo�bv
Z'o�n�6�=�̹X'j�U�¦|r	h� �xw���qh�d�I�!b��Si��b��#�6N�%yaT�6,���>�Ϧ���r/�EW"�ф�*�woD����#��|O�~�}��O��~A妥�vM�f�n֋�%�%�W���ƓBEj��6�c�',�����=g��xKl��U���;[���� JH�&}�����,9Ĥ+�V��14u֨P/�f>��I }�Ln�B)a��c&�1\�x�. ��>k�f!Z
x���@'��'nΝ��Z��x�kr�ˀ�z��m(����9��{�������ې���J�*�O������K��s��$�;d+L9���4F�̹fN}LzB2�8ˎ���F5#��*�b>cW��F��S���l��)�6�ǥ�*Ջ�vR�%̗%egRj�밆�mW����g%�!��f����Z��[�K��^��xůi6��S�U�Cu ����Ajb6��ջ;�_��ҿ��Kz{;��ޭ��\��{<-6����1�lZQҨɥ�6E2d��E @����C�1�]_]Ry=b�t�:gnI#X"��ox�gY&������3��Q�)N��_����X����..�\�D�'���|Y�U�L�������ߢ��x��M����*���R
"����Cٌ�2��&��4ө䕡L� �*S��UA!�X*��4Rr�և��Zp��tJ� ����L9BL�
��"�=���n���<Ng��������އ�ܬ��+��|5sb�L���kSs��i��P� ��o���ϧ�O��A$:�L�H;{*��V4�j�����y��9v�_}6I�/�UA�#���XZlW_�9��$�Q�}�̅6·)�0��BV��=Y��^d�
�~�v�X�U�s�ldg�a�,6��!е�{.�����)�:�.�4ܷ/�/G�ܲ/9������~�5�}G�m��}r�/�y�����q����T&#�3`d+O#�7��lW����^T�!`O���)���Y7*q!L}�IE�$��e�ot���L,�`�J�.0��/�����Ҽ,�{_:3Wg�oo)X�����q�j�����՚U�QZ�#��^b�|sK���������~��[��z�UoWr�R!��-=-7\E��u)8��R�&9�/�풸�Zޓ,X$�m.X[N>�%2��A�\h�;B2"����Ӛ�"Urrd����iW�)�ۯ�����B�;�<�0�"µ-�D�>�SCj����=}�t�.Y���$�d4�
Tf�,�ѷ�斱SLI�--���Ix�@ v9Z����n�3M��K�AA��00@-"&I~�9 ���S��������& ��~��[������?��_�*�,��b�����K�*�����7�Ǭ� ��+[�ѡ-[��{*�C�v�!��´���U���,�(H��I]H��]�y�r��B�}^�O��{�{@��!�:�J@%�cS^�\q�`� 8�%6y i��8�y�\@l���~����c��s_,סv���I�P�c}V�s��:�\�ٶ�_��$K��/�3r�&�='�C��i�/L~��>��i%�DN�X6����Ə+h�+i����eXk]?ظBB&RhI��E֊�0QV�R_.��5 ��bO/�Ol�>�k���c�i���l�|-N�">�ˋf� ��uXnB��B)T����������&�����0N T��f�O�K������Y 3��*Ka � )g�= �b�˅��E�Xh<�%���a/�o�<a���"��V����x�r��2�� � 2���rD���- �Mg,E1��8ِݎ�Q�ߤ	L� ��[ֽ� V��hd�l[a�t��g�ՂSQ9M�lp9-���u��bЩ>	��ڪ���.i�]��"�.�5)+-Je�(����_�	�����K�X/EY�hX]\]���Vd���K��M�=��_���`�9gn }A�EZY�%��}�F�8컃��|e>[�d#|��K *CB����[�L�ug;ġfq���E�@� �jG�4�΄n'�ཤ�f"�x��Nm}Ǔ �#0�N�v����@�/�1	�;���8�R��\wߩ�����{�����ږCl���x�_�����v�{ͭ����A7n�蕞[o�e��u2+�%w���<5x��2%����K1��*�g5��Ѧ���=�٨�L9���`>�*�;���R�������.��9��Po{��9�e3�ţ�����*��_��7\�51d�OU!�,���-�+.;�Z�\L��ww�����~�o��r�Ux��1�G�i�J!px� 2����;��~���J!�1R�/�-��:� �u b��Gzx�H[�v��<T5b,�NK,n�3�x�C��E�L�u�EP\B�;J!���ꊮ�oX|��+��B.�j���+ ���W�ʿ���(k��VDV�YB-7 Tl%�$G�:i� Ud�ӭgV���ւ���$Ķ@���#a0MHݜ@�b67䂃����Cm.d=>-�f��Pz>4� p~PPv	�X�u���P6b����w���0=�ƒ��ɇ#r�ǅ��M�)��@e���,8>PC�}�OFg�J�s���$3a�(�o�˟�N`���Y,�ܷ"R�����K�FA�V�d�.//%��de�����Y��o�A��:��_>������c��}n�����)�\���<w���fO�>w{^����!����K��%wc0�V{\ƨ����:Y�e�����ea(B���[\��ok�ހ��0sf�$`�H��ene~����!dň\��:2��� 7U4�{f���`i��>������o�웻�R�~���b�t�8�,|HZ$�HY%⚎[���^�xR��|��o�����kz�����[)D� ���j+�~���d��\n��L���R�$��� �f�0���Z.��ӧ�����݂sT�	�	�b�Jfl=3h`5���Iv|�=O�s!�� �[�3 ��~>�~.���S��2T���1�Tb¬D�Bs�)�77����A"`�V��P�\ nV��YY^:#G�Z�qPȀ�ZE (I)5�z�
`A4	Jo��q^^^�;4֚D�D�t� �F�������Y�S� �Y혗��+}��v��?��RTޝfp�����-ԫ�qp�s��GZw��`Z���;�������=`�傴"&�M{��a}�:�+{l�Ϭ�b�bv���Q���T��]A|�I���p����tDUuX�oLo�=����5��\{Ζ/�9��:f���̾��}.��2K�2V������jK����A�� �A�%ۆ��> �K��s�����un��rs
�J���w��i��3�9��(��ܔ��Ъ�)'��*�ss�1e��k�"ݵ2bxO܏RFH�W�qξK�|�̇EA�h5��u���+�&<�4�{ݱ��ba�1Oݏ#��)�C�._駋�u\T � 3���� t�����w|}C�7W��Xo$�,�[]�* �1��� �*6a�Y%*R�h��"B��{���J����|z
�\Q�kZo���A�9�J�z��iA�`�
�c��^HTO�R"i4�Ѯ��	�S�>b��o�"C�2tJ�鵬洢8#�&��m gk�b�<A�:f�8H�6�n�Rg��:�������J&$��3������M����/����n�$�ŞGcU�o"m����V��h���˙,xP����i���(..r���������������O����,Y5�mU�Ѩ��J�(�W��\|	�;���X��u�Cw��
R�E'��������y1�;����l l�
ؚFj�����M�.}��UⰒ,�N�r�Q��Ve��s��6��X��*s��kl���Ţ���s�������k<��wj[��c���������|�{s�����P[�+V�8�f柟z�c�kg,8G���b���{�*�ّ��_��+��$[��:��AtZX��x/x/
��!@��v���8;�D�gAp�1Ȑ�(U�B��X��I�p�R��|�1�_#�)�d��耴v\b�3u��t��2���ʤ�~���)x�oL�lkh|���k�'
iڲ�������o~����p�$Ak� 
׎ �7�,�0��
�9�R���z[�+0m�1��R���$�nn�]���zAO�t��gZ ��|R�������͵�lNJ��(܎SӚ��OB��4B����>q�:�,���j±����%�c
�RkpL�zq��(>�J-Hd".
�jFe����5���]Z�����4�L�/�m\,���O�dW7t{���~ ��-ko8-o$ߗ�5IS}y��L'�?<p ^�)��zF��3�V�u=w�ٔ~uq��˷��aE�7��B'ͤ��'�@�D��zS�0��߀����e}a;P~ߍ$2�{�m����l�TL��2Lt��N��X��Ƀ�x���eJ�������-b�W<���Wt]j]qv+�ˤj�/�n}�˶<��z�>�<��>�� ����Hǘ�}�;w;��&?���k��߇|����s��}����kǩ ��I�u>[�Ʃ.{�b�}Upϳ��0� �OZ0���,_ٞ*+$��f{"�8S�up|!N^���*@2�e�h����(w�U +,���'�
�=E�F����M�}�қ{p��B���|b�WDb< E�a#A�H>��qI7W3��z����zD�CD��`G���,G���#�Q�p U������-�Y�|`MQ蛎J܅;�a�%:]�c�UsJ���$����w�r�5����9U����D�SE�
���@��ns�[��?*4�V)� ���3�Lo"
��8�*6��)��9���r�%��֧:]�֜���1E^ 
b��[d �t�&��+�_^�ݛ/���;�!(�-��"k ��&�K|�By���;r�0���YJƬD�Yo?}�V�x[�|}I���z ���;z
����r��
�%��U �-9�����v�ي�>���+��Œ킯���I��]� �V�w������b�<��BT�#�f�s�[��ɩ�%�(u�h�5[V��@T��X�hk��e+;V6nT������1r��I�s��yJ��?��������۩,S���u��YNn�K�9�)�mϽ�;1|�}�l>|�q�ejl���[���9e�39�b8� y�Z�%��ؓ���0���[�O0�m���� 1�(��Gx��r��*l!���TlVa2��&s/l0��.v[��1��*+����������N�bެ��V�����h����)��eı���[�y74R�f0��Ք����zΙ�����>�#\�B�F�L�1tR���)It`��$ỲX~�-��j~qɉ��#-�?��6����wM�a�"�K��I�u�1�K�M��9�1	i�c�i�ߘd�Г���B�w}+sc�N�u??8�S�	c���m����}P�� @E^�ܪ~
-:]�`� o:e����]�!��& �9#c�t�t$O 
���U,�NA�=?�L� *���ʦ���
��BF�¯~ ���~�3}|��		x0���1pX�� �N�͈���6�<1i��q��}���CģdOS<f"�\�JϪ�E�_\!)��]���� /OY�>��	:��c0�YFeoPF�VzK�9Hui��^gK���z.Sp(��P�U�_;%p�%�ƾ�\��F�6�[w(��i��w����c�۷1N��Clԡ�=�����#���8� WJ=��o��3p������I^���RK�U?���d?|�B(�f��w.�8�Zm:.�Y��5E	�k߰�>/J�mA�΃lKҺ�2w�!N��Ӓ��=��$2>h�Q�q\$c��<d|Ca6��A���sj6�U{�׻��,��Dc�D���	G.���Մ�.u�j4�8����ӰsaR>�	 � ���K���*��N ��� jU ` jJh��DL��g^��~հ܂ -6�5�D����ʩ���?4Q�hX�:::�g ���'C��(�n>,����ʤ��;�{�����(��A��\h����18�i;l�ȯ��LAn��87+Z>=�C4�r�/+c�$e@ۯ C�������~���.U���rE�vÃ͕E|P[���@Vl��R��+��}���G����1e>朘�rr�e�ɡJ�8� ���5��H��wWѲۘo�n�RD�1"3h-�vg��ee�ʪ�{f(9H��	��ǡ��؟�Ix�v�Yzm�ol�?�M�ڮ��<�)��P|Y��}l_lX�=�'��������ܶ6Ӹj˾�cch����]���`�6y�x��|�����cfj[er9�=Y��_��`� ô�BU�������HbRQ���w�PdgA唐���	a+� lPу�#u�5�f Lc�+QH��1-m�(L�w�Գ�7 ڕ!�e�)�W���FI0�O����W�+���ÎZQL�C*��业ӗ_|A�޽�� �.�&�P"�D%���ֈ�����/�}���'�x(@�k���*��K��Z!�H��Zg��6�� � _�j�(:q�|޶�l��e���n^�Ǽ�U�
�P��.3f7Fw5�M�!Y�I�?nRE%l��y�u3�ځ�dp�[Г
g\߽�
�@�QG#�_�Fc����]���Q�L��Z;ę��w.I���P�HRi���C���,�w\�j��zLR�]���5+���Tf���VV�g��������@���f���eY@ݡ�v?ۺ�IЎߑ�h���^�(�7z[��rd�$f)#��xg+�6]��Z�d���/��hU�%``��t�z�O���^o��Ow"��{�����4����M���K1�7��!�U�=�7�����S��)۹�����l� ����s�|���>q٘�b����ڹ(�m�aA�����\,��(u�P��AP:ߊQ�B�\��8_j�q�Sԍ" 0A oR�۳e�X�z�`�M~����hl^�N�4���i��<�K6:sף~��\g9��u���<e8 ��3!$zgR��Z)D(�t-�{��/,��n ���NT
��{*ś���f8=�+ң���h;�+U�<����"ܴ1gn�J���������c�
��Jv�����u��K�^�e
���=T.z�"N����*�j԰^��z�7ś:p+9�xK�R�o[��K-X��S�#�9Eg�sN|�2�g���rǛ��� ��Y����t�m��#���;ԐQ���rFon.��bJ��X�l�jؕ	64�A����z��K?:p���f'O�>��E��G1l�(����� v�l"���Z얳�����o�I������.U`0���p�V?���z�F�)Nm�z\�IT��%�>��ǭ�$>c�� }�V*��d~��8�H��yNp��s��^�j��c�j���b��?1^�m�/�sE�6[u�e�����k���h���:�?����:���kZj�0�"�y����H�$U�����f�bk��8$��;j�������_�hb>�H��"F�6����y�5����g%�H<��5pc4r̨a.��z��}��3���n@���Y�Ri'	}�ό���߆�|�h�|Y_G������ahm�	��E�p�>h����@���Y<ýws}Gw7oh6-�{�X:����\�K�#[�ǒMva�5:�4���M�vJ�a *)��َ��ա]ۭ�;��m5欈��@�<r�Hka���^ܔO$���Z\9Keή��K�A�q�?ʆ��#�u�+��B�e~t��	/.��&�v: �]�e�4M]	 8��t�\dW�W����0�h��v1�Q\��� *'����a������zZ?�U�,j=�p�0�ژ������;}d̝m�X��@��F~�2D��e\~}����B��C�d�dKH�s�d�pb�wI�N_��S��*��)Q��&�]m��e,�9�{(��_ bؽm��ct_�����f�۷�O���v�����_�~�dߍ�8��<c{��(|.�8��9�.���qM��lh$;��N`�NQ�|���:���3��@X���z�����i��O�q�w���V�#�n��e�5���2��Z����@�.��]O&����q_n$��~������	�/�npYJmeԐ,�\XW��S�v�epڶ(T=U�Iϫ�&�K��s����{ �k=�G��)�o׭�ϵ�v���|ܒź�)�� �4M�*��˫�`+�lgS-�<V�4�^�1�%;���X�'M�Y�����gD���VX7��G�X"�P,*)X�~����!��cѽ{�>�w*ڳ��x�gh��x�J�`�,
;�bW4�80�ǁmcf�|Qt��l,D�-�i�M#���i������QX�6�uZ��Bv#���n�Y4q`�햼j�ᧀ�R�88C�`����]��0L�5+���]��P�(U�b�H��Lp8ɵ\������H@��;|�BXF,^�����R�q� i�z�U"�J�����Ma��^y���^�V*��V�\��$i�j��{I��y�P:��]_�}����a��}�9���\WU�h��9<�����{�qOu9m�2v� ̡}Ni�9m>��r��[��в��}����1�����n5MU�x����JkG�&�`l���wB����
xi�	g�O��مZb���k ��l` j��RVₜ��]^Л�;�kݮ��\sl-����Н�=��#/� R�xߕ]��������Y�Y�R�ܤPz��9��Ŏ"��k����l��90?zlz�Ѯ�
�z'ө��݇���.���VF
�1�0�ֱY�Ι�U�R�;��0��ݺ�T�?�]�$~�?N��:
A��+sDi7���S�~�"�����pE�� 2C����#.4��ū�2�Љ`�sE��&X�� �n U?}I�|I<S�~��B*fMj�w���z]9�՟��1��2"�GZ
<�B@x�{��l����{�u�:;�4�ע�ը��d��.��ǧD��	f+l�n�+��V�D�������B��ā�����uv=���k�O;C�+���ܦ���R�h���\�B7�1v��oC������ש�Ɩ�;���4 @=��覠$g�0׈���$����PYx��s��Q'��H�I �H`�+�=�^pɺ��=�ІY�`;F��O�@Թ(/��V��Φ�N����b�H]�%�l9�?@�Bt.߽����\z��Xwf7�"�,d,����g����<&b ρ8� �Ɠ1_������x��ocޥ�w�̈�w������`3�XQ���%*����_��|�����Oσ`�,�~��O��[wjݣR�-��2�I}�h/�?���ݑ#Շr��� 6G�����d�[�!gb�A�[��= `��7�MC~����ή8o���a%B�(��)H2���z�흾�A���XE��V��6�sv\|�H�R/�.I�ql�ڼMnp-J�"����x��2y�Ϯͥ�b����Y���X@��k�slqB�����/��p�� ��)�����������6����s:�s�Ͻ���<σ��m'5󒊩b�B�QÕOZ����J�3]�r4�UV�I�* ����gf4����]]^�����H�[�)�h	ܯ9 ��%��d(�����7�w����3�ˉ���|�QAg2�.�FDN1`9Y)vg��0A��� U�8ϳ��1�.7�̲�6,�!	u$�é�$�_������ W�t��xc#���)�vɞ83�>���-ԫN�4�ʁff��B��[j���20��b?$������3�T�gn`�xx�;喇��8���$0^|��Q}z�x�24�2�t�(RG��삛�����͘��py"�|�l_��&��{g�9�/���G��f�������R)��t�|^�ت���x�'��nO�kM ��O�q�}��u�cTzz,�����)�O+Ɉ���ǠƋ����x��KZp���06,��"]���"[���m�x�����/��~���ޯs�j�s��k�q������Z������v�L����`���f,�ُ�}�驵����	`>Na��he&2�h˼#]P��Tq��Dj�M/h�چ�0BVd ��A9���:|W[�S&%@W�_��^��F�#��$�H#y]�J�"q9��b<z���H��h���ͽ���f��E���a�P�qP��o�۫+�ԭ�P��ߘI��Pҋ聿}��<�=�1�d����vh6/8YhY�2�g�yJ	k9�������mOؾ���cf�	�vc���X-�2~E��Wi�4�FK'�e�N+�m�F��+���)6faV�U������q� $cK�H�lYm�+"+�ޏ����\XO��'��zud$lrr:H�9�wR.����x8�e;0�T+�h
V~F�&d�\���[>�D b<�{�l*e8Ux6�G7�� �[2^}���gn�����X�Nd����S���¶��[���n�#��v<��� ��Z�����{n�\��;�,�nyft2�V;�)��G�m�P��#�^Xv��^��?�8WI��W�ˎU�{QbWm�Ǽ֠�޶�9�Bm]b���
�Mf�
��/�ox��q�ڶ���f�M˓<*��P��r��]����-���β]�/ �T��|�Q��u-��5�j� YX�~�����R���P���t����2�+����V� �"'�kv(�$XL]�����;K��N٪A��s��I�Ä�*�F��]�wq�x�fH9WG7�qw�dG��}ꍠ����%�w�(`x4O5Y(N�:~�{�dS��f��LM�Ym(��~g�귽� �<9���w�Ee%�=T;K��-��ű�4:�飊�� �jK��3�w�{`�V���ɤ�+��s�0���,�{?P=�Z_�j8�-��q����3��9_�\ʄ�o���G����;o��ǟ+K1?�)�z�}���������ˮ��~�y˫�!p�2C�_p�y^Ӭ����e��@gYu�7��� �Ҏlq)��j#���z�\�eƠ�jIl���A_.�u@j�M��cMka�:��l���2_��B�UD[��^���R��&�{'�T��B&%���v��\��.�Dd?Zu�� �dDv�V�=�~��r �ww�;n��Iz���L�*�h'�r-^mx������d���i�QC#�j��v���k� AO ��-�5��R�@�8���7�~X��]g<�.;6N,A����Ԟ@]�v���`�',��y;G�[��_�#��?+ș^Z�a��B	��x<kgz��Ev}��(������$��li�Z��@�#TE,��o�8!����f��Y?�R��Y#�.j��I�ș��v�����w�.F�;�/9�?���d߱1Z}��X�W?��v����#m���f�����:�7��,���m�ǅ���ީ�<=�16�C�Ak`��X[Q�'���b4�9R�v�����Ym
�O��V�}]@��jj�#���Ge��`�P�c����>��LO$V6!85\��0���ނ9��}���v�9�4s�%x�=��n�W�ӹ�'��_���Ok/s�D�bRsN�0ְ��^���R�tj��֬P�Q=KN2� ��'�>R��gQԱ�^4�TO�� �񲚿�Z�=�'\G ���RL��l��y����x�f�#�_f̴I��_g�n�J���AK��S'�J�H6X�����wo�w�T�8A�tT#o��Y�w���#�jz�"J꼗�����:�+^Y��s҃��\/� �keV�K����i��$k7[�8�x�o)�Ѱ�N�,ź���wلg�O���|ـ=��܏�ktmCY��a}.�?�1P5��c��a�r0r*���Yw�]���'��������|�s���q�R&5���{�����'y�˂����ii1𵆾��6z]�Ҽ"�L�9�B��QV�Z$���|M���bTe2�';g�Þ�$un9��B����2.2����
�e��p�`�A�����W��-��B�(z23f�����vw���PH��T-㽅x$ٺ�K5i^�A�޼ |�!��J��k��d�b��{�E|�g"���}���S���	�2 #����0�l��V�_X��K�w��V�&}�����������M;"{	���l���4�d#d����i(2�R��yE�Y3.�=d���kZ��Z��i�a�6M~�	I5������n�dhW�+I�kg�)QAy٤���P=���\|�}|F1G�Z��gS�j���ِuTï�@����Q���
�bYʤS�o�OtI�D㓴E'�#g}~��w�.���>7������v^��ϴ����b ����i�T��aЗo���y?��S��<���EX8��P�و2�V���5x,���J%)��q�T��5�N��o4�L� q(��7<{J�\έ?׍&y5�$s9Y�"N�ch�q  �:!^S��Co���XǷ��>�(��^_�:�Ϻ�ơ�/	��<�/�^ R�R}E�m@�g��vP82���7��e 5�����cW�Dlt�ɉ���[����rm�S``�8�Od��ԷD�Bc�H�1�qq��OA%{�X��c�]��k�'�H	��'΢P19�i�+eD�J��P{���$������Z��ʧc��y||����M�d"�A��j���|��|�(5��d�߷	���Ӆ%6.vL�+�6�@JC9���}f&�d�1��l�{��I����V�\���&����i6L7��2�+6߹ǿ��Cf���`����mǘ���c�;�V���s ޹��sc�'��m=�1���y�u�� @俶,���m��q-k�~�������7�J�o7.+4A𼅮��F>�3�b:�>N��x�B �qc@p�kS���0ϗ
�����FIfټ�JԕT;�s�gAY�'�2N�7	�V��H�KQ��9خ�Zm�i�>8��>.�S���S����ĦD�4�T�q�V���F��#Y��E�����
Ϣ>f�@Y��
K�ˀy6�"��-6>�Lk�g♅ۈΥO�L@m��K]荴٫����)k��(���V�[#�]ОO�_�0�� J.m3�Ad*Ŏ�����`'����ϵ���9�ՙ�� !�2Ǚ+>}������)��:݉_���ץ�Ůp�Cc�޳���8p�����r8�;�5�%yZyR�|�~�ܕ��T�Xu�ժ�2![��ׇ��E�&g(qЪ�k��������r��^�aՉ��Ę��&�K��2�ū"0>���{(��m���9���9��v�}��s���s��9y��Ŀ����N��q��l��;��m)��9�,�H�y��fK㲊$A{�l^��oZ~5Z7Ҏ��hU"�j �6b-���[T;�kXl2Vg�% ��#J��Q�$4�^+\�E�
�Q�&G���o#��Xf�:�@���W���� ���1~EAb\�s�z� ��c��ΰ��d2f}5NrӲ�|g�m��*|�`�Z���H��E,��%�y���GHNȖ����ڮ�a���$�b�f$#�P;lX�^2>K���TF���1pm��U�pϊ3~7[�tvϠ�SD� L��7f��F �(j���0�i�:�e���W���(�R����l6�}�D Ƶ�J)�$?KN)j:�l��x��H+�Ԏ�@��~dM�A�.�@^$��o�j%��N���f������tĖӊ�s�B�-ǃ�B��dQ�x�+���������R����6>��U�q=���$CqĀ�{��~�i�_ӅxjLӡ6�}*st*������9[�o�@�������^t����?GtAv��o���������r*q��"���v<V�	�e�I���3c�6֨�d)L��
�%�
�� |J�R<��A,Z
eQ�/�>z|Y,���X�����D1�ʦ�Bm��Tʕ8�/��Kݙ��3��~z��l�F*G�S���	5�7�U U�A�	��i4���'�D{�x�(L^�TX��DϞS�hw�����3Vr��$Q
�_��\�X���gA;���:�f�T��Ci]\�,�H���9xu�g��|�x) c_iM&�������] bl���g@ح�8��*5�v��M���.|�v �N3�Д�!����h�|HC$.\�S}��Fc�Q|�`�&
���v��[��#S�V�E�~� .π$]�h҃��}[�v��c^>�����պJ��0�Y�4�1[M�@� ���ۍ�/�
��r���|9��m%�1�m;�����>��N3/������3�`�ª������|�9M�6t�>�3ǎq��R���㿄ɲ����ɝ��3�e����Y��l�b��F@@6qomEV�S\��|�PRդ4`��ރ��z���A�0$rN0jV�����b���R�{��p�p��Ȇ��Je2�[��߭	!e$�6G�>k�%x2&v��|ϳ{/S�G��&I�dg�vn��sfiL����[��:�$��dˏ��H�Kh�	��Aol<-��H�P����I,�Nt�P�_�#H�^�h�\�6�0��){���F+���\�����J ��ԃ�}u[ݪ�@I�R��7q��N1T��	~`����O)^���{Oo�k�d�C��1(��iqe58�9%�ϝv �1�h��/'��>�v�P7�&<���O���==<.�����C����Ͷ� �Lb7���F�d1L���,�M������C�Yr��h�Q���ky�QtV�w�v[wFf�YX��+������𪴂���v�Z`n�J@W'�RFMn��6 �$>b����S1���e��9�ٱx�}��s��^�{	�x~_���9�����=�vj�ع��\�y��Ǿ��*���>�NF�����b|4M�P�V9��<�
&))�,W)̘I�X�+��لc�d.l5VH�-<z��6
�m����,J����6&c�Qm�kK̡�6�f������)�5|3��UؤrDV>.��>�b6 �a@���+M�8���p��� f��R�B�3h�Z�;�(�1���@YM8��c�|���%>e���t�F�����.Y�]�& ��z�6�����L��b��ɥ�C�`�j����$֊�ָ3��.�	�Ui"0�T��2V�ݹ�����p-mX+��.�k-ٵ���_�����8K/����������������5�R��`� �n�&X ^���0}��D?���>�?p����� ::�����1�
H Vљd�WH-�	)� �)K#����#ˈ�VS�]�{�e �+�!��	:U��aB��-�k*bو��_��<�Q�t?4-cAS 0�D�C9�I_/�a	�"щ��:mܲ��w�qݕ���q)�]c��<������<7����1�t�r�c�>w�RdD\��sw٘�L�S��s�}@e_��q���9'����w���ڹ�"�ݵȾ��13џ�<�N|�L���d2a���2L(i1� dH�*	��nuOB������3e xb��Vps���#�[9�B� �9�e%��n���<�{��Я�yN��l4����1�r*�+���l�n��z>K���~���Bg���Je���;�e����iMKzZlh��C"�`L��H�xڲ^n�����޼���5�K[ �x�A|���|y�t�6�{�\�Z.�����
�P��ضɶ�����u\1�� ^4�ִ�/�+f�F�)���pb��E)@^�W7�~^e�{�U�A���7>�2�������jj4}=�����׌��d�ؠ��D\�����r�e�H������T���k[�
� ����ρ�������;~�?.i1BvF@���+�Ta�
4��O�)��%Er��tP�5��2�M�`_�]�~/o\�DPf���u~�ɨ��;��y+&+}\�գM���?�e7����k lV?�w�����j���i������>�(`]P>�Æ�%ũ�s@ܱv���}��%.�S�qh�CqR����`��9g�S�g�����5b���Yn6Ř&Jl||��5�<�>af�3�Y�5��&�v;�W�#/�B��#s7�}�vL^r|�֕dCL
dQ+�)s'z�v2?��k��z�.5Kי��C�J�_�Z�G:�'k|9��9)o�e��6^���x��N�MjMԣp�B
�����q�v������n���< ������,!�k�\S�Z2#&l4��j2�rPe9�E?g�}IJ�P %�-��,�Z.�xz�s�J!@YZl��|1�Ԇ�!$㦭ų�%qI�QC;��LB��r��`GnӋ���K�.���$�����0�A�*������J\��~ ,�%�z�}�[�x��X������V
�*��q�;I�� #��7���Y���3�af+�B�z�00?~z����?���'Z��b��p��:1a�Ϋ�FW����1�3��@���@��ƢJ,��B�@�nW�@TA-R�լN��+���<C�	�X֏��T�F��z[�>�Z8)3D��F�6��nD�|i�a,�����y*���Tt�1��#
����N[B���fz��U��L�ˍ��!W��W��k:��[?�?wݟ{�}��3z���9N�s��0l�w��������j�إ�ҹ8��Fe83;�z��i/~b�Y����7�����F�����L>��r�r5��5���O�ÂkLA��͙��#�� �Vr�5�h�U�FTq�z��+����l�(x z�RJ��w�]�CZ�}*�E$��g�����	{]���IE۶��~�@��9��k���^�5J4y���b㚼W�����~�[h��4�����[��~CE c|� �`��^Y�׫��D��iA������G���� ������=e�]r��$����߰�E%B�ƓMg,N&���ys��I�"h��m\>��1�ƹ d�+�ǆA�*µ�u���Qr�@*'+# �;��+��E��ͷ���=�)�a1�V�\A���6�vDg�
/2I��bE?����������T0J�|��͋o�0:��(1T.�Y�k^���iBh�@����
�Yf3Fr,������9{PlN�7]��l�cc��l}��]m갊؄~Z��͖&a_^���/�,~7"��l~A���'8���3��,��W��I2�-�;v�k ����t���h�@�A�w_�t��9%^��9�ېa����L�/�����\����k�7?߱�x�%;�k�/_��|N���o��z�����mf�lb3��w��ٲyP���༸�`�/>t���+��y�-�ԍ�R)	#Z	���I[6�Z<���u�5҅�S�' Q�U��}:64�y��>$�Pfi�`��8QQT9���kU�2�H��؍���������<\)nN'���Ъ�?>�ŏ������	��>���wCfc���;mVl?8���`WƓG*�	'Dpqt�7 +1�[y��-��rA�'~T��XI���#��V�����mܵQ7���UD��T���Q�?�j��8���c�2�>V"�92���T�%��
!���p� �*�|���N޴XO&EAI��(J2�_��9 ?���7���4+�z���*�
L�HC��Ѵ���X�7�+d;���@}��_o6�Ï����~��O��:�=��y8���h:�* \��Z�7>��肰��ڀ&�m��,a���A��k<u���E|��qD����ZpUH��{��|���$��H)ˮ��)�>U�j�׎�J"4m��9)��oo��v^�T%P x������^o8��c� eHg�u5�I(nʾ�
�2��g�t
��{-;���ϰ�3�/\��l}Û��싫z�;��/�s]�/��>���Z�?�NN��KغXG�}��m��Zc��VH\�%�(���a�0�#�
���]K�a>�|z��7�����:�_`b�� x���mkq��y� ѳ@d��@Y���x0��z�ȳcI�Ί f
�������?�W�������'��t6��7o����f��4+�>�p�~��˴,H�lM�#�J��_x�!o"�R^�e9M����S �?qg|��[��ODK�)�zdƉ��L���2	��s���O�.��b�(dP3�L���
|����]��`���p�Fe�+�r#�?F-bq=Zn_F9Pb 4ƍǊ@05���7Zt۲+Y�-�:D�����;�_\������B�>�r��')��P�Da���X/�툠{fo4��*�GfC{N�8Y�{���UA�x�ih2�`m)vu�0>Z�����u�"�O�q���̥)V��[}ߴ;W���|O���o��ex�B�Lt W�P�����B��dz���t�^�-�r�(j[���G���Q�������֧D6g� 0*��czy�6s���WjWtC8����V���?����.&oi>��>X)><-�C�L&-MWkc,�J*7��x���dT2)X��<cK-ƭ��,]{�Wgc�����r3�v�ס�~j0���O�������$p�
ǳ��㞚�q�۳}��} _[C9L���=����/gk��Dd����ґ2�-	�҂O��$�۳��-��� �����P�Q2�ZzX<��Â�l�)yD|֗��?�Y�F�]���.�@��[h�.|��"����w@��l��
 `d�3��@�7Wa^�oh��mYC�;�:r�Eg�����ј:h4���������������~�3�5�EWU�4�&b�݊�1�@�$��D���kM�Z��.1]k*��o�U��53^��� tT��8��A�*?�n�U��(��V?Ҩ�VCp��蘪���C�Z
�O�S3�*6�����d*��� ���W[8�: lb�k�`@��z�����%�:U�?�s���_5hH���^�������/����3���W��]X�2Н
��"e���'k�0�%(�	������'�����_к���'.��ڞ��t@��4��� 񹋓C$��$�h\"I���*����Р�g�T�H�lp�P��TC�ivD|hI�����$7e��V�򰑂TI<xZ����~�7W��o�
 �*<�+.|��cv�Ng4	�Tk�����1������2͂l#�O��:�K��C]��+���G��Y���6���9����g�������%��N}�yO?�fֶVe�����l�Ϧa��,�'�)+�ր�]\^��5��Z���.������~���O߆E)B4x�ںL9@�T�_#h� ˮ8����;\�GqR0=E���}�2���b���,Ev��sZ ¡5��4��(h�߭_Q�U�Y�')}�ڌ��"��M�h�P�����U�Y�
Ћ(����	�����>q���?�Ѧq�O�?�/��a��Hi�s;F,�& ��f3�13�Y\d$`��a��]���hr9��Vd�#����$�a1�V�P+���`^t�{��! a$�+�9���'%��c��d�Ւ�҉�����-�/%pͨ8C�<����l?�>���j��Z(%S�Z܏��3�*M_DA g����2���s�NC�Z=1H�Â̅I0��@��l.�X0Q�W��y��zI��2���������*J],���ϟ����/��o����J�����Z]���&��1H����Pۙ���;����D�Q�4N��ie4����M�+��iJ14n$j���5�V�5V2_�g���[]pz;���� -�*`�׷���yuy��$-�!����~�f3a/��(cҀｬ�t>ِ
���f�y��*�w�����V�qFɶ!cr(��`�_r�۶��\��%L�k�6sDi�;�=�b��m�2^���S���!��T&3?�_��<-B_��>��{+3`�`ꅖ!�I�a��J�9҇�uD ��5#LG�8,)D����+���~��O`�|�4D�G�L���`�� "�+� ���b �Ɉ*o��	���)H�`��jf��Ӱ���9}���!��NX.H�7R��p%�5M��b�� 
 �e������?��o?*�qG�Wc�� ��t)Sh�5G-��ɣ��6��@\�&�ƙ��ͫ�M���e�>qD����R�Nf���`u=�d�|P
b�G+6�T���ӂ���̈Mf��ˊ��U5����h=��gr�?��O�dI��E���EV!�ސ]��x�u�B��p�uX(h�A6A�`0�g����ۿ><�D9��`�onni�< �7
-����2;g/���Kԏa����A'�W[�������������< � ��)߃F�3
#jB2ͬ4�W&-�]Ҕ�3�忘�yNb�bH�&g	a`�{�Y �-��Ŕo4&�d��By�����+�Ѯw��z�6+�wc�%���0���?=<�߾������+��ݛD�@.+���2�����j�n[h��,�ZG�	�	P�2��0�����?	��Wާ���nt:�Q6V�����l٣q`��c�܀���|��0�s6|0��8��m�oy��*�j�X-�	O�a��   �[��V<��6	�V\z�4O���~��G�k������62̏���,�*t�v�
 �<��2���
%V���n�8���)b��ZMY�\�xUG����c� ���1S�J��$Y�pEJ7f�mf+�̛��GR��)	��*#Ē=F��EC_<�����HO�`��\������Y&��qV�QSG.��+ψ��H$���l�|6ѱ��=jT߭�$1J׉6��8a����A��m|���b����ȅ�Ո��e��`&������z|X�����[�����ے��� ^쬗\{b��u�tppl�j%�v:gq;�D!D��*l��4�z���[		S��̘&&�+�k������R�ɂ���<N�jY�΋����ZD�P�ܷt9��V`"3�����?����o��g���?і 5�L�YhӔ\ c�A6�/�}��M�plY�m�@-��|�Υ;M+����*��0p\C�fK�po���|��..��b���(��u�WH����:Pb��J�e͋Q�om�bR$�<q�8*K�X�7�ӇO���}n�u Ȑ�@� �zj���&��yL�;�x�G���&�?��W?�/����+ oǹqR[���='K�5�O��u���2���!��s�H�&�>{��1V���>�X�ک[?��u�"�o�~;�s�=RiݜǰL>�N�����`�R��m}�m����s�v�۷��J�-�#����cX��@����C0�53+пRr(..��Eg��ޖ��Δ�ߟ���6��1e�C�R�U�[Q�"Y��q _�f\\��ް�(&{e=�Sİz�{��c���삩��9���]�f1�='+H�G���ǅ����0dl�����1Zz�uBťɽ�����7����x@�s9��q�i�wƢ��0n@Q�,
�<s���M�1��@��i}"���S�Vq���������@쁕S�~�7�ZpY��ꉙ0߳���xB��A� �`5�����_k�C�ՒC�у9Ǫ��Jk+"�	�����B�.�8�t�>��O�Qj�Y0�H�`�(��1�쒌�.��Fg P|�D�ނ������?��ǟ����Ӧ	�, �`U�w~M��%�Q�87�צ�r<6��I"����tG�$����R|�㰒������MJ�7��==Ї�~��Ygd�o��;z{wMח4��i�AJL �nж���eZ=��N{��*U�~�T��W���Ϣ�U��3uMAa��?�g�������K�gPA~B���_`5+�썞f��Ҋ�v3�D��Qy���low���\<Pn`e�6\�c��i��j������sݠ�f�忿������^O���~��${��7� �(���A��ֹ:[�-v-�p�f@��vMU4�Ŵ=��l�FP3/�!؉����)�-�k��x���o|}@�
�/N{��j��G���h���.8����1�� p/��h�*��ǧG�� �L���'��q,x������͕�Ѱ/�8ć�8Ūz���)��R�,#�".W`�&�8�,9�ކFl�k�=��J��ҟ��sh���xO�|uK��/��-H�vZ,���(�0�Z�9cm�Gޱ��BU��!Q2�9�J��e��
���o��'�ش�1�edc�R��n�O�j��Aűz ��̨�gg-���&�6W��-�~`���o8Pl�:N|��Y�/�nG�^�ڬV�=NT��
�'�� 1��P���ZW��B��	_.W�X8��H�	3�s[�t(�PPJ7P�9�Z;�]����} [?����3 /�_���1�ꑀ/���~O�`�B���¸���Ȉ�ne��O�r�6Ź"e8�n��(���j�+��̀!�t��D�22]�pƨO�
سZ��{/�o{Or�)vC�����D �$n���k������wё9��IF仪��VK���,�X�������bqgF#����̈ ��cf���`䫪5�������;�������	������ll��G��ͱ�9�,�qd�c���q#���%GT�l���z\�'�{!Hx��\�_�<�����i~ɨ��x��{i[^e�#�v�s��U@Z`JV}W�27�09�D%W���^���辡�����ǸgUi�AܴR$/(�-�??L��3H������������������y7�����˯�X�HP23܇�#�� Vh;�0}*�T���q����4�,Ҧ��'����П	 ����@W�+�
2�u�� ;�X飢,Q����o=hm_��Hk3�%���$����� `RO@��Q!獘�>�ğ��#���n�&�\lk�#�^ Pۭ��~�s�b�h.���M_,��(����՛ΡʁX�cF)`*`VFTǆ�IW.��gl䀠?{��sI�]R�2=߃D��Z/�RX	>����+v�%=C�l�{�ZAY�/�C:s�.�6���5�ч��P|YR��F����� +����$�N���h�xE:\�KQ'���I�ҍV�b���VX0<,������ǟҿ�۟ӟ���	�}�4��i�t��k�>�a�� �eڞ_��������Zf�|��^`k),�⃚�͸�%�f��ۭ<[��.��u\ηHP{��yw��ޜk���C�z�F2 #��� q`&9YhB�& ��\�/�G_ �?��Q��������������L���?�߿�1�����#�}�p� ��Е�tr�S,7�V�-l����-X��?�:�`�ͨ<��K!�\G����/uh��_i�����^���D?t�<l9�I�R2sL�L�3���k`��od�! >+7�@n�O���y .WW���b�SkI�܉d������|}���Ⱦ�X�,ǃZF�$R
/�O�-��-�M}�X<�Qʈr�䆼Եʼ�G�.�/���p�M��ݷߦ�+��ms~&�"}�gi�U��!s�#gJ�d��+X�'�,QY0��H�RsZ�}�HA�_�}�SVdχ�}:�J�noӷo����ޤ￹I�N�n;������3u��,�bu�т��F���|�� C����@�@(�e&Y
%��0g&�_ʨ�+�	(LG��=T�5"�~�壀LV�т�����A�.b����h
�����������EY/�(="����=�vf{%'���`�4.�ՙ�ф�B�):ѐ*Q����,8��k��n��.=L@��`{��_�. �?&��׿H��Ņ$qH�Ś�Q��;���+i��%�:4G�6o(�d�7Nײ��桟)���*K
mĬ�Γ�x^L��:R����P�.6�B#M�M��y��K��L�*u���v�ӡ�qP�՞}�p+���0n��������b�$��#eE��)m������������<��n,�|d�4�\M��/�S �k��_��@�f��\ﵦ�g��G:u�5�)K����̬����ёO�����5|���3���?{Q`�*[�H�ִ7J�����
B�$C6�ͦۨ������58S���Ǐ �u�:�0����*��f�-�XURx��W��k+�ldwmD�eI 
y��A���T�w���� 
�D�Or�+�WRJ$AnOq��o|@�1k$+�\�Q�қ���?���e�v��<���^�/{�Y"�"?!m%�R#�RC�.���.���>��E�~�͕ ��{7�.�hQu�#|ҥ��E�nPQ7
�N)xge0�w���P	& 3�#��hd�Y�h�,�� ?�9��� ����F�\��~��=j�����+���h����s����(��f#]�=u6Mҡ=��k��^63q�G�B��!��a`eYR�$x�X����M6d;M1��FB:�/��K,�I?M��_~I��?�����&����������	,���{��9�]�E�Zd�=��{D�=�ձP�3��(>o�w��TX��pZ9-[4Ŵ	8$�_�e[,�pm��3�4�F����F���X�$�WH������q���m��m���%�������	`e"�Z���F ��6�������#}��1��_�2-���ݛkIЋ� �m�iD\����/cY���W��
f/j��l��� a|�k�ݾ�_�c��K��2"_z��>�Sf��ޫ��_�o����8o�s�)���󩶜j�S��x�c�ґ~�;�M�d]����~��,���"�Ĭ��� �{�}���ӵ% 2�LPww�\@�`�ˁ�=�"����wA_���*-c.[է�Q�#���*��槛Ij�,'4�Z`��v�r���Z״����*�gڣ��6rm�D��/���@6�k�͐m}V�|�%i�f��e L�6Y�V;Q��ʺU8�DjV�l{;r�~����8��M#4}�A�������"��&]�)RA%��@��������"�6�LR����1�*,�%����ɣ7u(�N��c�<l��o-%H&si.:��W�[��0*tfj�����4�?"���R`�~���t�M:?Т��
n����9��kj�[�;�h X�����j�,i��﹘Fsr�(7�G���X/�M�^?V ��L���&���BѦ�@~��IY��C�&���v�b�)��8]<�Ge�N�V�w�HܧN�+;�T7�.�_^���M�LaRIN�N�c�gm7-�>cB��26������0�Р6r�7Xoa8��̐m��5H�"�sfT�~A�������n���ד�vZ@��k���	�|���Mp�1�	�n��G�)�����Uad[g�)����A�3���zn��]#����6z��=��+T��w�>/���W�Q*{Gm,�t7�����/ϣ�$�S�V�� [|Ǚ����x�����{�����0S �;.�S�������g}�ً�_����+r��Mq׵=[E��	w�4��n�#o�7	�۰�<L���PdŠ��}O䓕��Z��a.̓1A��^��<�0�49Rq����v F��'Žt (�d+.�$� *�?���H6��t8��� K�� ``�z�|q��:F�-֟��-�,mzș%{�痠	~�(�=z�H��l��r3��swwc��<$����F�WJ��]aޱ��v�q���2"ٲ,��%��/�F�a"�f6�XC�1 &��d1��V��X�Zq���w��6���N�W �-ঌ�H�\F��R��p�i��R���z�i����WI�����T� ���P�آ`���6�σ%�'�[� ���v��dqj��Y{{��Bvv�]{��e2!�c7����Ն���"e䫚��a�	1i�����is������NQ�g�!��u��J6mK����,]��V��y��|;m(�oR{q��|�>?@��s�f3��2: $Q\��)D�d��%��lL�Q��h�i4�H�ŉ�%��5�A�אԞ�HG��S��4�[ltS���\��o��5"�l�h'5��:H��xM���3��5L\�_pD!�:%�����O��CO�m��~�����a䏰E��-�ss��`O�0n�|��̳s�;���������ζ/ۧe�����̞W:/�����V���z�Q/;�:�_V`Uϝ�M�A۷��󌩣b����8��Y[Ȭi���<O�����-�{]��z��;��J�:˓�)Sz1i�̈�5ȇ��!rp�f��`"�L�=p��� dP&�@��c�����}��Y�
C��WB�T��X�!L��p/���$�����������K����������AX⯾_��6�"A�^��8�lW�����rfgN���  W�NQ�o�܀Z�]F����>k��o�싶hZ2�q��y���η�������	���}5����<��{��)�@K<�:�3����\R2M������$׺�Kͪ0ͽ���N.�̭�T���P������٭��0 ���4�B��߉��@z�a�2���p�YhViEc-��,.qm��C����zq��E�,���E���C��cRn�z&�Ҥ�H���d�WN�o�P5��mz=���09|�K�L���w@��d��"�_�j��6�3����,=L ��n/Z��@�R�c�0�X�p�(C,��n/Z([�P�i4Y�>e�$��b�$w��Z�S�����L��0�O�����tq���k���o���K FӚ�Ј���{�~_Γ/9�O������瀔�E��bb���@繾@��z��sL���9�$(Ku�U�&��ٵ���e�*Y�\l�
\k��:ٶ���׋��o-�sЕN���#\�*�֝�{��elʀEѸr9��E���5��I�0��47*j�$�j�����C��a:H?4�\��nϲg3���A��/���n�A&ɼMX�P������-95��$���D�_O
�"��l������^�NL�Ţ�P��`���CR�4k���?���l���í1 �r?Z��Ӷ@ƛ��������s��9�k�lh��G]��pyd�}+J��,Sa9��� -;S���w!H�6����m��{���Fj��$P�媻���L0V?h�:�,�O�s�NR$��]�kzF��~k��H`D�b�:�:Y8��zkI����*h�4��!��@�R'!�luВ�7��7Һ�X<���AɨJp�&ǩS���N3�Z�)w/l�(K�8��K�Y���.��:p����|kEQ��PIM皽����;�ϦQg���w���j�מk��+$|�h��K1Ck_@��Tc�h��9ZԎӸIY��"s���$Pv�xzV$�E�����o��ƒ 6U���7��!���&��1j첰d)��裔
� �?�x����k�D���}�k��c ��c\�}�v��8��x
T�j�\yH&\_v������#+�+p�:4q=�(���ET|*C]���,��<`���$�H�$��(�I�9����i���~���ij��je?�yL��� �<Yt�O����H�F�p�R�*�j��Ո��xy�Mk`&�ps}�~������r�;Ϳ��H����������V#�!�pE�@ߒu���̾_�Uf?	H�XA���s�n�X���%�M|Mr
�F����e�ehZ0S�/N����9qD{B`C��@om:�Mzm�o�yUe}�-XcQ��~�=�RQ���}*51K�j���A� 8$�H��#��DJX l�{t����\Ce���k0�e�N^Y'"[o�WC���tm+���k(��>g���:MV�kT��ʳ�s��n��
��, l#��G�^�:��l����h�Oh~a��	��a��19����Q����V�P���^��H�|#�]K�ר�K6P�{j#V��6�b}<r�1~ �`�_*nZ�ӈ�a����"Cy�w߼Kח��S�����ue|�V;q�<��4<#��kг���3��Թp_�u��R���6�}u��;��6�	�������x��9�?�٩�>�{l�w1���W�o����-��pzZ���]EL܇"CD6%-ޏ�Yzϝdr�ިם}c�o�ع	��qٿ��<>�%���R6���S����*���;}��u�wװ�(0g��}�2$�<��<)���J�~Φ�_Y���P +���F}VͣeQ���o���)W�g^%�z`�n�һ�7��|+���r7�]��t��AL�c!�WSv�R;N�%��9��Sl�{�ᘬ�
@vV�imoG����(&G2VM�	����9��lu�Qs�ֹRjf|՗�w�%f`L�Becg���߼�HK1 ZN���K�k�
 H��"�Z!�D��|��n(��KHh��pқ�.���3�/��9LSp��T�^p�Z�z0�V�A�ٮ8�ոc�	�V�`�,{�l��Ż-n82Q�Zs��6x4�40�K4��ZAh˂��hLحECh����9���i������X[RL�P��ԋ������fP`��/�P�SM�vє*����X��QC�(�"
�8lD�\ ����z�o��ćŪӮ5_-y����6����|{}�~��w�_��O�|ۥ�����l�<6��q�Lc�(�_H��B��`��ƚq�ױ��5GI��=y�i���آEޮ:Bd��ms��g����zKi٩�{�������ض%(�m�kPC!5�k������/Q�}�D��-Oϫ��RP�{���XQ���8�q�V|_����S�s�~�:��NG���AY���6A�pפ��w�)�~��R�\$���=�ut�W�6G�d�β��f,�@�.5�k ؐT�R[dc�PR����tuy&���d���Gw.9:w5���(�k�?�*)	\F0hp=+($����ͩ2`t\�l7�� @�"g���l�d�߫�E�5)�9���<���9[���6�"{:G��;^O�P�$��wZ�����&��v�@�m3������ܙ�p~d��qO_��k7���U�G�}�����i0{�>(��.�#��;�+[�,���Y�շ��К��ug(&S��&����^��H�&�-��H'�47jq���E��¨�0���� �,���  ��IDAT�+ l9��u�m�6T���j�.9'b ���i�İ����l��
��(6��(S��F �+Z���j^���j�YX��KO2h���N�����?�A��}�MU;\�N����mZ�M[���/_�3�Jm��k����y��W���ߝ��4����̑�iֆٙ+߯@�X?|>�/TO�/��ǋ�^������G�Y{^*'��ڮ%ċ�g�� eks��?�s�gf)���x�f��U���`�t�i��a{M��K�vZ���C��y#�.~��n'� {���$�iU�.	��2�ŠZ)u���*U(O�{�������&ݼ�Io�\M{�:�jh
��)
��/jZ�7�35_Jr�p��#�+���-/'�{�M��-��ю	`���<{.�!��"��ݻ�n��x�7Ռyv_��2f+�?����{���!0Z]I?���.�X�d���qkV��C4 �=��wC��v��J��o$g���;��A3��$��~m�E��ma3ר`���
фp���iҲQ�8�M��e��PЦ��_ \(O�v��JAY��.D��ˇ(��$[5��[��-^��O��*���Jwz�1]X�ЛϜjU���q��Lہ ��`//D��^O�$Y_cQ�E#	�Fz����U�o��(�"�I��i������;o�麾�No޼Ѹ��F͈��Z�F�k��b�cݔ~=�5׻R�������&f�!�7��@�uN}>��� ]2�W���6��x |h���'�k1�����ؿ��k�Z*Q�m������\z�PڹM�8�/6�L�O/)�����1�j��|����ZJ��)q��*|��$��1�i�	�6�f}���8Hj&i�
vU��:@��v���ۛ���	|�sT��O��k�������0B9���4��ӝi��X�I ��尒�d��9��F,R�w��� �{ �C��6�0�0κ.B�4��q����CRB�R�u,�j+?Qc��U&�`���@;��k�
����d�������vW��V,����I�B�'�P�J�IȢ��4�ʕ�XsĪfP$XV�Yt �j�L��ꘋ��!�!��s^X����2|0����EcW[�Sg�)ir2Y#7`iF���G^-Y�ls�=��9�=�d3�����&^�Dw�1�k����O.a���%�H-*�i_��%���<�hm,��S�Wf�����7OB���Q 5D��ϵ�UQ�L��rgW������c�CJ)�n��tR���
2��%���P��~${od)u��ɭc����S�����%��k1O�uXwp�l�-�wy��h�kV���}�;��x��>������y�����3~���|}=�.\Í�,y���TA߮���S��1[T"��#�!"{+J%�jJ�����RaMn�`~(m��dc��4u��/�ȍ��̍L���R{-N�Y�f)	DY�
"H�p>}��j?} L�F���J��׬�i��9c�0�t�2f����kʣ}�
�t5�d�T����lXr���*K�rbT�xt��Ρ���y
�[�1{�i�s�g�F����.���k$ˣ�2p��3I�ىp"�&@��q#Y�7 ^e���:��ޫY�ojd	��o�nL),�,�b��%�H��}�(��_0O�԰�J"Oc��]��XؖB��͚���0s_�ޑt�t�[j��9��M��(�cẼ��3���L�+�ٰd�W�Ш�R��fpֵ�%�R|%�ғE$�T�S}�+��@I[�x�$ l���h^����r��M����N����e(f�ծ��0����s�r|�αЍd0K�k�(��o?���_�P?W�;��6F'��K̡QX�k�o��y�A��_�{y<�_��a�V�'�']��$�W���x߬�Q}Κz�if�4_�=�:��J9�W,�*���SsZZpU��n�2����C��E����X�=�#ɍ
�����L�b�QY$�G�6K2뛛�tu})�ر6mDV��v��w��<�����.��	��fjwVI/����k�~�C��j�3��?����|A�0'��V�v���L�I�Լ�y�O5�ɏ��\��3.`"�	y���,'�Ͳ���2��{e��/5��x��7:��񹾄P)L[4�Оre�ʤ�4�e+�TJi�#�V#�S�IǏ�L��Z�5��?�S$���rvG}"l�_�1憝VBg�H��Ո#c��܁{.��qt/k��L�,Xm�����Ĉ�"9�a����W)�q�G�,��ڦb���15�0���?|e&�k�!ĵ�붖�+���s>צ\��g���5ZNb�(j��̓���qt�D7�i���\c0��������_�f��#y,`���:,K�Y�@*��-�C���n̏	���9�'��:u���]�����U^��ꫯ����S ���LD��t޴�%�%�Z~����$(��Y�~��ۏ����s�Zm�t��)�cؓzOZ]�m���
.��ۺ�H|�U��O `s?Q����Wvs�Y�چ2����n'��V�R�>�.�)��=W3 tR8�3
���iZ�d�R͝ŀ��r 6�� � ��:͇����R �sX�7�-�i�G E�Y��%����+�k�j�Ɉ~r��5�*y�w�� a�fSJ�K�\T+fb�d�w]������5��]L��[��ɷ�A�\��\(0!��A���ҍiLl�0�	�G�tY	3Y����'����& �\�4@dEY����f�9[1v`���"IF#�Tg��=j>�qo�ǳ;��Q�zq�B�k�3F��T\&�Y���lnP
XR���6b��p���i�J}�z_���
"��*��`�f{Lt1��Oî���1�H?m\ R��N�M� ���I_c����z�}-�}�x&��g_L����O\䏙�^c�z�=��Gʿ���l�ژ|MS�Sר���R�����S��OW�O�)�3/���L[�$�:�2߇~�K�>j���������t�p/����Ӟ5�w�[�s��E	�D0591r�Z��U�#��9I�0"PhQ���&tE���ϟ���>]�o&9�O�6�{{�~�ݻ��oH��Y��t�>~����������Ǵw�/����ӈowe��Y]�U���͈��%���7�4�533����o�LX̌�>�g���r�O�����jv��TY��GAY}���S�Q�;:�%x�IUI��L�gG�
��1O�O����*���p�V���6�[U��Q[���*o�d�B���a�Wm�iȔU�͊�kOU4;?n0u�W��_��2+�"2
AU���QJ�U��J�%D�D�#�d�|��}�g�Z[��� �"�R�I�%�T��xc�Z�#���!�0�ѐ*�4SZ߆�VKi�P zR�Ѧm0-�`K�ku��"8��ΰ�r�}�������y����S�ʪ����0��VP�7/�-˶����Qf��z�G���)_l�{V+^v���T�������<Z*i���G=k�9���9�嘮&F�%vÕv�^y��rZB��!=[��e�ZI�� ��a_��ނ���"u�T�$��p�Ւr期Jݏ���BL�<J���s�iw��u���7�݈Br.��I�m����|?糋���n��O��g$b}�I̎%m���1���9+e8��Z����l���p{���������Tgq9�f��r��~�����G������9~�թ���Nt�%��b%�j���e���:Ϸ=�~�y>�8�7�ֲ�E{ T��Eѵ�8SK�����Ɂ�d�/��-�i]�r�:* �M�-"�V�6�d5U�p�ڏъ%
&GRf�8օ�r�犫c�gڽ#n�i��-���������>C�¹t�KS�� f�K
������,lH]�Vυ��hm��,�I��1i��^�4"Qu��������4�v���q��������,�x��Y��.�ɕ?09]���|�5^ˢ�0/K�9��=��⛅�y>ߟ����~@���><Qa����Y�
`O�a~��g�$�o�f#^- �����x<6گ	�xr=����/[�U�f����,i�Xȧ�wF���d�L�~����t9�D�+5W�����m���h1����L��]��m������>ߨ�F��[���=���`���I�U~�|���������~ק����7�Ӊ{�
,�#%�����s�|U�m�sO�����ج+�>6Lnn��Y�x��؆����g�1��>~5��W%p��A@:>x3ѐ�Q��-����O��'1u���X�ј1˝��d!��k��ۢf�h�A_����	�7�g����,����(���G�4s^ ��R�P��|)�X|p��IC�Ξ��b�l��*���� �4N�}^·J�½�[�dG�.�0�Oy��pj��� I�Z��J���Պ3)�x$�+Պ���a�_aج2��'���v`^���m8��O ��#j�!���0���UZ�m�R�4n�i��
G9�����H�|���	A�\���� �x��_?��O��������r����k����q����)��S��s�W���3?r^:q��}m�����x�Z[�N+e����*�~(d�%�"��J_W�w���
p�0��ڨ�W#	�G�+9���F�݄GF(0C�:���l9����)����w@E������!}��O?}�8��H=q#@���UU
�F�X��"5!s"��s�ZI�����
MiيVg��{�kɶ*�o�Z��z�����r����=5�\
 6�^Ы��%-tɕ)8C҈��.�	�5k�Үi��X��D������FĲ����l妟 A��a��E]��4�f9�ŕ�˵��ɴ�c��[6Kp\����ԂQ��Bq���(܄�L�26��9mˎs�"'O��@E~��%엁�рp�T][M��M�6h�
����4[�}����]���jo�cf���
�������pk&}%#Vʙ�Wþ7S[�S���t@
]*|,��h�����Ի. �����/9b{N1[%>G�y��O9s�f���G���K�ȯ�w�܃�W��ט��`f�:���ʩ���̤K�������uʼ��|��T�R����5e���aX�+d�����i]��T�5���MU����2�� ��H�{�����P�f*�,�g�et\��>Z�ݦ��W�/��y�]�ߐl�T�V0,̀��tw�$���S)���j�FY�G�7�Gz#�a����P�h٢�u�^��2r�h����r������^�)Gø��p/�R-*���q������1�Q9�,��\̛D)X�R�@<x�a��v^�X�i!�P)|�����D-&�-��o-��ﻃ5�����v|��rNj(��]AD�̆�Κ��i���K]24͙�l̂F�]��|�GQC03 5�ƣ�E'u��) �C�c�/I]ō�W��(>��-H������$��\c����5�.�@��� =��R�N�G��ãº��o��Ȉ.����K���?/��[���4��I\���t���qa,o��{56I��J�S�Lw�m[?榆z>�S�kͩ����,���f*���$�~��k�W�O'��z-��10���c�`ٮ�8�����A��0��鋃l��(ο}|�h�_��o��N�E2w���n���yH���:�2q0�	�����xuC��3c�x}襩k�a![]��N���]l��&24�A2����R���g��<F�@�L�z���Ŏt@��^��՟,LMK�M��a�ʫ~�ij���|X�����fB��;:���*(b��|�^�)G��l��Ɓ���qqB�MPH�PQ�<�|'o[T��=�Pm[�С*K"��:�*6��@8����������r�J�� ���es���U�7ͨ���p���+آQ.�K�$����+��ab��t����
Z�m�v�"��!�VT{IV5�G6꼕��Z�Z�Q`�z]`��<X�0M�ޗ����Ic�8�r�l�6�F��Q��KQ7=� ApC�%Q��!@�1����S�_v���ՙC�5>5�r��D9��-y���R��k�󫤙�Q�r�:o����������D��x�>�Q=U �[� �?K�V�zE�?�f��n��*H�����)����kר�,[��k0�g�.��C�2�F]�ט� �ҼHL2av��6�n�����(�r�f{XN��O��1s6T��{�Bp������3�#|���5�M��	�#�U͹��`�@"e��a�P�H{k`�.Dil1�0�(2��T|��yr�E�4xb�,�@������ݢ�_�"��9�7@��T�'Wg#�,���l��O�ɬ�½�����$m��e��=�����GM
���[Ax�8��q�7⊸]-�\���R����q��/'_�cΧ.�'�H�u��W���{dQ&����^9�D���5�Smt�3H�G��GTFp�Á�O@�N��`����@���	D���&�o:e�q���M��N��Q�3c9a���VjS��T�K���ZG�L}&. ��M�iS1-e�<_{7=
3�J.o5L��t��;�)�<�zg ^R�?���֖d~��*�M�p^�6��lv��ww�i7E���6Z�C�0��.,u��Dפ��'5s_a_���.��4�i��7Š�M�3�x�X��jY�>/�fVA����<��M��0w�Ǿ���9�۔�P��������Y��0h����Z�q����5֘/3	L���x�瞅�Ё������b��;��J�]����P�`��R�"yԯ&w���i`��u�#�o~:=���\��?E��dso�k����Q`�ť��8�Ƣ��}�HME�x0ߪ���vq}~na9W��S �)�>&y /5iy�YЛ�4�l3$�	&lg�/���Nl`"{)��H7�D�&�.�{�;k?4����x.��
����qhMb 7P·��k�\�Qx�<�&�>G�q'�'��~r�h� �֪.��B�|x~ta+ x�&Zo~F�>G{����z)j�6[���< 4�k��A� �CY[��
��U�����8�Jd4L�9shrm�v��f�T������PAg��%�bw�8�:L��̎��,���s�9��./��(�6�XbS���aJ�|靴,��-!�:��]�]�ϧu�K��%��Ç�_~I?|�N���b����"�z=<3r���N~��T&<�c�k�Ǧ�/9ƣb�������Hs���%�Vk��<yɕ�# &2$Ο>}�:u��B�����f�'X0|w��F��'����ymeEC����Me" � ���i���>���'�9l�8^j
]2n����N��L�<L���H)�����X�(b��o���q`�p �>�g2���n>���P�����'�Ɯ��Ƨ+*F��d���ߎ�z�%���#���  �Feױ'e��v�#�/��ɤ�����=���Ӿz%��r�3|�k�$
�D ��C�'S��k�,�~�UU�Wz�ʑ�Q�ɀ\ͧ�T�������N��!��d���YP�}�/�6+�rL!k5MQc�AV�j���|}�W�7L�Cy];$�\%w�����|�����s�+@6<Cv�5�_4�����-D4��8�I
,KԮk��-���ɆI�)� eV�]��w��*�J����M��������9\7 �DM"��!�K�O����k�p�e�/ލ9���s��~j���݋L�)uD���������a� ��2>ZRc#̗ܶU��A�Ӄ�R���&H�V�	h�q�J%Oe]IlX ��+$�&	����?���o��Ȋ`*X	�#���;��%���:'|	.-{�#���$6�W]�o�"�q���{�?�.0��?v�k��^jj���Y$c�� \ paޅ�����猀s�xZ�>T��<��������U,��7ZL�����{eT0F(!sw�n'�Ť��>�c�Ϝ�#��6>�:�R�v�Yc��4�=�U`�gy��k�;c<_y�#�Ahd�������o�_�����}��"ne����gȾv�2G��u�H0�b�B��%$� L�fٷC�5�@� �����4&Px^�{���
�L�VEܬ3�4��=���,�sL{G�+�2,�Y����>ޘ�ENV4���`�D��m�J�"�<19Vޜ�+ah��q���ݧ�u�>�z�9`�dh%kNU��ҍح�e�օ�P,&�z�釸Fk��8tf���2Xj���ces��Q�Ń����Y�9�*M7� �R�|~7κ7�y����K$l�=�4~�)�f���V��K�|�^�� ��?���(yhl������m�:=�#h�l�T�wfT�E'zIY�HI���4ˍ)W�^6�Q7 �4�v��6�ܜk5cq�c8Y&>�lT�Ĥ����p'�<��k[��*����<�D���:_ԗ��Xa��Tޛ��<�}ٲ*���Jc��2[������{̻����V��I>�i#|�+0'�+�C��l�ccH��p|��5�FD�9��>����5f��,�֋���{��9���Q����1Q�E�N�L��d\0��0`Ⱦ���2�����}��(/s}�%��.Eq��3͇lfF�/��c�T%��f��Il�q�2q�g�������9ѧ�f�<Ӗ_�R����>Tb�*�V3���G�qn��)8�ɘ�CI�>}���(B�?���ͭ�>����'o|�(��Jɢs-Ɲ�5�h���$�{ s���`�&�JcX��Ӣ_�4�i�rHn�פ�O{*����`�M�����R+�pkjߣ�8>��fmh�9T�ů�c:����I�c�<H-y��Q���,~#x���8j����1
0�v�n�k���|�(\&�sS#�^���O�����E;&�\;�A���8y8!�g_2B����򬓳u�M�9��<���!Y�O������zô� ���.��Q�YX�/"�F����d��d>3����g>_xI�r����H��-��i� � �M����?��c��yif/����P��Ṽ<��4N��L��]�8ѧ�="�������ߌ���Y=����5'��n��k%�Ǚ/�O�&����M����x1�6I�%�G9����*F�������AW��ٶW��	�}�����9��*ԏ�i@u��k������ɤ�������-_�(�� �k���L�e��X2J�(L��� �b�!5��>�٠O6a��͋��Н鸿��ɪ��/j����_x�#(��D����jv��kC�wp�x��:�E�L'�dl�I#��#�sM��l�0�.�(S*UA	Gw�*�#[�L������`.12�� ����>�l�i[��fz�n���{�b����3�u�c�e�}m�3��Y�j�� ��*i���,']v����?��V���&<���~�a�`1&'����ܰ��2
��a?n$K0Bm�Q:3gʬ�:%����d��İ��V��r�C���1�vR*�C�SnVI�\� `G�������F��pQ8pd��Y�!���+:۫��^���z��@k�$�0�A;��l:sl��5��(��̎���=ߦ�s��f�����-zc�
K���<:v]����A��Wg��vv��t�O�I=�A7��]q�s���h���n�_zd��dsb:����,��L�`MX-���j���8��D���\]]ɘ�gN*OL�0���K���ؤ�.��M���ܤ�����F�#Q@���m��V��D!=����1�׸X'��<7s������}`	�^��=�攂�z��8������Ĭ�$�L��Oc�1�u�� (�!l��3����ե�����'j����5��pL�̆/<b��$���Q��/_��!/ ��(�\��Q)Y^��O����T1�*K-Yy=+�W�4O}egES��	�㊿"FR*�C�d.>�Y���g�w&7�U&2��I��m���O}����g ��aH����Y����*>�&�<)g�1.
�y_�R���O���\��'��T̣|����>5����� �?�\��|\����	ּ�˨.C�R��Yگ.Ȳ<���4Y����R�#!r��k���I�����B.��
�*[��+[9�;�E�X�p�f��)�Z���8�~�<a���6:���`�YZ岕�Һ���3$�Z\k �Y".1hEhk�����p4LB��!p�T�i��~��Vɨo��0[�f�R���A~�9�S#��.��C
��}h���j�b��0u��6���xl�
�5'��I�O��F�������y�l��.9�����㠵�Z;m��7��[�d���n?~L�'@5��޽}+�G�8i����f�>X�� 20a0O�9=��T�|�O�����%�rb�^��5�U?<��b�������+���en�-�PQ���"�ݨ���Z�xT��%A������xOҳL�80[����͛tq~!e�����~S�YS*����:�틏��*��7�ڇ��\��h 	�3p� �x�V�V�}(e� ,�~��g��o&���LV9�CaM�)o|��3sN��/:��<,)0Hi<��ƌ�0���lu������<�T�j�q��{��&�&�-J;(�)�z�� ��.+6bL���M�����r�Ii^n�Rc�%E�ί�dkgM��T	��^�r}�E��
�;75d&G�W�bE2�d�DLN$x��Ʊ�냬 М8*�q*�����(⻣����t)�Kp��B162ǡZm�?�ڐ-�x�́�HΞɲ ��8}�S�Dec.D�n� *N���F���G��V⇙�%UŴp��V��}/�W�%i	�r�nUȔZe+��o�Ń 	�C��}M�X���h,j���g}���^m!�:�sI�=�_��P�X�x��������w������)���s�t{+_�-�4 �T�dP�Z�霿��o2`K~����Sti�b`�pq
@0�%�T����J1����$�_!��f�瀰�����z�6������b�YD#�#�	���רa������E�FƓѐ`� �����d������?����	�{D%| ��-�2H��*p��Ϗ�߼������ac��E�4#E ��QOM%9�īl���X ��?_L.-L����JG�7��2��@� ��VjB#���5��hF��m�g(�!�fb�Ǭ^���4R�A���1dKiB�� $qO�7�ڕ�o�!:J��o*���I�K�5u>'�k�ڗ����R,�Uߛ�]��q��4����Y�hU��s�^g͍2:F����%>��@?~dN�Ǘ�le� Ϭ�A�|����ƍ�g��"��Šau�j9<ؔ��PG?W4]{�����N�	�M�l�����`o���ߣ�0�1kKE���R"`��sg2��Py��:�_�_�/�V�e��8�X"���v�M�y-��Z�.؍�0�����؋�~�^�	�(���-{��%�M%�[�&��^h�V.���y�76��qQ���M�D��덉�}_�٧_r��E�c�`��i�
r����Y�ߞi>jj��ɼ_���7�䳦��B�%I���R�t�՛7�j�)��6��-�k�d�8�����y�˂���`��wn!��̆�_0(e����z-x��,4A�֔"aر�YD&ȍ�x{Q��P=}��7�痳��l ��a��
���Sd����w�C�߇B�-ua�v6�����Zc4�� Ȏ��7�@S<��QX�6�C�\4��H�yt�?#){*ƥ��� c�.�U�f
V�6ʙ��ĆbC���B��\�
i��5��Ϭ��`
���yX�=:��D2B�JQ��(�Y%Kiԋ���;䷂�K��!���A�B}
&x��n��Ĭ}��F�{qR�Fَ]�AX�˕�Y�?[��d��5"@y���'F�Û\,j9T��V�fK���K$�v�P+
%`S�^F������ n�	|��~n Đ|�7���l<;d�A�B?m��R(���ov�����k�A���G��8��oi'����D���ll(���&7��Ge(��#fv���F�|.���N|�$
N�	l�.7����n��O峋3٤�!��(˃U;ZT�{Q{1;�іj�n|��F���%�����ZRðmb��
� ff��Ӛ�'hdEk�=���e�bC�\�`�R,�v�TG_�1�S��׬�E��P�2a*�/�%*^����Yt#̑d�訏k *�CP�}�6}��w� צO��	��w�sG�G�Rя��\��?��ӗ����ϩ,{Td���'^|�Y�O���kJn;�/�s��`��Hl@�?� �D|��W����qø�s��2�{a?o��8xߘI.	����`���h�FN_� >�-O��W��c6���\��"�g�e�`���hL���>�������� �0J�K0�CI�[����ŉ ��^D7'KI1#*L���d�j�T�3����=y`�{Of�U�i#L\��y�([[�U��b�j�ZAez��䞻b_���^SftL1]`9�#e��f�9|epp�M�LP<}A����1��9����~7T�����V�:Go��(9�Z�M�X2�� D��|r]·� A..�� �	U� ll�M��Y7N?{	C��&�;���9k�������5��{��|bU����W����
&�w�#���~ٶR�{��O�tb�1M8�-��7����4 .��`�M��s�{{ݐ�rB��z�+�PkZ�f;��O�h,��,�v�@u��H�hf�@Y0�m��67j��ڄ�c�h,��s��d��n�s�u;y݃�sA�Cs`d���	=^kM���V-�~A����ƪ�&	~`6�W藵7���U�iqg�%��o|]^\N��&}�ͷ"�%@�ۈ�*`fhl�uɲ��mӺ�]
���+*�H��R㉟��+�'��죔TV�<��j���g��:�%�{�a���/�GG�� ��	\C����t�(b����{���w�[��& tЁ_-��d>1	����4[���Qu}=�U��뿏��8�ŀ.6�g*>й-��d��$��FO/7l�gS���bTd�%F86��y@��+&��*�8�O�(���1:fX�-Y�R>~1K��k
 sR+�ԟ,�4ˇ����V���h���h��q5i0��d@u�	�f�{���@ԭ*�j���ރ���|tV_�&��N)�_��z4bȝ�R����}�+��?\�X�k
1���?��V�G��HHI&�-���퍼r�"�܄<q�O3�,� @��Q��,90q5�%�oc�޽v�%y����������N�o�:AJZ_
�8��qS�W�@?h���h?���߃�"�0v�! �R�1�a�P	Ӡi�ݱ��]���X��x�@�rp�o/����fz4g]S�L���t ��t���&�޲�,*����F�}�=�;h1�^M ��ZB��Rs��ً��?~�K��I[����O�~u��|TXa�H���Q��ާO�u7�L@`���Ls��-|	���n��O�=�D�!~
��b�"k#I�T.l�1$xva$�< (���I#�W��ME")H��ñ���/�;Sf��5�Y��_��CH5��
3_����i
�F���t��mZD�	������K�D�s9�����e)(���5�߼�q.6�\M Z�C���f3�K������ag�Z�������~�EHj;���Zfr�\ߩ�3~ǧ:���?��\�(=c�0�	M�r`�K?5Y��A!�\X`�.�=L��:���\`��S�_��2� )9����~n:�,m��k �Q��r�z��(�g�~�{ʴ�zF{:�'yr�0��T�ZM�^,� esCI*��~����gL"�0GJ:<.����
��m�#�L}[T���jGV6��'5����1 g*ã�H� !��tJ�lR=+���¬�$��b���P�y����gF3&��P��� k�!m��J�T�������>� �yu�G�  �-���n��%Y�)�P��&M�Wޥ���y#�!�̎���	��`��̊:��B�%��7��+��ᏹ�M¾���
�
�%���_9I��r̡�\t���k��_V�f�-��i=qW�/���՘��` N���0��HE�� ��-RUle�e8�8^[v|0ge�r���яm���HW��)��RBc�A���o�޸cye�2s΂%Q209��:{V���k��ͳb>W���0�����Q��^��55��ց�hQrRbʘ��X1l�I4uM�(�34-������2�M���ozC�<uG���)32�s�|�qH~��'��+]�=�f�}7����A%�~�ùM�H"��	��6S1�P&6�,���AX��sI��-rqy�|���e�>��_�JD|��>L�o��Y������cH,��K9� �FK}�ά~��E��D� �����4�~��O=�|ڍ0`��c����qa[$P	�p��V� �JMk
�$���#��y���`݀[��ľ�$:�$\֍N�t)�O��0�tPQV���hLQ(� s�5Zު�~��h3�b��-�>?dI��|��t 3'��y����qcʬo�� _
`�l���HL��Fd��_���:��C���933A��ShCS�M�D�+]�K3�s4�!�A� �Xu-�]G�00���?��Z�|�y�d��-��n���)[8�]y�K=2r��?OB�va{�� �Љ1q\��f�5���9y	��3O[�FE���Q� @��q��5M5m� C�߼��(�k���KڣQ)�T�e_����P�R'r��u���2�t�Iss��ōe�W�Z���)`Ek�5?n-)jr���p�Wv�9�s�V_�j@��(�|2�3b#��I�px ��w���`��Ogg�e�}��Ӱ��l�I�R}7j^��E�~���GЖ�$�>g9���8d�H�d�\��C01��EK�$;��}gz�! ރ<H��{$m}mY���ߋА3��}L��@;vH8��P��28Dᆍ|& =�h�$x�<�#��ɳ�%}c߹c���8��=	��<���Х���#:��Z�A��fw�=q4g}Nx��`JN���\h9��+H�w�:}G����:�Ѫ��s��wwۣ_o�����9�50)�6߆469�{F1a��Hr+nj����5���t������K�K��a��{�ƀR��s�ilZ�����2%
v�ϑ���4N�  ��&�]��j�C{#�r:N }s& `3���J�� %R7
�j	:�U���y\����5�@+���8h�|�>�gg��0�M��܁�ce�:M����siYМU��Z��Fu� Ke?!�������̥G����ɗ{/e�!�є�S�BA����b�_I��6 �b����u#�D\J+�P)�נA��n��9���I�R`�h�$�$�DL'�a��I�ޤ����4g鰟�õ�yn�	Ly�����#�_�y��:�Ͱ�M������,3Q���T�Q 6��-�� ��>^KC�sz�&���t{�O��j�G�Ȋb΀l�G��:���n� c�bn�����'�o/@1���2�7MeJ0!r�L��2f�d��E�5�+��4����B�Ӵф�̌�sb7�H���*�e��-u�3��2<���
�EP�	8g�9��{x�R�Y|����Ϻ��R�r7&��4΄�>���a0܏���ڍ�Q�:�F]4�E@+���&�҃�.Mй @�KwwȠ��tyy!cx~q�Y���.WV9<zb�˫�]���:��x	j֙�c��炡�y��=��x�y�35�i=��:�DF@��Hf� ``D�����!�e|�>nk�O^o����P	V�i�sx�(w�f��������MoY �� ����x�/���h<�.��.l��ɶ(�4ti7ZV{W���
f��0W_���n��v�G�IZl���pX R�) �X�̗�/}a�֯ c�$`i�� Q
�k-��9��W�"=T!��L�M�ԉXh��"�`	����?;��l�p�y���+�X4J3��Z/@i���d���L�E�L-��[��b�aP&uh��|P���=�|0����^��̰^W}�:��Ae�~�ur�>lx�m8���X��x�Y1���`�w� Q<�n\R4@��!���XIc�:<D��R;!�M�J���~o��on�o~�m���V�0��qe���敌��ƈ��@~��O�[Q�� T�v�Qi?�P[rd��f.���.,c�J����e|gM��	#a��/�.}$6�������{����{��_~N�O;A�
 5��`p�,It�M ж`��dU&Y*�fB���l#�P�t�� \
rkm��no�U�,.I�ڊe�Z��|��"�wz��]4��hw+��J�P���8I6Y���P�*����^M��&��f�ͻ7�:;�dQ�\�y��]ۆ�g9e���S���7G�(i* �&�a�J�74-#J���W.U!D�I�i���}�DX�Ndǲ��ъ?�oN֝�0� ������Ï?���j Sl.��0��sA�\E){�~����W�R/���IS��}�AY��s���0W��D��k-��dѠ ��e)W��z�;)0����o�)��N��#�|T�$����m��W�e�ڽJ�K��dP���/rJ� ۄ�MVY��Xm���jK��vM4�Ygj;�����$��`���IԽ2��)�XY��dH1omR�`#�9����}�"<�WM�x��Jd�^0�4S�e����O����O�ߧ�ۏR�?��5�h����Y�\��)�T�˾&j�	ֻl�4S�$���_�! :��ڳ���U�u+�.�Ӟ�L2K����� ߆���Ԉ !��-l�R��`Q�⣬�Ŧg���{sbn���8�X�1���I��h��{�@KR�5�:�}|���xՂlk���8�}��pvΡtW� N��쾈t�{
�/�uڷ��A�"���Q�7bvVE��&��ö�|@��@�������W���.�}�fB����ք`!j���dq��*�"�u����|�53��$ayI,9\EҶ��i�Pk�eC}�č�f��Ƈ2 k�L�ٞ7��Fg�$�B���m/��i�������{Hno�_J����g��:��l7@�Zg�&��\P�0;+/d���] #�|=��yw�ڎm�:���x� B���|���>g�v6��9q������"�^#�����z�g�`yyإ��\�dp$�n�e��q�k��w��7���8��gIA��� �������v�xs���ij��9�$~<�.,TL��b�Fվ����"�)�&�g�H_0�ߏ��)D>N���O�0����I?����Iy:K��F��:#�{���{��zd����\�e΀���z�ͪ>l%�y=�x����u�h�V��>D�͓�?:�h , �b��V#�'N^[�~�'�iƈQ��^�P�'��1�M�n���L-ҁ���ng��:�s�2g�m���^��S���]�j�LX��h�%����
a�h�KS���C�/w����!-]�f�-R:M?v����<��_��I�HJ�i?��~�T>���l�L�����Q+�11��� Ӂ�ͭ&YRs��k��d\�~���%<�\��/�����I�g�D�������~@�$ۃ+�xh�����Y�.'�t&e&���i���+-����N�;<���¦]��[�0A�9 Oq�0��� oL���r�Y�����ޫ?>+�g��,X.%����,�7��:�����#���F
&��E�~��U���o�7o��ٶI��iP;�2Hx`�6|Ydd�j Xԟ���Fˋ"etF�3��p@�J8�9J��{��,�:�n
�����Bg�&�����xf���B`�Z�^JMVp����6�K�F��F0hl)�Բ��`t�T(
�$���[�+K g�_�/c��{К_�݁I��:(���hG-/�E��S_�<ͭ%�ٞ4��/��iQ?�b��5%�>RT [��$B�3#Ŋy��8�F4��7o�a��ﾗ�#�Ћ��=|`Z�6ȕ��{�F��q9n�q��G� $����~uʴ�s%
Θ�"�	�/��Y���<"PG`q�����T�sM|��/�z�Pj��Ⳕ�����k,|��_)��:hbݱ�eE�I�1�A���ج�Έ�戣��#2^/����g?Q&s���ON���,ǔ��a����s�c$��ۊ��9JMP�'T?��m�Ʃ ���s���r�aM3X#&�?_s�>�ң(�	)Ά�t4�1�v��K�B��R"L��Ca�w�#)����^n�y��EQ� zo{����ɴ)�U+Cp�2��Q�Z�-��%�f��_�$(�����ݴ��M?w���i�֜ng���\���}�����ɰHh��ր��1g_%0�ę�1��k�_��Hf�D�wZ>�rX���h�Q݇�ʥ�j	��Ӏ1qUٶ��KJ��ҷoߤ�o�K������s1�BH#1���7 a{M�ԫr��|�gק�Y��$�wߴMz�9�Q����%��"�OK�:�Y땠 �s۾.p�nt){~q%����Or/�(�� qtRk���O@l3�0A./PR57�@�{�╬��j��9D�HZ�TC�[��¨�������=�+>S��22)$Ӭi9BiV]֤��@�Ҧh�,��J�^U�C��b�j~��:��a� � ,���&����d��a~8X���|�L��@w�թs6��riH�%L�D����f�澍��cEM*��~ة�R����Pm���ڌvb#���&}�识z`���eZֻkZ���̼
3癘Uk��b;�h���g�D��_��7�HF,������\U:˪	����͚�io
0l���͐�t�0S����p4�e��``�$:�[�?��� �ˡ��0�>���50g$Ǐi���hީ1�@�1�`����u���c�}n{f�K�z����(VQ�l ��S�$�c.< `1�1���_p��t���5����٥��h��[Q�$}x{iKpr�Su慨D��z*�2SR� ��k�L��A���B�B"�q�K��t���Ϩ�A�5��xtS�ȳ<Z:$��d����U���ʞߨ)�c
�� �[Fd�����p{A��8.XI�j1`ʙƲ�Ӊ�Ϋ?*!�~-Lu�M�Z��D����U�����U�4KJ�͇�kl[uE����yzw�M���ߤ��� �M��N2y�Ģrlvn9�:��u'�!�.�~$��M�U�Q�HM߅[ϻ�o��=@��[	�콃������X� ���qV�2^�I.�]���7�=@��� N�0�V�:��Y\gR����!������5
=Ű�d�F�A��Zk% �����qq'8���t�m��1K\�j)2	��s���0a�����'mV欨m_盱{��K�6�,ml��Kp��vg�L+4(k%���E;S�a�M�VB�1M�u�q���&�\���jE�k"?-K��ǃ�D�	�8�!��\�r�����{�A��߉vF[�Q�60w�NT��〆vf7i�_�'�M����O�|��l�+�S(�s�N���q��YHaB�X�yM�/8f��X�Ϣjm�d���F�G&�YЋ�J�[�$o!�IML�E��'[+C�9a�22���&����t@;���/����&�2ov"�q���mt,���������>�y'嫺�1|����Y�3¤�1�5�E���h�����_,�*�Q�l��'�	 �P3Ԧ{���0��d��+�:���M�Z�����r����BK��Lؚ�{l�=�bl����6�:�@�+�t��	��Z] ��ࣩ��ٺ�b/z��m���6��?�n;݋7>&Q��������k�ǲ!�2�@�ΘH
�ZeyؽMg��p�)4R�C����>�k�r�4��� ,�"�1I%OH*a�h�c�h���,���x(߃�s��k�'Z<X��$�Ia#�� m��M�usަ�~�6����?��7;OW� m���#������������,��K��t$�,��	Z����,�</�sq��p �WWjVԽP}5X�7f:����:Z)�9~=�{D|�n�y��>}��K�����g�.��ٴ���1b$YF���e���r�J� E6 Un�G���?3/
yif���>Q�JU_bL)9H_1�8*+& ���6�1��߉�B���T�f��	?`_O�x7m���2@��68b��&lỬ�H��l�T#c���Xvr��9�RALhՃ�vp�X�mc��A���2��%ճ9�H�F|����&���65;
��*Z6�|��30;X�h��	�3Yڑ�`�7^:*�J��D���,����l.(�Vߤ�����M�q﹞0>�@������3y>��fF'���	��4lᬋ������q Gc����=�k���l����K��g�T�M#?g]�g��s|��Q�k��f
���`�4%�pg�Oj�C���Y���?1M��jt�6ވ���p+ƍ�q�o=Ō畳�C����F(Vd�(D�ڝ�Es��e��T���wǻ-�Rw���ܫ�L��ф�[��#d����� ȳvqq�AO���k(���^��a?��T<J:吶�Eq|o4M�A��������e�o�7>VNb)8?��Z��3j�` ��fz�� TF)�`� ���V��}ͧ42�`�2���7j���۳��Ј��l�s._xm���
��<��w�&���I��O?���杀6�.�Ϧ� ��d+�v��PΧ��_9'K�cN�fF�l=۪��0�);f��&oYj�����Z��(�ߝe)(����X�Ju�R�$�����������z(	�/:���g~x�X4<4�,9b�eP�E]����0,�	e]95"Ґ5����]����hf�Q#���A`O�"� =��.Q�
�\�m�(څ�,�TLf����G�D�5��f��[0jSX�`��$��%��2b�;��V�a���Ll���5O5�T!̎d`�~́�%{�I�Tc�	���h��k�����fG�O$Q"�{Q,{+�=�,6��o�G�j2;L��ajrCcc�꿷Ze���7��f�W3@hlC�?Z�&T~M���Pu�Ɨ�]fr���&,��ݠOP��/�cg��{c����@�m0 �R�����J>�	�b���?}�����jر˫K�|�pH���_I}�����C�����֠���̣�5~�cFa���L(��&{�K�|4�.�a��NsT���T�>�Z��	X�H�����
�>�y�1�Z�eO����5�0l���������c�E_�Y���5 �s�x��m���|o������ll��E�^eM+��]h+�������rf���>�Im���Z�@N+��QV�`��׊j�D�c;)>��G�A9�V�A#��N���A�L�b\�뛷Ӛ�������)1�<xVL�v�D����Z�g�๒�weU,ˢ��L~!�`n	����A���<7|����C����?�6��?���]��^���U4>���5�J4�� 	�+��I*P��ȏ�j�f31g�(x�f��PD3$�X�0%dϐ�-����W���0%i�:��D$+��6�����u�7ߤ���uZ�L�ܧ�	���S���pC�Dm2�留*�fI��:�\
N,���MI�O��6̪�D��v��	5�NԲ�/"5%�7	2Y<��U5r��kk7�gRxe�5%��5 n T#{�����K�t�c��-�y�<�W�XK5q0���0�6��ښi(7�����uF�ƾ���6<�����g�/rR)�T�͠��I"���l�����)4�E����fT�F�N�!�Z������c��+�:<��D��n����wuM�����3`�PMｷtx�7oߊ\k� b2SKZ�H�\�^���o�*Ɠ@�`�h�������u퀏��~r,	u�!��^�>�3�\��9�6���k���z��7��A��v�����_�a�@c|4/�ĨI���V�L��� �{�<*�ht10���dn$����?��G��-F�1�>�9f:�[��c_����.��u�����u���l��&�n� �	='�I��q�P�q'���%�x�$	�H
c��RL�L�n0�)�q?��o$Z\rAM�{�ij���L����N�f(ao�~�./�dm�W��~/ѫ�'��b�{��^���c��2�j���ۨ�UwS�ՍHq�h� \dָY"�/��%@�M83���1����'�M��H�$15w���pU]Sս;K�#����)�����UP8���h���f��
�G��Jd~�)*�*��<;��y,��|������t�	��!���u�	r�dn��7&6�Y�6��~Y�S1`��S|�����ބ��by�~d����^���P�vL.���E���X�Ro���F!�����D��U�bV�k(o0�o�T
��pY ~���X��@���^%RE��f�K�z1L1�
 T��>����5 ��ao��(NN��E� k�F�'��K�Q#ݯ�u��h��P��=3GC��T�Ѯ�C#KY(P�CU�<�3_X(�֖�/H��"���uѷ�B;c�4�d��u���P_�cV�;[+k���Rc�7�m+�.�����J
���yU���Q�g�px��m@�Q�~�#�2�얯�~\Nsǟ�E�Tl�bO��}�!R[$<~��9����o宴�;LV+���#�������9tvv �j|A��3���f2�e��|9C}��<��!����Zc ���;�_�^��,>{P�@5�mY�pmd���Ct���h��M�>�ޗƏ�z������Y,�3J`x���Q�sЎh�ׯߔ�_a��^\@Y�J�N�{���Zf68 �Á�h��h�`��Ϫݧ��,���W/��50Yuʒ����b��z{\�u�:s�u�.�Ϣ�Ҙ�����݆_�H�vl8NX�G3z�Hd����T�����A*�U ��F޽}��k�Cl��������1|I�$łmY{����nW����~Q�~��i�g�����԰RS��3\o�}(}��2�Qf�5�H�%��u1�;��2K1#��m׽�̔]«�3��w�8�d�a�F���RV�}5�s{K��L0�'yxy.��÷��) �<</�;ܪb��C֪��źb-�A<��2��0Q��c��.���k�+VrQ���\���\.m��A߮t�x��A�̜B�"�L�V�v<��0�G_h{�\T��r��퍼y���W��QW��2מ41�E�p�?�]uy%/^|���ƪ�l�q����vt�%2��dLV�������H&�fH��c���c#գ�;�ry��g�u���f����X-���f���XT�
�������+��"�{��Nc���t��J�S;�
e���j桘�rX{��-l�ZԘ/�T`�<���S�YwO�ȚiAoCӰ�͙/�n�VOY+�MzS]���͠��'J!�a�c���n�>�iO3=����C%��Vc��N�Y�}�v���0��7�WA�w�N\��Z��Y�}g�����ke��:�1� ��K(ړʶ�`�-�1!�Y}P_��j�k�Ν����yS ����\K��Q`Tn�t�d�GY�Oky�d����3�����k����׼_��{�:T� s�믯K�X�ύ��Çt={�d/��W�7ǊD��݁���]ɘ3�-猲[e��嗲Yэ �{�� g�/��N�gS�v�7���v�����*s0=�s7�����	�s����'��4�ug���qM2ςf�g���0����-�\�|�ѽS�B��1S�H�W��w�^
�3��Q�.�w����i}Gğ9�,�#y�g�P���ꝗk�y�V�\��Ѷ�:�[�n��/J( �cB�;���WI�=���Z����yck��&�u.	�n@����S2Q��2�/�Ow[�::Q�ɵ�"�M����W��1��0b�]��c�`cg�M�
�?yV�g��P����:�S���d2�oB��z*�ӵ���ܼO�fe�n6�N�]=z�D�>&W��ȦLRП(y�؃�@+m��ֲ`]d)���\�'A� OZ�VLkg��fWbJ��˨�� ؠs� |ds,���HPI���:'O��6�LNP����}�ƥʁ�����ݨr��/�M��֚�Z_����4���9��w+fRe�6d9�eօ�* �~.*�A�뭩p�A���T�1f*Yߥ��Ɖm���Y��7-3e���0~��Ю���{��\��92,���:��� �9G&b�O��ǉ��Z>.t�_�G6��7����O
�����?+ #�X0��[ $�?GM��O����kΊ�n�"ɼ�W�9{�����k����&/_�Rׇz�G���w+�2q���{R��F�ZQS�_7�c��/e�>�Xt�)��[�ڗ�g2�����>��vg�.@��3�`� �~���}@��12)k9/�>�
.*��%��4>��B��Np(e  ��}]���� bl��
w�,b�
\&�ZX��1 ʹ�/ZV�_�0VJ���f��g	>��͔{��@`]"D��*������Ũ��^�krL�}������-���r�m��egT�3�ڷ�3�z�ao���S}�NA4~3��7 ��&��Y�`���S)��T4Z,�x�:�~�	&��;e�H<�o���6�����tu��O���<���w����[Y��=�X��1Hsx��]9�M�S}�A�M�����s]�!������5������`����a/,cC�DA�V�9Wƒ^-�\J.��vu`�6�����4��N���5��y���G���L��CP0�o��"ճ� ��"���#yP&(�9�ܨu���+��%�����Vu�9����Aa=�}s�.!�:�;R�{jh��
!`�Ga��@�%2���ج4�J�Xّ�R2�0��>ƔTX�S9[��ו�`��,���^���0�JZ��iv���"f�3��M�E����L��ԙ˚`���D�H( 3u��'k2��%л���V�����s�A ��Bf2*��B��7�j �y�kn\0Aa��@���LBc��n���#yƟ�LHa��砬T�c�b��� ��l�84&lb���e��P@���ңGe^���R�^�4c��`�,S�A�H x���`b�#����O?�����B:�@� ���o"}#���K�1v�>��t�{_���1w�Ǯ�[G,kr�u�v��d��(��j �z�� �V�K�"|V�����^��l\ ,��`c�|�C0�Z��\a&�b�߼�F�={�c
﹀p�N��i]��7*nZ�=/ْ�vm� �������d�����37b��]e�V��`=$��k�x�S����e��׽}��XV14�v���8 [���s  �5��5{R<C��=@7���i
�����]�`��Fs��b��]Y>_�s�A�O�>�	v{��ɣKy�`��3U����u�
D���&2S�&Q��U7|. ��Y�؋�/5������Q9'�Eh�����J���޺=0�sL���C�N���F�@L�U9&b��a��,T� y�Od<n�XJ� �W���u~����U­>��:TO��d_m��׷L���e\6�3-�<Ġ�m�f�����jSنV]51�M�栵��ep���k� ��e�m\��gI���	�3Af� &�A���\覅E��j�Y#���$IRS�9`UZ!Y�H�w(�9����~$��"؞,��z����z�|)c���;����:5�W6h<^n����
rOV�Ճ�k���qc�|�>��j���j6z^�AA�������kT�V�]����}����*M���J¦��T��I�K1�#�<I�Y+���Ҍ/���ln8�m���;�>%S,�+����!*:��g��l�{cY&X�����qt!�T� M��|�]i c?��������WW�
�VM� ���:X��w���҄����[���?�T	6~ee
0��|���f��ŉ�������P��s��f�����6�T���1l����Ę-۳�p?�6A�WW?k?`������w0N4��,��������Ϙgg*_@��p�eM{��z����[XD�~�ٸ�N�~5���ӿٮ�����?�p߄Ĝ��T�콅�t���d�Z��Y�K��kR;t��s�I+oWfg���a
[gL��+��}��Y�Fb�Q���T��BM�I]t��]0�J�b��ҿ$OE�WM��.o#��/w�y;�����Y�I���G	���@➨se_z0_���O+{�݇2n��5/�t���5)��+�݆ͅ|��o��򑂗���jh�ק�<=+�� ��.�Ո�+k��N�		���  ��2S��v�����"�-�4i��Ë�Qp~ .��:;+k|y-���`s�};<���P��VKDw;0���M�pڹ�mj)���t�[���%a����,Se��G�jL��}s�?[X	`��,�(3���eӥ�)��у��u�v;���B�\g����z��B�{B/s�
�;�TҴP"V�0�
���IW��� ��.��8x��*5ͭ 
�%tAO���#���ƃYM��`⏽Ŋ9p�1`_ itL�U���3Y���q���չU��|�lR��Ήt8�1��b#pye\Z�_���5�p����|q��|���3��'w�����穮�|�R�m��&��_X��z�<K���9����`�
p�@n��O�^W��Ȓ�Y��0 > 7~?D��Çz-M�(���xmR ��n� s^ؙ��پ �gɵ�I���/]a�r���1���a$!H]����{_�}���6�_��-۵����M�����:��U�
��	��&�ڕ�s�����X^�P|�K�x�Y�x�xF[���� n)D���~��/�X(7��uf���|�f8%�`���#�?��k��Q�5��U����2^)��LmEv*�������euui�:k��T�+��az���t�呉k�Z4�)��\Iu��� ��^Oy��\��M-�D�[5�1�P��Ie(�>~$O=(�6���"^>Ю�u~}j���������*�!Vg��R���}K�����{��[�g�{���me>�I�/�5�=�7t�?u�2K�OH�5�.5��B0�qtA��z��7pv�7����Mhsm-JP36�������h3}��f5q��y��r�ƪU��:'�;Q>�(wy�P�ְ�
$�Q�_�F_����� �w
.6+��V̔���<�0�L<h�m95����b����8�U�5w��w쪼�� \k8�Ί[O��8x�y����/_�Ɋ!͒�m��9Fz;���-\ݾ3�����/ҳp{r�U7���`v�и�f�i]H�
�1V�aS�+�U�ag��Yl��A*��8����T 6M���m�b�b��%�K�K�kV�B��%{�I՚as�nh�	�@[0P/^��F\� 赩���|�|��5�l��ǽo�����H��C7ucH �@���~��^������Rgߝ�\�m���0W���ɀ%C���4���s�'ٴ��~���u���C|�R1�����];.F����z��	<<�>��Bԇ{`���:��
��1���,���u��G뒌x	��i�0Z�wu�S�:�̝���{�iA߈�5�s�`+Ѡ}�+�خek�F?�`���^��7��Bڠ�g��z��#"k������N�k���J�u�:����ғ�LvB�2�1@������-� �P@�y�
F���r���e��a{�@����g��,�Db�I�Zq@�;�k��[��
=�>�eￔ�j�jr�>O�E�	���i��b��|@�G1X��}�x���t���@�b�f%�陽X=�
��&$�m
�,��Z+�Va̑���"��MAv��)��C�B��dt��Y�?0�-�o��g٨ڔ�`0�H�/!Ht�wv	��e*�ҰH�E�� �L��Uـ����U�{ǒ-P��L>I�J���di��t�4�;&^�(ĄVO�ڶ�s�}����kr���,R���V��L-���E�4��<Q��+mi���j&v)J�P#�PݎS6�(���k�3n�R��8�~G�	��
����@�Kθ��օ�83���LvM�W0� ����$N�Ū����|͵BBW/�c����}�x�Ԗ1.���uc�7���fe����mm6G͜� ���_s��9��9���_���}�j�Qw_]X���+U೼W���|?+��eƐ�c�c�q�3Z�X��g>~N��쵯� p߹��Im�.6\Ct�I0�������8�*�x��ok�z�����Ŀ��܅��Y�p=�AõO���~5�D�֩�'n�:���}}��ڴ��9�,9x����xLX
)�Gw26~0�+��� ;��.��)�K�!v����ʊ��}0^��W�kS�]�̞�ǰ��~�8�������,V�/-��#���+�f���{���2'WL��ȗln��*�Lf���}��+��,��s_��e?;�����Z V���+9�(f�cL�~�Z1n簇��փ|�g�S�_�/Vv�<yi��4�\�T�g��g7 (����W�w�:6'��S7��Al��?����Ҡ��F��/�*��Y��W�?X'��|���h@�wP#�nǻ���n��rL�A<z"���Y�v�U�	�j�.�*]0&8�*����^]��?S��.d�u�  (����s
F�b�b�Rkc�Jd��@�s�/�$�ꪬ���nnUwm��ف�ŋmL�Zu��s�5�/�7�J��S���x1X[���:lo��-�F�� ����`-AƋyP*ۆ��cBY�2�wK��`��gt�}-:�4qv��\��0o{>Տs*��_~T�N�8ܽ�g�k�I�zr��HKW���i��^�Ļ Dn����I�6S�wlp!�* �� `��6`��ݔ|(����v�CZ7te5@-V�7���0ՕP�~�aGV��}r��{-P[��ٿ�ǧ����1iK0���=�e�~� ����:	��"e��"S���<�u���*�Ivye�?sy�h]'R`za+/�.2˔n۹��6����ڡ�(���4�<JN�����.(�Tt����cxسXU >B�rgMi<�����9&�.��,����e~n��n"������xt��J%�!��Lh���1��Z,�h<�{�����=�R&ge��~8�>��-����5�&���I�]�#lN����O,?���Ա<Qzie]�Z�;��#��zl,i��[�#{p�uU~.��\%��1��\#O3R��	\.��E���t���kM���z��q1P8o@��Ɓ��k��	u�p{���!���ݩ��I$�E�LJ+ YP��'���x�O��>[���A��C� ��C�b>���T�]���8�h���P0@\���� \�	����R#S��&�k�p�����1��
� ��֣�^�Y-���-m&b��\3��3�o#Z\E'����A�h������u�5}���R��b�zS:���84E�'�5����mJ?�)Mm��CA:�NY��_�-�4���@}�C	a<օ4yܯgv�� ٯ�p��cSA	�<5�}Lf�1W1�4u�z�����/�u�h��?�&�S��;�����3$�H�o4�Yz�X\�A��ɓx�{,���d,��Yg]��8\$8 ���o8>��/l�|tGm6븧<�f6U�O�Ԃ�%H�W��X�S�Y��T��h�T@�),�}.ה���̜�������|����@�ދ�O�;�w��e롪�?$�nK���!~�I$~��4-c��9f�٩�j�N�n�zsPƾ�S����1��� #Ӳ�M��7f�Ln&�y�uU �B�e�xbzqƐQ�»3Z�2]a�ks ��֮�T���#�w��MX���\fU�×մOmoo k�{��m�9y6?��Y�d�����\���<p|�MI����S�WU�W �yQ��2�K`�:*#8�g�˛��\gEj�vҾX��4�q?���z� �z]�5�B��+I��N�3hR��WJyr�����Ff��0 ~�ي��5������j�%g�����gZvb���fklWz�~���ܨb�2_�<e������l��޽I0�0�xe�� `(~;"LE�E�ݪ˦���<e,[@)�@�	��8����e����lU���ب��^3cQm�� ���x�{k�PХZnA��^��xν�+��5�+e	�S�P|���]T�DSj������VMGA�>�K�
�
�*m�����`!{J�Yrl��k�,��U���HB�L��:_�ڡ������)��{�U|��;cQ�˲-`��r��������-��Ŷ�M�.��n�tVv�-��5�qA8"��Ɔ�6��2�Z������#v_�v�����ƀ3@�r�ܵ����{�\/��ގ[��p������������k���g�б2����;�p���Zz�3��y�aX��F�ﯭy9ZҊ�R���U�0����Cl��2�u-NZy��8�o8˭�_�z2.�aD�X]H��;`�wN�xE <�Qa[�)����0x�n�ߟL�z�bO#�,�3�=kϓ�F�D{?���#��P�<�\�_� Ҭq2_�|E�U��!g�V��ˬ�܆���lX�~8�ߩߨ�]P�$"�b����D�Se�4)���r�Ww���3��}O��;"��E۝�f���)��fP���x�n� 1��_�F�dQ{#�i�J�L���pF�.�����ss"�h?>�ą�l�q��:�ep�{01��P����
�����W�P'%)�Ś�>�H�ƕǃ���X��ִHgB2����9]o�XGe�'s?QQ�e��4�z.�ʉ?U&j�7�k���Q���3����nَ3�.���I}���>E�vUw�] FV���l�Of�
�����n86�|������+X���`�*��2g�F|���p9|�-}.�b`����rͦM4|�̠Hr�Ս��1s���FT6%+�l���5��*�J�	�������H�ˋg�r�#԰0�&�Vl>4gZ2}K7�om�K���?�9z�����5OŻ���$��1쯳2����)�R���pט�����=��8�Nbc��M�� $��֝��v���ձ �Q�v��~�#y��G�'^�3����J[[<Q���X{W���M��^���P!�dƹ�Ø��97��!���,��[)�$!@.�<�:�m�:�Cua	�F��z89Q7��z����^�������0�ߊ|=�$��C�������lk�l1Wi�~��F]y�FY�d�-C�����R�a3�2��PTx��)����]ki����>� 9�C]�V� �_ ;P��S6�7�(����tbE�u���7�wf��5@�y&ki$
l�ab��`�aS:�\V����R���+�$��T�>ՕDtbn�d��G�?�n��'�Y����8�Y}���?K��-cÁ��d�'��6�({�|yl�h~pg�t�Zu5�����*�Q��Z+��X*}�xtSG`6 ��|���(SXe @��� �%y�1��T��$���[��2z�e4��������2��Ef;��Պ*�ʃ��r�[~���%�5��ظ�V�r`���IK�"����-���1%�h�*�Ȍ-��4��,Cw)j���gvLĘ4=}��_�������
ܫ&�Gg��6��C�w�-�`^���Y�:@�`�j��w6N3w~�`��o���8� a	Ėל�N�Y׺����F1JXu�c�]\
����u#[_�`������h��Ǒ˖xA�΁�լ\u�4P6��-7,<�ߍ�%��3��;�2b���k��5�ɟ�U���s����u���ZZK%U��X{<���������,ufo�D-*�����Y�\7��y0b�^���;���Ў\�Z�Y08���h�a"��y�a"��5әZW��f�s��2j�u0׿�+r��C3�;{��K��RͰ!]&U�;@��� �!�3��OqO9��14$σG�u���)������S��M��e~)SG\��j\&���c۽j���냤j)�,��~���m/� �����z�Z{����`w�Q�� ]�x/-���A�>�&4�a ��0�,�=;�)����N��	B��'{`+S��vѴ���@C2bn�x���1�b��x]/M^C�$R6�?�v�*����Igf�ƙA����a9���{1p���"�YL�u��Dj��ݨٙ��h�b<o�
�6��{�U�Y7g�W�٩.k_uA��6�Eyѡ��g2]�b�����cC���P�'�4lD^�9G6�&�]T�ޅ�fcCe���S���|#^������̴rP���.�x�f��!��O4Nf�aÀ��?�/�Rv���?�[���9�3Ki�ֵ���kN������)�>;-��K�.]g�v	�pP\�f3�`��l�'��a�k�Z�6������ۮ�ε������h�l��ޘrg9�Ԯ 3-�ͩx/7"�������T�(ͼs��r�}�O���4�\³��i�%U����\�%Re��k��Z����e��	�������}vѦ4ީ�N餦��J� ���^�l�+��Ծ�f�8����Z���a�Ś|\t~O�d�x�Rb�Rg�����z)�ҟ���m�ſ�$j���{b�k~q��uw*!���9��!��IVت�h��IZius�:#��T�!=�|�ҧ�y�j���($�� :9:?:��,^��XZ��Vk��4[��0t~/�d:�N������A]my���bÏ����w�Ж���e ��u�j�l9�����%-z]D�,CMY�r��D��� �&U1Yqd�]�����l���`ޙ\�vgnGޏ
��[ԙ,,N�p��, ��k��Må>�V	�Jl`���72��d�eX<����Ă1�U!�v��m�#��/0�w�����ͺ]$<��.Н���U�Ni��yR�LZ��:J��j�R3�� ��%0@/�A �9�����Ϭ>(Y�\e
�额��c\��j+wP��\� ��P�:�[���>�~�}�a�s�u�w�܋��w'��ߍ����o���h������md��w{���3���șC8<��u	�n�9<��ץIp�v���c�6q���3�v>, y+���0���~�ѹm���
k�*͡I=Lp�����}{����2����j<:L\��ˡ������Y{��d1o�X������ފ�#�|�@,���+�Aۍ&�]vJMR�Xa�j�eM%�9��f��g�4�g�1��+��Ɏ�y &.�L�kF,����z�H��}�0��)�*T��6#<ni=W��B@�<Ôٛ�T�P�{�f�Z����=�o|`ک�(��qO߸8rnp�:�kZ)�"�u����T5���h�W�c]�Bhέ��WА�>�[-�z��p�Ec�H��O,#�]K�ōu|��Zټ%{�W#;��2J{a~�n�	�3�2|6��'�[���"�Z[�y�2� �i{sg�Fc+�(i4X���c��k�-^̙���3t�k]��Ւ�L�_��\6��NV��]�1)sâ�L~l����	�t=.�����Z��6X�Y{Ff����,%�@�i6D��Ϗ�|苵���,��⻼�m�)�N�Hsc84b��T�g�P�����E�.T񵾚-��H�nJ\��g֥ڶ�mk7���e��v�7u�?9�z{���y�ǎ��>�����-v�ǥG V��f�q�84�V�n�h��٫�jv�)pC��	k^k��M�uW���)�k���'m�z�ύ1�����<Ⱦj��[]yzT�����ű���R��3`���~���:O�ʊ��&�h#����:�T���OY�N3��O문���[`d�G�Np����tV��W�L�u-pc�{55�mh���pԀ����a�1U���m3�jls�ٞ���,�����X�F��KF0��U�T:6���~���XT��|/���ώ?�����M���T����;���) ��Y7Tb���.�Ё����˷��� _pS�`���D���f��o���Z�QZgSPhLF�ז[oj�h0���̳�K5Ѡ�"XU��:��H���s�r�		���o�[ha���IZg�w�E��JMTW7|~o�{c��5!M�ubY"���.dHM��2�	��XQ�(k�fօ�S]�(},�c`��F�"��~{|��@q���۝..�/�َ8��7�I�3q]�[�� Z}:V�S6��9��n���^D<�-�
���!{ω��4s�cqX�)7�s�瀲�P��qŅ	�nX�<S2+�-v��68�(����0sg��;����&�����ιab<���Y	���3���3ִ�g�3�ÿ�) ��wgn1��|���-��>&nyx|U�ژ7��d.��n�(�� 2�����L���W� �q������w@�	R2�n�����_k(�j�,��ʞ���T���	
#�E:��lL�ϧ���5��8A��˦m�,Ȗ#L�W�������g�&��j@�,����a���qs��Z��u���6#�c1�tN6%�N����n}~�t����>�@�pV&\��{��Z/�no������AW�ō�$A���1b.����٘:�q��?�nR�cS�T�T������C�^m�|���o�R�;�% c�|��"%ۃWʂ��k��)Z�䎇�0)"u��頫�';���G���Kpr���V9^ S�)�d��6`:�� �lJ��P�ųU���ნ`��>��v.������2!�4�F�����:��~)�h'G`
���	0��`��[e�r�����M�i�앁=��z�[f���u [1o�����X"�:k����َ��jnW��XMH��~���lqj
���KX�̲v�]��-�}Mw_NaƩ�,��ړ�i��$�����Y+����y�B�o��֛�]l7�����Z�6�֍4��X6M�@9;`>f.g�\mu~qޤ���e��1b \m���7C$v1�+�
v�%�E��Λ;�
P/AZ�f����?y�]����^�{	�!��q�s��6�����j�mSF�cӯn�>\�+�ޡ[z`I(�
�;�H�c��>�Ċ}��3����0q0`�z�l���AeW�u�Y�:7g��Y��E�W��(�y��%a���.��l�3,�����$�˻��#�[����9ڙW������Ï�'p�&��c�涉���\���[Y<ZM�a;rm�9�]���\k�@Ju��^�SY�t�{�Ht<�.���yQ��X�SW%Bzȫ0TI�vHZAҨb+�>Wvy~�58�Y��&8,��L�Z�I������D��I� �m��Y�o��������.���FiY j=!�ǜ-�h��9ܠ ����*�[�n��B�u2���o���OT��Mg�c6V{��q�.������b�+ǿ|���=�(����/-�����u���ӥ�5�7��#b�w����E�.�Z�q~���7
�a cv[ �^c����9U�>�l�~U����\�e��Hu��2�OǢ�(u#̰�Z�X���"�LaNA�"�nQ<��LsSD7�?޴�w����}���85'�etL��tn�^�^�,O������lj`��%K����?(�;c�5�&
����7��\��m���{�͛��
��y��q9�#�-��+�-w�?m�?� dA��:G�����:�h�����;�c�N���������)����Y𼹔�f��@�EqC�V���l����2	�]rW�_1B�e�"���B=K���$�Ԑg �}8����5�>�Z�БCs���k㼾ylX^�F��k{e����-ݯ]�J�k1ٝ�����Y �>�l���&��AR������ײ��~�F޼/�������v�1hU�&�Y�IP��-�0)b<9��F@����\��B7�����O5Uy~Bx�͍��P�� n3���L:�f��XP9Y�$��l�#^��B�����2�6��8fo�´��1`)ͼ�:��"�ꟗ��|�/�;u2�q����^i3}�4Y��H�=�k��;}�4{�ar�:�ypkdTw8�&�=cS�ţ�zW VY�e�뼹O�
Ζ]ch9�#u����.�K����0�&3���΄(�q�`�,�V�E�XMcf��5@�>Cg�k��rI.,��bMI�õWF���ؠ�\cj� H����bc2�� ��\�i�ā����;��x��d�?]�&�lS�hm�2���� BX��MՒ᯳f��i5g��R���9��Z�({��l�,�<e���&6ɗ/_jB]�-e�6�'O��`y��=��.,c</�HZ�����f����zw:~�g�
���y��c���6���^y,%0.�N�����c��M�?8��[�O����kv�]�T�ْqkٲ��_��sON��ꋕ��9���{eR4�OĊl�Y��p�;�q��bS�9��v}�A�3����9*�1#���&�O�]/s�k���d����g߼}����ؤL/�sQ@�~<�ԓ,`�ѣ��@kO�C��r�To���i����s]S4{B�x�=���nS���0=�rd;���g�����ُHh�`V�b�+g�V���,�bUP�0�]�h�S���lb�3gc��?��VޢڗZP���kZ�������9���h�J�u��Ie��0����Fϻ�����'5cդ��o(���4�P.��G��	��<�%�'���(���sF��oǢ67lW�����_y����wi��-Y6`����A�E�������A��� /q9��[��x|w3爵���Y��V��x@Q��X1��AL2Qxw�ܒH�j|>�{��,�M-���Mҥ��l�fu��ߜ�p0�.2XkeS���a��`�o
�Vn����b^��`\O��$�]�a&*^�!o��Zh��2�8�x�L��N��`Th��j��Yr�~�x�G��~�Z}����(�@�M��yҬ/��ل�3���?ʯ����
�w_�������q��H�ک�M�~�u2g���;'�u�G��ǀ׃�q���r���}��i��>{�L���[��(��J�`a�FLf1pu���p��.�ܸ����+�_�Z��c>N��u��j,�1=
}���//�y�,,|���9c�Ԅ��c]��i�\�߬ɺW�͘�;�����ܬ�.	 �ӆ����=�@�_��1��;X�	Έ1����s�o��_˸yR^@��$b�z�����Ys�kNlߞbX���
�ؤ4�(c��>�zP��w0�(�<�:�(��������Ok+Z�&3��u���'��>�sy�19;��~60���XNj�� �x�5�*pG�ǁ�T��b�s�PR�n�=���{g�}��9D�S$��}� v+k��ط��؇&f�Oj��u�hxL������ݏs�94<��O4 �
���t��κ$Ꭾ�G�4��@,[��ν��XG��<�/n���e���r:�4�x�?�A����Q�~:x��|}j��>X�w���	�l�Y0<��5fW����ٶ��7X����.6xݨS:jI�EY�+�Y�٫��n��rD�,��V&���X3Ѿ��+[�	�3W��u�6�ƹ�uh�w�Q��k#��tb`���$����f�z�Ru�4�����e�l��h�h*�b�������^��W��ǟ~�������>�&ֺ2��z����좴Mr�3�ؼDB<S��Uيi��j�z9'�#l�0]�o��`��A�o�Q��J˹�Z���q�q��n�r������q��}�8h�w
.�׽�P������9��O?�,��?��_�H��� �J7eM���M�3 cVj��1��m��K��8�M��D�a�hƠg�ec�B �k��FdVu�Z����L)X��ke����{e�4�zM��ǿ�V�bn��k��v,�rm/�=2~Y��|NG��h�S�h���Y<�+�u��D,n�)�;r����S�����q?���پѧ�&��I� �3�c"cO��Q571e��!Y	4�gBQ担[H;�*���hkiƶ���!g�j,�+�kq�r{s����7a�`D�9�����t��9�j��5`�C�x����k4X,�-���n�0ϓ6�M��b_��|��=ӧ!�j�4 ܞ��|F���tqp?n�٤��a�N���}� O�V�r��m������{Q~���׌�q��7«��e  fڧꎈ,L����5�S�x�4YMJ�D$L:[PP�p��� 25h~U�Q ���P�	��S�ng��^��tkݻv�׭Cs����6IP�:/Ȏ F�����
�{W6!�j�Ň }ַ�����5;���|<�7��I��a�,~�ş�/(��`�Q-.���/�ʿ���-����(�z���2�E<��z#�
 ��.�z��ʋ��� �{0b����q�LW��4�e^��Ҋ�81�t��^]�q�a[]�϶����E�%ܙ������!؛-X�����#�>�e��|ܮ��c	�����ڱ)$��;p�5��3�?�ǟ������?�8Ѡ�ɅR7p	�������&m��!krCb�
v��)U'�H�<�р���U�����_���F�� ��t�z� ���?�/�Oe��������^���0����`��h,%*>���?npd7�m��d3�p��#�3F)4�<Dcb��M��Le�D��CV�J�ΣW�0�F�����ݴ�yEk8�-���c�g�xda
��Lם'9Ѐ� �n����@k��Bg�a�il-��!j��\�V���'Jy��p =q.�'p�!�}�N��&cb�����I�����(Ӟ�Z��t|5�F۩]���+����4{��}w�۸�ja6������4tU_��蒦����Y6b��U��|������q�Я%N$u�������������Jj��߰6�/��n���C�Ԋ��c�r��V�������xJ���7ަ^�?i��l�>ũ�4m�R��rvyj����c�s��X�hc��Q��.DT������E�x]�EY�QC��q�����۝\l��.v^����re?(R�)�^u�������c�36d��J׋�b�p�0 b���F���O�����/��"Ƈ��k�)YEɐ��/��"���:H���ђ��ް8�ZQKh�M�3��J���&q���z����n�gϞ*3�/�����;Y��25}�dc�q7�t�/�.���>���:��;��~����w�wTȨؚ�x��bv�m˦�������o򺌛��u1Gg�;�A�둷�c~
�=/�� ��ϔ9��d�Vط�[�Z���o�Xo"�0P�~R�
�#�{F2	�s����B��kӺ�y��Yw����5��]�]�}u�2���� v�9�K.�@�n�
Z`p��]m�u�,'+?Ĺ�ڐu�W����q���������)�@�{�Ѥ�H5��^?�LAKhKpFN&����l�Ρ~�6#L��
n���0�ִnfX����U�.�rr�?����7����5�fB�I+ؘ$�fA�;���:�d�8|M����O9��f�H��cb;��B	"���8@[N��L�)^������^�Iy�����m'ir��u�I�z����	�7�'\tq��k�k��rZק�6�d]�aUim�5�w�A��][%V�?ʱB����:��v%P0;j=6�6�� �4��-)n�}ǎ�E����)Y�}N^4��ky���e�Z�i %,ta�2KL}yy��+�}P��`{����d�%�:_�gQ�uGa�[d�����i�	��@��T�7,O���n`�������|x;���Z�=y�� p�+^��OM��.�[C4����$�q� 6V����_dqbG)d��^V�J7���w�n���M~y�k�䶪��4��=����6Ǧv�g檌~TW��\�Y�]ͧ������2�e�9�an���S��]����ȶ�aTN���7����ט��WZ��� �J���NZ5�׬M���ԾH�e�^��MG;���������P9�צ�=�r��;\�8�z���>� [�������W�p}C�>�XW�>�O���L*	c0��8�e�௹G�_���׶�1��X�s#�����$6��V���k t���?�߿�q2�Y�r���{1\����!��g,�!���o��oS��L�������-_?��s���g�W��W}��zUֽ�����J�X�C1���q�'�t�?�ud�2E#�»�VZ�'���T�'i�)����1l�n�nλ���{E�e�V��ޔ ��hQ�f�|����jRρ��=E�CV&��Gyo?1����g�3d����NA',�UiGT��ݵ�z�A���e�Bx��fȫ���ƿ�������j˕�� =E��T��m�=��Db� �kve�߿{S���\^�=pM�a=ib��Ī�ʀjU��ݐ�:�g�������MM�&�*@�z��h�1`�c��_�m)��J-R���yf����?�u�OuNl� `����;p�|��ɏ�f	��j^~�onvǩ�W��3ˏ e��5����8���������S|Ӵ�Zb�������n-�H����â��q=����e��>�A'"&'Y~Y� ^���b՟G��oood[,@lΡ�m��h
 vFU~�T��P|�%�R.�@L´�G�.L�o J�(>p�H�TkhJ�O�ڏ-��k62�R�{B�f/���˗�
�zU�d�������nv��|xr�d����`ngtk5:̭D�T�����31�g6D��]�R�=�Υ@��I#��d(��H��DL\�=����˳[ٔES��&��k0�F�%�ԀfY�_.��j��y;�����(L�;LO,@B7�����T
a�^��X��k'*11�k���M F�ag1�}_�Q�9�9�������zƒ�[�0m��u
C�4C���� ��Ÿ���֝Ʒ��o�( �J.�/5�l$Z&O�Ɍ�u&Ƕ�&��KPY����u޵��|�N��/�D̮�	0d,��
�b#�(���wM����9�G~VAaY77�Ju(wqJ����&X�:�=�w�Y��+�,�s��XЉ��!=�	eb�g�P�\���+��Jt��d�6E�)� S�OA��P����>ȯo�I���*B���)�Lݤ�L��~w�PWjߙ@�Y���;t�|�����	%
�ȧ����
����*�=�6(��Y��XPO�]e/,{b��a͵ԭ$�Eb�����?o���U����Iw�iD܀���������*����E�	�� ��x�~e&�
��-$o[{*?�l�6kOn�?�3�8���B�3U���f����={�ӐⱈJ�+[���{k�������Go��s�~���
�:�7��6�Cyu���8-��RL��Xݐ���6��	�ZN�/1�w������� ���0��V��'[$��j���q�nM��:����;�����A�����۷o�}�ԭ�K0�5&05`���06��ț�{Zz���Բ?��̥AK*7O�E����%�������$x&<;2����1���e��f�G2�<;�-]�K�澮�'�ݮQ�]��Ygr"|q����ⵯ9IɀN�;���_�c��q"ܘ#3���8�
��� �awݙ�?���TW�yV�p;�o�s�x5lX�F������y2�H\3�k͢��lk��A~��'9?��/��O0��W��y-����z{���{�#VϪ����L(�����9�1�j
x��L��W����́-����RV�[ n���<F����L�\eͨ)�!
}���2��}�vA���\̐�������,i
.Q���j.�b��4�@L��yf���Ԯ����Y������m�R-'�Y�+H�L�`i��ʯ�ޖ�*d��@��pa�E{��;��T��ݭ��C.t(�ꀶ�e�*������Hcv��Je))q�k� �Պ�{��wF8X|���y₁�2.4i/3��_WÖӐ�|g��\�rbweA}\�1dGp&�uȜҋ��M�%4�1/t�T)� ~n"3�%6�I���|s�I�L�Լ꯸��ɉ�~/t�D�_cSZe~f�Uf�K�XU�ѣż)�3�ul��?�\�R,���"ă���.���)1#G]�L�@��+�# ��$,�{Fbo�bk9[3^Le*�%(kv��ָ�����υ!ن���eJfm�=o������O8��/D�l�b��R�4�MwQ�\lsM�x��\�&P/˴x�ǎ5����.��{<Rn�����
m�W�<g�=����:�<��;`���{�q�^�����jDH;o~{n�3�?������qp�lv�S�w@W81�����={&��ql�oK[���
�@�p(��g$[�b���5J�.Z����� ��	Su%Z���h�s�����6YS+�ӵf8���q X/��C���Z�k݇q63H��k��G�w�M77�Xe2��q��5�AD���J�;��e��PJ����F\�(h0���ט�Z�FOR�7fM�鶸���ke�ih�^i�в�&��bȊɜ`/�,�_fV|<���ce�*�Q�ѩ�7��Fv� 5���L���3�����ܝ2Jh���"e_y��F^�� ����&�z�t\{��^�u4Z r��ps����\:$ٵ��v{|����0�6��@<t٧n�a������V���-r�,8(�OS��d���]f%���}����s p�/3�-t¬$=~�x���~��X�0��gȨ1W�Q����~%|"s{���לd�:��K���?����kL!��q3N���;( ��g�n�u�>i�	���Y�q2���=G�h���nnc�`_,��N/���܊���O��(o���g=GꃩNX��{pY��rW,�ҩ���[��\��젰f�9U,f��|Xn�)_�~��n&�e�j�m�L�ѩ�׫W��s%q/����m���A4��}F�AZB�c�3�, �T�f�깣�{��lc��i^������xg��Z��"J�k��| ��Os<����l|K���ZͤO��??��9���|��~�3(��.�K��k�(��w0��5���:3���&㼱�Y���-�We3�Ή��������<c�>u�71�:�����[g�5����A�����ھ
<�wt�d���G��ъS^r������U�E��G��<�|�Ϣi���2;�*� ��[���7y�⛙�?4��ϟ�����E�Mͦݷ&�#���}g�s�3��Av$X�KY��+���2dJC�ƒ�t#�v,N����\U���!�Wb�Gu�)�a�]�m-0Y�c4Ǧ�>M�Q�H�6�BQ7x�m�E��V�ge'lCh�VU�������wW�i�7w���S>X����=w&�ÌP�c��Һ<۶<���/eU@���i,��:ז��=#�W8p���5[�=[y"���n˺�V�uq~N��L�q���lRx��E����V&�+�����^������J�Q����+��u��c��5-�I�*�����j����U��l��-F4vp�q�ݠ��3h)y�`���`�n����XA���gQ��p|�-�A�����|tʃ�j�3ic�����ڗ� �k�h��k�T{���Q�o�£k�G���Hq���x�T꘎ޛ0�i����l���B�oo���\�pj6����4$d5Z�c2�/�M���b�B�B�/;���,$�}�z�� m���ۊc7�U�T��s�d��1^��ZV����ߛ�8#���3���|J�xr��?�F[�Eg�d�ۻFBa~�s���]'䧵��S��C���S����.^��{��4믏�7�*��l�6�ǽm�:4�ԇ6�a�ծ�-�[��)��K�R���{�DI]�s6A�؜M]�}O�����1P�X�X�nz&l|(��4T�o��[������`�u����W �Ճ��ￓ���*l�����&<xx%�����_^�*o?��Ͷ��^K�L$��f��2S!4 -`eE�ziL�sݨ�iRU�j�bi�Z�5��xʝWfɪ@�+��I�Z`6ΰ�gj����:�������܎���Ì���P�%���6���ǟ�����x�H�$���a��U"�c��7Z=D�ט�5l�Ȃx�Y���]��Bi���4>{���5?�9OG�xb��@%s�{�Kc�2]� `�A"rڕs�P����4��濞 �a�8��x�Ն= ڱ��Ju�q��6�;}�m�ԓҡS,�Z� �0v���-�y��l�˕erW`G���V2����uAIl�Q�#����t� ̩�vW��Ǝ��%$>��٬Rc54��G�!� ��@��}�]x{�8!C�X`�>ܰ����9��lOw۰Y�������@/X�m�������@��2E3Xֺ���uaNdyt��)�+�n%�*�[��ܯ������hFdu�j�v��}q֡9�a�:bѱ�X �[K�#\%�q��}�ȅ�\�u��,K������4j��p�t7�̍����@J�{i�����D�}s�}ґO��G:��r�s�u���5(]l3�e���H��)��k2�X����s��e�IɌNϮ��'7�[rus��q<s6c�x� 2����y�e��\Ǹg���|i���n^�����ӹ���:��HPoN�6��>T S�m���o��v)/^<��~y)��O����� �;Q�V��x�̕�w�' u����� �aB��I݅ʚN��A2����`T�s j�Ig�0:�0��Ѡ�3k2��gԸ>sGj]L+*�IB�I�������չ��m5܌1Wx�����qn�K���?�E����� v!�$2�n��M渴���������;y���\^=* �t��S3.#x�L:(�-�����Z��=��/<����$�W�5q6��Z��SZRX�y�ve��i8��m�Dm�X�R�R6<�tH���6���o�1՟��k��j�_����ذ�� O͞�o��|��|�&���I�U�����EL���fY���P�ȁe�$S��%��s�-��&�fюE:7W�������Et�b��_�_N��;~�SLLA�if͚���U�����!�Ej�j�ZG41�T��k�|m�|��j椺�:���X��E��-�����1E�����ޘU������vG,�-���qf�f���S����i7�vc�{s�C����7��s\+����hA�8s��ud僥���x�܃e災� 䚬3_���ɗ��;;���1V-�w���*K�ޒQ<�{�[YF�-Y�%��_���F�!R��IMuw%A�3`n�E��1�+K���:���f�˳y�*k���fJ� ��I˰��'ҬSȸ�ì��>#�6{wf�~�1��b\N�� ���᚝�����؝�&�����&�@�P�rq�Vuw���%����\[�0^��Q��
�4�/��+���)Y�^�Ϯ/{�����<����9�������xgIL�a� ,!���t�R��X�f�za�����p'+��j�0�H7�S��^��/�^���Y��y�`S��drD�'C7-�����o����
^&��a�ֺǩgȐ�jHh_-۵ոdx2�no�`?:+�d��,�x��T �f� ?�q�+���S= ����مf�zazaֲF��讖׉y�����p�	�zNt9�;R}RSD�[��c�@����+y+g�qϯF���Hkq!�g���5���������e���f�����\���6�)s��>_���dN�A�A9x�����!��lI*��r�����ә����&5+=�4E�3=��.G������ż�/��|wwS��ڔ����+��z��:q�nX�l�VqO{�\�5k��'a`��H��WY��B���mai�*������Mh�������EQ���,�����"���6���g�k�Z ��fЦ��s��sч� Q�5���^|�U����̯��)G�t>۲4��^��i�^2`K v߽�|���Ɖ&�f�����_�e���Y��P������>f��5kK���Z���KY�K53�e���Ml�kEf	�������R���_�,�r��H_4{�Z���k�h$Ea��H�GZP8) Ҁ�1��n����@��&�QCl��;f6Ȕc}{py.?|��#ă��pm �I����;K����3f�o���1�vRF���b�X��fXە@'��J�Z��JeDC"t۴��JT0&�;��hLXg1��1���נ�\p����ȶ�M�Sͬ��]��#�J�������]����{Y�]��Kq�I�^��Qvw
�x_~|p��
�V����Z]�n0����͵��o�dT�7W��e���!��D����4�)�l}�&�Q?�Zx��T�ݭ��7�F�Tί�w�6Vs(�r9*��V������1�^SV�rE��r���#�K�����S���V�U�N���Mi��jc*�5nb>3����3q����D���%S#LP��@�0f.bΈٽf�F��y�K�����n'��.A�rS�@4- ]2x9�vT�H$U��i��H0�1's"���*��Y���Tip�,w��9S��S4�/�E���+y��J���c� S�n� ���F�%��۹��E���'��pT���\�~�M[JS�+��.�`%�X�~^���|s�8���a'*���I\'>+����Í �o�]��6�S�_͆� ���/�o*��ʳ���.3X�m�Ά��D���>0�a����w ��a}.5����$�T��Uz�c�
-��c�݋����O�g��<��-�}�}J��2^
�l����#=ݾ��G]�����{V��L��^ЀP�'�
S�fƺ�������ɔ�{�c�ǵ��#����z�|SֶGT���Wo��~��$����_F��x�L&���΋��Iu�^"��ہeq ��C�!+3�"��]�u8p��������~ػ�9����9�N�������L��]T4��P��WW���n�����s'��<P0tu�+�W^k���V�q��?ww]@Ν|x70� �S�����Iդ2�O���F�@��y� n�����Fw��A��f��/�k�,�rHdQ�'2�r�"��희n����FCy�����X����Z���u8��� ���0a��g�M`���|Æ�ŭ���>d�A�N@��uv~�@?~�V�o�R��ȱ�P0*@���B��������y�
�yftf��s����Jn�+�P�"��Eyy�Jp �,3�Z�͋��jyX`�][���v3]Z�:S����������Y�Z���M#le�&�5���kn݋2������O�+��Bٰ�����%�󵾠�;*�酫�-80ik�h��v��:G}v�f��1<��)n˕���q @���sK�W�)6�|-㾖�_��I���X�e2W�k�N}͂tP8Z��9��ߴN�O�hs��{�����1�3�N��#hg֩�h�;z�i��LL�;�Uŉdø����`q��F�ٻ�u�@a`ucĵ��c��ƒ���Hn�vc�rn�6���;�-�wr�/��&=%�%,�~���8nޗ^� �l�Ȋ�o$�0K�}��t��ݪ���+#N�b�������NY�����Do�� v��9Y��({����r!{� �q��d�k���k"C7�˸Q43]��������,U�;�uk�h�aġ.�Zc�����;��!6�\L7{����'����h.��EO5�/��F�d��\����W�Ϭ�{��%�@���|�* ��(~���low��=��ԥ�W�$���:�vO���u<�O�<~$>�+�J>����g��d���f4��C=/�~8G�Y��f�1��:�(;nм�7o_k,���5��6�
HF�ӊ����ᱪ/c�j��P�e��T��=���mz��f�0�Q&՘�'�E|�q���<����twsS�إ�Qg����ks���5�T�[ƥ�_���EM�� iM'�	2v�xt��]8�R��S����&�zX�О�I�f,�ؐ���tz��k�F� l���LR�Y��MN�U�jݳ[��j�y=Ic ����rV#Y����Oe�<���Z޾����4����Q��IU�K�^�8{�Յ�K�9�m7���\�wN�s��?��k�u4}/�����ڲ^n(J��ʑ�i�Y��Շ<I|/[���25V��୏\�}>|a�~��Ɂ�|%�}��4NN�k�pr?��o�[^��@\=w��ԲBs���}L�kЀ�1�㫛�x��z�P��^����P�L��:�����E����0�`~7+x�-�q�F8j��>l�F�}#��?���ǲ�r����k��,bw9�M�@ri/��0��F$O��ը�P�gp�
c�����o���a�W�_ˇk��qM5iFû��WǲE�"M���@q���J:�\����hF��:�7�[|N�|i�B��yn,<b ���\@T�Zc&3"���g��TV(���){�#�9���T���[y�v+��/�_��W�J���/�?Y�6Z�]h�x;�YF�'ȁl�K��;
���������5�a����ۺ<���!/3j%������e�<�J��g %�����qO� `�y>��
�z{�
��M�!S�d��L�H�`i�����4��i��}������a�I}S��*����Yf ��퍼~�����Ս,أG���ӧ�������NLE� ߩ;�@�4>	�J�`]��a=�����Id���ڐ�N>�F��BW��8�2��]���r�e��AR����js��$�@���:5�(��`���tl�����3�V�ֲ���B�W�8jm�$h�� 6���A�����D`Fdo1�Ĳ8}�W����#���n��A,6�/:�l�~��0^sWc ��v#�M�eI��>aUγ�B�KǛm�
�j)!o/�l<�0'_��<~��J��f��!`�lP*�{qa�����.6�ʬ5��>L���� ̦NZ�S���k����#.w8��������WZ�)'���,&� �� �����|�pKX��>n]�)yܗ���V�%���	E�X��7�۬E��������
݅{���m�_ggT+�f��r;����;@��ր
��L�2�5k����e�p-@�/��B��c�j:�U������G�w�Ғ<�Λ� ��@�\�#�UΏX��v��0�X��de~h�=A!���M�C��Ί��c"X�8��۽�n��MoN��j��dL�߻F��-�:�ćN���r��§Cw!�ۃ��?~.@�Nk���V��ۧ���$�X3��*m��������f�3Fu��C6j���UxXz�SB�Z	#�k�
�z<�c�������ƈ_3;E��K�� � �c/�q]�O"���������Ъ����%�݂��.A4�����Ϡ 1@��p(�3b�0U�d�R5F���2�h�`cڱH�������K7�.������k�������;T�y����\��,�h�,S��P*x�#@����8��|K��c6[GâL]k7S3��{�[�M����k:�8�?�]���dV����-���o�j����=�:�'�.��9+����Z3OԷ^�Ϭ��;�fXj���-�I��i�_��{�����1�~hj����ז���Z0\v�d���G�:�F���rN���^Z�>�1i�v��.ZM���M�:�`���: ��b=�X�Qn�"���{�>k���y���}�N)��̌-�@�1/�h�o�2`�}�����S��E�I���?��'&���/&"��G��ɏ:mL��k�cԢ���|�]�M=��c��u����b�H�:O_������z��NqoL���πx�~`�[uUu��{�aOɃ��M��s�F���ˋ3�}V@���\&�LTZRƫ�d�rLpH���h�rC	;�h�-��x�d(}�Γ�Āsc5���	b�2��J�r��0ۗ(S!�txֶΔ��K��y�R1H�3I��u�-�~s[�F~W@�O����y�P.��]��Fg��*���a|�9�q���|����F��W�ѹ�������p�ՠi�r�͌����lb㼴a�u['sÚ����>�$	�xn����S7&����Z�-2�����y��1��A3�~*��S}&�#]�d�)ƺ0y�v��2F9X#��,G�S(�>�M������1c��w���k���M�=Ǧ���^�e�Ym�nd�w�
�s:�&�wP�CLrd<����|�9��ģ���N�E��iT�~�v�>^E�(��_xU��T$�U�fe�����
g���;]k3��^S��ҡl�+y�������<;y��\x/�߽��
��x�a�ζ�����`9��&^�h���>�h;�m�d@�b]��GVo_Y(��g�-��8���������1�cd���h�(�@`!�o�(��Q�6;��H�kcI������:;�X�<����ysnƻ����{���J��#�	�:'���@���(eϨ
�k0VT���N�[ք�������cşi�;�4i6���ə��藦�ڠ��Rg��{��h{�-Y��J��#2K���sp���w��ka�8C�hud�~��6���:����TVdf��6-0�q�Z�Ę���ު�8���1[~78��/<N�*%���c�F���Ж@s�0�;�p��0��Њ�I�bh��LB��4���	�/_<��n���\��LUo{{v����φh$��1��$D��9t}v!�7�?��u��]�A���>�H�X����06D�)V|/d�!��(^@�(;&�7�
����,}��u?X�뎮��~Cx7-���o��l��o��Voz��-����������M<�*�Uʇ��2y�Ɋ�,e�R��&�l���:d! <Q1��2�?�0֌\˖� �F}Q�{ %$ʙLE��d�{����w77�^���]N�4�ݼ v���ߌ��>!ca�ٍ�1��N�5����bŬ'��Ы)�7{�j4r�pT�olFm]��=ۜ��x� �Tpehe�ެDp۾y.�4����6���<4a�	�~6/qJH����\�\��<ͽ(Y ���FR�=R+u��_}1K-�k��dN �G``y}*��b/�l�)���;U�ŪFĞ��_~N�� ���R��L�}�8��^U�!��[8���Ǟ�r�a�6�����a���ň���s��* y���Bx�Æt� ª�R�!.%��,h^@^��*8���"5�� t� sz�Y10�|��Zް��!�_Kb"v�����@|�\�P�a���_z����ծŊ[�뙴�bEW8 (N����-��^��n��%@Vf����W�(H$m�BTP�H$�o6�70�ˤ�ܟ4��)�̙�;�۸ʣO�yɏ�*�rU���^ ���=����Js3j���C���u�h�P}yAW��t{��B3��^�|��'J$�W�|����
)�:XJA����{��&k���̡�r �l���F����}p�a� �ڬ���a�UJ��1��>���9���;����|�1�G����(� �r�@�[}�{�p����^�/����۪`Lzh��i�X�0�#b���Q�TT�cO�6v/��`����X��(�3��k��[����E���Ю��yn>������޼���+�'qL�}�m8�����3q^0���((�}���I�V���)��Q�sk�@*@�T�#5���fUA���Z�`���\����yZ��>Y�9� 񘊷��J,<�\S� _������$wsa��\'#%��X��!��˹u�$�E��/����?��l�q���P�镢�,��;�J�4	!��Щ���W�<��>G_~�)}��]��ɼ2����a�H�tqq%c/䟆��^��7�/������U��2�p8����@��ɫ�̋@fX�{�㈜-�M��_׺MqRi"��~4���a�Px��j����NJu@qՅb�U����C����;�Y$KD��ի���'�����`ȸ�N-�yN	ζXOyO)�_2�X�O����1���=��	`��Z�3��O>��no����^sy�s���'�CuC$�0�S�q�舯9!��
�щN��!����Y�M�R����B�;H>�*Y5��u4w��W�yM���f
�dLu�*a4Ʀ5�_���b��	b��Ψ�'o�̯� �<�hd��*�Z���&L７yi�VOƀegQ�"�?�لB�Ǜ��Mٸ^���uĹYFN �电��U\���n�]���5�j�_�ni�J��<d��B�Yà2��S�$�K���y'���j0J4)�a�ȠVQ.M�"���g��;N����,���;z���>��}��s����O_��l��8����q�v���n�"j��i@nZ����
��A>Eyʨ*Xd�����<��k2������qC���^��r�{
jGI�G��68r�ە�aA�J���
�!5L�υ"d
����ԼeI�:S=H<�+$�����*^Ƭ��AK��� 0��RE��I����Q��@K۶���3�����H��ŐrZ� lF��a,xMV��Sx�Tl�s����MQ���%�����c �JV��yXϮ/�zA/�_�#�S8T%+�� �W@]�j�	���g,�e���ظϧ��Ͽ����������w4�>B�kK�R��A���6N�c��{�� �j�o%�<H�yJ�Y��nn���!�'�σ~�Uy�8�=9�~�)�|�B���c�p�������Tf�*	\���=/�qO��F��WAXﺎ{}���$�K���-�Un]���k������JΟ!tg�gJ�Ai��o:o{�{-��0�z.�5M�Kj���k�����h���1�8�k2�]�k_�WM��	W��sTK��O��O/
V�ZE����|���^��|������y]�C�(׼�J��A3:Oz9��r�pT� ��U�s���:�h3�A��ӜC�W��J�����u0O� 26�n�<8�/Sk>���@�s���϶��7�&�|�&�*D��D-�Z%n߸��߼��o?Лw����U{��z�L�l��B�_0 �WN�PXk	�r����&�Z�E� �hk�A��{�Ș-�|���O� ����4����~�wts�2Z.� �߽y��NBF�݃�4�]�x��~���Ӂ�W��~�\���އхQ��`L#��Z݃��L���������D�B���M#Ӂ�bA�r� IeF�����G���3 Z�e��`��2�u(2�t����-�ͬ���P;~�" �k�A(?+��~�]x�������*B�̩ƍU_�xFϟ_J����B'"T�8����������5Q*�י�$�(a�0sC��}�����:����o7Z"�U𳱷�����͗��t� LvKQ+��Wfc��k��]��K{�U�j}�(*f�	�P{jte�>}���o�\$_
�^�?��?�?��?H�s �̖'2�5\VoZ���}�>2���^��	�S�|o��:qO�$���ޑP!}p�ëW��y���~K?��Z��xN���߫U��T95D���&���#y�v]N�9�=�$g�+*)�|�y�'�C��X�{��K�O��:�@֊�8�\x�2��{�]��œ���q�����Z~m�.u��]f]H��*��Şi�3΃�\0��E@��l��U�b�Ѥ�A��/�����s��S�t=dOϨ$�KK�:W#Yզ٪��{�ϷF����y^��i��E0����֐&
�%�C˴qް�2�ǹ�R�^�p�m��?DUx̍�(�Q&�i�'a/8h�$�}���NX�z8���{�p���_~�����.�G)���n�H3ҊFXg���e��K[éW�F���@��s�D;��Q�c�������h3��w8��u�~�K2gN3 �?<HK������ƀ��(��W�]��_b�1P��6�ݑ�T�B������� P�>��k��ox?�m@��j��/��&j��Q1t��8�'؊/q��`��gF�(=2 c�x�J�[4��M_]瞘X��@��z�Y�M��&�SP@��i�+(?����m��ۈ�1^>���/�%�=T͏�0��2��A��� 4ϵr��x��J�Jy�>�(��l�M���M!� :Hz����1x ��U�q��R�EH�mW�Rݻ4A�O�Ϟ�i�Q_ ��ԠХ
���G��^�eOק�~F���o�����_j����bG����� ��J�!��<������Ŧj��[���R��G�Đ��	U�&os#n�~������%�4�	`%��}�
���N�U{��<�W�T�E�����`� ��9~9Hji�S����7�M�}��[ȑm���7�/�-ɥr���ze��Q�Rd%�lF�' U������ū��u��#��UL���������3cgp�k����[�j;�! �T�qJ�ѨDYUK�iV� l����?#W�Y��t3`����-�YG%g��%g#9����ʚ�j�'tu2`����ż�I�[�$	G��#-:�4�C34ճ�Md�R�8�� .���  �ӒX>� )Z�Z	"7<tv_	��ָ7�s� ���⸤�RP�@��5���Ò�vg�7���pg4l:(+a�`6ʂ9c��� ��9�©�mS��*s�~����6W�ϭ̥�w�VpL��$%}G��pZQ 0�O1%��&��g_�N+�40UV���M=9�`�����0�{�M֭�/v��VJ�˰�A�/PJ�1ZȎ$�l8Z(�|��)�qK֥y N��c�<?>Cٻ���G�s�"�|y6J�য়<� ��6)Ը�b7q��ä���z�¢0PfL�n-�l�#��@8{��X+������J��H�y�L���L�)����濻�6���0{M1 c7.[᧲Ji������	�g��j�~����O�W�>/��nWWW,���D��g��׿�/��B���@�+�u�i�`k�h67V���B��Ǡ*���-Ч��c^��̞��^k���)���!���!����^�����N�	�x�[G��`�?	����x-�A��'<�,�ʤd������Sn�5�Z�mW�j:{�a��m>��������sZ��9�d�������˫�����|�~x�9h���I���ݞ>����o�w���V��yUJd�šI'��Oi�/*�S.�σ�k�Vos�$])�pq��Cѓ��)x�&S97�����4HD:����ːs3$��Q!�� c*_���g `����V9=�[T�󱈗k ��Z���#�(�V�a�g����s�=�=	������|c��$ߣ=W�5�C���\��ԃ�5�����ӳV#q׎��ܶA��̈��|����Dٱ�o���'cfwf��M�(�E�վN����B�rI]�}pl�,C+��@�M%U����,����(��&6C9�
;e#��l��~F��I���Sn8�*I!W�����~,L��e��E����&���kzBLj�%<��s,��ڢ�Ž����'_���`�Ū;�~��J(�oNN�g��ų+���D����vg*޿������}��skGKA��ު�.�3���k��p��������`x%T��K��ڍCC
����5 ��֡/(>��;Kn���r	?��og#U��I�Wϱ0���s1P��˯x��1���.aGX�k �ILH�5����g��G��b6Nw
 ��h��~�ۂ��D&#�Խ���HU�<v�?���d���o�v��
V�~����xto��X���p#�"�s��>fk��m��� �X4�����Ǹ!�j5��8y�8Ο+EL
'�8�ބ����[h�}�g ��`�����8ɜp����ͣ	�S�b��6�)[�b��<ӣ�,�D�%#h���]C�K�N�A��Z֊5>����z8Vp��A /PϹҽO��#�g4����\N(�:۽�sQ���Ƌ�����@�-X�9C�#F�3�?';�������Njdp+:�;�8"���hƤ�KK�D�W�܍(*�!�(���4\�/�g�W�TUV�J��<�p�~��;c�� `��'�p!��qQ�4�Z�*�A�����O��ʠ뜆�%mΞ�������L��V��KX����R�	ax��T<��O���B\�,H�䥥���Sĝ*]P`
��`�}-t3��N�O�#�Aތ�[a�*�U�Q��Ę<a�{�Е F�9�ѱY*'6,�&�'N�}B���D�6���@q^l���������Й��p�邉Xϵ���o���޼}C�|�g	e���������}�"����T�^^��Kڝ��eXoy��������6��{�/��JϡUf�V���@�^*�A>���A�>-�����Hڄ��z�a���(�3��ʟ=R̰�7�1
�9�j�3	�]__�O�жF2.���U�����AL�81֧�)���\��T�������5x:�	3���5��N��Vq9U�^+"?�����ݕ�zFY��pC�߿��`��ڝ��97�_T��sR8�߳��{n�,ǪB���K��//�]l(�{x�-�%�cv� �bm��A���b;��+X��J�����~>?<� �q㜆����sΞp��>��oNH[��? h5�
x�ԙaCm�����(FZ��+"�tqh��)~�^�� �&��T	�1]fa�2	�f���|�eZ�1 �k��2.GK%1.B�J� �c�{���� ���fe*��sEn�C��3�Qp�����g�ϣ�MV�6���P!leM[g��I_�jI�M+�������֒���SE��][$�S*�s�������S ��_�5�r�g.
�d{��S�W�Y|���abB^9��i)ƾ�y���G�(ab�&��GA��A9r"\����^�����
G�$� 
 �ӂ5~���9�9�h[�=`��'�Ea�d
$>�ئG���JI!���Dv���lה�ɍZ���߇�u�*���@?�tK�o����n&B�؜$A��YI�Ɋ�J+Y�2b��uA;P�(�ZZ�����>�Z�K~�G�;*f�p���%����d��o�z���؅݅���}����������W��si�
�!�$ȫ�i,Ċ:�2�������*���Ri�`Ƞ��Z�8,�ǜѦYh�(�Q<�$��?���Rr�>�V\ϸ��6�UХd� _�pm��.����K�ZT��s�)�-��0��
vS�ݚ/�!��G@��8A{|��k���ս_8�GT@s�#��@8��={�߽{+�j�f0(������q�[���^
;��D���o��9��M����A�������d�!�^�%�{�k�A�S��Eֺt'@��y�p�d3`����k�`�F�v�����.��O�%o��A1�5@���D�3iG4Y�|F�*ya[��C:��H<"�(d2Ϗޫ��bt�U�CJ��vy��J$��
Fv t�]*@��ɳ�c��	6ɸX�H��,囿݋߰�[���=���[���g���e���a��Q�k�}>)�94m7�8�+D�s�ÝF���*R������#m��Y� �M�x����ߗ�M�>�m�qR70T�+�����VHA$��hy�cD�ћ�r<v�7����w?��;��}��I3-��S�PT�o1Ņ�Ő�qR%��JM���fɀ��l�`r�੒sۄU�l2���J����HLm�p�Kp�Ѫ>ɶ?;u� v��.��h$�6�i��뱗 H���!
���s��G��.BO��R9u/�7Wx媕GׅgQ�Au�V��9ʦ���J����;z�ʅ���ne���'����Zr�������篤[=~��fc��7��3�r��U�2Sr٫�ao��C�9A�ɱR�����+�bX���m�I%ǃ������x�_�W���yY\����2����"D�C����
��
B]�do��Du�*�����z��X\ٸ�cZR�O��S@�t2��1e�C������� �"���X��#w�|�z�«զiٳPA��BMG���/�͇[�����?|O����_��c��<���lNk�B�1��Pl&!�s�~QQո������|�wf���.�,�f��`J�>�?u9����Ez�ם���-Z�p)�T�U�8��Y�����hZ�?��fҊbai���t��͙T�1�fl�B�1�l�y_�f)?I�F�yZYƊ�m>H[ū��1������G"_��ߒ�6%�dk�Ĩ�nxf�ll?;5p��v��)��%�<o��?�֑3�d��C���YĤ	>��S�4t�0�vb����

)Y��	~"�nu
�P��)��VJ�I��=�Wr4�{&����F�fyM��) Ca�8��+�F:��sbkf�(�h?}�
lY͍@��R�Ęc [�~��ڐ���%�>P��:��EVK�� ���&���zl�Tk߱��⨣����/qɂ�U�ö�P����O���M�џ����ba������� -���[������K��|�ʺK�5`|D*��#Wyi����q{��o_ӛ7?�r`R����t�� ���+��w_�?���?��zv}���+�F̚&����i;�/Jc:��;Y�#�>���l� (�/��
�m�V|W���3N����G�SB�#���_��!L� ^k!s*���딧g	hs��|cy-���$�P�~~j��^W��g�c>ߏ>��@Xzߓ;6�Ҽ^i�a46:��Q�O-�^�3��� <Y�c/�*��춃����t�����{�u�k��}ʤt?��3����K�nz�������10.�I�� j����h��̺�k_a:�g/�<���޾yK����J��o�& �����h���y���7�LƐ)�2����k�p���Z\�'@����<{���EF���f�Q#�F�K�ٓ���6
$��,'�F�R���1�����-�E��B�Ej����cަ���6���:�?8X���Vq��Fhn�rx���$����Z�z�)<Cz���l&�淟���\`���{c����{��*Gx�t�=���\["�[����sܦ�z�S�(}o�A��F��T/����g#��f����᠀�O Ւ�2���Tx@����	�	��(�E@i����G���TuΩ/C3�{�?���x��c�}h�`��Mp5f2�qG�g�حp����i,���������e�/B��T�I�O�)�����E��A�3���qI4�v۳B����MW0���z��������7?ЎC+�ط�\�޾/����+����ě�?~�?���V+���7��n��x����)7:c�s��;Y� OZ��]	�7��k����#��^A�}��'�����G��%���3q�w5W'.����K^y-e@���58A�l���ầ<`k�������<ZO}���ɏ}�;��g�5dU�2���7��S�Ns��a��,zU�-��%��U�O��o: ��o��
K~������O��~��'?��e�x��S��H8.{O��;��A�%$'9j�=k��i��x-����С#�c��Y��`�������>V��Q�����~9���<n�A`�ۂW�
���PM1�dp4��KU�꫒y�s*
z��ig�)+�����߲��¡���p�]��>�H�]���uU�P����<�uPH؈��H��d0�*�"5�yR~Q��b:{�E ŝ����� i)�(9Z�����ߜ�?������5ĕ̈́}Қ��������w1�z��牣#G���3�y�( T�'�?�f����&���%/���B��������~_��7S�tws 新mH�v�k�t1��V���QeУ��HKv��~������xүZ����Qbg�DjvJ�v�Һel�Wc�Ee�S��e����W�� `��V��#�<	L>�ǔ<�'�( I<e����/���
e���ao�����Y�`j��t ����qG���������K�R� �������J^W�.��@�t?J��=�l{�s��jʛ��x5Q�oTk1�~���k���O����������mg�����޸��i�""(���(��=�{V�v��z�,�'��4�����=^�0�z��%<X���TK$)��wI�\��0^�x��B��W_�u�;��0�/�bG��r�K}���ȟ?��P��0��Rt\jo��\�����Q=�/Ι������ͷ߈�Q;��DB��{�y؋a����M��7����zl�F�@���A�\#�3i�L�%ט�]��Pm�f:�,��Y��ە W�)H���9���ޤ�&2Wss�joA����  r6`�2�K0V�80�+b�af0�+�B�2��X���Jx��8��+������7�/�{ �ꄸ�z�23��)Z�3X(r�0x#`���N?�	�D�0��A�=W�l�Ҭ̖�??��ü��A���ѧ��a�Ņf��Hp'Jzn%�ܷc|!�4������K"��/)� �1Ư��|=�?��}ɹ��[��8�l�6Q�
���>[k"��f^���/y�2WJ����_�,�����f�o��O^��q��yZ���%G�۩ty�=y�������������M��W��)�÷l���#�_�x�� ڥ,��~�)��Vfl�ٕ���x���d��RI�hH����s#�=�*(2������T?��l������-�'�źjI��W�ɾ���́;��ڹb���ɻ�"'N����- X	o�S!�_����K_���O-饧-���~d�V���#��`�m-�نp���D���k��D/���s�OW��ׯ߈熓�o,ɟ��c>Q�6�m���)#^��ʻ�=��˟�B
+�ј�@��+��n(�p�ҩH�\�3���[`>|�or��W\�͹y�f���_�8R�h0�K��8��ܫ���3�;�D����Tn��F�g�/E��8�H�SZ�|~�� f%T��s�ɔu3����7�fr� !�I�YaB�!/
+D#�����1ĺFU.�R�S�r�#	9���&`ĺ)^�Z@�P`���Ѹ6%_{�!��f�<U F��Z	�QK�.�!�{FIw�R^�L҇��kk�(�6nuS�>+ض2���l _�<�&^!��׶/,܏3��n�ƙ������LEq�|?���7����;����b�B+˷�� ������=���d&b�#>�) `��g.v!߫�� h@��a($�j���-*��40G%Νu^x/'#\��WŗA�F��
��S0���iP�����f��E"䴄�+�X \\TeO��s�!����&�V�%���i���$�s8෿����v[��RG���_�*���&�rLcE�y�.iN��'9U���Ek(T�82  �=������!'A�pwKS#����p�l�rͣ�:�5�
� .IЕX�-���x�{��+u�ﯟ'���'*?�)���|U&�h�i`�������_N=��֬�J�UI >� b�pO���o���'�n�4t���	e��rJ��<y� �"?99�1N&T�C�U�]��gtJs��^��CVs(!�.��t��^0dhUt)�VL4&	K;�)��h�B�<L���
PhwX�2��I����`�R=�G���5g��G�%}�9F�hfCI�FsіV`�����4���\'�o8L�������Ϸ�N��W!����������b�T��=��5�4�y���U�2s�S�UJs��r-"���	��V�s����3�!�"�6�V׏m�N�L���_���$��Tǋ~�FXz�M|g��ݞs�����Hx�bq��M���jij	Fϯ���'�C�\[JhkX��-欵�$�E^�8Z���eދ��!���})󳸀�5C�p��������}�j(�f:-��n_ x��6F��ȑW ,�	�dE���S��o��}pw����:pxF�W�'�c�p��X��E�m��n94B�:�s�[�������	�+���2�]����T���c��s'�%J�5���?�!�ɾM�#���*~�b����~�������#�#���ų<������YVW�Ņ��~Zc�G��G��H���v�����7�>���(h^N���y��%�
W�6��{ZQ��i^�䧎au�@��0�dtD����3�ꫯ��~�sι�8��B#�h(�%)(���l����`�����"}�\ə�U�5:�����Q�Nc?$��Wr��nE�K�����oݫ�H5�r�i>�%�%%k�_wH������Kօ�?i�fN7�ƾ��̖�L'�$Tu���3�G�S��[����w#���eT�" ��0����D㾢���D�3qNv� 9Ն2���ʐ	��b`�f�$g_�Ř�c��W�sq����ʲk��~�۲x�����)�n�����<ijls��f�s|'�?ht@��\��E �$o幒���;���*�N�$a�l�vS _6�d?��+�!�0pE�� ��#�6���N�V��H���$ ������8��b�:�7�z��p0��2&��c����:��ŻN�|����EN��b���ŕ�`�MI�l�5��Md��.W.k�v ����`^��ZW5%,�Мp�4�9����av�s���݃�dc3�Z}��a���ī-~,��p���%ݲ��T�U�?�O�2�a���!�O�R�Z����9_��ƭ����#SPHB��G��|n��q�i���$�E��q.<8f�䵗��c� =<��	Sx Wwtb:Kz�|��R��m��rh�g&M���!T���D\��M�-"5ؖ�?����`P�@����-漘�=���K�C�M+��\s����֞A�,�>����~&gc?(=�q�)���O�����<+ǥ�4=�/\�����>%�=3'�W��y�܀{�9ƔDL���ȸ	����e;���Y�� E�pLm�PEZ��wDU�����'��{�:@�ļ8�ftO���z�*��.d?�oŹ�q���XdIV�V1�<���/�L���c�/�@��r��&�%&{�I	��,`8Sx����Ț	���>F����m��ҷ�⿎m��vm���ޔ3��j��A���<wBR�`bz����'�����J0'���\K��T�����N(Kz�̾.�SC��qh1�����B�e��ԏE<�.�͛E���2)R.�9���%u��i�f��ܿ�P!Lhw3�@rEV#N��M��ToJ�	�<��I�N���E�F @����4�I
BYɒ'Π�=*+�j�ؒ��i�u�f]�qU�V�G��.����ܗns�1�%�����(&i+�:�yj�IHz�?Z)ޓypz�;�8�r��~)��%hē�Jm��@�J��bPE���m�=�w�  ��IDAT�/fq�`�&Q�4S/Y���� [�7p���HK�ܿ�_-�2�*�u���Yh?zAa��b!�Ņ�3�y<�0@ͣ�ԓ��a�y�}��f<m����t�8�lv��<GG�tj�5���C����� ��V�V��H���e,���h�3��WW��ó��5a�bc���ۆ�f���/����
���&��Z5�X��j��b��5+¦��qZ�'��>��]x��#y��#s�m�k�C�¸���o�Fǭ���`S��F�>�5x���P�5�U��������qVORQ1��")wO�P�aUʺ��k�ж��٨b��w�F�Dn�׃��7
�8x���֋�Lwȡ�A"�t�lTsG i4�є!mvn��4oN�����wN��K7Y�%�k��c��)�z�>s������?^V�;s0Nd�\1Y���

�����Ǆ���o�+:��e|2S���	h����U�K�#T���DW���w �@�j5�M���ȗA���L����Xh�0������kh}�s�������~��$U෎�Y��$�����%e{%/
��t�5���x ��4K�`[���Ul����D�KK�)-���3��7�l+���� �I�����`�����c���"m��ذm�5xT�G3y���j�Bk� ��&W@����&�uj������G���<D�E
7X�X;b�/��*�yv0�𲆥�HhB-f�*���z�-�A��IX�Ǐm��<�G�J����S����k �T,x�kX��1�<�)�N�\�[�Zs�$�2o��^��,G/hM�<Cn�2w+<���I
r1F�	(�|��E>g>C��������}A
����w�~{.� ��W?�)82OEq��K��ilD'4��#,�m��%�\)��������X�d���(.�+nU�4�������w��A�`[=�gGr�AU������R�,�N M��� �u=K�L�]q�9�B!sq=�ywƺP08� �����u^�}����8���H�����Dc6�6n��X82CUϏr��q�&?�L�C�s�9Ɯʺ�]z�K�J����L#c�����̋�(΃��Q����!�|��*��0��y�*E��YR��}J^�I���j�Օ2k�V��u�jS���J��t�(͗
	?��tS7��K���F�E/�f���dt��A[霟��7��;GpY)�=�Ż�j�Yd�O���N�2����.'=�4���h�˒�t� -�´o��5�0DE���O�d<��9,!�R����˸�u�.���_���޼���[�|��F�E�C00�b��(Nʯ�R�+����Em�C�haԻ[��Tt">��{(F>�����N �mFcヵ���4U��X���*s��M�җ͕�`������/�~�#:4賠3D�P'<�Rr�8�P�� 0�����"W'���[�k��4���z� 0�dE�w*�h��Uf���ٸ; 7�Ӆ�ϟ	y�$�^�z���.K!*R��I��ZS*�4ԣs���A�����i�ǅ��Z��S�2�Y�s�z�q`όQPQ`���gN=�н�+���_+�V��"7�� ����	!;���&Ş%N	�א;W,"�����?S+�b�T� =�X����a~ի��X�Kˮ��!Tj�QdT3�1U�d���5c㌻�G�� �WB�f��tUI��س[����쇹��.���M���<�os"��0�����y�T��o6�Er}/�Z�y�N5��v�~��Ѝ������-3#!q�\��97���5�Q�i˵��'dh������˟��|��U��X_LU5���r�7Ν�<=���ժ'���`fWD�+P�Y�Ӂ��9�����#����1h�g+ި�*��NBB���8X�ɲ�!m7����ϝ/%��x���AAW��C��d���Ô��Ά7�e ��%l�Ǔ�+@i��r1�b[4_�E�J!(�e�����J���e%�#𴤏�4�`з�[�X[�o���
`c.~f�>�� ���%&$�O�v0b_x:`sx���'��6�~�,����b#�����\T�!�8�hK�$7,�V��)n�-���;�zH`�Ew&���tQ�N�T`x�,n�c�}�<��ͩe�V�K13���	Q<g6F�Z����9l<�b��9۷�A#`$9?R�#�w�P���b�����!q�p^߇%M��&��fiά�����vaT�$3q��&R��Qr*��0��2y����fs�tLav#�T�&-'�ǈ,$c7+�(,
���?5�����L������h�J����Ώ6Z��B&rx2�J�F��¼�!��F�������} ��SR�*�I�K�E�K�ָ-���"�Es{6Fd�k���{�K>!����呴Ë%�o�8-.�6t�����|x+-���o��_~JWϥ��y����"f$|�^�Q����� l�#�3��ECe*n6@|l����q%�y9�_i\T7pW���S�c�)@ج�	�tcE��%$������>c�(����: �M�O(\ճOt\��Q���')ɵh�{bחX���+VΎ��6�:{ �":s�%�<�g��޴�&I����ч�����i��˗/���K3'ڻ;A��2Revd�d!:��}��ڲ�G���9%x�B-[�x���c�_j���_p�,�]�@�=�0��5��hӐ�~��[� �l�o\��p{���xB�G�O�}6&#����g;;N�vF�a�VO���OU�8��[p�L|�"��RQƳ6l� ŧ:X�-B;���V��ٹX��]�p>��QWw%�˿�%,�j�ǰ��9zsυq�	G��x��@�	��<.��r��+�jZ��MЋ�||m��-]��0s���[Fn֪'�'pF^Q�3݆Y����EEb�ߦ�̅U�B+�N`�P!�d��X�iΖр��ϴ8/@*U~���� ��X�5܇���]�d2�jՐI������,�'@��ax�g3��:��s'}d�s�p~.JW-։$���XjP�sCU�BZ����W��Ps�7�'M�߸g/b<�1����Rϴ�O�����5�:��n�I2u#tg�q!��j������dl�~�{��ha�d�����q�L�</�����i�����r�AX�&����w����þ���+���W��_��~���Au<���Gί-�(��/�_x�5S�Ƀ=�D��tA��A%���� b'^�#��L�KN��wj{�ɕ�VZIqJ�Єۍsȥ+Ar!���8�ԓ*撬�Ƽ�E3���S<a���$o=��`�g��PB��cT��Y�1�0���*��JF�OQ^����� �����ڷ{z�pG7�����A�g���.������� �o�yϔe�IiyM))����e�<G``���$P>�Trz����-��ɍ�)]���T�le���L�=]�ϱi�J��B��Jݠ�]&J|�����{�����3�W;����W�w�C��\7�� y/GM��V[_L.�W�b�ظ�=�՜Y����������s�8&dV��x �!0x�!�8U(`�W0wyI�iL��   ���Ѫ�๭���,�9#i|�� T��C�xW��=Ք�A
(�h� T��t^� �A�g�Њ!U��[-#or��m���l
�C�����/xB�8j�c�YA���
mR�L�ne�u
��p�I�s.�ѣ�=��	E���-�˥e����z��nR�w�u�ī,[�}�:!���z���'��4�v������hۨ�a��C�� 5bL�^>���R��u S<�	l��n��(0�Ii����=��%�Q#�J;��xq��3���t��@wo���?h�݃�TzvyI��@��q��f��{M�ꪆ���h�'<_�Y �����������ǜ�o��`����M,�o���C#��k�)����l(FV�Hk�d���N>"�[~��p�B`�dBXv���6�<�XVřv���;��"1��=�BXY5AJaG�
V�$�Zʮ�Ͷ���l����St�����n�����J_\_�5�>�z�O�����ݞ�����v���جn��K��\�%����T%����b�,�@����)�^�K+<OPs+D�ĝ��5t�=�I�f�W}��"|߿c��[������I������4�������/?�j˖��k��^#G��k���C$�*���A���b�����A��>c�M�,����Ԅ1^� ��F�Ph-=�r�๠�jP��;K�c��>

��Kq��T+AP��@1�y���n%B���E�vN�&�G{����߻����.Y�x�ve�	a���rc�D%�nn�J@��)��s�;`F+(IЮ��d��r~v��1����(�
���7�����=cq<�i��9�!<h�����F�Y��N��vN-��^��ϥՂ����sr�u\��o�vH*7�ۧ���6" k9�xxJ<i�64�kٗ��_?�����Y9�R���TR�"|g��6���9���݀��rդ�t������&�wn��@
�Ր�F�qN�+���(3���`@+Ә<�+9OX?���B��!��<���Q��3��͞��+���m�<&	G�A�H�^�y���n�Yv~\\li~P�2"1���K]���@�@�SD1Z�,V�z����G�����ad���� �?W�2�:�p}��ڌL�T�l�Vu`��������RR�ְx���u�VpY��z��R^#�����S�F%���l�7��i��K��i�ހim^Y4Kן��9��F�:;����B��$;�4�Q�����B+%���j7�sc� ,+�B+@�唼˜��<?�RZ(h6����Gsd���]��2a&�� �s��{l�h�B"pg��{A�=��~��W ����Dw ��+nm��o�GI`�7�'�O>�}�R�����HV�@'K[�2FnW�!$�T	�'	�B��xv��6#?:n�]��Ŝ=���Q����2H4ݛGk�sNW���\8+�1"O�'��R�	ɺE��C��Bŝ��&�2&K@��]r룆��'��`{�����
0�(��Ņv-6F�9ʵ9GV��9�K7ܤ����jI����X�>���}�"�$�J!����V^V!}<6_3��`��r-�0��f��Jc=QR����`� �a��H�9�G� ��
�}��D���������O��m�2�5�O��e����~��L�7���.�Vh��t�k�%IY��R�N���<�c9�Ш򼚶-{'� �̋(t�� ��q��k%N��U�LI~��Yߏ�T�������a'�j#�J���F�p���}_{)���d YvN��%:�{��3�P1��D�F�Vyq��w5��7=}��W�g��Cl�ŞA=�F��;e/rz	�"+�� ޹
���d��e"��ꤠ|�7�PT����4�.�[<�b}A	`#-��0x�|8
@�9�09���;���R~0�Dl����k6}���'�>�ˋK��p+m���k:���[F�~��Κ�Y�^���Ñ�ީUίZ'+#��eq�c��$�O ���s�\��71�=���=\�bG���Ɠ��
>�d��fBr��' �h��;n���[J����+�X~���t����x`�����*-��&�*�i�"P��̸�Q�9�ps#��e�"e�G#b�[��CJ)�_�%���:ߎ��4�Ζ?UlӇ�ɝO�������%�Y��������ݽx����~gU<�@��$�m��ynSX�_�	��oZ����k�w)��{�
@f�#���f�=>��`�0�6�fy��A���CK�cB���.IFW�ǂ�EyܒgzeT���3����vcU���&+�j�������{����1�f4��[����JU��G���^�ܙ��+o��C�Lv�4icp������󪉷��m��![��,	p_�������s��]�|��7��?(�0],�`�X�n��|���X�{��"���6GT�h6s(&��Zݐ�����Jx
# h�J"������wO���C/�p�����z��(���!��N�����dr�� ���<K/���Ie*�3�:K� ��2i�q~��M�9�����^f�Z(&�0_��B�D�Qț��~��Ic\|-����V9��	I�!%���-S�vܲkvA�>�D�(���瑏l��l*ӷ��7@|2�����J�/�4v\)sT�!��b��e�j*�M�� �&���ZO�X<&sb,� �h��#��[|ู�ߏ�Ƴ��P�-wJs�6��XQ��'S���D���X�r̨(U������ �q;n����`̈́��$�7n��F?N'W$
�$w��&Ù��@�`��ޘ�HccK�'��rB���2I��ϖ-
-���%+�P4'�_����t%8m~����!�� F<�=4WE�w0�s��=P<�����2�պ�\�q�|�10 ��� ��	6k�D�.@3���b��z�c��"(��G�T�m@H�`[]s��4kWc���p��N�!5Y��{<��g����Wh�O�o���ތ�r�E��\������%��'�#Ƶ���a����J;C��O��8�B�4@)�q�|+&j}����D����"F�ƀ6������jm�RG��z��~'7�z�qx���������;����P*ˈ�¡��,ͅ��0��I�$�� ��2�B(�,�K�v49�A2h�u����,�3�s�M��y3��^��V��t~uM��$�?5]��>�Wϟ��Gz��JWt4�3;x�� �!�k��B�	������8��G�s�:}�Asͯ2ޠ�M���!�_}mU�$f<�|7���-PgYN�d��@>�D�������j �i�x{����������v�;��o߾���]���+�s!`��㸺� �&�>J[��K�/�����|dE�C��ܑ B+���y�pH�_�4T�%k`�����H�w���R�ٚfP�yN�r�~��ƭ�$j��`����|+���|#��^Jmjy�ə��m�ґƻ]��s��͝( �);Z~Wk^_]	���������a�����H����M�GI�wPN`����S�V?�ʴɒ�Gy6n���x��]\�˵���Vo�-���zm���݅��V �U�{Q����s�|��y�q��Z�1��hk��w}l�q�},��+��<�H�}b ^gkPBD������͋�c�-L�&;�#��DJ8�׷�J�o�yU�i�{�^����^r�лP���t;3/�:��iEJpJR�˞Q^I0&����K���c̀�ז���G� *�&����d��E����u�D���oN|~��g^c�z\x����ş�-$� S����X �x����̲�dw���އM<O��e����IK-�g���3;O��k��r���ǜ������A��J5 "�������M����g~��'��.4�#om
0g[���=mʾZ�W!��8�L΀��&j`�[� ����+øe���!���:��Q��=��V�0Q8���l^?IC+��}�辯�����W�ҋO>��ե�N���Ⱥ5� Xe�:*xU�6���V
(�Z���'�{@��xE��G�C�z\�C5�\�K�_�o��HA�`��,[��fQ�	�e�m�)�,6/�,ð�C
�c,�b��ă�X�#�հ8���4PEq������3!{���Aԁ�?<�]^��EIu�z���'zǡ�����
���~WuNu���T=��G(�\j����sǤ�"+a�����\�����-�p�����#� j�-9v]���`�=L�=��:�=(�ꗪ	ļx�;����ŵ(��/��B��x^���M�s$��L���0`�q+��A�g��kaO[�Z����?9�	�Z}�I��h�\��~1Wη4g��>K��pSB�q<+�o��V������̠yv�E�%oi����%���E��(7�w���[�*��?��>��S��Ot��D
��w����rUUh�͹7[�ܖ�eVb��q	 6Z VE�wRCD`�Wʊ9�M]?<��so ���bu�����(z�RP�"�A����{t�E6SxT��������J��d���v�5\�4���'S!��;��"�<"y^r*���9-���р��{�8ٜ��I}�᾿'7��h��U^���<��M�rB[!YXǼ,��s��+�AI9��˷�$��E��J���V{Z��;�޲[�'U�u.������tܨ����x������������޼~��|o��H7�ݙ�	4<��qN3�@/��H�єr� ���"��m������$�=�58hI~/�����o8o��Aք���_��Q��c V4�m����/h�6N��1��:�zF�~̞=�L�֦T*�y#/��y\Яd��ȸH����Ci)uO��B�t`��-�WY��,���gqfZ����!���XF�b�%�[Q�7X���jV"*
�@Ia"��	�$�j�h�������?���[��yG�9�=���e �ۢȥ��Q��h����4_������������� rE���X��)���Q{d2��*-��A9~�R���p�a`�x�%�=�@���I�΃F!�Oܒ*�����\��g�4�~���
���H[Ql��'����-5Q�Q<����p�y����f�l6 ��?�g����K����(E��	��&��3�o��ܛ�b�^r�vN+��O�Y燽#I������G֧�,���faF:
�EPK .�f�K���a/��'�����c�=;��3 ��g�{�3RɃsQV���� ��-9Q�ؽ�p�n�O�e���mԯ�5������B���A7L��|���b"��9���P�l��s��q2/�U����i:8h��&����{R�8��^K,�����)9z�{�ڄV2

��V�u�hv�� �Vƛ��O;X����ZW�f �C\�|�-}�A{b8��s4e��/�˺�&�"o�,��o�-t4g��g���t��yQ T�e���l]<Ms�Jn�>y-M�V�)��fl�{P/���9�{�s�;��3 ��l/����}` �Ix[�^Y����+L~��x�3���퍬�R7:��� I����^��6"�y��b�@�+�T��=8X���}c��m{���~��SŻ4�&#��E�&�k�]{/C�����uK � ���2huJygkJ��Z��E�VS1Z+�ڡ��d0"�_v5��B��%]_\���IJ��/���Mؓz����[@�G���
��E�{�d\�Q��-2\��]I����>�)�֙9���/e�Ⳇc�;G�<
]�Qн<H����s��/�:�)��G�mZ���/`$�RC�L��C�2'����}����@^�P�L���->S�e����4M��d$J�(���1I%d�]yl�0�B�QN�m�3b���_&!dݙ�5��}��B�}��΁��"?!wgwe��Ox�j��n�L�#��q+��x���!$��W4T���i����2�Y��Ɗ ě*k��"56�B|Nno��+C�}���IְV]YЬ����Y����z7搇zn�ڀ��� D )�(T�5/�&��0je ��(����\F�}TCF�}���w����~����&��
�X�0 ���|Wv���,��Ãϝ�D�s(J�EQ�^��0h�x}��  N`~��-�I~�z��]��A��\=>��� �UAy��7[�$1i%�ø�	�g�Y����9��hU����rA)����ab=�),xx,�y-G[C��C��E#xɓ3 ���K��:�U��arm����<^l@��/����?��=7 ��:"�Qx�yN��Z�M�OlZ�a�Jr��s�y5��|�ى�z-�" Xg��iU���!����F�Cm�����A�V�$��K���HN�!��7!(U 6���FU�;�뺟-w���xg�9�}ќ1>������{�uU	y�8������N���m��U�`���ɫ�����@�� �/���P(�6Π `Z ��q5K]��vص��e]�������|=j*Ͼ0���/�n.%R ��FAԫ���\��Ç�O��9��+[��r��~�K�3�9�e5|���G���Ԏ⟁��
X��aI,G����a�_�|���Iւ	s9��9���*���W5�-9�,^��� �ң��{����h
�������ޚ-���h�k5�
,�K���C�
d9�Lyl�{��2 ;H�(b'˕3�o=y �9��d.�=��˗�b�y�z�򮅕���{�jXI��;n!]��; WKkD���2bէ����u'!V�l�
[��V���"�d6��K���V>r/,��"�7�����./��Q�6!�VBXG��%�B`����'�8 4%�BF{�MS��6� �竉!��܉``�V ��K�c��ҫk�4�RAq�k$��;<�L@i��)��EX5*¾{0z��{��B�r
r4D�a�����|����ˋQ��޽}���k�᧟�I>G5~#V�hg3�L���� @�d����xҲ4��g�Rx������;Z(P=8A�BC([����4�`z��>���ځ�H�}�d}����8\��s����d���6��+�{ 4'�#�W8G�a��kh	��4�š:�u����%�˼(�䅶�i�G����i���� ��=N�7���d`�O��o����P����ժ�z������B.��WG�qp�)'Y�E�e��j��d�;�g�e+�P��+����z�F# �mS�;�����:��}�x�bP4�s�Ӧ�S�܆�
�imD+�-:jd�,���ֹ,��E�H�	�\̋�'�ɸ��, �|_����4{�$��� Y���m�� �-�fK��r;1�,?o>ZԄ�Q"*�'B�����O�x*����-��g1!+��e੼��Fo�����8��g����sH��i�&b-�̀�1q�9�f��-�{&w�; _Y���29͟`ap�Paĸ��sp��"4  ~@i�-`�gm���K&��'�T̫���HY� �rA7A�R%	�Q�8�E�s�86-x2A���/���e��"�\�Hq����s��Z���R;�gS���s�s�gK*�ThO;Y�����Ҵ����=[�m�jI� a�9�����$�C�қ��:{=8�D-ϑ����W��Lɘ�/��\�n��'jပ�����iӰ!+W�\�� #�h�UO��bS ��� ���^ի��P\(5�7�z�S�)� k"R�8x�,c��J�9�>�����|N��ks>�.X��<+��U�.-��4�x�Рx���%1����G�����U�8����n��0�f��&�h��(�����4o{ͮ��;�pr6��\���{��rX�[ 	=��9ɛ;�ݻ5�a��!�1��)r� Y.{��U�Hh&��`k�(4�{�`o���7���3��&;f�4��&�����od�b�w���g&��Iݰ�5D��M��YZ�>�&�Ug@��)�3ڬ��X��z��+y���x��!������)�s�c�Axo��\1�bx=�>������C�Q�� ����L����@
/��D=P��0�tH��p�y��/��E�{k��� Idlu�'&����v<�jZ�y,7��ye�x�c)�%���2S[�9��&�M#�v��F������u�v�b�[츂CMſW����Iֶ?��Y��T8M��y�1ꨄ�⯲g��Ȃ�u�0c�Ő'��w�����;��G9ƅ���QM��̱b�8a����/mO �l��OʄD��)��2+�x�.����}Vĥ=���-�i=��Vu1_�l9_po������C�r��O-�� �0.�U�|}�\o ���tѠ�/����-�4�I�X�& k���}h7� �l�4��X��n}��gM�'ɛ�5�+�ثX��po�
�Y��ai��
��0��G�i[�}Wp�n�û�n�H7+Go��=�A�	�%`�}M�e�$4�����9���3��y��Ĺ
ꢢ�M�����`��\���,��\�(��Y��f�!�I@�
�U��'� ���>�8���A�����Ԃ%o�����(�X^����ك M~V��ozڞ�O�?!yL�lB�������Dz�I5��Cu�ܬ��F�̒`>�ڃWQ�Hp�P����D΀;��d���_���u�ȣ�y�޽�\ ���nF���xuVt-<bp���|.^�L*��X���s�n��kH�<�k���gr<+j�54P'm�8_d��J�D�<�50�q�l���挄on��y\�y.������=�.�aAr/��z`�����s���$
����=�S0�50<�fC�iJ�,̫yd�%O��1PMs��w���&Uo���ݧ���7) ޾�� 5���P5y��mw�p���n��`	�r�1t�O�*��ȃjd�Ib����^����PY	*�=	�oG^��L���3��)��3�,.��s˗��.q���y�ё@>�a@�:$�8�_' s��ֳ�Z��(�8;$]�5�lm����U�#
z 7�@[�. Ԍ����qId^� d}�}�|+���A�3u~��٬�X�pb����G���G�Ǜ-���[,虅#��+=�<t�Օ(+��]��"�*�>�cWE_�ES�H�`Y�oH����k���Q�M�*�-8/*��eu%}�|�CX�a�S2�V=V�~Vר�G�TL�f	���z���NY!�?{|=���doUY�j�)+a>���Bz �Z+���cJEq@���U]�GI���3��3�Dn��o�_�a��v�;��YhZf̖�%rM��\�"U�p�R�wӁ��7$_���WK��s�������̠kk}�8D#<RE=alI�d^���VI^` ���K����1�k�3����z�|�������Η�<l�k(�-DrO͞�="R�y�u���E�����%�G���X�I��A1@R�4x��ZS�RT��+߃��Dm	�"�t��������a��J��-���հ���5��fV%��9o����Rs�Xְ�[��,V�x׸:jP�� ��)�|�ªJG�p<|��PT�*���A�P�ճ�C���a�͠�VxZ��	����ރ�D�}�O�wR��sa��o%r�cxW�ǲ�]����p��J�dLƯg`���E0��	Y�m�l�a����RZ]ՀA�9��	`���y�[5���
��|���=m�^ͼ��p���'m)ȴ�u�[��TY���m1�\S�Fɼ�&?r�������c"����奏3</��L����(}������_�d>+%�I3���i'k-�@��➠�f��P�,��M�v,���$ߙ�^|�T����{�م$e��cP�:�4;\���_Y��ٳE��Zm64�=~MZޡ���բ_�y�yp/?��nk�����=q�٦�=B}�~�8v�:o�N�=�e�Ȟ*��h[�}��VDZV���>���w|qOģy�$!��]�d��P�uăq���<`3<<6�ɧ��������xd�zM�q��;o���}���-��<ؚ��<Ӥ.E���,k��mF� y)i� M�m.V�����"6iK�7-؜ߥ�\�+����"@N�XZ���{��ꇼq���ۍp��aO/���\�����t�{�>Y}N�b�8�� G9���S����R��_���^�^7���_g���AX�hv=����בs[.�������m-�d���>*��q԰+�,4Q�6j%�����]�j����xT�
�M9d2g���r��"A��L (���~@Cp��2�J�@!G&{�]���#��-�/Η�����W����]v�
ؒP�=�ђ� ��/VX .'훧^@��NH�"��ܺnV�]ܓB��P%k�Yސ�i�1������O
%9�i�GkT��7���7k�*�E�d=w{X����2�<���u��=� 
Ϭﴷ+r�4����a��#H���R�I~���A�VY��:��H �� �`�$<Fѳ�`�,��r3J�: -��x������Y7�4��V ;�P�w#���!U/}�����7O�&|�K��x�M���/)�1�ou?M�I>�Z�&��#wH��Tc=��|ޣ��k��F�8{��$�RC۳�|���� M���~^
p�-��p#;����)E����N��ܱNpM	��Ɵ~��3�0p��w/�����.F��nd���=X*��s��{DG�{Q�gs��uh;�h8�B,��X�]:�:Y�����r�Zh[���3@�vǎ��h����U�Y׳��g���Һ�E���:�k�,=��f�<{�B�`o�ts�ʵ�?�5W��Q�8�H1�[L �a�H��Y>�٤�f\[X$@��=�g3�����Q��yCNt�K��`�sxj�4CȈu[rd�ɚ�g����Q�:ca	T�L}c�����HX���Sx�"ɯ�Ǖ.�v�Wڔnլ��+�}:���{���Յ��^�pTz�|h�x�6�}Ъ2v���3�IHQ����1b�S3�@�>r,���Xd>�}j�\�qJ�����b��j ��xZے��g�<*�	�� v��+)���:y�I"��N�{���2�j5�##�߼_�����
��������;>?��ּ��hJ^����ͣ�Xă`����������C�ܜ+�w^��돜}�h�i<'�\�Z]w4p9,�b��g��DPA����/�GSk"����GK�-e���<���?�G�?�{`o�N<y�؛y�@i���	J�&FW���(<(��㨉��.��U�7	'��c�{ x�CXS ��3%3e�(aw{�AZ-m� �
q�z���oS볭U���N����[�԰7�y���b;wY��S��dՕ���}�j�	U���2WGW��EP�IM�����H�g��t�p����b���_^�ӳ�K�fa� ��9d�b���y`��m���l_�f(j�(��}d�?����L�]�*� �Ae��Wެ�s ���*�_����`9��+E�U^Sq��c��
�-`J�em�+5W�v�ŀ�=_e~}1�n��*�k������4$^�:�s��#�I�T_M�MVt1�y���ط�֊�qԼ�I0W=�󏖞Uq��Ȏ&����S��
$;T�E���U,��,\�뾟����}^�*��<K|��F��z/����˹;R�p��F����������7F8�4�LB;�}hv�N�1��s��3������g
7fb�,�W�i�� `\B)�R�-�N�֤�����dW�!R�V-�~䐳��9�a�����bI�SW�mQ]:eD`a��@du_�1Y}��2# �`nn>:�8�
��7�=�����cŏ��� �*�B��w�(�#���,`XG�#�8:%�[}������)X?<>��,Jk�F�ؐ�Һ8;e��i�#���tv@7o0&`(�
��U#�Z�8�2����8�eZ�k��j�>>T��A�Q�-K4���u�*V��B�Ma�#��B��죦���N�ە�km<�cS�z`���`�l�+~V0[��򓵃���w���8X�u��Ue]��6��Bh��r�XcT��U���>#�H8�kͷ����^��i"���X�ۿ�
���B�<�Z�s�(s1��XƱ[�`����٭n"��% -��hFw��D������M�0m-X��6��$:���v�9��aS��a��vf��f @�do���Z5`��*L�b����!j:sC��x�Qcm��E�i���n�J�g�6�W`�Bf�2Ѓ�v|x��Y.�|jc���9nk)Ǘl��|0r�S��Ie�֔�FS���9 V�FuY�ƺ$tƀ�U�+Dyo��ִ�ݖ5�QE����3i+�N�����U�ǲ��^�ĝZu��E`��`�A����2�Vu,����Q�9	i�
�1%fYgP��p`�ّ-�~�Gg�Y��crB�9�A������8�����P���e�ǚ	� �x��kO��V/`\�L'�Cɠ 5tKY>�%��M�tcN�F�d��>��w;���d'�$0�����56f��Li��+v)�m&���t��� �$���Y�J�jk�v�4n��{���;�*�~�gIq��`�L�V&�*}���i�ɬJ�|�˼�y��v��ic�M�
0#dw�@k(b6E�~�2LVE��U��Ì��
�V)^�E��Qn����e[��z|���?m0�4�X���&P�Ɉ��^5�S������ �l2	����w�)��Soq�%�_�-L_�����^���/�re%	�����ps���l'�͎]�X�A�CJWS�x@�N���L�h�C�狃�L�)�U�������ff**�e�4U��q��`�����o	O}g%zP�O�X� +&p��`t�o��`��`�HO)e��4e�,� :�ST?$! �~���c�j��T���1q�Y���%d�,�e�y�g��ٲ �瀔M��u���Z��U�7;@�ө
�U{��S6��HN��S#< Ƅ��:��^S�;�T;hN��M�s��Ȯ�riN��4v��<����:�	/����k5�S���B*��1�X<g;4ј4Z!�Ժ�[�z#��`Eni�������h�[\�,M�;P��Ƀv�|W�P���`׫��1�g���YYX��0�ƺX�P���,�7���Y��h}������W4Kݣ&� �?�j�H�jd�㟙8�g�Ɔ�?��wޑ`6����UuVΐ���Uk�Y�|B2ۜY�B�8U.�S}���ʿ���k�fo���i�6�����?�.��9�Ǐ�d,�Ģ��`O\�_����N@��l;6i?Kj���=$����4��MTE�s�\L;`�t��Im�t�V�WtٞT��2�R�k��:g� +���qz	�gU]2 u��
U��(���٪�
i�	�$�l�49�LY	�M���'�����B���y��H����|�Rӂ���֓�o�Ne�x�7S���ug�Ij�ov�5�t���VZ}%�;
��j~�VS�������	���򮁋#Y2�B3��"b �|��E&���y:c?�&����<�ae&�q���
ɯ3f,��c'��$i��ٗ�积?���́��S[���-D��pʧ�N���&�6���U�V��96��LҊ�OO˴�-���9�S{�	�qc�I�f�'r��i���s����©�ڜ҃����R��ά�+[d,ǘ�nj5��߫����<�z`d�����R�,�Z�1&d0p�X��\ݘ/�{y�9PZp#�Eח�*3�?n?1��r�4tJ�4�0�/w�no�y�X����*����Y�$�y���C�_3X	�6�����B��t�Sy%��k�2q!�3�/˩�*Fȏp�
=�*�m`�X]]kCy؋�M���/n�Q����ʪ�YE��Fi>@F�T���$��w�{e����#M9*����z��t��_�VK�����`K_�'�
�{���v`E�\Ōt��=�k)]S�)+��7j/��|��w!n���m�.��W�)u�Q[Zu����j�3�����(��T�E#^hB��z��2�	�'�)����^
���.��
�P�=����9��@���x�ty�Ƙj�6O�ɕ���r�C�oó=����/�W��c��A��4���8'�Jc�`"xT9V����_8�DW̫�R�O���*=��A���L��J�	7�͖�IP�A��ZʡU����蟛�|��/^���w�����\�a��5�� ����Ԏc��h�9�
�Z;V`L:���^<���l�,�*����XL��*���e�iu�������KR���a�`Je�Ha��̨�5�� �O�q��A�#aDJ�LX)��$@��� � �k�!�A����=�1��q�y�ayg#���������r2o�償����Z3
�'�8z��2q�����DW��_�{��O*�����~�������i:[�G�d�&�X?�]�Y%�	N��"�4�#���^Y{���xd�J	�-O?S��[YO[n��I#�I���G�cp��T�&Ԡִ`�Ҝ�)���H�!�-oę�J�����>`褴�A�
�?R~{'k?EE����gkr� ���hs?U��@'��s��I�o�hU��|�f�m?�:(w�.�ٙ��l�g)�jTi�-�bZ�(��싓�Aa|@���<9�Ve�-��8>t�����w�s����`O���ռ׻.��n��߯I�*>t�Z�Tu��|\��ƸcF0��DɛxѼ��Qe����8.�����<��j�4%L�4�����:��3�Z��gmm�}XW��jč��A��A� ��7۟�g��p]�����ދ�+{�����ؿ�u3�D5m�,�$/�꼳C��}�uN��c��v���_�l]�1����)���}��c1����w�7ܧO[���`��`k]L��V:ƕ�=��j�L�o�:Nc�u+����!�����#>���W�?d���=9����` G��Q��Ȁ��Iۯ`)A�k�L�b��JY�j�� ���Ϙb�ѡ���,R����E�x���3�VO���U���z�{g}�W��	�`�T~o]_�V:^�tdf�Z�k4We�k�v� '������b�e>m�� ��
���f��}�v3�� kU��M@d���bf�T+�At��5����P5���b�.&���I���ߣh9~��ݠ���"f�Cj�)��Az�d`<|�B�4H�S���^bi3H��J/TU�O,�񕉹A͏���WYd�h��I�|#/��gg�����\,��}�A����� l�����bӰ���y7�y.s		�4�6=7a�۴)ߠ�����4���� �Ȟ�G�bަ��:D��-N!mp��<Tm�o��6}��`�P��J�!�i�n�"�D��2V�p�δ� �zp�~~�����H��Y�
�Re8n��t�t��*)B❲]��'C`�	�힪���MlYu���)���耞[���;�d�&���q�I�p���[cJ�]A洦��p�=�Z�@�kq7pgr�'ptV���~i�xֵ`���̏1h�����n��r��@)���׍S��_?�GkX����@�e�/�����V݈�M��S� '��T�s�I�AX�V�F�[�OY+!��$�Cn ��c��to�ta��d5�'4`�t`[q/��� E��� Y�RL9�qB����O�[C��ro��5�"\/��Œ��T�����z�Ɩ��ҹ�Ř���{���4��e@��&R�;^��}��ξ���XY��S��L����d����\�s�a�;7d0��D�v*�1Cdo�Ҏ�e{VcW}�U�-�
�wP�h��8bcW�#G�rǙ�ڗ;�r_tʳ
�b����7ON���k����sE�P�#�ڮY�`{�wM�l���,@X� \	�����\^�SS|�G��'�`bET9-l�YSVR�pĎ�3�6���:g��*>E�@ �����[��!XT�'w�k����N����_~�M޽��lxz]�?kErC�2- ;�*�uz4u
^�49X�`:��8��2@��))m�J��V�R�=7��'~�L� 7e-��H�VOK&� ����w�ӈB��;�4��j2z\�#��d�%�J�0��M��0���ʊ�t�I��ܲ$G,���R��s�秠��e��p@WN�ϗ�ݮ���_h_c���S�QS�M�h!	n��l%��萶5ňpW2?$T7���VCA[����`!T舯	�`�jJ��R��2M�`s�@��Co%�s/�D�ۧ�P����wM��B��r���V?�4'�#�@��+h�<6�P�� ;8S�"�N�դlg��|ʠc$;c�b�i�.����L��H^��>gn�UYW�>U^/��y�78��J�h��4X��f�5I.�w`�� �)6
�mc��J���{�s1�dc��E�4[�p�07|����� �3�w���O��8���E
��h�!�Κ5;#�>x��P�[*����ΌW��eP����Q��1��PO�㢈R�����{c*�3b�Զ8�4ςُ`n��=/U�>�����UWl�8U���L�Ʋ����N�����������'�ڲ�-�K��$�V�2fū!�������'
��X�����,8`�d%ٻr�F*G����ъ� ���g{�ٲh�ۆ��We�5E&�kh��(���[6ܼ���0�_e�F�����/^��_�cW!�tpnڞ��ٻ�h� �L0�i��H(,��-q0G�z��f��[''���'|����A���	����"m1�m�\z�)�A��g���۹Φn�qpD�b �6�P�.a�����of-�p �	�����	Y���*ž������cO����N�<�����	腇�P�������Ld6�Ǆk9�#�b��}��.ZlMj0�s��B���)������N��sm�O��=<,e��	��]
t�Y� ��v�ʗH)͝�AT�U7:���e��U8Q\�YR-���Fg��.� �S.Y�8j�J��'��ƘS��7al!�^��mh�g�*�9�܂�b��Q��R���=��A#c���5`û�oe�� �7����MEzA�� ���t�9<H'Ճ���V�V��F�h[s���go�������lc���n�&ǭ�a:M��&�E+��V�!(�'k���;�Q�B��~]�}I7���5N�c��:��ZO�sb�혊���Uec�*K��;��_�+
�-r�|M{�mCMM��3�N��� ���W��I��gL��ȜS+�&,�ǭg��Juc�p?���+�۩������(�Lg-�z:�7{s�J*m�:�'0z0���YĮ�!��g?���z^�"��7��w�+ ��2����H��L0k6��Q�n7�<�� ��+g�� �?�3���􏎏�`���,��mLо�
�5?�.+�Ll��H�tWd���bܼ:7��G���1v�9|��
�ߞr>Ao���)�s�z�6M�����Vۍz���a��=�@��Sb�
|�l.D�m,x�`Z�$}�|@�y��,y�T!IȚX���,���J��v�P���߲Q��>��3k7
>�����f���jv�qI��t�Lӡm�M�]��~�1y���*��L�_*�rу����5c���2��ߘ$#��|vm�W�/�D�/�}�Y�Q�{1�j�T�YİŖC����A
�k�f�NE���-���U� �\~����}�B^\����� �Q�fT�a�2J�`q�5�� �.b�����)kװٵG� ��â�6��%�[�����{�e>�3��zb{�H`�be�.*�{�ioᡓ&!����L.�^q�nW;� �ë��rIK�|�����	vqU�K[�
 s�OS"Eo�`#d�]��A�/+IGpzJ>ۥ$���R��:���ͽ�=�eE������8U�لb���)د��2W��S�ʊ{~���#j��ag޾�x�.����@z��
���s���{�?z������4X%�Z�"��?>:���C���0tL� ���$��ۣ�9/�.A�"j�lǄ�`>pr�(����S(
�	S��荡i�d���<���)��!,F��+RF�Ҵ�rIЁk�������������:kڻ��?�өA� L-Y,.�ތX{$6�?�BN���0ā�ߔ�m�H(q]�|h}�u0�ujIK�Fۧ̀yզX��kj�q�^�M93kCM���w����v��F�+��7��ͼ+������D*��� ������z�JOؚ���sZ ��J�:NX�����M�9f^FA[3)��m�.x������y�X=�<иQ$���O�z�N�)x x|Gcb0�84>>����]#^��~�0<��p��ެ�߬�1������Z�K�:@��C�7{�Q�����zʺ�{<�D�����wb(=k+RA������L��Ѵ�m�t`m���Gi�g��w#��}��)èA�l��^D�H-ցb�� '��3x.!����d��@|�ݶZ�ҥ1�jq������!�V��ue/;K���Z�a�~�.��H�B0��d��2�8!���U�m�
#�l�䘣�I�*�g���������O��F :@a����Ȯ)��9���6��&��Cy}u!��y� ��خc9N{(�cϰ���ǼQn0o��>�=O�ߴ���ጒ�rj�*�G�-�˾�z��A[�� 2I�`RQ��m�E"l���=&��d.�g� e+�v(pң�c���$mgrq�Z�^�N�� @gB�B�fh�f#�y�`��x+�Io'^��iݽW�&������#V���Ƀ[���c
��?\������_~���}J@l��8GG�v�@�B8
��Y���6��&�0�is�sxƂ�	��=_" ��ȗ@����%@{�z^��n���c���㰗�)����"�gv L��<�/W�L$�/;�`�f��^K�/.�Ӝ��}:}����:�^�wK��zʀsv�6��Rԓ&����7ě�;��=�� �	[Ơ�b����z/L!pB ����/^�˫K9�q�Y����sp-�w��G����G����3�a].�	��.��9��AG��qj;K�WW����jŴ���d��"k�GJ+
�L� �(�)�s/0�*D@�<>9&������� e��:���J���+��K�>;;c�J����� �|�=��zo�] ��R��+�X��j�Q���zq]��_`���T5�4!8^^^�?|��;�����)��|�����Y?6"���E ����i�����C��_�[ƣ���/�fg�_�P1fWW/�����#�������k-������i��䍛E�T�� ��<�'�NhGA�sCO<�6�X�����@WVQJ6�������P������V���& �	��}��}ü�࢏� ;+�p����u���{�kj�=���_�幾������-���^�q�����\f`|z�O��2�0Q��zpС�`f����t�ڥ�Fe$�*7��]U���� �������4-��<�[X��b>5�{=DC��c�F��Ӛ��$��p�0w+c��� `�w�*��0xel���^ǉEgGy��)�?�)9�^qL��1`/r��Z,z�A�/U��c ��m+����dwWd���2��W@!�n�^2K��թ��?��|��+꽎�^�޼mC��d��:b�lX�k��J
���3�S��7�l�4���4j����[���X|}���(���~�3`��i>L��D��?��2'�ve�{�W�x������rx|�b&[4��q��7vOX�Y�0Fa��D�j�1�A{�y�`�߃�aU~�}&F&�{$�����*��d�8;?��A:I�M���Ҧy��V�6:�7i�Lt@Y� �C��t-X��εb�`�����g�#O~�M�"dݛ��N�^K,�^y�iJj�E]�wt����'��B�l�P��7a�e�ROt�r�^60���t���Z��aWx+�E��Fwx�N=iG���q�j[T� - �m|���)<M{"e�R�,>���� ���A
��W�NZ�4'�O�Z��FI󜛷;�5A6���y��57���7���OJ c�#�n5����<���7o��i:i�
�TcM�;��7�`���O�����m`�m]NR�Lc�t��k�J@��������Mf�r�X/����Yqc��&�����~���b�z��z����W��9Y �S���L zl�W���/�y��_�|����O���� sj�V��׎�R����W�^��<& �Ё�<O����Qno��{��e2��r`�̣��L�a@�������{�O@�M.Q� 0$�ҵ\�=ҟϽ�ׯ_���o7�[��0 ����/���|j�(ʘ�%����_m� �Kٽ��o���Y��o�\�}@�B�����{����4�17�Vv&q��28@ŭ��-����s��o���<����5�h̎��� �s�.��=�7o�� ��cڣ�	��ݾFzt`��2��	�`�� �6�YO`�*�&����i��+^rQ��\��P4��xQ�oƾ/�p{PGto�s��T�d@���}$�<G۶�?��g�����ſ}��es��O����)��%�p��8ú� �	�Ct�}���q���k)M��<���W����o�����zq�*GvH1�K�a�cܙqqחJ�/}��2\�m�-��Q�+����XA�5��>3m�?�='��ݟ�㓬Og�zL�5*9�I�0�4�_t�aiN.�=����٤	Y-3���s9K����*����Z���%�[�9j)�jnSՅ��1�����ƥ9��7�[��1*0��:������#h�ˋ���כ7��۴���ן������o�_�mڌ���Xu�7��P��7���&pֵ9�g��s����ט)���W�����i���r_��P VgGw�ht���ֈB]�3�c�Y��q����$��Z�|��Kw;�ôy'�ˤR�/z�������o��:b�����;�W4��OR08�ڋc��1/7	�znڪ�@�um�W�4�S]s��,�'x��/^�bp��s8I��� 7ן,�C�xL�"��y
N`- J^&`��7oe�����;�.��x�&�f����`�"�o��.ܗ�#���ݲ��|���������	�`�$����0�~����Z�����AA�2]�Q�Ԏ�T[6gG�Q��)�?U�{X{ >?gP|��EZ�������� �ӯ��Jv�ifPj
L�����?������L��|��.  �g�'L1��j��P_$���U#a��x/�� |�p�½y��}���<���0�>m��}�����odan?�H��3� b�i�O�����JK� c�G� �M���� �XB�xx8'�d���}�K�.7���g>g�#vrr���U�w^�VJj��<�/�W�|�ǇG�7�AM~��:O���7z��-gi#�����)�W[+�Ҕ�ꕴ�)�Zz �s�?�(߇.�igc���N�Á���"]�k��b�9��k�o�7�f��"�����~Hs�*�����k �� k����G�[�`��8V`�����q���8?0�&��z]�;�����ZS���������ځx10G�&��2�4��\L�p�j��G0���J�TA%X���m���*m�������a����Ƈt��Y�[Sx���f�]FdR��,rɫdL�Y����d)#���C�� d,���ʶⓠ�j�
�t�_�ǝԁqv�&���@q-��F�}�B������߾R��Z��U�P�^�4*�;�Û���l��}!$�XY��\A+/�&��Q
(��,��h�S��<��{�c]Z���&�?`�q��2}�0��\����OuM�i6]�5���1;"[t��e
��t"�Iz��ҭ�,4-uR�fEE�~�z̪�0X�֨C�BC��ԣ65VC>�v2��W�( �j+����^J@�X��{�F���D�h�������ߥlB�ݒ�����<���ۖ����& �5[!1�"�$+"y$F�<�5����_��F��tP��Gz4��Y
d��B�1sW��!��>c����y6	[�Y�����z��	� �.Df���	��>����~b-&+R	Ե���e����
L_���k�X58z0+��pĚ�<�L%N�Q���B*r����q@��iڐ[�9v��UZ')p�p��N�9���i��yX=f�X XGǪ=(� ;�M�/�ϱ)�j�]
R �/_�`P���7����=���x��u3��%���\��	�;��ظ�Bc�tnը����҆#��Buc hT��@,��|}.)O��d�5���sMb����Zˉ
�3N�VP�3ά��	���3ڇ�OО>�4>��?�;�t��8��C
[�"v�MUq�p]�i���C�+��S��7LZ�����ԣ`�qϑzľ�q�ZԽ���&]��q��p�R0��|��G�\�i\P�5=,-K�O�t}a�:�}�zѢ̧��c����}֔1M�5�ۂLԁ1�gi�Dݦ�M��杤9��Em.R�[�7����6V�P�� py�VN�!������l�/�R��!1�cu�q�����J�V�*���z6���Z�[��X�#̛�df���e��"�<.L߅�c�7nl�oTw9֓���ؿ���$�1��A��&��L;s�fӐXOW�9,� <X�����$�í�U�a�ZX����J9�6�(�%�6���8eq�����,�K�R�S8^9M���d
�	�Z�z��`��5�������k价/�~�N~�����:����k���^>�Mg����i>��6��U5�z��b��
�OT�Ģ��}m8��H��1�>v���zM�y��� |P�*�#&�AZ�4��g���Q(���a/��ū�L`�ƭ����q����`c�� $���%nԠ7��,��1�<~8�G�	V��-f���_���%(�u� ���dUD���ZO�dP�<<:�F��-?�"w^���L~��\���u:-�����_�ۇ'R��CM�A<�KK�zQI[[*2�F�C5n�S4o~�J�~>�H�E��ZE}1;�r��xZ�}ȴ�A'S�����g�\!���Ҝ�4&1;��B룋��Nf�&�"�;bEJ��i�@X��*_L{���UՄ�d�ԡ[7!|,�d�80:��/A�m�+�2�zH���X	�4	��cxZ�)��	������JA>7��sq��Ҙ�A�4���xе_5h28������xr0��� �j�oJ� [۬��(7e5���}���������V�	A��Ǝ~�x/�@�
��r���x�,�OM$ 
��C����P�v1���APj*^/[}�h׍j<0S��`7Ўپ_'���ْ�A�h�=|���[6�n��p%��Y�M[���i���[��5�A�:o�k��hpa/9�;0��k���J�:ը&��RػP	�T�c���
Yp�����V�z��Uf�57|@"��:=�sF�}���HO��=�"�H�6~��B���7��i�� �g�оj跼���7X��v�
" 4�ru�
Kh�{�0��Pd�*�\լ
��a���g�����ឩ�)|����"s��Yz�%+�6*¾��,�59�l����0 c��s�utxzµ^#%���]�T�T�����_����C�>���l�k����59��zf�HW�34Wn��P_���R�S�>*���f��d�c���:a�����iQ
tvƪ��%��Lnǵ�bq����b��f�B����!�V�U��P�\���Y1���ɂ{����9�0�ʿ���Ʒ���Ǘt@��Cz1A�4_����(�}q1@�`O�v<:��wo.���_�"���72O��v��*��/<�k�I��׼H�����qc�\z⍊�Ӟ�{tlv�xv nU�_Y��P3:��Wɹa�Y0�FǢOsF���^����ƽ����xA��A3pnLA��*h�{�^\I;Sc��W�(�=���$�N C����`bU�M>Q&�1;� ��hg˛JN��M�,�f�Y�W6�h�t���p�&�7��M0�B����*�5�c�X9M�j<hV)�`"�ǟ���t��D�i�ki���EATcjm��+�R���{ �٤1+��c6{�1{j��8ٽw*q�m��u���#��9'�s���%-�_�>�F��H�����	mc�[Q[��~���z�EJL��p��K�P-�F�*/6�B��L�9�v�x���T����z������ˤMq�U�z�5V-�� 6!�2�X�0�'�h����Qec��9���oh�iD����U�)5�
�1�3h�4%�Z��T+���m�:�����^p��L��V<�yC�U��"o��`�x�fBX��P����B�n-n�� 4{�T����s[��(X0MƉ�v�
Ź��֦![VhqF��g����B50#x��[�@+����5#zB�J��G6��~����a����:�8�9�� ��0�ߍ���<��١�d�5��v.9�榾�ܓ�1F�Q�`ͮ�Lհ��ҾM�?�+���U�u^d��l�9��
NgG`�T�����S����+�����A��ӑk��Lek���̺��ZqA.��g������> ��@`\�u`��	�Ӣ�:6s�=e%����ʬ�3��=ġ�0��8��}z\j�U�֣�ܠ�mX3��w��b,����<�t�Sw�d��V$SY������oPĶ�i�tvwQ��Y�X��`�9Y�;
�!��7��_Ҁcg�ܲ"��g{�����>�;���������h ��k�!cL����i���#��k��-=9c��7/�������o���3�ϣ�GVk�0���A����S2eZo��y��C�:�~�\��H�my�̬!��]�qN��"��/�f��)g��#�CҾzx�b�1�����枋�j�Z��������z�i

���:���gjF���F�M*g\�!g��¬F���Y�Xr�]F�� ��w�6��%�A���6�/���+!gsz��Y>�9��(�/ ��j��������ك�~>�M�
����V�I)� ���.� �������Ƣ�����
`�"Ȭɒ��2r�^)��*m�G�^��C���W�O���ú�I�3w|���ߴ�$�\�]�S��ۛ�&rv�6�IM�2X�t�+v�S[z�G�0�)�E�q�',ۮ���dJ�s�����j ���rq;.r^2�d�w�+���Ȃ~k��iALۅ�&�'��Fյ�5��[k��@����f+��<n�V.��u�����2q�?E�\@w͌����PƃO�8pt�}=�I���@NOΨU���
J�Y衙��_]�+�.�R��)3	]۸h�������6p��Ȓ�i���c�mm�5�7\���Ֆ���~�Sa%������)�q7����c�����
8��S'7��ܽ2�5�z���s� �R"u���U�<���o�N}�ԄVT�������i�*�}Z;kz��4e�Nu4�~��*�5Os^&�x�5�Ui��2�T���I�~P���d�U�0��*��{��F
4=��[��Q�_���p��KB���D�6��M]�.[= ̨]�f`��Jh'%���z����~�{��Z�c���B����-S�d:{��{X��8V}��i�[�i�R������������K���v��ux ¼�Զ��ݓ���2V����-%��L�X�EV
���N��|�jԂ�ݐ�Uܜ��r��"�1c�!��ꍁ��6����N���00��^�'ڄ��O�_��?�?�􍜝.�F�iCP�5LTC�^?�4��'��2K`f����z�*�d��3��v��0n�5�[�
]S���Z��A祈�x+�tK����l�U��.��A���3'K� �-��!]����j޼���\�kuF��T�*U�@1�z�DJ�����]�,γv���?��6�{¹�CǓ	J�#�h�sV�Q.U��'��Ȉ��I ��p_k%E���\�bq�|q���x}Å�翿g��l�6�r	��j;��dU�6��x2T�(���<�?��M{��%��`�Wvi7�ܾk��y#Q���r�&�_^�����N@�ϧ�z{� 秇rt�N�����4�:�@�E�����l�U;�کtJh�i7��v��� �[;�JR�
P�}���of���B�٨hDʃ��,&6O,�6�a��*�����`�.IP�}@\����5=�6�6u�g��{ݼ�N�ގ�"y���T�T���u���7榬���EZ2}�9���Z�h��ߴ������T��Q{B�}2{�,f�*��� j,`[k
:'߃��S@� ��|+��B��n`��[ec�����-ҍ��kO�麃v=P�����O�����U�;H�	��� C�Wvۋ 0 }���%utM�E�4ӥ���gn�<h�]�Lq�ŭ�Ϭg�eV=�2��������O[�Y��{� cA�����J;�hJM�w�S��.��e,�}]:N�m�~`�j�Jx��UT]�9*)O�9�;��A��c�H��Z���W[gu��	eʢ5��W����Ւ�[�'k��7[��}H��S�m%d�$Z�<u��A`S+���ښh�}�B��7 d]3#s �1Ø/����AN3�g��=��ay�Ki`c;NC�|��[3A�aJ�S��H�4]�³|�{��^��ڵpA����w��nz2亟��Yz2��hȖ�(���VΏ�^�?����}s����.���N	jm������B��L5���� �B�
���:�7�t�yJ��S	T�G�2�\t:�q>Ln<G�2���K��,�N�cl��O
`j����,Vp-�r��^�`(f7q�8���'}z7Uec�I��L3)�RA2Sԙp���rȹv�CMA���AfBߕc�zq�����'�F?Tf���6�^�>����X���Oa"!���������k
�3��}���M�L�ؒ	� ,��:�C���MjV����<���8����V8^��
�q��2<��"�rz��W>�q���ǸR*�����TU� �G�'mP�u�Eܳ^�V;�Z�#l���7 o�SL?�1A#l����\�j��X	8�8�Z�v[6���yv�V�.͍{���\��R��S�L����F�W�k���\����L���at^U�X{ �^����ڧ�-�~���1=6�%O� &h���U��D�^7,nl�`a6�*A�wpcS$�\��U�*;WOf�za`{�t�2m�[ܴZ����V>& ���J�.��H/K�ai.���d������t�\��z:���?@č*�N�Np~zƍ����7'�'r�B�o�c��J7�8ݿ����OuU�Ԛ���䂥k���� ��t0׮G�-��8`���mڊf�Bn6���A��䉦c7w��f��O�D�Z�`���,��N��?����LK��|��'v���Q��p+�ɨL�1bL�N̼�׶?�ժ�	��δ6�����b��-7f|-�+�2C�f'����k���l��`筛�0u�Z���= ^$صjG�I��q�;M�[Am�j�����9���+yq~���^���'8؋�g�Z��{o�t�8XLճk:!#��s����A�S�U_ W��v38d� �j��R�a\;�������!�pxQ���2(���h�zeљ�4�qh�����]i7ƃ/8�����$ծ1�H�PhpK�H�?�	���H;�XP�}xf%[d��{c�=�5Zq��x������ l�����K��;z�L;b?f��"l��44�/������O?���)��g���Ɗ�	��e���`�Z���ɹLQ8�8r�h�ˉ1ͶjJ��ӳ��Y��ja�!+�M\�n_!W���֮̋h��~�NL�R�e��������
g	4VJ�� X���1�S�I�t���@4����R8hz[Ć��A����s2 �~���Rqѳف����Ʌ����M^,�L�7(�|��A�Ϻ����u#����T� @꿐��o�j���7�(�������fZE�n����;ǂ�=�٪��x>Y��*����4�����5��� ��R { ��)ji�7Oa( *>(�n��;� ;	�\ �i�e)���R68ٕ���z�桚��pcS'|(3�z���C,��[���bϣG�t�YnR�W e%�أgOnl��כ�&�O����cu�^�����&i3P�t�0��` ��S(��C�h`oG�~J�0-,P��,Jm���9��*������(�5����N�X�C6R�����x����I�E������! J�w2Шv1?�GZ[h8�55`�Z;���LBN{j�B[FH���TY�`��^#4:�<Y��M��Z6I��8X��e.�G�f[�^��X�v�@�&��U�ߋ7�VϬ�������@k�t�����փV�Vs~�9�,��U�����ڶ�spt��M��*Cf,���DUd�>F%�:�?UX�w`�P�b�F+l���Brk4�g�fV��5��2ͩa�ȮV��w2�}���'��b�i���v�ς=l���N���C���=��h�Z�v%�)��hy�E3&(�9L�}�����'_4�ŀ��`sM�ZM��dIįY�f>.d�&����?�*��b��VFX�GZ)�x����vY4u���;'���}����4K��<���p���C�qg�2f���/c�_��L�$��CN%<�M�Y����4� ax��2ypФ��r|0��˿��R~��m�gi�l�ߨ�\�~D "����*����X�`���6�Ͳ�7f��|���{�e�� f�7
��W���<�>�Lˊ�,<pt!-�EK鐗�(�%�_�&f���W�"�F�o'!�*hY����N�!}�iy�;�zI�T;ʎ���d�<jz����uNN.���XE��l��V�Z��,n)>-�х�b7b .K�!����8���}vv,o^]�m`7�V5�!AW4 V�Ņ�P��[�0qc`��nb<�Q���i�h���I�2Jl�8�����|eA�3C(�"b�<�������3s���~�"�9tz�7�)=��sH��FC�
,�eAo@tR�[U��պV�}�6��F>���t
��zmփ�'�w��.��hil�������f���ҽB��Ǐ�F�'��rڳTn�N�c�ڕ6!>�����I?4�'V�l6"�8M�~ �/�)����^�+Z�r����;zѫ1��IOV�ZӁ�|�9��x�`HP�^m��j�Ra���o �N���6L�WZ�=��]h؊��Z eR:VE���5�5R�n��4�\E���Ji�u��k�ֆf�Z��4����7���X*\ ��C���s����Fnn>������n�[�4TM��қ>�X��tY�挧�\���%�)�}zД�D3�����tiڈU��*���G�� X"�R�:n`7//.��<Η�H�h��Γ`� �R�-�>Ѝܗ�h�ksZ?��n�.7�� L�h�*s8�E
[��Gv����;�𔦺Yb���#����V�	��֏r�;��m�QA{rt�1�5���7C>CG�TkM��  �Nh�<O��Lp�L�b)r;488��p\�D�Z��L4Q�W�>Nv8�+��y
�t�qEۻ�'h�pH����aǲ���T��%\��/���ƅ\>��*;�K��<�R�{��*�GZ��L��Ew�A����q��ɮ؂b���Zϩ��:���?�wo/�h��w)
���'�=C����uՓ��,���吻pT!�����"+����lL8O`�3ӨF�E���trt�,4�(�Y0��AQ3c�l�55�f4[����N�G^�E��5<5(`m4_ZK>�R-Ft!�I�u*UL;�m���&��-D��K�\IX[�heFmXH�ő,��)b�W~���|e�'�4uʩې��h"�\��@�Z���ĺ��T޼~���r�N6	L�T�υ*��ͩ���P���0X���� (�5"N\AݲOS�k��a��g�̵㯲��b��F+vM#1O���¬@W�]dg��������)�U�����順X���I���Hţa4�'0�c������'��� %��B�=����g�A�ǓQEc��+J����������͊��s.:?��"��"r�< ��{"�����Q��6�v
`�*Tl�DUS�՜�:	�����˨�Pتs��8z�0�I+ڽ�Ze��!(�l(rW/�����.5VQ�Z_�% �Z��U�NR��o�,L�Y�
�z3��i�mq��ȇ�`�M�>�&j��N�i�F5�,<0`�y���t�2���R�OKP|,
魤�1���u�ן�~l��.�~��u������K�3������̘64�рLPn]Bnl���40G��i��w.�*S�5��6�9J���A��90a�Y��qzrªO�VR���d}�_�T�f��ܮ�5�\�0�A�J���=@�lhT��ϕ�1�U�A��L7j'�4XJ��=����m��k�gh ^��|+��
�S:^�U�UF*[���0��6�]������Lk������?|�K������JC�y5ڜ��r�*g�������d���!!W~�7����a���+��+K�P ����w���"�X�eed�{}���=+��N���MV߼L{y����Q2��v8���M@r�Ɂ4`�V�C��B��2-�����ڸp/��;��ב+E�K7^�^K)��8����
��MiC�R[V�cS��}��c0r�{�T��1q��*&Gr_(^�t.`�v�(׎�t��Hag��篡�I0T���m3�׌]`�jr�����I���:8�lBBC�x/��n�ٕ��*7�����������kh�R�UL���S��'L3�܋*>{H���5J�g�e�ʇ�ˆa�k,��#��l��WޣЩA\���15O}�ދD�N�����������E'?�˟���矾%����N#����iv�����`�$��.�I톍���]5c/�U:�����h�t$��*��S�3�=�阪���M=@6띓p2���`�j�5�D�+<�Ea5�� `!5�@x�q�W꜍�>=����4E�aol!��&�f�ZiY=5�@�~n *ʳ�
��Ό�X9���.S�u�2��4;�Ӡ��5�Z�A[-Ώr�x�J��n���e64nr�n�H�=-V|��z�U��y���u�G���vw�~J7���m]Z+6�ه:��]��l�ҳ)�����앶�I���r=C�D�ۘ�8��H9lv[j��~�}�A{U��`)������6ml��Sg-�tgL�bL��`~h������{�'3���8��|���F�n3U;k	�6�/��>[�`[��Y�`MNs! j�Ĕl-X�`�L-;�-�ĺj���`[����1��1���V�� �žS�uh�9��{oP��>��(V!iՆ�D.�0.���՝�:�=4����<}���}�?{�1���]P1Pv/��C��zY�9Zͬ��`qL5B�6NGF2c��	$�v+vWy��6�7g�Ff��B�������;������Pz���7��=s���Z�Q4,��݀�<
�4�Z�!�V�e��a�� J�mF��~�	�@�y|���o�RL���9��5%�ణ6�~��4�OV�вg��tgu>XD�!_س�ѕ��$z�>3���>	�waH��H�3����`H�$X+����C�B:=H����_��G��P>�ޤ��A����>B�L�y�PX�yrE��T�-kn�$�}^?`}���/9����V�W֣�b��,\�>X_��BU�"^_��$x���!0P�Ӗ基)�+�����/��<<��׍3`�b��l�>R��>�ڿ*]K�|����/R#����;Fo���^U���6���lVˋ�s
a'R�ńJ�(w�]�Ԧd��f��"Պ��T0]��
ZP��V�d�E�(��8G��%��Tj+��!��=[���ԟjJ;���i�` "�
����T��	�ߙ>�zu�ΠV�C�8�ɨ��*�LC�&*���]3Xg�P�@���̘����0�G�����,�4��,�f��5X3���WM$ �� �'�	��P��E�̡IH�[�.��+ع��D-Z��۫(��X����`�<5;i\0�k���@ �
�&�}k-�p*��~�U=iz���C� Mv
L�ڸ��Lg�5Z�Ё-��a�+���jZd@;�-�����LM�9��}�p=w�A<� �ދQ�oM�����2~԰�b�!b~ij抴��i���אL~��$8z�t�kJ��*��c�2Z�H��ͼY�y�EUe~]�[cq���SL��Ӂ�0�s/������D�� J�Ҿ���-��̵~ș>%�1���T��&�z�#�����,��x8�z<UL�_~������)]K�~ʰ���tu���0�8�<ގ��(���0d����9�<��������mR�i�cl�0@�,8�L�~;����,�XL�彑��4�i�  {yu!W��l1��d]iq��m�b(ѰB�� S�f�k�|C^��H�Q<�>R{����o�	���VV�Њ��\c�6R�&!Ke{τ�Mk6j��󪼊M2��y�:}��f�`��r4��c��wmHg<E� �������t�� ̦�8e����.� `�BDp�Sso�g��&��l*:�в�@R'E�Y���4B�Z�̞)R�WV[@8�`�999LT� C��ѻ5�6 �r��(&\*`I!���yx��"���	���r���:޺��O
~��X�J����>_���[X3`�R�ʫbm�K?4}��=ɦd�>|����o^��鑜c,�[lP�T%0;�~��#
�Qe��J`!�00��TY�Z����s��uC����F]����ʵ
�m�k5��[�U�+����"��郱�Q��bz]�-U}`�`Dyz~!��	��Չ��I�Ӣ�6��Z3t�Sm��f�h��"gBڠ��ڸ5�4��zɈH������[�J>�@'@�6`��>M��5%��\�9 @%�26�	,>bNfXE�^��0����4@Ņ�*�c��:L�nԠ3�k������Aգ�N̰2�i�tܭE˵�Bkt���8��"5���ސ)z@!e�" �F��x_��Df�׽AS)���=B<�+tQ (�P
|�0E3����!k&)^˖ ZK-�nba��Χ����m
�����H�[j�q)RØ;j�������t�^8w�*ǍYh�Բ�Xd���櫶VP(��h�V�t�[0�dCk@`o�e�.E��'v�o�wX`3�s�3�B�P�⒙q���H՟_^hUe;1+����iKd���S56�,p�����,-Az~n6.�Ne>Ӿ�ZQ۳�?���a�kk�-�
��*��#%U�+=���*�i���Z޽�,��=���گ.֜4鴸�����@:�\�A>�G��ʱ�ƪ�xa��\��� =b�9
����L��`��uq�Ê��&�H雭T��v�ek�9���\��� ��Z�)����ř�fJ͗t�CQ)�Y��C��1UT�W�
_{�0bP�rv!=��֜�b�bg&����ll^�ء<,���	�x��oUW{ȱ\F, ���[,/?z���i����K�q�Z)&ah�F�E*�����y�to�*�V�=���
����Wa�T>G���_Od+�g��RɰZ��.h�(i���L�%���Y���FF��?�ʚ�0F~z�$��+O%�ęy��>s����n��k䴱))м�G��{3K�8�⭗B����k7zӽ�6���Nxg�Vh��\u1��u͆�+ljd@A?�sj��W�HS�媓���,7p��J� 8�*�*�K--�S|:��Q�`Ƞ��)��f�ғ1
+�瘬Vs�SfDc����9�S�bVcBl�r�� ]����7���-�)��Fw]��;c��i��U�"`��cK愄8���?��`�Y���_�� 0V�M:�߱*U�2
��尙"��?���v�f��@�F, }��2լ��`=Ze��k�|{��zУ���%���Ӓz�N�nj��M<���&����Z�����%�e �Y��F������D�6 ��e�8j����)E���z�T/5�d�W��� �Nl<�n (D k�x�T6���Ě5�QSX`�zK&s��{�^��	C����G��C>�ܤy���� A�l̳�z
��g-@��<��hT�Sx�`ݟiab��v<����R��CE1�]���=R���=w��IV$��Z=�xA[Z����oP@���	BO�GZzt5cS�&qF�kM��w�ֻA���_p6�:"=���?(���Ԏ�n	��^yŧڠk�j�E��[`��d����yo��7x���9(p��K��݇������f_a��H��.V(���W&֎�]�l�X<��;C��8�-2m�M�=d���Zai���imB�ѨƳi�\`���ZA9�q�}�E{�V�V)��M�YE�]5<�*�HvB��f��);�j� ���G3�I,��>�Ĳ�f��VF��=Ğ�����b�a��Ӟ�v�-�Q��z��(͡�������,�m����f����5��(&G)��z��i&�É��"��Ӂʞ���i���v��IF��}c����đ�f��@#p��/G�`�)b7d�tv�V�M@�l�>��U{����vy�2�#�=^�ElBa񙇒3}1��Y٬�bu��/��� ��Zhg�f:>�����lW�P���OP��	���J߭�8�������ޓ����k
��D=�O�Au���qC�!I'�X=�"�<�=[oC
RO�~F_�u�ձ`F�	�9�������cz9��������I��|F�u��$�����^ִBz��Z�L�{��Vm1����7�|��ᑰ���U�� t?/^]�7߾�W�_0�����!�ϟ��<I�
��V�_�f�����O���(X��{�vH�q	�u�@��˗r~yI���~c����[�閕i��ܟ�o�DIw��H;�h����_~���!��%}� �qO,؇�G��]�H`)��!劃�C
���{����θn܂� ��>%��c@��`�36_�g�OϋrM � �|z�����Z� ��"%Y��3�����k �;��A	׉�\0M�� 7ޠ�@ ��&���}��9ݻ�,�S�&���v��	�}�7����l.4L�^YA�����@;�c��	����K+ V�왁���v��!�V�
�{�Adc��HT2�`Oq��g���R�ߟ���S�����M�In���5��Nρ��S��+ ���,6�:ߋe5�أQ��Ƥ�.�����Zh�ޮx/qmG<(D�z�^�t}�4�~w�7�66�� D�b}[�!�Z���,�	�T�����j�����N*l�� �{����.��ؕ0B��DK�*�W�Ѯ���S^��_�����g�_�t��M�r\�N�1�>ڹ0k�::8�LEΪpks��vч��<<ū�^�����,a���ӽ���UJ���R����0��a����v��P���;k97�mAsm�TLO�+/�"y�b�G��!��5�G��ENA�v��X����Z��`��<Am��^Ր���X�UИ2�4��N2��_�P�v�
9T@X������u�=4�_�2�j�-0 H�S ���C�G��*`V\�Q��4/����g����D7Y�-+M'���J��Y�����`:y����"���hw|3�<��?�O=������k�j�B[;=9|�Z={8]�x �1W�xMOG`�f5ߜa����]�S&�:[4%���F~;�(���� ��Wq6�OsF*Zg�M�`�ZmW\������q���^7��]�a�6�K+�#tTm�B�y��UOo��=g������t2P�- ��̴:H�D��f��E�fzb��i�/�Ŵ��`��@���y����Lg���zVm�:��L��S6Ϡ+�P�j��S$�1��Rp=<9M�u�6~m���`si40` -����*:��-з,>OI�4����y�XlC�����_%#5�-�J��b@��'��w�2n�g3q-ӑ�^i�7\���A`�&iS�
Rm�iϚMmm팀�)M���!�a(���FjV2i��>j�s��A��@��9�;0����5"b��ʂ�M��6g�%I��&�HW��UiNi���y4���8�����Vx��������w��V���"�B5��j-w�h�:k�^A@�V�i���t���	j��F��P�{�5+Z�,װ��4�eԴ��|Ě`!D�>�\���)f%�	�r�2A6pvo�ӝ�M#	p�@� �6dL����{�K��LT��ׁ}�6Z��s�s��2@�c�3Gj?L#�h#��M����7����������5��o��3�Z��_܏�bb/掶z�ς[~���^Ir�G����_0�5�/��um="�5%{Zi���^�H��͈��γ�WEI�
��gk;�k5�j�2����q�.�D���c�#���;t�^���(�:����o�&��{z��in��L$�[���*	hm66?��IF���k���X��_�E�Rv�����hD�h���)�o���:=Ye�R�ka�-r+	��R:��Y΄ʗrs]@a�s��W�1�v��5>#t-(�lk-g߻\I5�/�Q� í7�.�G��кdЛ'S&����h�9����0����?~eV��W��c�tK'�xY�Y�,Tf�A�5���L�����mB�K'���}���?�3���w�#�dGv�b5��1<u`l�`�"��AW���i�dBq��[���]�V1~}�`��+u��B�{��?ȟ��'�`�H�䓣c��O?���%O�>|H'�[���.��l�J<8��39?�bp�����|�S6ټ��1�HG��ӥ�:a�+�?��n���߃u;Ls
�./��"=P4 /5:�[cpT��B�0.8���|�F.�.��n�u�gHu���:���݇��wKA�S���Nz��|�����?���)��k�6�X<��}�S�.�Xa��7V���P�����7���� "�F�X?77w�ujۿ��6�����@uy�RNN��P�*��!yH�
��w�?��Ӛ�k�A%
#../�g�>]�	+��<~�� 
���{2u󧍜�\y��΋�|�����狅�y�RP�u}�)��Z�W�8��v�TC�5�=��ѩ��]�{�f0��H��`;�X��~���Gi���i@N�K����鷚���a���n����;��_i�6
uM��bƼ� 
��U�#�S'ggt���|�Lq'�5uydi{�*��s����,��57=]�{�4����+�t{"?���\\�ӳ��AׇT�qZ�`ݼhcޚ���W��>�׼M�m�,RWi�?̀��K�1ӂͼ�� J����g�����t�߾y��d1;��Z]� ;��)X�~x& �(XL��<ы����>}~�$Y0d��)����@� ɜ���7��Q��x;���^�}��7�m�m��2,�6
�M<'�U�&�жZSv��kŰb�	���QJ���)i"L*T����`�cuio%V�0��`��a�&��;li�B�n�*|5��L��F<�x�sS����jz���t*q�P���"���|��y��/���
҅�#o����W���7���	��^a�B�d�A��:aǕ�e��_0^R�%��\F;pb�;7],�'k��w�6���F�� ���J�Q)@*��ot46�_���:)��0!��F�\��P熡��J:M����F��6��5�Ĉ�i0����86?k��&�xŚH{����������D��6G{����@Kg��Ni1n��yX���.mp���l��fS�oSi�G'3Ք _��i,��h���\�l$j+���8�I�vƴ7 N�*e�.�����\a�	��y#0N�_��#�ҔM�&U`.��Ѫ�Y��2���5�6l�3g����������s2:U���0S=�Ī ~���y
�	 �{�� L��j�4��������7
����`��bq$'�=���Nb�xڜ+�'�b���n��8ī��
a�/..��7���Ɂ���^�g#�_(��H�&:��fѱH`�-�N�D��)����?��t�9��ag����o�����4�GǇL�~{���ۻ�L6�*����U��3���bڐucR���]иޚ�׌^#��s>�0��Q�8�a��9g � �����i�w�il��mЇ�7�&�,�F��)<��`A��ԼW���;h�T�I���߬>e�h=��L��@An���HX� ���c���\�>J�W1<�>S�;YQ
�4/`H ���w�"�0�:K� x���{p`F���t��RƎ����,�2&�j�
txpצ��]�3���� �g��'��\�R���Ր�M���z+1�t ��~F��4x��>���a$�c�W���u�/�0�����k�a|ԃ���(�A@��qNZ���S��!��*P�fͽī�9��!_�(�i����K���7.�M�\�=���PE�T�e��c$�1`Q��,�}>EJ8-������_��x��������o�uR�ZA��޲` Y
r�g -�^'�5��|Q#0] �FU^[�4�Gv�Í�;>�o�;��j����*�7���#��o�=~��By�}��weq���"���Zu����va��IM���6�犚��Q����,9�q`&Y_%y�2�㕡#t���;�cV��}�tQ�
��+��Z�ͥۼN�^��<-�v�����z�R�S�'$�Цf������ BL��E!z�H7�9�@�}�������߲g��}&x���c����>|�_~� �?ko�$ɑd��{�y_u���������+��P(��i]�:�"3.w���T�ܳ��ΐLttVeEz�a��T���w���-�ia�˲=�:�U���x���v+�ڧ��@��%!XV��UBC���k�R8�&�¹jc��%D8 -v���Y=cf zO p� �����T��^^�L):�p;;;��@� Q3�����Qr��C�%J���ұ[�E�+r�v���Ό��*�5��J"l�Q_�<�����qg�/��:9��d�?���&���f��- @��0d�Eǭ�`�@������qFl��P�#�h4��q�"zd$G$d�J���v��T���C��NIP ��{�5�♺�n����斥J�⢌|�;��m��<�?��_*)�f�Q�\G���E�|��x�lS�D����K����ew�8͓�@�(ҽ����81��Ժ�̘%����Z����TȒ[�T�l�y�������J�nҵaP�-������C�x,T�'�g?Mk��F	B��n�
RO�<�z�f�@����R�0eG�ʘhv�P(�c���"S�^�(��ǳI`3�/J!`䜍[R��"�L��J�X*@k��U9�Uq$�+��(�1�UY�������7r�����徿��.=tlO���3&��5��Ӛ��,�M.5��z��R˙�b)�l��X1��E����Cj�޻n[K��h:��lX�����ؽ%���{�R!��~6��0{�rN*�V���
�m�zOk���u��G�2%њ2p�ʍ�	�*7K�u?�dt��p�y_�/砗��s)_A�]�����|iVC��_�[_�3��x@\`S-���샰��¿�3��*��_�����.��֐����ɞ�#�������U$�����u��H]~ȿw��fyE2��X��h���` ұ���>��t�@�u(�w�=�)
�1?�2�fz�
�<s�K����Uv�.ksʷ�Ŏĩ��i��}n��S++:�Ys���H�1r �ReX�(��AW3@_h�WQM- }?O����rr|�2�v���iS�����A~�x*�N/�<E� �#�� ~鸐M#]�Z��8��*�����P�m2������2~�H4��t
�D��C�9㭃��b SG�Ȩ�8��P�|Ha���k��E�>�hU,SĿ���	���@��H j�7=nſW�~8�go' ���D]��P�QPb:|�l�&����26�]G
;��yo1jgai��8ߡ��������ڜ!ș�S�<�T�ų�1��&�P��KŹ�S1�1N�5%�����sݰ[E��|��cNT�	���p��� @�nXl���l�E8G ���P�n�`����a�	�ꔢHyF�>l9����&�I�������`<t���`>�<@:4�ʠ:u��d�Xg;n'@�� /2H**�ZUʭ��c�����ӹ�,9S��;��
��"��Hq��a�j%'�0{׶F�,w���+>;TR�5
cr��(y�����v>0mY�ct\��\Ҍf���e�� ���g�ӫ�ͼ���55�Ɨ��ߦ�3e�Ȅ{Y����f@u�㒍#w����RuM� ]� ^���������^����1�����=���?VWh~�s_Z~A0��h�NO(��B���vb}��Y>63�Q�nL.��3o�p
�7����a�Vl�RN�'a�),���"'c�E�����u��P���ҿ�ѨG�����[Կ{Y؞����pRW�z��$�3f�Ѱ� �G�~�&;-1���so%O?�CH��7k#E��b��pF_��O��s4F���,����4V���?
�q�JkNL#���+t4E����Q��tج:
��7���P�jG��J���X:�܎��U��[��g�HO��R�L#�E�hY0�2�j����BϹi9��|d�pc6��0~�i�Lg6`I�q�ȇ������Gy������䆰�.��d �ڂ�����'���D_LI@�*h*G�l����6t8*��i�cG��Xf�4�nKd3P^�"���/�R�f?�J���5k^c9Вi<cjcqr�^�ީ��� �cg��i��jC^�ы�/�
wa|1>3{��,G�D1��[0
	�mg{Ǯ�v�=g���s�I�5I�6hY3;TG�ȇ O�yð�\��ej��yHc�,�/M�ʮ�i�]���bG/5���#�|6;SCu�@i�rڮX.��k[,��#�����8v�(��a<���Z���f��hr!����\�G����D��n��6y��wH\����Jm�3<�h,��������]����ܗ�G;��7p砓���|���%��������>f�  |���kd��t/'�7M�?G�
�:l��`���v�0�(����|�y_�M��u�]���=NuX�<�I�ss���[���1TX��
ff�3Uֈ~��l��&�vS�@��z��z� ��i���⾈o���Z;<u�����*��h�gѶЅ�����._��:�&�U)&��º���=[���t]+�iC@�`n�Y�C�U�O>c��Ikbզ'�������Wf1a׃�hK�����FM5�����]E>�H$(6�^ѡ��B��U&}�\3O���H_��?�
O�1��<�ǝ�mX�4b���<��6,t������`�x�1����������o���~������xIͫ��ԮYP���.�CC��v�v��y4�?*�ѳ`O�t�	�O��_!V��dt#�s�z�������\��fZȭ����"ŘV��M��뛬P��s�������oԒ��yk����0�K3�UY;v]��4Br4�lRsݐs�⠨�Rۮ[Շ۴���P;�7�\s���=x-�Q�D��� \)�ǿ�����x�b@�ߢ���4�>	8q��Tհ�c�Cf�;ܴ���T�ͦk�✭j�!rGW� 'Ϊ�*����(jIk���"���
��M�m��nOL���U�؇�I&�g���}$Zh}-�����?���6�]�@u����:�
�R�k�h�����/b���6��z/���h��G9q4��=*ĕX��l?+=��LCe�:@��0��h��h�����ǃ�f}zTl���GK�G�{��NR�K'�7YP��c
+%R�C�c�Vu�saU���� 9[�-W<���b��`��p\�y� ��/���@gJ��/s�m!�7́|�u�`��< ^\Á����U;��Ui�$vk^XW������S�<�a����6���g�#�l���&��35ehT�C��Z������Ps�?`Y��M���ۜ_�*s{N{Ӛ�]���rb�T�{�.�+�G�,��m��w:P��߅��C~>}Q�iɘt�ƺ`5[��tjB�f���Z�3
�4���~�-�Sb+�S[��J�gJ�C0/��+�Vˢ^-�7*�N�aBkUp_T�π�Bk�Ճ����^��uջ<����~�A��g���>EE|��gc���}C{K��B�DP�ye\��驧�=� �����ד�����֪��Fǈ-�dK3��^�����}
��yr������_Ԡ�h�H4S�'�4E�vG9�2b�z`�ˮ����J"x�Et:��4Zb�� IB��k#��R�-F/�S���y��E����ֿ\<�e:>���t5����� {�f��F�Ũ<3�a��O����^e�����z�L�U�&�m	h�R����L?_0>Z�����MĈ|.�2;ĜS�ȭPa��``�J�3��{�����\aϷ$�����t[�-��m�l����#o732gv��̰>�v�?����JaQkӴ����0�F�o��S��l����0����Rn�.ٱ�� �;7  ���Dv�5m��� 
8�>h�lpsYj٦b�M.��g�Ɣă����6�FA��K]�X�J��9�����f���ݬ�t� �f��.���Q,U�]{�Aen������'[�����Ŝ
��P�\o|跈+|C^b��ԅ� �_t�w������X�26,AY|`��"�x�M��N'8m��=����6� ��t+�[�	����4����
:{� f�R�)5(-b�ZmG'�����
�rx::҂�r����
���r>�06����^ `��tʢ����2�%ߏ�Y����fD}
\K~��អ��wv�������D���!J�Cd\�rA]�E9e�{G`��FM�},�\9�(����P�
`���1�o,z	a������2U�<8qi
�jgy%�%�%l��f�Ħа��P|)k-���)m�e����@x:w�sH�4,�J��@h�y�z�����C��`o�u�k��6�Gi��	Յ#f��Q�#�cz�T�TST_L�7-o����R���/ݨ��'�?����N������d�5K�HF��rQ���FJ�a�G91��ӳ�*7���T	��Q{������\��l8�4�&g�=9��(���{�\ӓ_�����?3ޡ���m�E(��ݚРXYHED����L��v=���A�Ě.��ܜiqTgQfV���n�1�:�=���7J �앂�$��,C�(xD{�m�%�6*)�(����|̱h�nU�2�P�4��o@��cr���Z���4A����^��KF�;��A�����g-3Q(�P�eהNa0"|Y�Q�����s�cU`�ݟ�ٳa�:[��O��{ :�k�����<-_���J�P�����g�4��/�p�<>�)�s�d7a|��B��ϋ$f7b@k0��9Gs� +'�2�)c�(('���t��f��jm8P�� �	r72;�r���-�![��� G��DW"G"��ٍ��X�e���Խ���P���T���iw�ކ�|��X�yf�(s뾊7ʏ�'�KT։��1���bh�q����)	�}�G ��Q�df�J���V��,����t�s\�<H[��ByI���S#��a @�j��mՁX�]�y���:��r$O��_p���K���@��$���ު�Ԁz��gA)<p6a�u�p�RJ���w��B��ۃ�(�|��o�����"5�ށ,��>z.��d3H��Sș�.���AgDz,f[k�Qo5slFm��4�3նP�+�������&��d��wѩ@EE�];2w�3ޯ��D����M7s��>�e<�+�����K���pmw4�����օ/�������(�g|E���V=Z��M�BF��� ����C���V�U�zϼ{�������_ ��2X�d�����:b�h٤�rNˌBdtLȎW��_�M�[���;���;D�J9F�_�E �"t�w�x���ץsi�#Of�ll�,�-@��5I�/F)�N+��g4�z/d����h�=�Di
�ra������Qu�3AV+��@�n��I�0V$��o`cIԙ����C���ܡ�k~hm^��3�`Lc���2�dJ���x�9G��V����*��u�`��FD���Su�4��92� ��t��.��Hg�L\T��-��G�V^e�OP@��1�٧�l@�Y�<ZF��@��=�Xe�+�]�2;s�6з���� [0 LԖV��w�r������R�e��U���D�<)�y���B���-]P�w���[�f��6��E��z���V�M����W=3�,��A�nk�4x���*�c��<�R/3bO@�{B���\'���lLs�r�ā� 0nf�I�AG'
-����"�vp���`:\�<x�ôn@�Gwf�Q���6ZX�L�yŌ����֞[�xIZ���	f!�
��.=�{̀���Zې��s�3�.0�!��}����-�B��jv�j��U�pdf ����l�(�(���A�Z�oTD9`�6����������	@S@�z��R�h)s�&[cߢ���o��L"�	��}�Qff$BrFϯ�6W�xY&�ٖ��k�R�+^mm����s�U���߭i���~L�ͮ�^hi��)h�/t��4����H�`��5� s��5�`7k���a �����k���l@�	��ݭQ�,���*�?W�p?���vic6���6<ߢ��(,|
����]�T��7�������+;��U�E�U>�Vq�X� (�E}L4g�VбKkA� t������td������.~g��eq��n��#��v�sB{(������WY���uO��ί����I�ʯiT�1�h, æ6F@fx��n����m�1.��_�P����1qW�1�{��)��"�����; &v��L�]9k~�r]�(��l9E ��R��ж�����w+U^�x�]ya�1�YA}$���=�`u����rh����x�`�rT,9 �Zf�Ȍ���
�:�P_���l�f�<B�(�_�nD���� � ����TxZguc|����ћ�p'�����l�6�_�."--+1:�w��ٞ�{<�{�5�c��z�/6�����d��j�{f��L�%���r�q@.�F�<$0����t[�b{ N$�f�֙�.���/��ZTEz-����Q�ڢp#���B�wEʹ��,�Z![;�lÉ^�;�qxwwϹ�$q`��PU@w�c���l�Xޡ��i��#�0�>*-��Y�d��(
j��lP�����-�� ���a1��ކ���=�JAc#A�#5�m���S�W ��	T;�9���g�90���5�ϰ�C� �7�I�Z��jZ_�B	ɡ�A��6X�n+]G�ު	�!����\���'`�dc��t��>� ꋶS�Oָk"�3_F�S�,�x,c<�Z̝�js�~��l-�t:_N	�r9������^�uMG��&viV6��d�W^�Ժ���<\��43��I�|?�n��a1�v$r��fC͗�8����4\ں��8d�%7�>|~�n�⡐��k�ߙ���}��
ժ�(����zS�4��غN`%�k����g��P�Y�#�3w&N��Y,X�0��	�=�F2��'��3`��j�C�ݷ�������g:�U����9�(��)1U���>��J��#FuԊ�yi�~˂HN�g�����S��5�
���h �IS�:\�C��nM�ĵ�Dr�hY_M΄8��KʥI:m�M�d��n��{UZ[���!U�5�xv,�ə+3�A#T8���K�p^ќ;fZn0������XC�	 )|����=����-�����2}��g��2���T�^��� �0�g�(��"�' 	
Z��[�����:m��Z->9��F�m!;iSl�K��V~��b�ߠ;.\�%c����A@b��1î4"� ���W�t�Wk�"Cm���C� ��o�5_�/G����]D��OG�yh�\*[m��&�r4�5�陭�t�ٍ��n$r���HȚ�����I`
�mԥ������k�3�r�0�;}���}�y� ���Vij�qQ:�Z�ie�Xv���tdz
��>�S�# r0/��������r �?�qv���L��C�q���:����
ǅd���=��#:`x&h���::zV��-[1�C����p~��}0� \F����X�ϣR�(|,J���$�u'Wio����{I��Y�5I�
�j+a8���͍/�S�"[Y*P½Cf�E-'�m�3w?��`��V�ôf�������e>6��l�c�$W`��[f���%|���hD�ڠ�>��̶e��,�q���3��㠠�Z �s�庸���u��*� 4�]Ե6�hU��e��B����^hp�B��J��k�	�hH43f��Z�.��>ݻ��6Ѹ�e�Z������hR�ea ��u��>+X�)y ����ִ렁u�k( ���Bf�M`��q�,M�?-�.���z�
B@���E+8"b����;��E:Neԍ�����OX�Ǵ���#N�3� ��d���6,5:�����i��4�6�˷X2%>6��cy�;z��tM�X~Ҁ��@��K�JA�
�U�4kh L���+h���Wa�/��M	�"�Y� �-����qX�}�O�V®���}�p���
5,Ťi��� GwB�X�Sp��w��-E������+��2wY��g�@EC���y���!`mG�8���>�ʤXP��h���C;5���+�r2�JED+��(ʯ#g�:�����ݸ<0N��[ƣ7�32b�?��S̰�F�j���j���l2�����b-h�a��{���Q��#��*H�W]&׀5�1dP�;�͚ʘUa���B0R�l�sF
ˏ��E~z?c�DI?ʖ���^kd<[婕�K;bU�f �jI��V� �������单�@,^�V�MC�V"�d+t(2�Q�F	�^ߘ�f�8˶��j+.7�*�������	�����mU���YP.i��6���l�>=����[�|4�JN|��<�F��}���F��_Ȅ��
Kt: ��6��3��j�X�=|Ƽ �,���˙��e�q� 	C��Yz4^8k�^@Bu�R�; �1xn��	�r?*��z�IK�ps� �����+h�@��.>������{~��dc@y�vp}�λ�J�wr�ދ�tm�ǘL Јi7�s�T��&gY�o¸���>����s�@l�
�j�uuqu�L�����|&gײ�@,����N��a�K�,@l�f&�f�I��#�����-�-Əb�)�����y�>��l:�/x�?�Y"�A`��U�EΕ�����"��a��MDvo�v��Fy���tG���6��lkiY�'.D} A�h@��9`+C��d�
Nm6��bu)�_%ht�)8P!S����ZY�c���!`޹�=��|�\��2K��=�M�����ָ��i���ۘ�=���k*�*��>��B3dX�|6���9bma�]BkA�e��7j���a���lr>�����oo�����7V�ZA^���e��T�<�h� P\������+�,ד�Lp���� Qn�k�|6mm �隫ⓣؚiT�>�Z��rVZϿ���Տ�'K���	��-���jt f�i�	�!6ڥU���ۥ����^qm�>���xpUO�u���,Mݶ���p� 9.��� �g�l��s,�%]&��wt� ��mn����������*gŔ�L [�-�zʹ��55j�;Ⱥ��	��!����"��HZ��T7�&�G �jY�J�T=�e�2r 1Hׅ���{�2Z̼��2xd�~�N��-�j��}\�$�y��k-*{��g��&���QIڠ��Î�K������ ������E��:B��ǳQGH����L���A��%Į�"[�aD���;4!�<�[��1q�`���$ �UBi�Fx�P�L�ë��q���<��0�p,�$�� �~������9 �qCB�NA�)�������\������yP2[���Ò�5W	�`�1�����ë;^�����?��B����xk��ɩ{3Q#t� �d1�$�e�T�
?��L��/ӽ�tz�����Qn��r�@Fټ��\\�(�P����kf� 9zf���|��:,������$��V:#�l#>|!��ų#/��3!U�%%����s����eV+(��6� �+����@dg6�%�׌����3;������t��[�8ܫ_����۱��7iF/�ݦ����TΒ��?��,8 �����SJ/����O��l�;���O��R0�&��а�{�u��T��/������L��$@�3)���[j��f�+����mͬ#K�2H�`�&CPj�@bͮX6e4�	�@����*��3^����H��ME1b������z��*���tZ,�(����\b�v��Q�ۨ� �{Np�w�u��Y���8Fa�UJ�IDs�V[�N�=�M	�8@�h�R+*'V>t���3�������6mzOzV!��5&����%�1����+n��e�d1�T���.�h�V\G7{G��r�������n����6��aa�kU��E�<0�fD�eS6�uɢ��^2���ЍC����X�I�RvP�@���2`�01�n�d	���&g�����3��I��I����o���̗���j��	kkp��[�"�RNkQQnVƫ洣��H�yc���o�hiAi�\k��U���d��n�H��f��0�3`������k����E�lA���1�a�{,<�\21Phm�<�w��`�o�꨿�ܢF��SBYm-���%�r&�$}Py��R ]��k���H
�²�X3A����ݤ�[ ���j��k��}H��6��ɏ�gj$Q
B����@q$US]ܻˊ�D��Ƒ�yf�6J�EUw�l
��V�|�;N�@E)	�0��R3oQE:qI��E�Qp;�XZA�>��%� �u��*f� !)�;���ه3�n勵kw/  �X��O�K�G��{���Q;.1���R>~�����`Z���ҵ��.䗷����Љ�ظ�#fgg~H�������	�(����/�7,�_L�>X&�yIQNྐྵ_����������ށs���2���Sx���#�;WV������H޿����<��c��Q'0rFݠ���%>�s~X<��ߑ�5�\�Y`�8��S�]��C�' �A����C�g>�����<}��sF�*�Zt)�g����c]]\% R��fs�p8W7 #�rw�T�Ѱ塚����h����Zo~��گ�k�H/.n�ҩ���=�	����o	��R:q����C6�:���&�E&�#s�2�"�.Ι��M ��p����P����Tq�J�h���&�C�_�8����Y���/��Q,�<L��g�%��qPEE�iT�;ݚfU}dy�(��s�M ��L�7�5>�P� -�մ��#�d���	J�G	�Z_i}#@Z2[�5f�g��HP1 �1IvjȀ�JX��4c�$��k�/�? 0<��"K���O`9ك>LXG�3p(�|��{	R�ׁ{B���{��=�;�N�=K�w��`��h�	p�e��7�v�:��cˌ����ݽ�?�)�@��?�jNk �%�p�����A� nҚ��N�� �y:�L��h�}��Ç�j%af֐�Zr,����s�;����'��(v/,�I'�' p)Ӭ�����L�1w�]�-�#��(6bL�_���H���r<���΀��;v�b����M��D�5a)�T��NǇEjr�x�B�������w���{0�{����4qR��<�����wzv#�S��贰A���Z*�t5bs� ��@s� $�MEQM|����h���T�܈J�oyO*8�ɃjU���.a�t�YU��ƍ���j�pv��*n\L���D���3���Q�cCn��e�Y8p��qE��b�$A�P�h�l�i��������yzÒ���!��B5��f�|(%��ąu�!�G���NQT3I�l��ad$z��C�����IWƳ��Ua��|%�w7��M��A���/.��}�f���O9�Ϟ3��� �:�N4�/�P�B���O����.���PǠ�Ͻ����~w_���������sf�\�[��ˏ��FKk��
�����Y.a�f�!jP/����O�%9�b��R$��98'Y���Z'��J�Q��â����A�}�̬%��|~�NJr��&�UC�\�xJ_y3U���&�������Iw){�qT8Qdl���o \��0+)�b���g�0�9�s~\>��N��P�5����\���C�(V�m8�����o���@!�
n�<�(��6���!q=ݏ���
� ޻�-'��'� ��뭖H Bi>}G��K�%����ߛz� �vX�6�q��9/����`*�z����⃌>~N�1Pm�,�a#{PB_�ǛZ;�8pr.���\&���)��y��%����%A%��[���B�)�#iu�@ʤ�E�q<�k2s�hp�~��Z��;� ��/	��J�P����<��1����4�s�@���rעf�*�O��%�=���K�a .d��l�9Q�_�,��8��#D`y�������o4��.����>VF�p�-*��`���w�Y�}�IN7׼�!��۰���c9<ؕ�/���a�xA��)�o,}L�Yȇt�R�ί�����G�?;����j,#��A,�K�̓ţvg����g��vd�oSp#�9�V0}��˗���Me��F+Km��!�������Lvf��;��mz>���S��2��Z�yu"߾y���V�E�]��%g<�S0W��svMG&�lOTH�[�k�JWÌ���!�8�����_��W��M$e��m�F�jF�6dZK�T�V�ށ�M�E��YR*�wX���<��y�Y�F#���b�����[$kج�t���e}�ݿuZ�wo���?�,���iNd[@>G�U�Q&{��{F�hU�n�u�q�]e�;��.B"3�|a�K��� ��W+������P.Xa��*�����iC�`�Ul�xJZKj�V4��РѴ_-�C���t�)�<I�i�z�M�Ե�vYj�4 JcmkI3a�
��D�Fŭ�Æ�;�K�f��B��wwv5�fC �FBp�(m)ɹ�R�r ��Q��A��5���iFQ��7���c��Lfr��Ŝ��I���/�?��}���]����\�2֨���/7��m����G�v�3����[�{�0���F��A�	�$W�u2�#��]��������`�@Xv� ���X[�ӛ	(\\\�</�1P%E�,���.?�z8լ ڷ� _��Vk��*�f8]�-I�t�(�=��zI��n��Ŝ��̴5NP�Y'˞�?��w>O��R O�⃥�����p|h��OeA@�<��Λen�����[�\��R��p� �?�&����,7��ڥ���+�C1�$O MCp��j��l(EQ�D� J��K#���=�UX=$�v��F�,FCn\��k�14d�s-��%��[%��!p�
M��}��t t A�Ռ�4��ߖ�l�g�J���\�>q�h�V*�A�Z�Z��$J�?	��r1��	�p�u�'�C����i �^c��525����9��2�g ��ٔ6#X0��
	�����ݗ�t��طf���Z��h��#����_�oE�ղ72�ؿ��P�t4�gǻ��ٱ�iv�4�
� �s/�yi&)�=�QH*^
�җ�k9Kv�J�p N�U8F�;Syu�'��L��v�F�<�\Np��+�ӳKY?�K�jL4Yyy��"k_^<?J�<d�����J%�	}3{�jI����p$�S sz������,�f�&�'���L���@Y壔�s��r)�dS�r~vE[|������[J�,�R��� A�&qT�G�D�J��P���} ߊA�ξu(C���l�W�#��?k�UoV̙3e�W�E^nqQ*�r׬g=���-.�g8Wv�97R����4�eI���O,~����ܣ�����j!��l4 ��H[�JP����"K�q���x��p8eא���V�V�K���=��@��:{?S��Q	� �>��?�*���>E�?���U]~�Uģe/@0��Хq`��1y��8m��JΏ�Yn�W"��pH0D?��ڴȸ����}��W�tͦL��^3n�4R?h�� ���8�9@��W�^���hf�Tk��������Q��F���h.j64�X��~�NXe���Y5KF�8���=yv�>������QrD�I�,K\^^�H�"��Ψ��Ǧ�����N���d���<K羓-�!���Z�U��-�0b��\���/��,��[��29��k� C]���2�Ɏ�\B�-
���C�h
�N�TM�Q5�s���,%�3�c�%cچ/6ܠ�/�-jW�J��CQ��C#����|+���1�T �J6ϲ1@� ���Q��ĉv>^U�F�G�mzmU5a��nTo(���TvA3�J�.���D� �3!�wK��b�1�!T6�
6Z�_ԑ�k�Rj���X�<��&}ތ������̭k�
�آMJ�fVe�HNi�Y͢*s�8;�R�\���f[ҳi�u�D�M�۠���BrV�U�*F����Un�;,u6�,��YұT�6�v��X�/hGfYz;��>��Eh��`��h�`��}�����#��5�~�X\�(�4�`"���OҦd����C�� 8h���������y-��Q���`�_���hي�;t�
����C~�q�+?��g9>~fݺ��&��wR�	+ڐӽ7���)�lՓ�c���t$��}����rx�)#�0㾢6]���r����cp^Y�j%�������<uf�@����q5ώw���N�����*������}ؚ���ݰ�<֫�Sy��2S�]��l�Ky~�'�_��	�}QI�"v]��}B-l�f���mJ�n�����)�n�op�������,5�Sx���˲��Z���ѐ�	�#|'J�x���^\�u�y
Bo�������Y�W��C�j�l�&���&���{k{�t��ev�:�N��f��dH�R���N�V�y��wɢ�ܐIND/C����V�F��r D�Ǔ������,6�JĘ?�)��ʌ��3��8KB�� l�DJV�~���ҿ�tv��t&�	҄�I�̜@�d���������5�����������v%���ſ���� a�ίO��r���0�%?6��^@��rnr���P�N,���೴;�Q�v�d�@�^��9�4(~a8k��� (�6>	�Q�U�{yL���<��xS"Do��+ ���8���F���/�͛����30ͮ�|�����&�G7b��ϐ�ߐ���z^붵���L�})��+�g�D�;��"�7���7�_����`�l�E ��ζ�����	b� �c�:��BZ��o��?����{!S���'Њv��o�D4.i]p��|���vpݯү,��39�l��(,m���в�-�S'Ù��" �uS��h4`p�	~/=8����\��H3��h`y6uc��'j�k �c���^Bԙk�E{��ui��6p�P=S�W`p���*;ܘ��7l[ǵҐ[���"T���"�ֲn�@�A74����>l�v;V�
�	 �ҳŚܞN�^�=<�R�a�Ѯ���杂��'�q�m�1<�!�I܎1@)u�g5�6�LuP�M]�h�mԌ�f�4|ӽmov�t��i�m�Qb9{�f�]�T"x��Z�P��޵��+k�w.��+�9��K���	W�-4}/W��ϸpm��,ҳ)[m<ea��3�v�N0d�5Q�ZR T���`���qh� PRC*�l^a?�9b�Xr��n�Q3�YYA�rR��D���ŋ�6^�����}.�ʩ�M%-���t���f`��$J�w�]�-ӄ�@?>ܕ��)m�D� ��ae�\R���U6��,����RW���p���}y��ɗ��dwg�>��Ώ�$�ḃ�p�U��\ov�==I������%��RL�l�(ݟ	�_���T?L:�j�2�ډ� �9g[�{����wa�2`�
"�ȌZtޚ�e��xlmt,��w�u�nUI~�,d		��v���$g�q��JEV]C���V4�!s�F���MBx�Ff�]RE����B��������=��(t�ؤ�f��$�d�Ι�\2��x�D@�'�j�����r���J
������H�#��0�h���B
)DpX`�P @h�(���1�9��y+����3di��z�g�:?K�y�d2�ۻ��@��DN�����y�G�f[��(�3��h�_�f9p��.��"o?|���6Q#⒳�L}��N�_���9Y�f
�X��JnP4݋q�����勣�Y{tp(-��7�&���V��o/��	�����䘮e0�J�m��*��"�+��8C9J�r{2�Q���Ǉ�w���z��))Q�B9d	w'��dW�M��/?�*���Ȯ���BTy^���O�lZ�c�*d��+��Ry$��t�C�b�p�� �g=��$�'�wRt7�O�[���b�H��Ȏ�(��(�ʋ-�O.u_��ӗjZ���@�8Q����y�2M��K$w�~�$Y{2���:I���54��J��RC��Buv�|zNDL�-g��c���t`�j%�̴'���k��,@'�e�R"�2+$h�/�Ge��K��Y��:yè�#�lD\3:���ȺbB�0(��%��Im�cy�,kW �g�lGlY��I5-	r{�d	��$9���>��ճc9��%����~{'������'�[$C�T�R��PZf{�R����o^�H�}7َA�l�6�ۍ1��UZo��"3��"ff�<o &�Kɚ}j�79 m�ܢu�z3�[�ؙ�h&�-������
Ŧ���{��h]���C��B��,�ɵ���}e���޵��+>�2��S�`&U�i�%����Ո��U�8���R�YCs��u ���zT	
�k�Y�%��vw�ͫg�6=��(&�p�f��O^�LX~o���`���^Z����T��_~����"2��z8E�K���V���s����5AV��}΁ݖQnŻ�kVo����N')G �Q�.�[,��= �m�!G0�����=�Q�NOɟ$UݎЏDً�:+Z&���J�$����\u2�&�w�GJ/��X�s��q���,���k�m����]b�j����:�J�#�S�֐O��������?���\������}�O����J�� �U
�������>J-�Y�cE���x��*q.�4Od�Y� C�q�������ڼ�L,7 7`p��,������'�w��7���]�N�ρc�ө�Q!`�,����ͱ�P�&:�f6	|��@Nt�F�7��hs��ո����2ԋެ�k��e�n�~D�P9eh���tƋ ���H���M��Iu+ެ��&������r~��[���KJ4V�X�t
|͔P�h�D:�o�� ��EL���%���P�f��_�������H��˹s�J��h'Ek��H��6S�9O�mNT=�m'06� �D̝C��˫�{�)���w�{�4�
�="�<I�g=.eog��ۄ�x�rz)7P _�R8xF
8=�� �Qn;���w��#�c��ͫ�ߞ)!;��d�H;��	���!zK�]d ��&0�ݯ�!���c���h���:���Z�h�.l(�K2y���z��v����9�8dY�u8Us���|�����i�D�E5:�R<��y��������f�w��H�U�Y��H5B�~P3
 �-�A��J-r9�I�jp��4,#x�&�s�\/[����js�<�#�t���H�ln���I�;�d^:�-��7�_$ ����6[���C������="�F;oE��)J����ￓ?��MZ�3�׼�%~Y��$����g�vbl�#[p�i��^k�¾��f�<�e�w��,���#G��m�{���v�Mto����H�5d%�2��i�e�ܱVu�$�=�)���#�=��e�bQ��Ԋ���~5{i�5>�vh��zi���ь����(��䈩=׊�h���s��u+)K�j���A
^��A
b�v�S�����L��b�)6: 2]/��'���l��o�❵�{M>fLF�$z�ݤ�:R �h�\��J�ʩ̸���~�j�6L��ˇ�?{������G��.����Ȧ�l��{Z�މ6��dFh�u�lr)�d��w�xw��P�r#�I��|��{�^,�� "N!� ����/�����TN,�'x��HE������<����4j�ݟ�Wr�����lQ�@IK�e�,]?Բ�\�^"т�r��|)��d�,�������ңڄ�����;���΍pt���;�1e��9_�ϝ��q�`4*̀�J������]��)��|z������]�,�]:7_^�R=�;�|G����^��a
�b��CR�C�X�VG���/����Bwq!��t�a6�"I�i������t�d<��	�i9x5�((/�`�� ���̘�aT�*��\,���k���;���I�>�&$�7J�i0Ml� ߄)Cl��ˀ��ƴjht��$Q�.M����1��+�H
}�Z�j���F3<Lw+�o������]GH�Nj���d ?���.E�ߤh� E�	[ɨB�M�V��v[V1�hq��6�������������_���_�I��aQX7� P�c�yy"?��&Eu���<�s�Z���0���,M!"L�ut�#ۻ�����.��������̦�^BXV�$@�j8Q"�� �:)�b�K�0l �{{{���+f�nn�x�	5 ��-�g�fqTju.ka�ԝ���dT}^�S��g@$o�`\-�!�0v�#�kM������N�ٟ�v��d��F|ce�|O�d�e�=�ssia0��\�iG=퀂m��g/wEK�q܏�X%���ҎZ�Y.�� �?Mk��3 �o���Pf��2�.$���g;^\%g����V�\)t}-sF�/���/��[y��X3ԍKNr��=7���6.�܁²���K'��~[��%_6�\��������:��s:�u8�#�N�Y$��RI���>���4���CZN	Q�#�t��2f���#�C�ʞS��M"D�qJ��u)Ш�F�@�1FS�o[_n˄ZV�٦a���I/������(M�rE�U�hbV\�d[��`�͚�V	�\a}$�N>j������3�q
B�x��Lu����5/I���+��K6v�u2�&&����p������>&	"���ro�=?ry��b�mƳh���N����]��h����Pk�Э����Ǔ}o��߀�B����@�����	1(���ܒ���H'5h3P��I��N�E���r����#;=� ��`O�7��A�ส,nk%���{��Ç3������qop}�ހ6������صV�>}�I6�'�������<?�g��'G�_�@�x$�ɱ�,bH�4��1�)��O4P��6�Y3H���;�����.�h���^ų�c�I��2�?�= ��zΖ��=�6����N�3U�(��U�O�P1`E��ǹv4��+FÌ����&�'�舥C=]��#�k�N��9�aF#:�U���X�v��n�2׆�
l�hL���~����M��6�������w�嗷���UZ4+n�j ����J�k�L���Z{�ʥ.L*� 1{<Эc|�\V�5���qpV���c�ݴ�R:��J/�"]�.	|kt��s�ܗ7/���?%P�"�|(T쏒 �8�J?��:[��YrL���E��:K��[vHnt\J�;�����������-bhq6ΞQ�h�_jN`ob�Y���3!Ժ�����5��/.�׿�iD�*���1�t:$��$�Z�ek�����bUS�m��������!7�:٥h�Sc�%�~���=+�t/q�8b��ň��,tX`��;U�&���������`P�>t��J1�%%���"t �_3�^�Kg��m��yb����)��E)������;��}�R^�<&�H�\
H�+��n�@z
�f�JKT��.5̀N����^~��O��B�K��D�ǉ��G���!���!���i_R�u�X��4��t�(���su6d1J#�igT�|v�F���8�N�vlϖ��	��3��NK�;���qZ��-@�u�NA�����ks.�E0�|8���2 D�N6�� ��{�i�a|G	����-��K�F�XD��ʇl<�L�D�p��������珔e'�<����*��y>y��e��8j�	�#Q�*�7��l�,+�Ϲ8�B��R�ͥ��&�h(�Na#/�]��}�L�����K��Qe%�.�����k��|��2^�;���� 8�l9C�Ҳ](��_�)Yd�h���|� ��W	<��xX�5��_�NC�|�y���xL�����%�ɛ#�F�J��@�l�:���>}��l�o���Y��{j!�^���ú�����x_3gG�s�Or��H�}ò�"��"�C�}�`�b��@�f�qC ��Ym�W�@c2B�q��/z`ղҺ���n;����kcg>��Z��e�qs���c J�{��� a{��iZ��l��W����e�������]�*�7k�Q��X4]�o��Ƭ�i��w��.MmL�0�a��c��k4��" �i����A��,�4K͌��FK��	6���b�6���{�����Y�����?�(=����� jㅲ�q�ę�@�6z�!�h}Fd�2(e/L��И֚�>�(˴�{�� 	݃���lņaA���W/y�ۛ�t��k`��(�̳�`�m���FL��I��$\_]�ĉz9������XV��Q�"kO^�:a6cP�ҽ��:��=�ۑ	 P�|	 ���+�%(	Մ��@7���!Ql6zy6����h�O���3j)L���g'���~�^^&#ylF���Ez�y��_ȪAZ��hu�h�X���`)�_�
�z�)S^ސ�~�\6�lDG?4�%^�2~^�uh��8�ɮäU}Y�+�9���n�������W��Q�>�/^���ze��ˁu��ʝ=b$�X������w���^%��'y�옥����^�~=D�HV���mY��6�sFw�����g������߼�d˽f��0�����҃w� j 2""�&E�W�Y6a,?��I��@�{a`@���j���5y ��~@�Y��}Ϡ���:��~֍6	�i�m������g�rQ9��nʪ6��KǼv�����E�l�(�f�A9�ɢ|�`�u��6�Ӕ�4�#���^���غk,{�§�9f3lJm���JPރ���͍���An�o�:ڦ�.]=�ɳ�wr,Ӳ��(CN&� @������1A��x
�#��HwY�=<����i
/�F��j�Z�[�l���t�mV-�&{$ߣk��Gdh�1I8f�z��  ��IDAT��� ��Ǉ�N�^\�Nk����`E(ԣ��ri�N=8#?4�y
`o�o����5�1�|j�=h�!@E����w�B�W���E��ɞ"0ğaw7�9��)�d �{t"��>|x/o���]RTx]�j`[u�v4z��ǖ�Q�{jJb@���^���-o^�ο|~(�)��6zn�Z	����H%7pʢ�A��j|����b����v��Ս]�{��Y�.�ۻأ�^'���i�����,!&��Ky����󗯤ټX-�H�ݬ���E�9�C)�bUJ�|�i�8����A?Q<���bϊg^�[t���L;�D�F��B����r�� ��q.����ӡ�.U/�,�|� ����������^�:M�x�/�e(T#T��ި������ܸ������a�.G��W-��	�Б�������/�5<{~Bc�tʥ��������u �g�T뇞��dD��^����9�^� ږb��`"��SD7���d��ó#��2��8m�ݝ��NNY�E���?	i��YzMY�d��%7	��a��-g�!��#w6��@�L��o���
���#���_(/����K�!�-�����	I�H�Ci{��ӳ3y����.7ZN�Sf�6�\Pv������҂9\Y,K�;�3=_+}0c@+��"��WpGhr���{u�E���
�: �s�|�fɴ[/J�_�S`��{�z�,t6��� �w�=�� �����ٚx�^��]�>3�hPF������o�ẟ |�����[��jr@7V���3��u��E �*�㴞P�Bp��xе�N��#�K�:y����D �q
�vw��E2��w��_��n�	��z\]��ק�7��ݠ��b�ٮ+�Ղcϐ���9 ���B���a��o�u��g`CQ�,A p�Y��GS!o6ۿ�K��&��һ��L ���9���ma)΁��f�U���v�0�4�Ł�x/u6��5�85��3�O����A~Z!\�f�M>Ac��t+ʔ8��{
�%j���Z.g�538UV��u�H��A�)�N������1��\JNA�`j�������w�#p��AX�.�����6a�����<&�����+4��Hh&�8I@nw�T�B|����fL� T����x���6��M�v��Zk�w�,��)��8��v�0�	�B���C�a�Zu���0	��b���}!�07�
��pt�'�;�
�����Ge�Y5�4��T��c�(@�--1�-Y�����G�/�K�	�e����_?�Lk�u�|)*:(������sd�v�����s�{(R o4<J�h��eDRL}:���ؚH�\���'������3r�x��H��� 'G|�F�]a����!��O��;�E���<��|�z�����;��1"K^�eC�����ǖT�)��+���Ӈ��`�7؅�ƚڧ�}�:�4�ߤ�q&���Gj���_���L��%��4��cV~�.Y'Є)�G���C{M�8����@�۷�ɯ�����9��3ZN7�y�������oK٣�j�L:[_$�,dH.���GqR��58 �g���9=�dvQ�3�V�L&g���0s�MC��7��&�PƠ��1[�H��T	�~�B������Ä��|?�y��[�/Rq4	�]I>H�a�)���F��q_x_��}�x��k\k$d���@�ob]�iD��I�Eș�{[={ut%���p���5��g�|��Xפ�#����@��݊
�\��?8���	�@�r6c���\�M�y;��o^?��w?�M&vq�#Y�L	�stp8������g���Ǝ�Od'���ƫ=����Y��0�E�r����kUU9kYS{�d����6�,�1 ��K�Ys��-�KSKqɅ|z�/5�Oz K$W����{$�S�O$9'd��?'�l��8�̫
��e�jfZּ���N1���Sn���1!_����XP��w��$��������lj�q��[t0�gW�x��Ϛ���s;r�����nYt:��L,`"�b�t�L`ǆ��}Cfh�T|�#p�y�$��yǺC	�nPQ9����IBo��߿y)�8z�m�����ە�h"����~nH��$����������O�X�kH��n�!��6P���t0\��ONN(���7�K��[�^��:j���������>�&�(a�䖠`s��pz�jP�p��.�V���)�M�L��2�o�j�E��WW,�:XƜ�8��j��H|:��D�w>q���W���d_v��R?�m��O,t`95ٌ?�{�B��va��s�#��<�ؓȻ��|��[e����e}���dA��`έTn#ʩ^��n�N��31�C9Q"�l��9%����i�ea��x�"� k�����+�z���G�f<,���Q��?�J�qC�yK�3�ga��mr⒄���}/�~��3� >Z�Y��#ހ��`*�p�6ۈ�nT#J�?U�I}��`'��G���X�K��D:�˫X�n�`Т:K�ߡ� ����������L��`l'��7����/e6�d�3j͟O�X^�5�>&`��1,<��t���^��-s�YÙeȂ��" �M�ur|�6(�J���A������]`&�b�B0�ty;�<>:Jv&;,!VL��R4xtp�a���Q'�î!%�R�1��f�Z�A7���dKp2�V;�O��SQL�pL�j�ค2����k�]=�s&V^r�7�,hו�A��/�`'��V�m���TXJ�zN{Gs\��&�@�� *T�r�U��30���hγt�K�Dɿ�ߏ}�}�o=>��O�!���p>���! �NN����s�ƅP%�AЮg*��Q��Z�zNRj�Xk�|c)�Yrj�EI�T^�k0�!������S\��j�����H����9���3Z���|y�#���Q��$�~��E�goQg�b{��2�϶����z�߳�bb��#�OP9�6�@�նF�@G[��=+� Z|DKw/|Ԗ^�fy��<2�,<�]t�p0��,GCdA����od:��AR Y|d������af���m@f��ꜣp��pY��X���ʖ�,@zP�d2*�(Tl5T:n����M6�d���\'��ȷ ts�қ����&]XP��)x@	H�&-���EI�x�0�ߺ{|�ͣ.]�ݑ�j�j�TD+.��lM@����� TX1��:����t��^_����떜j<[�5�F&L%T��2��2@�{dA�k�Vȧ�4m%�)b���1��� ��9����G�fӞ�ٝ��� �����R�5����K��R�.I�ٲ�Lu�:�t�)��߅Xz��@2�T�5т�`z��g���=p���Ɩ9� ����:E�T�Υ��N�B�Sf´�7[�Q4$�9t�@�Yy#���"�@�Ѻ�.���rk]=v��4Gg�����v��}���έ[E�����"}D)�@�j��,9�F)�����-JP �L P+񲶨#�I��@B ���[��ڴxZ�;��~���ù�3���@����3y���l40��*�������0!>;9�����ß����L<2O��-8Q��H�Z���Z�퐪�(�@�1]���׋�'�IH��i]��S��]�!&������=F@�0�0��>��W-��r��ň@Hˣex�����;y��T�f[]�و�d'������u�.�@�Դi��Li��ZR�m�%c�GC�g�hp4�9�x��칛�ȸ��@ި�{���T�$dǷL�U@J�P�l<ɛו�sw��G�d�j �����]��,�q�"fE�+�a}��pc�@P�R׵�����ww���z`�Iݞ)�����{����E��#׺:�s�Ü�hYǝ�1߼�F޼~#��L�}Qņ���9�m�m�{2�T��1׮<�+���Q�At2����^V.� @\/OK/Γr��5Ǝ-���}A���KLR���g���X=�̎$[&�;���])�QXwl�����{{�8��������C�wk�;��Ѿt	>��%Λew�I����!J�Y��&s�3]�@�� L�yep �OT/��<G!Q}�!	?Yb���F��ve�����Gc��z��  8�v@W�TrH52�(��~� ޾��d?o/�y"�齏�~���L0�Nd�� (�;�E5o�<�л�dO':��e�
)(=e�7���(ٽi�.F��=��IcZ�a�����O8J���Z.�nR�~�.�
�iU�4�&�wr'K���r��:֌�F��
z����6�TQК
4 >R�վ@��4����Pj�JI��P+FV� /�Q�?l��]�D�r_��q�`�h$V
�?$ ��↝��Z�B?�L`�z:?<�!����Af	���\���#�F���ߏQcg{��Uv���9�!��� o�k��QqX�|�6��h5�>)(E�F�i�lȭku��d�E�E��b�����]���N,3���lhWM��/=�S����po�;���R#�2�;ҳmK"$"�n��	|]��م|>�JN�e���f	m;��h:BzbF>�'���U��6J����Irk�����o�a�,V'� [;��f/^������;�ã#9>>&S&k�an��Ņ����c_H7�K�r�癦�^��)f�]����7@�#ӹ�|E�5���+9����Zu�����j��r��ॳ�ts��j͌��ĝTӴ)�C�T�G e��F��]�����NǢq(�����#h�g��\@Ȯ6�UK����Y:���k� h�1����f ���$P��*@�u0N	89M m9��T՝ĺ#m��J��G3t�ma�9��jF٥m�X����J��᳧���z�qX�l#i��}H�;u7f(��Q0�0�;��B��(8w�O�����9\ұ�X��E�[r)5r}K��xح�l�9dBv�G�$9�`G�E��ܧVK��-�����\���+sV���*;�3 �$�'�Z3A��Z�t���SOԱ�p�e�rֱ���{��vu*�Fː��/�_��������0;��$&=����`^���So׮2��ۺ Y�R����ٍ��Px�]�gFt^ ��B�E�,��uh��΁c�0�nheOͼ���˹��Д�����r�-�H�.�V!=,�&kVrs-�-����k4#��
�k��b�B��v�U�:��9.NC(����������d��UY��~I~�N������x����K[Oe�>&)@�&�9�[�dw_�ۗ��Y�N]��P��9��(���ך�1OyjF���(�]`K�dvۣ]�(�B�Qǲi����|�O2IM��RY9N;�����u�s�����&��X��1*��0�oAb�Vp�� `*�1�9�!X3\�k �.Ȣ����ɶguy��Չ c.>j��*rѣp�;f�,�s�Ub��d����WD��|6y�"����C��Z334�!�P$,Z���|���������ںb$��J��q��֝H�bl<9�-օ�0e�nD�q���:�~]��e�W�u�h<�*�ME�_�.�;�2�ms������R8��sAZ��N�&i��/jzS	��){�$C�d!{��	�ΘQČ3D"���B%"��й�d�������z��:�$k,���<���EQj�L�g����>����g�|����"R\A���jI��U�z�>h���{UY�7"n�؂Ό���0��A�A�c�ؐ�Pw,0�l�&�dx��_���������&����`?��=n(�a:��j::�.�ә\�cp�Jf]�xS��M:�s�� O0\-ז�	���I�c� ��]0�ݬ��w�O`�1J�Fj��>��y����'��@�x���H�a�㯝sVB{;�5���M$�dj�UȎK���@K##�]aK���N	�
����,H�[��=
��w�c�i��5��u��F���*���<�� �	����+:�
^V�\�E�ҷ�d�g,h5�N��3>N���y�˟�`wF!D��r ���s����m�E�m�}�~x�������@�}����Lk�����˛��ɥ����9�L?��&=s������=�%fPK�(d�� �3�u���_��NxW��YAy1g_�����̲E7��_��$�Ѳ����߿�B0JaKk�6\UMW���G��h��`�ǃݲ�Z� �~����A3̔�~~�y�J�,���:<��B��e(���
�o~��|x��#�н��� ���`ǿ*�C���ƻU��^�l��A�,��8�'�K��j���<�(�'���� �ד��GlL�]��!K8��@�N�T�2٠��v1fkG���A޽}GZlg�2Sy�p�S]>� ��ZM�֔l�_ ��b~��d?GM����a�8k�WӯӶ���i�6d{0��d���K@�M�]�s�]��FDP*��&��ڠ��t�QՔ���gQ税�m´�lN�	�ˑ�l�ltodqc=Yz'�٦e`�,�{���������V����X�Fl�$�3���k��n#��M�+��WT���w��^	V��2@YȲIQl�NN2XW�k�2���U�6��H3�,�1�� ��I�h�3�\zB#3�>\H5��iZ�����N���u�\�`�l'�^� 3����Ȉ%���M뭮��pǤ��v�5�E��-Y��(U��n�� ��T5�<�W=������,)U8V�z��"��+�wэ��?�@��ح>���(�H��9+zX4�Ш���^��2��j�w%�0^V�� ��%ʜgS���4]Wc37Z��
$<���Z�} pj�Lm]��)��g»h� �1��|����YIWͤFIi���'���E�@�7�|#O�_�\C1����+��	ޑ�K�?(D�0�ۯLY���9v�rƨ?�Nj��1���g���P]�Ì�r����0���3s�;2/�%6	����Y0'�J�eÃw2DG���D���ӥ\_]��YԥkU�M/�Y����F���� &�\3��Z�C�VZlU�FN�~s{ˠ�3�T�8�ҹ���q{{J��"�S�m��xi3zR�zƟ�L���n/�s��]l��`=솔���d����d)��/������V��������$��u�Zm����i�*C���������|<�vG�@����x�\���XW|Os�hձ�d�@z��ta`���M~���"�d� pb筓�zl��>��<1�f�Lğ�/�$�*N�bݦ׭�גՒ�R���>Pb�$�_�\ɇO�^����1Y|W�������4hoR�~���?e�5v@s�:#���j�3d�"��S�H���jx�Uz헴&��+�Nr	�@i)(����%ƽ�'��|d� ��:p��Txܬ�pB�sT-��> SA�1ӓ�.h��N;j����)%�s&*���m�Z�ЭXd`d��vď��]O9�'z!���C��Ϟ��a��d�P��;��BPK�ܑU�*�_f���YS=o�6�h���MS��M-/�8x�@��~�r��C�5I�L�����z���Z�/F��#xi�d^����U�����;�t���J�}�7H�Sn�Q05J�yd�HM�HFD�dՈ=Р��Z
��N�v�lu����hxy�t=#a��o��ܸQ���ɤ�e�βnxOD" �$Py���ڈ�v_��d �l�"��{;{Lǿ�p.��&ۚ.��䘀�Hi!Wh2MTsQ#2��TA<s\��S⣕Uۨ��ps��~iA�x��gd�:Y�P�s*+j��&Q�ٵ�W�a0���~��h��c�a ��S�d�������xM&�JϺ��K%WO�fO9v�0-b�5p:(G�4�#�J�F�g�+:Bk��,�8R����짂CE�9l�m	G�����˓As4A��f�2�Tٚ�r �<�u�yy�2{�K�����d�9������h쏢a
-�	��	�r�V�3�0� ��� �4 �s����!!�?,����>JN�:P�m
��SQkji�L�qe���0� ��(��1�;W^��$��TY/,�UX�,�EFmJ�75��,B����2��������7�t�����t�y*V¾�/	��#3䋺�|&.�+�_�������ݳǬ��J��ã�|^�")u|�_�hP#a�Dj��B��`��`c� >
�o�:�Wp��o���;����|�����L^��Z�=}l��g�����)A�vI���� �r�s�내w����V�Ae�A������X5T~����g���Lf#�N�S��O�?ɇ�o)�2���|Gv�;l��pl�Ec�>s�rJ�G��;(��Շc��t$Ͽ\������ ��yd��wƟ���2����ӵ��-�����e����ny��(�$�XV*�^�� �+�ۃ�٢������h�D�G9�s�����J����� ϥd�j��������2N�� )*�=xP*�#�%щ�Vj�3�����w}�$T����Z�$���Z��Ҹ����F����1�l��]���C�n���M_B�m	C٥�ڕD� �Y�J� �Q:`�#�Ҕ��Uu҄R3^n]2љ��З9�3(W>��?��"Tx��hs��2�TxQ;4#�lϬY&K��K,�U�՗O�=;�Rq�,EY4�r����g������b������&��fW��25�ONN�q���;� iT�L��V���4tEΠ����jy�!�d�F�XBc2J����Z7.\�te�L�Zc}����G�)���f���S ��Dg�R�	 �LN�ȣGG��h�_�F��������ƨ�YHnu�=e6��hk�R�в]#ZB�J�5�Z���Q���;�h��0�E�=��b�ved�2�ۀ$ɻE�a	lN���@��`�]\����3.A{9ʇzتoS�̹)�@���ģ�=�;F>���]�]	����` x����@ 0�����aFb�%��!UU2L���r��Dg-�Ć�d�(��?v~��%�p$;�i����r@~��o�x�3i�6���(�� X�)�,4�b�1�� ������ŴL� I�&�5�����*#>_�̦�e��Ƽo6�.a�f<�(ڈ]Y�[z��VY����4�_�]�j�[�ﴖnM�Y�by�7\س/�2ng��4ki�@�\�9��7�[<�b�?x i7q�P���_9B���Rv��d���]���A����R'jW!!�����Y*�`9<k����7w��m4�'$%:��QmA��Aw�QAQ4T=:9H6{_���+�t�_ɇw���W��B� 6�J_	����$� ꁀ�i�����P�& ������Z>|��
'HD���;T�t
H�Z$ۀ!�u�9�YA|\'� �K��6�^��?�ȑL�)�^�xDr�tυ���y��~&Z)��]j �͇y���U��8�� �gK����bX�9s��_Yȿ��?��=|t�	��XSRtnóQ�ն�V� ����B�]���\ld3VkU伦�m��H��ᨒo0�ƛB�v��=�Qz��w_uE�sM�x˞����:�
���HQ�� ZW(�9���q�Om��d��H�!#�3�t�PWN4��c�������h�'��U	�:i�_٭��1bb.Y#l��F	?jr���/�7��.�u#z��$EA�K1�4c���/^XgM+��6�͵tR�dbb`��K =o �~��VT����O*��(��2R��`mooo���R��q��:=m� �A�8.F�Fii�����:?�����W/�o�@��N�chߠtِ�i� (k��7�d�Jf�Z��Բ�*r���a��L��u��&��d��T;�,�gQ�����D�H=�b�R�c�p�	čg��W�O�:�;���@�:���M��Bg2*."lJ>*��D�֚B�c;���FG'�W�Lkm�S�I���l]XCAv��-W���D�J&�@]鼰̵��֞��8�����e�7�,0D��%=�gC�)�;�4
*��s�Aͮ�L;�T1^�O8����)�����ic��L��Ѭ=�Dg`�c��$x�ʚݵ�Y*�#f��ǡ��������m�/���B�췺���AfS�P?��#�(^��,�f�43�,)���6���Y����'�K��:om��k���5���������0_*��e���Z�g9��N:寱�j��J�_y+��/�B�X:?~�P�J�L�R�~]~ 7��s�LW��<<g�_ǼҎs�R�����W���yA}Kۋ,�c���l6NA�|��c��F�:W�,n8�}������ʣ���t��rqq�%�tQ�jj����;��0��n�kj��Z��ސ��OA-|ƙ!����X�~���l@�b��#��F��om�	���0=�%\(�u+�zA�ٛ%���f��s�=K�Č�a%���XIir���`��m�kl��r"���g����-D���\�yӳ�
xi�Z�2BG�$yZ���X�Hl���.ֱ�ֵJ�T:"E��n�q�V����eZ�5�?:�m XK�]9t\�=���
�l<2 3SS8@��B�79�/fܰ���ck�H�wSjzCpș,�����"��c��y 1���P�!��Sߚ�ˉ}v�:�?��hNչA&���ԙw4�Q�B,�4��i���ײ�, 8X�sdF�Z1���S��� �jw!�+S(	��ʣ�U��-�]��͂�'}MdD-�	�XCԒ��J�م�H�7T8>==�V���n~>�����;��m\u�Qci¾�M댁�ON�R�w����a�U� ����h���d�@������ťԏ�す �[.��K�Kk���$�u颜�FtҰ�CKN!�o���8�*v���m㒹S�a�����p�F���������p�jT'��z�)�l�^�3�}��:��k���� �\��H�/r1���c��1�P�.x�'߻S�Mޝv��$��F�ʗ�6�~1((m�3u!�ڷkv`�vN��R��Ā��j�F�ԄɈ���ɳK�-:�JǏ�;^���k[;��Iݴ�&��o�vƩb^Sk�e�\���6�6P5tm:�3��W��*Z����~��������C�{A�m6�4���7q���gv�)� ��
�jô�o�f�7���3���u����ڐSXG'�3x>-��T��B����neЎr� ����=�ޒM[���3��f���_d?ټ"hg�z�o���mU���Tnnnigʲ췯]S���z�	�rAↂ�"o���Z��r֡( GS ?����U]8ם��}��,�Yu΁�˅R/T����WCF}���n������hՉ�(9�>���ѯ����?�U�hϲ��.Ĭ'��i�q�ZR��'���q+9�Q3��ߓ�Du�MkQÎ�.sh�k��+M���m�܄WH"�B<�a^�V��������{�s{�e��_�{�X~^%��^��*c�͜�`�7;wBɫχ��
���uT(=�k�HG%�Xd<�҆�Agi��[d�6h��H�u��ɡ��{��H1 �ϻJ��J��Gy>�`6~`�g�%HD����!�T�1S����Wa]�t���jךw��6�S���n���� #7Y��0�΍E[h�<(�������M���2������û����]|��s�*�	�%�s�Y��IMҁtt(�\g�a���с�^~��08�_?|��;��
�	Fa_���8���K�!b�P�O� ��_~!0�� %����[T��!x�&O��eWdg{�f,=��Gr�7���D�f�L���:X/o��U�0�{�_W�N��5�̅f��9�5,66 ���i�� �mV��J��cYt�B�c�Yk�k8� ��J��A��넝����g(�&�T�<���a(C>�H�k���`�`	Q�oF�4��Etax��� 5R�E�Q7�;f��S^��Q,�y�r�䌖�{�D�B�{Vë��?G����й�e`T��r0��U�𱔦r8ȇk
"��4ѐy�Z�z�N�Q�B��Du>.��wJv��h�}]�s�!��U��j73�H�p�Ȑؐ_��h�Ơ���̦!��ۧ�h�$�u��uj�e�+�.� ���Y�O��0������3�E	u\\�%�!jyV5�����gS��U�>R[�h�1(�����{V<� ��9��U5��M.R��^�R~v�r(f��-;���\��s@;��7O�e�2ҹ�Ԍ��d�����?��O���Z0�D0甆\�B0 {���ŭ\\]rtYU�*2#�U�<Uf!�Iv6�� ��PZH!P��ٓO���_��Uy��{���ڎPɇ�ľ��a�T"v  P@�9e�� �J 3k���i��_3�1�_f��B�]�]��ݞhNϦ�6]��m���)�2�9Ө��^��Ti)s��2鬢)�f%F+��Oeyߺuh� r-I`�ڽ�-���2W=�ɳ�2,��nFy�s(^���_����*M︣��h�ؽ	>łb�..؊i0̀U�ڻ�ט�#��@Z�v�"�[����uS�;��lv���r��j����`�{4ڃ�����?�%V'�Y��hܢr�j�(�cu؈� ����J����:=��'�s��}����U%5�����A�!�C���e�	��u��[���K��,��n�D�b����}Fo���̘�)��M�5�ȓGG����xq8�e�eխ�Nȣ�=�v�.2�.�=�A<VD��g�2�N�ۗ/�8�}:v�[�x},߾xFg���.�S��G5���9߽|.�~�þ�wY�P�Vˇ�C@ ��vp4U�⺝��[ ���e� L�5�Qb�B۶c3%<[�/�t��h�d�~o ��#r���gD�Bi۱�5��9���G8���Ur��X���;��% �r���\�҂��g��նjl�Q�W�u�e�7�WZqƱZJ�lL�@1��ޘh�'j��Y�"�cԄ��[7�6��X����?�-.�'2х�E���u�8�O�k����_��ZZWtK��'����2��/��=]+�0�
 l�����4�> ��k��>��y0�'.��,��U�ky���e����δ�l(?#�B�W���I�0���<G�D���?��$(<d(�"�*?���3��J5�*Hz�ژh�;�W,��Er�e� '�]�*w�L �
Yc�ձu.�~qus'�>a7$��s4f	�=�yB��q~y����k�;�Z����$��_���s���v$E�h�oBڨ����5���W3ٚ�)�Tҡ����i���H��}�=zt�/ ��f�gEyo�J׍�O�7�3�T�N���R�E�JA�a�wȷ`���ҿ�a7-�a{��X�ة���=�}칀b3?�����G�9�h>���@&i��O�kB�g9�p�	;�/���~���D�x��+V�-ə�|�7|�L�t���(z�4�7�=��o� O��]P.{��e¸�C��O��(*m�F;�Q�b�V1�����:+@xcM�2c�Ng�=*��$�D,e}E�c:�-Hg�Ʊ�wr��:��H,�7�Q�tU����xas��4P�����H���Yp�����G��}�~~׿FQ�E�7�����@@T�s�lBɟ�@?a6�7S��_�w����u�<h����ad���8:B��N�t*�ܮW/_���(��∭�s��?Ju/��9a���4*��(���pخttц�v��*�
��{c��T��3 �=y,/_~+��	��G,�\k9aI�\+6|����� 3���/72�҆�u�յi��2OZW����e�v�b /��JNFٳkt����:A�<�L�����F�le\�V;�$�:]pN�Аho��#�H� DTl���a�cZ�U2b���i�Э����  �X��y�]D���)�P�׍)��_�Kd	�0��,�{��Y��3I���Y�� �]�Y��0���3���x����NY�-�u�h��cۻ�ա�̞�7ߔ��m�.�������~Q��q/��9��:�q�����_�o�%N+� ���C��KS2 �����y�F�%٥@u��k�Q[)���0�j�GA\Pڠe�����b�5m��DeLXUM&d�{��C)��n�h��Y*�z����G�j�L" ����T)Nc���0��l���ƚ��dM�@o&6��G��?�Q5��?Y�)(۰�#sQn%J� P��%�o�q����i����˅�Cۥ�nI�����<}��`m���s�tת?��Xn��y���v���c���&�Mˬ��*}�&Q D� Mh�ٛOe'�
��XF�B9�m�`��W�t:�_�z���N<�r!7�az���i���!���cN	��b^ea��j�h ���+��w+y�}����z�]������9= �&P+8/U��XOH�|��lSuyO1h"b�/�>2C:I��X���H�wJ�!ۗ�ʈʭ�u�w�~��k3x��f?q�E���j���=������� �v�J+�k0])����)����u�$7Y���gVW���	5(�PV�yE�~vc����g�����2
h�i��t[g�� ���	9�CC��
�B��<D3�9@U+�?-�jG>�ƷH7_4uB K��� h���%��'�8�]�)~y�C�,׭����f����wr�@	�,������'O�*�>I�z\�uq���'g6Q�=<;%8 �����c:���9�RR��~%O/do�<E�[**��g���GG�uJ�$�A\�v2&�9���B�88;����9=�J�yN#�n�#EnE���h���c��������kJ��)��]/侴
P�R�Ò�YN8�8 B�ʈe�������fِ׀��Ȩj���0C�l�Z�o5��5�e�L���fA���������(��h5��~Aw�w=�k�����St�m41��x	:���r�s|\wg���iϔi�'��<J����n]Į��˕֧ I���)���D��0}&�S���Dtn�3�<3(AA#��KUfB�g[\H?S�זچl��._��zeg��\R�e\AL�SV��lA22y�N!�M�V���3��Zf�A'�TM�מ_��	5�Q������@_�mԍ�ou,	�w'#-+s������Q-Q��N5�1�S]J�@�Ԝ�hD ����Ip7��Ŝ]�:k|qi!vЦ�3>`! k,�������/r��yV����n�0�'��r��p�me՘�tK������~6�D  d6.�yA���O��}ͼ#@M���F��vl�uE;quM!�KV+N�؞���kۙM�,؁��<�{�N7�z��|v-?^ʗ�[
�:��u
���^�M�'F�t�F�E�,��F���	<��]'��L׾�T$�k'�ڐ"=���u��EZ�5�8h��Nk�\ic�W#���Y��DEN���ZZ�Z�����Xo?z_쩯�O=�h�����/���o^3�'<�������F��si� LB^Mp��T~H�D(Q:��)�-����.g@�����D{w�XKC�Du^�0����ː�<��������%*���w��ܢ�2d�U�M��2�i�>�1�Tc,n~8_=�Ч7���|��(J���b�a���X�iV���qw�w���G�q]k��P2?�x 1NX�uw$�T��nu���SD�5}t�,ם\�,�z��`�
�,��Z%j"k�����}S�0̶�t @���� qU|�0B����]'c�c��/Rt�o?����5���4�+'��A�8�8\���7����T�X�� :;������y�᳜���tP��%(6*��n��
L(@�c���VO���3��hR3#��&��"1��Z(賬X3
E�h3�D�^��h5n}DW�\ \�
�)�����C�ԑ���KE*H��J���R;�`���d�7��fPp�ˎݲ�B���*�m��!��{�֌Qi�3��Ap� �۴2�͈�s"E��%�.R�H���qw��ﺦް�4(��F���jÆe�Iv��n�.6鿷��U:�\�C�r$SU�.Ֆ,��ݥ�ߏ���u���qUL�X�`��4�����5 �!l��koo�u�vE�����(��:��"~/牊����*��HGGYyƬ�Y�C�)�ZJ��!�� e���.˧��L��kY��W��dɞ����|!�*�u�D�u�����8J��	�����J�mR�#M�S[[}0�*��u�>p���H����e3Dl�NM8��)�X#��d	V� LADA��ٲ�I�{���Qk�4���R�y���Ãz���ѐ��ҝ�6	D,X2�Jv��Ԑlɗ�M��w�u�l��`KO�#��EV�6�\�m�|�v(�E9=��?����l_�<�������4���3c��OQaaw���F���7��ʻ�)H���Q6	"���,�߭A�����̶'YG����[ʲdf�S�f� l�k�������� +� }
I�d�nӹ;�����my#��E��W�`�2ʚ���aS2�LH�	&�T����a�8�)���g�3���rL�0U��o?������-�	���=[-bэeG��}���>��]-E|�ATOT���MD�TUa79�8b{%#�κ �iD94��h�w����߳p���p��+u�����w��Ha��^�CI2����-�:-�Vo��k�V	B�~l�D2�r~���`��w��FG��:Y��i�nWɈW��U��='�{pD� R�O�r�z������օ�@
����r��, D/8DPbFsz~ͮDL�׮0u  �Ͷ��kiT�f�V��k��ݲ���$�~N����� *ZL	*�W���|A���w�}����lϸ_�ҡ�I 
ژ���9I�m�>Dt{zv%o�}����Y���la0�TAN�Dn�C��B�-4x�ؼJFb���NPP?j6I�)9��_K}�1�}=1�:����r��h�5!C
 �^�X���,�p��V2�h%G�9GAmM��:���g��!.LY��<vi��^�1V,붊Ţ��ƙ �"�3 �8L�S1U�(��)J4�����}��s���m��>���h,u�!a�f�ikx0�,=!.'`5
3H�a����;�ҾB�C�Ud3�\&#�3)���6Ӝ���`��%y4���J�}�����eIaw ��q��B:eoo������_��������]�ur�p�:2~.z�N1�V�@A�ɢ,��eh� ׸��,9�-� 1�|U��V�t�^[�J/�/*U���ydL�ϐt�'Pj�Y��mJI@�l���i����ٞR�f;�[ ����0��f��f�G,�f}�Y���` �#�? G:�+� Z{�#n9��5��hَ^�B3�zZ��2����O��J޿�����Հ���/_(C�F
M��SCj�R.��x��v�>:�e ��V	��Ò��c�U�ư��/&Obt�Φ;DK
����D���b
˽>#�5���$[zi�*������oUiy�5:Fi«5m�6�\^߳4�!�܋
�3�l�Ӌk��Ǔ��{����uC��I�.�����nŨA`�����o�%���iM����V������W�Ǽ��3��&B}�A����mT��3�r4�Ｑ��	��`Y[�}�]����������Djo���}t���[4�J��~�g���1K���y�F,�l9'+8���ܲa�����DgA�n��
Ě:d˵��(F�m��b�T�B�FD��Å�_d������[Hu�z����70̐�E�c�7S0�巳�^s��YÇ�y���W�}5����{.��
f� Ho����,��z;En\�y�&.Z+�)i ��c�A�(��`����s���'�����' �@��	@�Ȟ^�����h�`����x��-����������My���}>���ۣ1R�҂̾j���+����O4`E��#W*b�?�G)�@����!lD������_������7�@$@�&s6K����ő�ծ���Ka��
�ޥ����5?���\���%�p�{�,MhE�KWyWq�ݔ1�\��Cd'$���05�fk-�3��nrb���ׁ<9>Jk:�a�M��T'�#ɪ�κT>Ԫߧg���֒G�E�\�w��R��g����<E��	LO�I�����v�;3���o�hWk: �f��ޢ8
~��b����IxG �Y&Rt|V�RscG(�FK�0�L��X�@�Q˿Сc���6��T��Ǽw8Yt(j��j�k�%�3������&��3Ct�y�FW���	'�R���T΅|Ŏ����_��۷����:9�0b�7��lDZi��L�g�� 7�9�n��b3������8}���(t�"�����ӕe�J�Hk`d��5�6Fs�I�5����..�����%��xm0�'���aՐ���o�ȳ�'�a��9rM�BK읍tj�3m<<G��Xf[�|�* �M�K:{{���R9r&�Ia��A��~F������:���"�'�j����2':A�L e@p�p2ٕ*:S �.�˟���r��邍E;P+�/�ү���Ԏ=��<��|!��QBe�I�`��A�|�s1���M[Ӧ]c�}+7��R(����Ħ>e�8O{|:-�s��G�[�{����X��
� a��A� �3�ί��?�"��{��$��ҵ#𸽾!J��Ǩ#TR*���H���+5 ��?�>���F�(�귧c^�G � ����s���BT� ���U��;W���q�qzZMcr��S]Nv�o��7 E����(NI
YO d?�Kk_��x��a}Ƌ�ϧ%�,`�#��2�޺>1�}J��Xoة���߫ ��>��ˍ}�uA�?�T���`��ۓ{ 6̂I>�g�
y �����g�/F4R��?KC*h�E���C聚�����w�s�]� M#�u_˛���{�S8�8<D�0(���?�V&��z�#VD�����tz��ѝ�,�%��W�9�u���E�.Rt�;�f�O�����w�D�-[�m���b#>�ɛ��ɠ޲�A�k�G� ��@
M��m{pJ��oҡG��+���./6�0��`�& ������[Fw�w,�N�a��V� �G��U���~��i�!�Cڹחg�� )��bĎ,�)		�F �u���A��Ú���9�a���TG�Az���\�ʫ���,��G�a��n�4Ƒq`^hw�F��A�-t:�����e� �z���Z�鈘�? k�mU��d_?9����^�$�G��> 
��7�ᚖ��*�Ɂ���@p^�%ú��%�wY��Fi0�x�2R���*�}�D��PgD��蔛�?�L�V6�.�t���)k��P~�Uӳ���������U�I�ΒGnV��	 ń���h<Mk�^8S8�p>ggg�.9�_���v(?
��r�J���clY΄���BP�&�³����ҽb�����ﾑW/��7O%�8����3��]ړԻ��ܵ���/'�t|���J���{�nqO�l�g[8��TRƅ������W���sy��I%[�^*�`�0�"�a�nx�`cHj���gn��95��ͽ���:=74���\Ed\�̚l����R"�Ȱ��^�7)0\��$X�.m9a�&�.�N:�J��gЩp�� �ڭ9b��a��}���ܭ�kn�, VP�����b]~k�H0?cc����o5����{�C�s�w��iޮ�Cd:�HE@� �U�_R�ى@@��u�a6����R������
ϧ�3Mg���`��l�&	6<h���?�t}�� i��m�,Ȯ Spz8v���\��N~��~U�]�g�����yY׸�4S8n�=lM�2Tr�EH��U�C�ςeΕ������g���Y��.j�̇�S������J����17��Nr2������w�Y5f�z#���44�X��VU��l<���������x9og -��� ���d�*8��"mO]�"���C���=���#��Z���t���w`�~v<�QFj]#7�Կ��h5E�ӊ�ג�m��Β�&E�����̫V5���M�R��:�����E��uZ�O�)2N�	�OatAz��fy����	����3�����0d��F��W2�]2���N���C�n�t�C����oߝ&�u-;�P�Y�(s�$�a.PY�@���%'�L��g�3�X7�2W�7t6���WZ���"m��/��|z�����r�(
\����9 )8�ؓ��,3a�l�:� �l��P��!r,0ܶa����O�=�����<=�.,&��~
�v��i�i�v�r�K�6kY�i)g���>�ۨ��- �W�:ڙ�w�<�?���ͳ'x��t����N��� ��r�j�_i:w�M�����i�l�s}��1�Ñ��
�z7�(��D��UeXS�^B�'.��i�1et�B�&�����h�Ϛ��i� ����M{�~}M�FJ@w:#�K���"�����gٞ?!eht}�+Q�l	����)?��_��G� a,֓�ͦ�@��x��� ������0�1���tm��s�S�M���1:�dw,ӴO:���4cF���%����:�*�S/�^�x�@`'9�1A������$�������ȶ�9i�������( C�&��Q~T�s�D�bQ:����n�<'��/��3�?}:�U
* ��9���|��[�*`��{k�E�%]P[�od}��H���b鶍y�i���pu�8� ��>þ雪�;�C�#Ga�Ԧ��U�QH�� �d�7P0��`�ѐ#�J�X&����l:g�j������Z���r�4o~Vi=��\C)��B�����,L��(�w
�1�ràE�2]o���״xNȶ!Ajj�},���ؐ�kۛ:eD�@?���)��3@*q��7�X�6� ��6n�I�/��:���� ��]�B�m��ܑ��^A�}z�Ne���=h_��q�(��|���U鉩�Q�R��A3���/4���ʑ�{��5]�q.xy��k(#_�0/w�5[z�dËv�e�U�qJ�i�5�k_c��{`٧(�7��덿}A��aC��&�l ����j%�7���6(@��zy�,Q�cq`8�.F�Ҭ���f1w����x�|,��;�C*��dh�͂F dh0�{bܯ���~������%3 a��H6.t`h���q3{�lR�iW��ɨ�Kf��� �(S�5�싒���h	�R]���ł%�M�j�Z���mh�b��'"Q
�,��"�d,�vH23
])d�0�>p�8�+�n��<���������=V�R��P��&#�5ٖ�ޖ<=>�ׯ^���ȋ�XwӚԫֆ?�w����y�<^�&F���`�3Bp֬�q@jNg&��Y!
ƫ���G���@�A�(�(�;jW���*��H��Nu�$�S���FL�W���\3G� ��W�*U�ZY{��\��~Ng��"�`6I�PXjZ���ڨʂ��P�d9������-��-(d�>|�(�W:/o��������K�K�9��ɓ}_t|�r��a*\T_|�t������y��m:+�_�M�Ni���eD�dX#��|� �x�;��)�Lv����������zkf,6�3U!�5Ǚu�[N`�x���	�cK Ҝ�)��ξ�%�z��)�����V�3��Z�w�/a����L>m��J wK�\��0�����Ay�a �b��
KZ�9�F&��:kM3�]p˦#�W�3�,��΀M�1ܥ�S�3�y�??jMZ3����^%i�5��l4�:�3�h�Ɯekw�5XTY����o� {A�����&��]�b (6�
�2�c���d�Ag�@o��]��܌M� F�^:�[sǌ���~� :_\k��T}�@�^)x]-T���t�j��f]�܏

ʂC�H�̄���$'�� /6�,C�w�ͱ%�R;[w���:�z�J�M�,p�صN��˵v��q��Ri.���KqN�޻w�η���g�]��kY�������� �庌�<I�I�!��;�ۋ�^`��-��Y)��X�]�TL7��A^O=������7�{Ȁ�_��w��8	�ߧn�W���s�rY�=��Ix.�-Xo�٧:0}C���7�ע��r@��]��";���h�5m�qT�";��
:�S��PH7'G]G�N:<3�X��K'c�]I�4�d� q��I�Iè�����x��Ҿ�TlW���׌�Ӂ�[�(�����3v�;���>H{�)#�����`c�:�q����(c����	�R�{���)߲��z����v��=Xt�Ԥ&Z��GB ��uwR&�XMS$K��)#/ �v�Y�N�i�"�m`W2X(�� �Ff�ģ�}������|��D�v8�N� �����S�	 �Z�X"�G�Z5�h+y��@Q�S5�@2����Pg-�*]�=��M ��w�22�9����?�LgpZƸ�9u�Ո���}���5�I�J���ÅU �Er(;�~�RY��l���^�L%�0�1o�wXi�X��� �����g��@��?E��Ņ\^ ����N��R!��^\�ɿ�뿤�\��o�L�&�'����!@X2��9�7���.�Y@�7�ь�'�����c+�qm@9�ƣdI.�K�Y� ��u�zAUw�~B� xy}s���{�@<�^`2�L�)��P�_�&H�]A� �F�6�~��dk����E%�B>�9�]i�~N�ho>�ˎ�쥳 � �p�J�^` `ڝo'��X�?.�^}�A�+=h�v��P���J�v�e�;G����,��`!�=�E݆�Eh��A	��Rmr�,�s�ZӴcp+��]��>�����bW䈲rVn/����i{�a�P:���c�q��Q��k�i����D�lM
H�7����p��adܻ���ٝ 'w<�B�����Kv�c��Ǝ�66�]���4b@���ӧ��O,衹��˕�{���
���)��S�l����92X3��g\�$%� M�^������P�dT��f��F��_�`��v������=$���Ϡ���K���a�'�o�O�C���+�+b|ؘXE���Ė�/�Zt�y.��Hx������b���u��ړ�W�ǩ�1��P`-~��^������0�����B��=���DV+}JT#��Zk�˸��� �/F�	�t����}
���k�\�-՟�@��L�I����N;-`���'�,�u9|>)Zxmը~;�t��(h��R��G*��ƍ��`4��s*A`T�VcM�_��$±Uc8��>MGm=�L�s�Tb9�_���a�Y����jI�g��LI# �3�u�������?�3�4$gI�3!FQFJ�T��٣#y��Ic;����H�W���{vqEqHl��@H  ����DY#��'�^��������V̠���u�\%0�)���w�I���Y��Rm.�{v����9��j��wtٝ�"9�翞����^��D��Q��1����bE+���U�s�M�f�Vx�X���r��I�R�D��M���g���q�B��g��ֱ���X�7a`�g�`����씜�u�X'$P�̬K�6a�$(���l��L�����sH=%/�zb]�`PEm�)h�]^]ɛw���/o��/	^� LT�B�N�G�%Y4P,�[�*%$:���J}-�ՃK��~p\6Wr���Y(�C�} 6��!ɀi>B�{=��C����3��+4���^��1�V��k ���x�+I�&��̖�񡞛V�҆��6h�S���.Ȼ�������>^A�f`���0��v��R+��`�֌AQl`�vѰ$�g,6��ݩN��lvc��st2�Xv����XXQ��zyF��"jr� 0��QBl!�*=��%:��������<}����>�pDQ�_�ߦ3���[�����8e�MOV��c5�_D;�~/�L���:Ψ#5u�R��:�ӧV8�r��,1� �����{��8⡟�\A\�1���5��Q{���\�W|�kW$��8�VG<�&���.(p�H�ZS��J�Ik������z�Q�py���L�tp�Or*�7�V)��;�n,-�e�ˇ��}QT��!/�_�\�LD��
�8$
��eih�JC��f h��8��
�PV�V���#M���D��F��*��� �9K}c��wT/v"3<J�T�ǐ�Έ����H0��185Bp�nJNfǨ(�:�:�`YdgwW�f3�M�i�M��Y7
�a�*s ��űZ�+N t;�)�e���kYVthuk���� }M�f+����ۤJ}��~.�
�'���]N(03`J�Q��b��՛i�,"�"���;sF��\{�H���Z>�(��_R���"��h�w���4�'͂Yy��#�Yk)�৬Y���ܩ1/-k�L�����O ~��ǭu|�2֯5n&��
B��rDy�����?�,��ݩ<�49׻t=K�+�D��$D�ǜ�0���4���uϠ��~���*ك5��-�����Kr�B���Q���GT�Ǵ��݆2w��P.C$�,��	�*�:���r'	?Jmk?>9� lr� Հ�&� Zր"��'������)��X�1ҡi�J�Ť�w BU��QQ+ ��O����7o�/g�	�-8��M�^1�:�N�h�����}�A��Oi���N��*��B�+m� �f�c�l;�1`����$�Dt����I��8�+8=g+�or3֢d�Wx�[+���ӧٞ��뻵<B�W�,Q��@�>�����%���]���b�Bе�*u��OiPK\2���E=�9�U��nCJ�E��;��F4di�DT���wf�K��\�j����v�nT,`nh5����sϚL΅���Z��T��T�b��J`�V�/�_�L�X+f_��x:��T.,yYmK{�,W|�����,6��8/JA��6|ȏ�7O�ʓd0�@v�����=;KA���{�5�dK�%�	��h%I\x��{ ��s�t�)�o�Kچ���d2e�ǭ@���mT.cgv�v�+_2�U�i__�l����w2\�?�^~_�B~o��~Ʈ�ZI�E�X~O˂��%�/`���R'2�2dρ��y�5 ��!���7��/Z&�������O��i�B�}��	4;,��!o['���&B�l�;J΄��@�;3����~�Z�q�9R]#%|�n��5b�G�Qo+J"e�q<Ճ	QD�Z�}D�/�M��H�LB:H��}�J;;��"m�D���w�Si"xŬބ.���(�����S���X�'�8k��
ȰE�L����t���LAn��/��U�F�P�/t�(�X9�@a3G��C;�	=��T��H5��(/�������Y9�SA�Y����m9��&��3��d����^�嗿ɻ�ry�`t|�"S ��1��8��f`�2xp�Ś@�6�$�(�>h��	�����ZM�pլ�Δ�՘��l2(��:b�"��
���?�T�5O ��D�K��׶�=���O�P�knN 8�L�]5�N^����+��b)��c�C����4̞NF
��	�A<�q�	IT�a^���YV-4s�3�d/	�b̤"��'35�Υ�A�0��kNNN��n��&3\�,K� �7:��ׇl�E�~^`V���͆ �˗3m&H_?�rM �Pj"R9^	�Ƞ��@���O�뻏9�9�T7�~����y�q���f۩�:��Ȟ(8a9�6/�*̊���	,�Fˇ����Gьs�<������#qU}�A����������t(3ϭ�#��nGC�C,���Y]���W� L�̚��6��' �Sk�7��Z�݊��~M&�C���D��2�.�� �/p���Bѿ
��� �5ղ�;�<���*{�u��ӛӬܚ�oO�aA�U�l�WP��N��2_�\/}���3��00���K�3�)^<�o�y*���,G��TN'&�{�#O����=W(KBX��4G<�v�8��;�gE|&k�|M�LQg%��$�W]���#����[����}�=�+<�%^X���`$󥆿��?;g�2�+�zR�����hB����Tk-�i����d����XzM���m������0X����ɀ��]�|��,J��+�
��kƱ?���~WS�j���]G~��'"|�{�:{���;oyڻ	F�?Rula�>C7
�۬���Z�-�2^i#�B-e�=v�]|�Q�����i��y�.��Q.+Fu�i��п��Y\�R��t�����K��i���vm����8$ԋ���/��i �ց)�Qe�	6K��
7	�Zfjɋې�Qc�&���$Ԩ�p��s��'�XF61"'�XHMTS�0���h�v��#F)����O� ?�z�A��a4������������%�J�3%�+�+m�WӘ��R �b�3B9��u��%�Z>֥^�߫�HS���k��28�|����H��is���$5�:;%g�\0t��P�==a�����k}��Tvw���_���_|�����7N#98ضl�IY-��i�� ʷ�Ke��r0m��@�)%����8�?�Q�O�)5R�5(uL�&���������������SѪL�v���!*�lp�0J��UE����-k�P��k�}]���U��Sx�����9&L�~���ʾ�^����lU�_�Pk��9j��b��,t�qe3!k=1[�ya�NI�.���28f�����im���G`��@@ea\:�>��N�Q�#�l�'A(:EK՝=D�L��6�5��6�p�Q
�0G�R4/�n�w�M5�7�3��/���\���ח��W�s���%śWr�����"��Ƞ{565"���j��k��m ����P6��#�"�o���&�(r')�N:,܄l��>�E����I*�����\;��cf���#�tu6���z!�i���p���߿��~�^~��<{r"[[c��@i5*�{27�~��w������d���BC9Q
Bg\-�僙$())j�A|�Ih-ߢ"�!���&`��U�X:��u�/!�j���a@�7)3X�����i���hƳ3!c
���1��=(���Z��+U�E���R묚U5͛ml�q-<�em��
_���\~�������HON��>O�:�5y�	A�إ 
G�����5C�?X���2iu�q�����d�FI��cw{"����Va%S�5F@,���nW.//��o���NӒ�E�N�l,�����)�_U��5��jF�k�$U���:&إ$w��ƚEg�*�:�X*�ܔ�5*&����ۈkX�]^)��a��l�B����n����e�%�1�@��ꕣ�]#�I�T ��`xX�f��l�G �	�S��H�cEH؍��%[��pG~������jV���P���ЉBB�(�#��i�����щK$�:rm��s%π�o�dR7"٦�.;��c��x��bx�"��Y��\�Z�(N'�1[;��¬�u�\�,
#�L�`����O���oؙ{{I��G�=9"Y{b�M�T�B�,��l�mv�f�Y�I��g��9k+�0;��EK^�Pk�O�F�E�[S�.zm���@y��z�<ϫ	׭���r�iU�3A^��lIfKf�ʰK!�Ʃ:��(�P�# �|��,�#0R��G�6�ƚ$��6�Z�� ��m1(�QI�V>�v��H��q�!�_�^u�.�Y0�E����tֱh��=��~�oĲ`��c�mEڏ.���UY�G�3Lb�U�R~$З:kgA���G� |q�s\-4�6w?8�K�Ҟ�x��A��f� �l�c�o����C�@��B���t��	K�
�Zq�X��-T9�Y�"�y�"2c�@4�*L�V݈�� �c��ڼK��޳_�E��'|N��V&�k��Ùg��&*D{�N\ҢM놌��ޡ�x�T~��y��<~|";;s�4uz��V�nࣣ#�15����~��T.�n�*L%A�jpu��6 0�gg����9�3n/��`"!P�vj�����qm��rv|��,�N@��#Dze��_���S�_1�c<���	���)����}E�0̆���W��>aޗ��J\�t>_G��h�v�v�)>?`�G�;������6u?
S�τ�����<�ĥE�C��b��0��W+%k
�d���Lk������,�w��y\��	�,8�$�J!�������S�D�آ#�pȊ��?ȿ���W������B��e.�˱���@lP��uN�HޥҨ�dj�k���1Q0�a�k��1��h��^�Q�P��oR'�16ɑ�@C2�:��J���7�1�đ~��&��T7~�6��k^h{Yf�0�i�	Z����;�|y��,:�	fϝ�-�[ ��4dT*G���ه%} s�2�$�Ҁ�����<E���3�?�N@eƶr�� _sљW�G�eAv-�I�L붷M�YJgg u�+F�߿��B�,��*���O���UH�\��ԋ��� `G�:��n�U����M������|���svX���(H�lQ�� xJ�0�� �Xw�s�����}��[�S><�2�(���sC�ͅ���s����^�f]ۨ��fg�t��a�d�n-)O������0��wj���l���
�f���i�>�V�p�m��xf��y[�z?kV˜󂝍k��r��i2�[��
4P1}��r��v*:��H��DW�£�g�G���o��$Ω銱W�F9�c�T�'p��Z*��R��l��<@��3;��1�jNj��}xʱٚb��6˪S-��:b������w��|F�V�W6�zI"�m�8�(���4Zd���xW�����Y��_Am*���S5 꼳���"�����^��w��Ͻ���?��'���+y���������^�6��;bXHz�`���%࿾y'>�rl��3:e���C(��
>��ekH�ؗH�h�CG[R*)���T�s����DgɆau�0c�´�iĵiCK���e�ր�q`I�������O��{y��9����t�4H^�g�E��[)X����%x,Ǐ�ɟ~���?��J��Y7����$OͲ��>g��m@#��0)�{��	`�� u�i�*�M�*�7i�~�N�i�i�3 �� J��i���L]���� |O��r
�c����ƚ�
�7�qI���H��@-�EP���5"�pb��<��I�������4g����e��?_D�+���?�y�w���G;(�q�^�p�F+�𪦢���8�Cqn�(�[����O�ӣL��ڟO���z�D^~�(9�=3��P���h2[ӂ)wv��u��\����[H\�p�=���qg�<�H��Z	�|���U�G�s�҇�B�X#68#2��d�L�TAYzdÖ+է�r��G�hZ�kf��bB���6�Þ-��Љ����|J�QF��1ERAEd��9<1����χ3Ő���+���9�Y�d�R�D����"�Ih\&�����v��F#Q���u-�����0*�8=Sh�!R�(�TQ�����K�(�D-;E����/�	�2�g��L��� �N� d%���n�ߺ��0��eSp�,L ������eآv#>J������� �TD�2u�_>S�s�1�X�� |���Z��hl�q;a>���٠3%(�ic��9�D�aY,���:/O�yk`����q�TkB�̬I���zf�9[��l��.��ʓ0��r� 5�gY��֚v}�Py�9888��''r��LJt�"#��$2�]h!F�ز��<�ҨT�wЍ�^�u��' h��$�:�a��YE:Hݵ�3;��0�f���� �t>OXAF�`#v��|nww�r{��ɲ3.�J��6U�K����K1�v���,�Z��S)q�6]�g�h)5�� X �p6Va\dt�f%M
����5Kj�����ﾑ�'P�^���Q��S Ͳ*����%�m�;�� {a<�i!m󷴧�LkL�D��y�{�ܨ��bP�®*��O$OF*w��#1��.�D��5E-Gm�*M��
2*��}���m���l�+ϟ?!��ݏ�'�u@*�v�v���%U�������3:Ok��m��(���/j6iFK����׮b�ʩ�\7���mv��~���VdE �Aۀ�h啵�s}c�O/sY5�̹��g�\�ޫ/N9R|c^}P��Lbv���B�w�������&�Ln�pK����'䷩1Zk6N�8A�n�JŅ�Z��C��(o�\��MY8M�kb"\�Y-E����w�m�ACl�����7��Gч/��L��e��f���F4��HX����.���"Uj��ښ����@��x-ϟq��zq���*�k��F�����O�c�
2�z+?��by��!��W���LR�Ά�i+(
�2�3F�O��A0�M50 J��9�q��M��#�,��HVK#�k�|�dF6��~/hW��u��g��S�%�"d+�&�*g���g��o��<��|0�&�?2	��{|�7�NJ���n�B��$��?'�p����{S��׫vb2��).�͑>�ʣG���� ��j�*��n;N@����Rr8��'����g	d�3p��_�m)��<"�����zCǿ�RF�\ȩE��A�󢍔��ݕ�/����]k�����h���� fu/�_Xz8<<L��OЁ=����l�8�R���q����q�X-��5������_~yC�0��Eռ���'e`�DyU:,<��<������\�q��y$�9���x0�૵���C ֵY�������s�@��7�G�r����T#y�&x;>~$��?�M&[�J��Vf���X
^��³�c�'��>��Vg�6K� d����ؓI
�^�!�T@ ������~�YrɎ���������w����Qr�Sf1i�Ç̒,����y�(�0bdրe��^�Mh� 5�R8Ea��x2E��Q�1V��h�3������ .�j
��m����f �B{x���^ɏ?~'����w��A� ??�Uvְ-V�9	�(��99=�(5���ly�h6CF��-�!:!��A~�9]ާEg X4�J��KoD���3:�~���u�2��%SI�}���[�ޏ8���G������oI%W�M-�oبc��-[�YoVf���3�T�V���ٓ��[
po	�����TZ�m�bIQ�S��8?4X)�&>�_B҆�!�ֲ�JU`�dZSic�F�7�S��V|�b�2UMCm�[���(�	����B��>^��mMJ�m��B�8��5�k�!�J�||,�ʄ���Dޑ�����!=���z�"��\� 	�����=��͸)�f�le�����Z����/���aݷ�J$��x9³Ö�O��W�2q�*Wzљo a����Lɋg'��`����mx����QN�)(�`��aף	ˑ�JA�p�Ttms7�"g�P��T�HG`x������qëΌa��f(�stDa���cK�|h9Au��yFUī�.;�~�i����dA����m���~�����������j�@����^~Odh�I?������t�K"��ײ\5�6_�\����u���9p ��%�31� @��ސ���,�� 	��(E�pq��#��I`�������t_p���V��Z�cm���y���R<��~�/m��}	v�.Fp��5��.�@��d=v��8V1S-=���l5S�ٞS�L�^ ���y����O  +K�DkspE�sZ���k0���S��QI���ˮ���jЍg�ԛ]���J�-K����^2�Y�+Sb?c�iӞ��1J�M�C� �ՁS&�;�"�=�L�
݂��_���ҜF�`NK0�<@�¹ lß����霥uE�
�[���^}��Ϗ�B�@�߳S,��H��j�!�x!�R�ӓCy��Yr���^����[U����h3׮����:k�/4�l^dGo�"�Xg��5��ٯ�tKu�F
�pߍ�~�$ئڨ,�叁��b����� z�A������ ���y�6U��c(�'  ��!�hk=;:b��8_[��l�y��\]�RM�[n��F{�V)� �������eA$Wl�g�]��?ֲ>�&x	�|d���9���(3��`~��J�&��|+��	��b@���;]�@���V-4r��Z�ĳ��?��CI�$I3��8���L� ��;��� w���n��{�=Z�%�����GdU���%����n�f��f���[	���>��|�-G;�ūV�taԜ�m���l��U_R�t���h��v��$��[�Yz�L7�2Z�<:�K�JU�ӹ�����i6�(_X�;%Ca�7d_��M^�k��@�V�XO�f�`ql�3V[�b���؊�
�]��B$w ��T�KՅj����6D�9�� '�i����~����^��O�r�2�X����Sh�.���c��
��2��I��o{��[��Rb�}����
�ʍr""Wj�AZAVR����;�?"}s�b�O#�¹h[wxJ=(���ݕ��O���C��?����|��_��f�I20)��SUa�y�p_�L�������4�;��,����4J�,4�]�Kd��Ǣ�i~�����?��:��
���)�1>+~���O���?ɟ���;�x� ���Q��A��%H��뿹�EGs g���^����_�o���\0 7��6@ݒiCX���T�t�2�&#I�H����N����@Q�AvN��#~��H��:Lꌲk�w95ͲI�+�TZj4���\U���En~�c����f��V���5˒^�	>X�2�������&����KF��J��J#I�XQZ�R����E��<3�f�$k��r"���"CY��ʀ�n:���a�
R�G��M�r�m����ɿ�nK�q5W��WQ�3�Hi(�w&.M��|P��rb�kft�����D&�1�?��Ȣv�[�p*GưK.0sA�y�GG�|����,�S�1�����Ջg��������������_/���M��6H{�2⾖����	�0�
�h1�8|T�&P?M�/��{ruu� 4��@"K�l�E�M���������0�2�X������O�,.�A+��%�����Y 'LހGC���"��vS"%�
#t�r�w��
���dt�PB���G�*�nyl,��[��lE��0[�z{s+���Skk���éʩt:V���3/��/�$�V�&-���M���_�\�e�C~Mop��X��~'Z�ډN<��Na���{�����W鞀k���y���C`�
W�eP��(,d}i�K�%�cm" �Y��#�5�Y��{h�|�t����Q�!Q~���Z�.�/������ւz��Z����� #�he��̿(E
\8���K�a�lh�~���ڽ)<�N�"�f.��'_�����%5���|���t،��YI�2���ajx��/�_�*Pa���uY}�b�@XJX�!G*Q����b7 H���whqH�˖WdMo¾���.3āP�Fv�I��H!~�#�Z∼?�ug��qqY��s.���`NGT爋��l�gU42��=M�b_���hu�v(��	�ˑEr��Ѭ6[M�!A��U��LQǑu̃��� �s�!�����d�ς�ԇ��w ��S���_��WҌ�tN9�`0pcvލ�gc����M�{����.Fk���&��Y�w_!_~�3��O�#^XT�n���B7���X���N ���?���S&�d���VSU�D8\肩�����(��&E�/��Ӟ��cQ%@"E|��`�}����3NuȰ:MЬ�4v��5Ƹ(a�lc�B�#p;|ˡ|�����(k0�^�)B$g�R�3X皆�*�`�e��ڵX�Ho��������������_�5�ՙ��N�뵇�G���������(;�J2���|K�z\]_+-}.�]a��(5CE�2��������5������Y��z Ӈ=(����[�Am ?�K�%B<����2��Ud}Ѕ�L8pS��Tv�v�՛ײ�����%A�C�/����|�ի�X:F���E)hH�PD�ળN^��ivZ�5g�^m��Ƶ�ٞq���on�DH��B�����y�CcHȎG����_�u������V�'3� �B���
\`��c�~0-&τ��݂�^ ��J�,���	���"�|���^
J7S� ��Zvk���S(0,F�-v��fVU^����K�ڠ)�0igg�,��p*m?��6�Dg:�Ȧ��:���A��W� &9å��Y�?�X�k�}TN#��3�&��!���JrYw6�=ޢ|AEk�i��ߪ�-�JnM��5{��+���C���9#���آ�
�̫D�P�L2���{b`�����z��`�V�a��٥Tk0nG.�;�3Q�����iH~�h��~����{=L�x��r�
ޢ]�k;@
�՞Su:NrSE����<�>Ѧ��E�;n0�����v�d�9F�=>�5�9�U��xT��HQ��V�<#��cٷ����-�q)s��1����Y��.J(F �).d�$|��_��s�Au���*� ��f�t}��f��lB��J�hɹ��C(�n@i�ʈ,���4<��I�����|���0j�����Ӆ\�5��U*`�0:]�k�M�(�R���b��kل�Ƭ�c�n��ś1y��p2�N� ��a�"��AY��	�Ȉ��u=i����I�3����O������d�v�ewF�EEW�֮6dy?K�7��k�L�}���x��^,$G���'G���]���m���ez�[�Zi�grD����l��ag�/a���v���C����fS����Q~��x{��Wʅ+��=�N>d]�Vz?� ���Ś,s�w�YW�e� u�"E���T�V،��St���Ճ8��Y��ZCJ�@ɟ��!e�������W�S����J�}����'�;��O,K��1�m������嫯�b��kDm�1��S�-�nYSaO ���\޽}'��3:��-�zd��
kb�z{����_�^�|�\Ȍ�����;���q�(�I �b�N����Z�{�횀��Q���	��l��}�RU�K�C�48��jL�~��z��]�Rn�:�<��iM��׆��t�חruq���6�P���{�� M��,l�,��K�����-YJ �k�n�B��p]�s�ڒY�>h�@Y�����p���7���������-����$���=�b�F5U���3�/D�S�sEv�3pA��/��Ǐ�X3���1�cM!3�nP����=[�u���	�aF(�����38�����7����2�g�<3�)�[�f�A���#���'��Q��X��)Qџ�2rd��2h#YiOo�茮_B�$W8
�ӳ�DP���.�(���z0 ������U�L�r����\��݋NՇ� o�1��z�(dn���E|�6��߲�n�tO�a�ikRq���L���tR�&,������b�m?}ˈ�ؼA�S���������Q���[�o�J���7\X+%��`�j���f	!�%�8�R�KU�����E�V6��~��������G^�nu(p�8����Ȩ�x!l.�6�܉C��r��p.�����.v_��xy���5��RaՎ���t��B�
͛��|6Е�@Ѷ�eGEm��( Zh�NÝ[�̉#'�$���}���WD�+8��Zn�Gbj=�4,R� ��P>6��h�+%�:�Dy1w�5VV����1�ZPi�4
P�lX�38 �{tޥ�2j�����q����"�a��|)�gd�6鞡{���Y�4� E�F2G�5��l��K��ƚ���kp ��d�ĳ�
���!hrqT��R��xS�;����#	�U�#�L���`�)��M��*��2^��t�i*���b�K�.UF ����X��x��Y0���!���9����j`��+3�4�'�� ��/��R޼yMp���-���� ��������7���mo/	����o�XOC�.[h\d�ey+�AV���h���f& 3!qQ� ̀���~7G�f���\��T����<ɋ�3�,��Ψ�̴ ��q 1��Z*�-�˓Z]�˘�Ъ�D�Ǝ�fN7&pz�l!�F������l{� Y=��=�f�B0g,pU�|cN�e�\����5sρ�.�a�>d��	\�\�0c>��4M�Pж��/,�c��;��I��4���9�	kt:q�#�����}%s��
�U]p"�+�CR|�6���͵�����Ď�����,�h�����@�m�nU1�9���� d���W�N�2C��K� ,�S�n�<ū0n��b��8�[D�O���U�|�7P�BQhV��%�j6Β\��!J��R	�����W����J��&��RT���C&mB�\���8���)C��HY���<��(ب�踏��LA)/��NA ��	�3��+�w
�T�s� 0�E�Nf����9�W�s�zT��9�Q9 -ը��*.��X�����K��&�	/�ɧ�T2����@�P F�q���}����ɗ�|����g���@�[0F�j�2�Z�S
����V��P���e#�h6�Oi��ƍ�gg�qD0��K����-�N�(���2}7�}WX�����,EKas����H���X��������`�2�b �W��^����#MȕY�R�?쬀��4��S�<*�܉�[k�B���޸�-����%-��(dZiu�����Y�'H���6�W	��{�Pg�1�AUgoG�1��ӎl�sI�Ǝm���
����H-�����|8,Ʈ��S�$ul�䦑�e�:�Y�����O���QypTw.հ�$R��=����j�;�J#C�\��4��J��U�Sm3�9F#rtw�w����k��t�6��	 ��vF���~���,>�E���YB¾�`feČG�{K;��Yc�'�:���W?��R���iQ�>�:�e�� `�ɹ򹵽��� :hh���"H�SG''�)��j0vG����k���{+(�=�y�v,�/k�{�!���7t{w�����#���M��(\{�3de@T.��em�̫���5�B�"��֦�%����r5O@7��!ˈL
�|��ϭ����FK�m��R'��Z�k��� A��GV
f�i�E�3c�B,S�\<Ry�����+̯�t���}cS�D�O5&�Fm� ����!��gc�VԌ�d���b�KNX�MO|65G�b--ȣ����"�
ԦsZ�{��Q��m���sy����� k�#�v:�3���>?����{9;��{�u��wgw��ֵ�����t	\YH�@�E5�l�53���Y�
�j�U:<�&�vP��e%+
�� v~�����O�ã0������t[�$+x�u�v� �A΂�N� WкD��[	�3;�1���-y���v�<K��h�=�|�J��߮Z`��q�c�`�(��m�
�C���������T��ȠS�#Ŋ3��7f��ف�L~eQd�O?|����kY$�z?��f���<�!FSŘ�&o��~�1?��V�Aj_��7�d�V�F�QlD�t�a�c��j�!�F���4�-&4*d�*��Y1�Y!������"$�S��M�-h�D�j��%Cɋ�8�p�X5-��������rm*���ǖ{��*����
5-��4�K����13��pm��7-G��X�.EN��HH.�a֫4`15�����<;ؖ��5Dc��ѓ��p�v9/Xr����njm�U�"I��] �]Z����d$�V������.�P���M��R2�K�4ath��¼$�o��\�[� �NɻH���eSy}��Ȏ����>'e�TՒ ;M��N%jL�ՙf�\.����n:�[1�\Y�?��Ri��a+�U:;��\�������^ ��M<rk�@k$��kT��F�§�%�༨75���M�,�h�*���z�^ф����4�N��8؛� ͤ����>�%�ʬ��+]�Ӂ�b<.�Q1ӥC�UU��!?�<�1xf����Աp�|��/_���a`���P|����s7y}!c��5#��߇�:y G�`FL���up�'���YR��-C&.w�bvj��p2Գz��VrU\G���pк56�5��;��@X��=M�{�V �2���(C�;��j���W���%[(��4_qh6:�s��gZ�9Q�txp�yI,!�P3������|�Қ��B(������1��\;?�܉Z��hs���Rp�.�1}��:U�%gF*��n7P6��Tm�Rf�`@Z�;�\ ���
�M�D�3k��ܜ�)�R�j9�ٳA�a �(���ȱC6h��)����8c�Pm_tHx�]��̮!�O]M����y��5+f{{`#g�@i&�P�ղj��s�&v�G��*��>Q*�5��\�rW�\��T��ƺ�ΰE�*��t�Vn�A�)m8iJ:��5ώ��g�<H�彜-dݣn��A����0��s�Nٌ6���~�/G��~}� ��2��{���]��s^Kt&օ�6���)�uT�4���s��̇'��'I
��yg,k�	�=��t]Ng�VZk[څf�
f��M�dv�I��J']��/�"�ӋƘ:_c\@��]�N������9n|����'����=kf��0r.6!���Qh*��P�F��f���ce
�d$Z%�S,��85G/��,l��ޫ������![�_'&y����yĆ|/�U�xl�6���|~ �;3`�Z�\���cA�o9e�4��|.��½�i�A��p(Ӎ��6�I`E��m�����f�Ԓ/%6,��<�h�d	Y.�Bݾ�T�4�����w�Q�Ƈ�+r&�x�&%��_S����1�����O�!Ŝ�:�8���v���,�o8ND��U�ph�ܒ񸺺����U�� x#��W
(��\�<-eiD!�h��)M��27p�ggrz����pk�ܠ��ҡj�9Y�::����y����_�_��y�� t3G:�
G<� ��q!��(���ɷ�%>��k���������ɭ�t]ǞQ5�h���w+���o3"���qssE@�Ǌ��6+�k��|G�4������v����������ְ�(�a>�� �=�U�W��{_��4����_ij�z_͒�4ޭ�� �X�6b8��*;������9/�"��?2|(7��E����g�6�c:���5� �Y�r`�T�Gv�Nn%g��i����^��ȭ�}<�O/q��Mؔ��;��Kuњ��~��xx�}���P����$����kJ4�ݧ��x���_�Ç������ymo2��W:���� Р؏�!�u��B��TK��H�k��1J{�B$O4g�M������>���4S�}�`k���*SL��5!����$�٩�{�>�S��p{.0o�ՂRaԌ�2��DKA:	�K�MPO�f�"���M�e�'�2>�V:��0(iٞ��_�$���M̈́�A� Y�2�� e�-ȇ����6�ų��3>���b61j	�#Gt�����2 �^.�z�5��2�3�Rkyɀ ��4�&�3�b������T�
��)�4x�*���K0���^n���Gu��^p![�#9���-��n��SPssK�1�7�7�AE�لQ*W��A��0�ZV^|��K�9� �p�U0��e��Ul�Q�> -%)Z���,�H�9�� fO,��HF���6Sd�V��L�����F�V���#�.m]v���d���{�K?�Z}Jp1C��t�m���	9�
���BSq�P�JF`�=���������u�ZM:`�-� �9Fk7S�����-yq����$�#���#m��U�CQ��cp�_�2��0E\�``��Lsh,���	�lp4]���nM��;�Z� �L����#a@"�������h���y��������������-TN�UC���O,mx6������Y*�J�X6fc9��a
�E8:|�����D��=��Z��7Գ/D�t,t%XCi�"�
]iu?�������9�r9�
 ���.�������/2ѕ`�����₂�6����ۀ�w(���N��I����k���d�idD��~�w a0ݸf������hؒS����K�L�~v��&���G2� b#]t�_�5� � x�@����Ut�u�(�͝�맆���:X�S�����)+,;D��R] �~�<6qL��yBڢ̘��0{E�O�q��H��s���j��� ��s��E�ο3[C	�B�N]'�3`,ɭԙ��r��R�k� �uyD霯,ˍ{Xut4p|(Eߦ�����0��V˪	T\�{�i���f.ߟʻ��	ֺX�Kҕ:S���WFB�l��ŵ���;��Љ	W�� Y�c�h,�!a��<
����w�ޑ_�5"�0�vQi�@ǘi�6�a��:;�+�ؿө���9�3�(��V�f�VhvX@�,Ra�Lv��bFл�o�9�r��� �L��2�P�q��f{9� c��� YǆT��@9�oh{ЏzA�gI
��"�����3+�g��&Z�@5������{I߳!?�V*t��RM�Ǫ,x��%�MO_7̢vZ.c���bJ��Җ��ȑoK^�ګ]a�2�gsħ���jV�`����S=Ш��T�;�I�CJ�.�d3zhLc��?5{��6`b�~�+��V~l�k"���>�6w5,�ޤ����8�g��؆�l@<�����cV)h����)K~��*MR'h�E�k<z"�!=v�%�9�bt�JǗ�٦2s��̨��^�$V��% �N49�(>}=��Ҧā�{\1�Fہ��cH��\%�[�c�j�1!}�%��4F���ܱ֜���0m����_�ߴi�a�g��U��,9���<D��^�ثZ%V�u��Pr+}zQS�9�p_�趀`b���F��67�rt�+�;����r�F*��Q �ݻ�l�U��d:~*H�7��͒<�!���4�����90U��2*N�u��*�v��JF�}���N�E��3'��C;ʧmzJs�s Zj��1\p��=�Ʃ���-[�� i��Q�D��vD���/��Ay�M�|���ru5�N6J
0���ͫ��w�"���3oL�F�� �%Y�*���+��2Gz�-`Y/�s8�S�Ip{V���s��*9�@ JA�T��J��.9	 H0,Qz���C4�1v�����>sw�_e�/G����t6�ãc�QA�k �<���¡b#�l�q�m<0���eU�CqH����� ���	�@������%�3��kS#?M���t(K�(�%
��Z��f��3����c7Mh��R+��A<�^��M&'�2�� �����Di����:{�Y�4��J���)z�ҳz�ϊ��9���E����(��+��<=;%ge��Yp'��W�፪ʮS��Q��t{E� ����XA����5tw�@��=Axw�tL�L�qI�,��Y���o%����|<�`3
��U �^g`66B�ʊ���m�P�����0h�ٞ�Xו�'f�:oX����Kv'C"B?Kgs"K��h5���rI{	�tϦ���r2'���1a��|+�P�q}�ԿZ�{��Z���	���ځ.��CK�����2��N�p,�ࣉ4sN>��D�f`w�b�����(:��?'e
���}\���l˜�ۺ�K㠷����� �jUUE?�k���ޭ�ql�ә������ۯ��#�o�����{.VЫ���k�u��#�#8�JEl�Bps� Q9"�_�5ݯO�W�!�?�s? ���<v�Wk�f�mf�'r<�Q�>��s��$�:j	f�:��CԹ��&M������9���`y��ίD�s �~'��YH:OR�z�6��V�w��v��T���^��ք_����w�����mTY��F��D	����H
�Q�'�_X�XT���Y�"�u��&t��.}& ��2�'GEj=آdޑ��5��Ws����E=0Myf�E_�]H�!kE�y�TwL��:�?���2�0�v:��=�O���xS����G2��@�jwg�����R�Qؾj)M`�xoZ&R�ԕt�ݪ<]��S����u��G�t���i�a���%�7�~2��̠
��@ǒ��'���(,V.^�f1K��.fV!���/��^x8n8ݕ;q�m�HtF9 \l���m�Z�LS��B�]k�_U@g֣�(�1����s.n<T�=9�0֨�2_,�qM��h�s�$"���A	��ߥ�;���c�N�e�x��QbBI�m.5B.���
��ՀX}�t��v��&2�\*�:��ap�J7��7u��3�>>^�F�X|��b��csb9�"�Oʚٯ��K�kjY]�uc+E��?�u�{@�݃�#o�6Ά�m,	� ����l����Y��P�P���Z���+�3�@�م9��~�E��r�\p�j�@{���l�Ǳ�*a������z�9��x26�}��w�k˸�]�g�ץ;p���a���p=�����\�O	��RjȺ S����.�9z���R��}��VK~���Or>��ʴ���A��ŎH�O�-)�����{���_'0x���4�T���#��$;����[A0��D�h�(.�f0��5���%� 72� &}pH��`�	۴1�L6aLۇ�p}���<�����s�"s0���h��%����C�"�[-��X�D���$�:�`�)�q`P.3:�4'��+���-�v/��i�pw�g� �W]-�z�)%_���?_�6���"�>�LT�g�4[]XРC��b���L��xJ���S`�M�?-��ͼ�<�����P��%Ĥ�bg3��}��H"�Fa ���S��N�������2[�6� cw�i�Wڪ��b4M+{��8�/���kZ���.��'6@�	�ywwfr�|��U��~�����D������!�������S��J�WdN;V�_1fE�Z���%|H�oMKѺĉML�Y�t�wRЌky�L��S��UTT09�B��v��(����SA�d�N X�FA̚t6��҈n<�O�W��8@+%��tTߟx�]�Z��y�a�(�W��z��r�f:z�"�y�S�1Z�.�_gd�� �(�Y�3לuF�4f͔p>M�po�n�ώ�x��� Q�P�)j�U���$g�\rB�&k��1�V�_�N�)B:���ж��q�o�F1�A��?����LFSQI�Kk����6�5V*�����K��\��J�cr�>�̀�S�tb13�Ь�Th�o�p>}���N��w����˗�ZFFP0C�����fS�a�GNOSd6_��Zg !�O��A"���� {}r�-{;[\kP���?���^�����@н���=U�q=O��H��=u �Z��AY��e�mt���R��/�/Q2k�zr���Ҹh>�S� d ��L�����k�vpb>��?� ��_aɉd������A2��� s2	fZ�U� 1�I|D��u���,an>��ń9�5��r�$6����lF���B�M�4�;m~UX�A����D�R��;m�v��q�[u�����R+������ao�}���*؟�Ɩ��ѳ����y3#��P}09_��mhV�a柃=�u|}ugr1AϯS�fT% G�+kf�p(���]�����v19 �)�+����UV��Z�	�ϱfX��Hn
�Ԩ���-h&H{����b�5��ks4%_��?���R�W�\'����;������ў������oo��p|�� @a&�q��T�����ץa� ��*{��F'IL�� �foG~_|-�߼��j� �_FfL�լ�m]e�GQ�&��m'�� �����cT�"���u]��g�C�KV�#��;�yAm��昝����=�E��������ܷb�6��Iұ�>J��[�� e�gώ��/�������*�������D�I��("@��u�2 �9�ܹ�������O�@$��9lɳ��w���Ǭ��+�E8���t���_����S� l���
������/	�Z� ��
B�ȡ�T/Up:��zߤ��U���5������rA�8�c�C�|�a!��S�͋�>lmDZ(�4��r�Mދg�r�0�2�rY��Ѥ)gFk+�c]k�)3p�Ld#%��CZ�1A	��ު��Cӗ�
LT�g������ƚ<��EP�!�(�֦MRM��LPuz4����1��G�F�l�8��𔥺X��j�U��]����hd��-p��6<9��/�4~�KΈ<X�v�]_E���?�0��(���ጶ�`P��$�y��W�b�9̠��U�#���Ɖ�˂<��VK��_�����j0Co��0%���i6�&�ÆQ/M��� "��Р��ɍ��]����62~2��}�qg�<�=� `w�P�lȕ�Ey��#��*?���&�rc��ER���a�-xp�H���"��-�U?U�F0TW
r���Qu�jkL kLlu��&p�Q@Mc�l��-3bKM��J�R��Ǣ��4���DC�n10�tb�y����ﳡ��>���˟��ș0ə9_����=� Gsb��X[8αLpȚhb`?*�/s�Ei]ʚ5��[���Ѡ̋�9�-��.����W>�n�6&���MoAnX�bC�Чϛ"Ù@+�{�6l�f7�G��AǢ���9{�2�Z�_Z�X��?���,ى	J�e����6�v��]4NT��м�©�8y�@��{#E���i�+��o�jX����ę�X��D�����C�}!�7W촜�����}��|��e
~egd��Bc�x�Y��2��^�a૰`Nm
�UmA9�&��>��B��eAs�-��V��lR�r M�Yb�}^���z6�T���#W�&@��u�4f����	���A�1)�T�5���&(�6�C�ڄ8��<�N\NJ�Zi���� @Z���ݝd_�־��;
2S��4�4�Ҝk�F;�WL�,	�V�+*2�϶���S۲���@�fa�2��>����0��5��r�x�@�dw{Kp�K<�uձE����YY�eC� ld��àv���ew^�4��<��r\# 7��;�G	b]�fe��L3p1X�%?c��`s{���F]yI ���s>�	sFKm�1&Y�6�4�M]18�E�L�[�s��8f���Ѵz�:���$���a�����S�W7�/ȥXA��H���J=�4��`�U�ry7�nԒ�
߱��-_�R�|�B޼>�C, |b�_���!�!ˬ�|w��w �̩�SDgMcYB�0L�|� at
�Ls2`(��3�k�������w1��ހ��I�Y��!�s�hF�q�"O�)��YP�kP2C1�`�/�"��M�z�!֊aC+t���E���o�a�hY��?��������c*��������rҬD�{���j&Aa���S�G6�C��~I %t8ܯ4X����wN�1�L�KF��Ҳ��Dr���eU�$\����:�6��MXR3F\�N�f�b�:P��o���cű�}������	l~d$���p8�o~�;��]����g�ż���
Yv������d�Ţ��_`�8�\{Y/�54������u�R)\2}��vk��;V�oON��U+��Ep-g����65x�YL��h h�Pp�����W�	`�Ks?�����&����(ٚ9�	%st�b_�V��3�(&�� �/Ӛ}��B���(N/�b��;ĖI_C���x�Ex��v�"K�z楦�D���q}0�%P��"�zT�:@|����fU�������rI�wvVr|t��_��0��� ������\,�����?���&ߦ={��:'���A�X��U[Z��q��7Ǆ��g�<�:BM���F(tm�hp��s��."����m�l�{��R�>9z���>/����P�PH���[��d�y�JNa���N���i�*�j Q��}V>>��b�lxV���{PGF�6N�L�o"w�)�t6p�3��2|������6��ki7��3���/�H���I\����¤س�$!\\��'r�B>O�(�pJG��5��%*��> ��7�L��~�&'WR���fQrm��.]��US���;���=66n�3̣����o�Z*� !m?�dooON��dZ�Ð;��ц�Q.�E5�K\u�.���)��"��4�b#�U�Z=-L�#�s꼼&���ڥ�ՌSi ���+9><���s���tv-�N����`{�B��tb�`�{P��2Tr:���~�L�����pa�2$�$�!�	���wh��m&虵{��_��D�\�[��z18��Ţ�7�p'�:L����vڂ�õ�n�={�g�k3{�^#�Z���'b7�d���*�X��f�pC`��Aw�`I�e�i\�`&����G�U	Zg�v9�U�Q�v���r�aė4 <�<���H���~��Sؔ l2�� �	� Wi�l�������Or~u+�rz�}��Z.�O��4�T��/�m�@OR���fr��)��y��,�Ԣ�Lm#1pM���h�7x��8�������~��x�|'����u�
%�NLP6��2�.�D���uϦ�������A꜇|�\�N~� b �-Ϝ�RCi%�%�E/�_�����e���#��8�Z��q�~�e�1�:_2�[��si�u:'p
w�3H�I6��hb��
����ٜm���N��

��˴&�ݧK���(~��RZ�\�h��@2H��RIߣq��	t=K�����p0n��~\�.�5��4<^dOg*����y_G��,�}:��M๠����Cb����������{������o��B��Q
{�e�[yJ��V�R���5�`�����]��(�l߀a#��v)�4K��aJ�Fd�}��.���'�}��^{������6�O����b�ol�'�����'$�c��9���o����: ��lB���,ٲkv
c�m����C�":�i��t��5��YZ_�H��W18>����#�Ub���
Bc�B�*��^j����N\�>�^�ź���Iؼʚ��r�+����I45�(>�ύ�v	{��xJ��5VqBQ������@�@S�RO��@4��u(�4���a���&4�AM/��s�D��:�.@v�E�~sXF�Jf%k�J�C��,��I*�a�R��Y"�����,C^]�ʻ����"?��N~M__߂���E����Ä�&9�ŕ�Q+��ܟ�ț�G�</�A(yIM��5��6�g�N��F����̼o�w˪�>-މ��Wb�<��OA',���{<>C����snA����"o��� 뱁Z{[��ix����� ޼~�u2�|qA��H�T�g%QZ ����|>tnB�}�����Qr�[����i�����/&�4V�v����;<���s���'�5xvuG�����ls��{�0Ub��joal�ɳc�����/^��:N�K��í�:��q-t�6����"9@-A �L�'��ʸ�n<
 @�˲��_�J��!QՖ�㭉9JJ�D<��N^m8Fi�F��T��0ù����4���k��>���Y0`����
/��>8�<�І�������+�}$j6d:�L�t�
��i���u�;[�λۛԦ����N�5�h���d��2�-�G�z�>�R��h�MP�0�B�6�IV��w)�O�p�.������g��w_%�vr$��1V�cWW�1�K[�6�������!���ڕU/�8l�{�drA�1A<d3�˙�v���q�Q�M[k\h�ay{�ڱ&"p�6F�mJ1̄��l�վ�%���m.��@@?����y���=}ʖ>|�:�����w��8������Ï��R@�Ў>��0��	�w�87�*����k���w�}�S�D�k�KӋ,[9H���'�e�N��dcV+KC���UҞY�L�z��^�}���r���
��zo]7"2��8����ƭf�4�����e�J���$>ے7[��9��>l*��m��-d�4^��5�����c�m�%G0��zd���F9.LhPk�E��!�H��i�~R�&wy��j����u����r�!�z	!/����U�k2��mU3k#^X�o���L�D����Ù��_�����K�U�X���W��^2V�{;�=�x��
4�Y����p#�(�S�}��و�����	����)?�e�l�5+��#>�U\ϐ����΃�;҆F��.
�s�6o��5+��A��!���u^b��F�Y3@㽉\�,��x~y�,�>�kY��e�JNOO�	����� ��6���s��Z�S���(mG�=x�)N�iZc�AF�m��X��4?��&\S��t]�(�1A�v*/w��_��o���|��e������a.�m2/O����#W��{I�S�UѴ侀3���fcf����"�c`�����s�:S0_�7��������E�ֽ��LY���օ��4�����={O�N4��#Kb��`��s�XfC����=;�"G!����39><�J����[#4����Y���Q�#� V����*��еY����&B�N�����<�B;�! Z��![{��+��5�DI�J�����Ե
A F`�����n]`�7t>�^6l�
\'�����z��1��A>G�|E���T��ڜ�J�+m��,�d�``�A@a��u�3�)k��ǽ)�AW| ��pz��k����8���<~<|]�����/��G迠�������b�G���Xv#v����� #��GG�v��\���$V=S3�a�h:Y��W�� �H���y��X��m>a(>�Yed�'AKjT�Sa�����}b+�l���Q�Z����JK�yY���؃0���/��}�УǞ�}I�ߨ��i���B��cP�0�\3��2B\o�e��_2���9|�\6��x ��_]�C۪3���,f@%�$�wz��3��[̓ݭ)It�7���އ7&��S�;���/�qZ�E�i����R��Ï�����䗷���q$���WA��(/�/X���2i��k�����b͈�~?k/,n��X���X��g�9ˣ�k��o���?��@��p�c|����D6n����y�?�߃��~iZ;�\���\9j�mPF�nު�v����� ���hHs���l����;{��� �0��&��y�)���ӌ.� ��Txs��~=��l�h*�����n���X����_d%�Z���G��ӟ䏿�B^��'�6�����O�����z#��?E�-��W�vrrL��s�YQ"B�d����)�����Kfc�
ηd:��@��	�vs�} ��ñ�Q� ����0ҷq�b�C �+�2��Q]g�!=�0��,7�;j߹�kN8;hX1����ۢҲg(�Q���
���z���47���"��o~���y�Bvw6�zI��H='hHhǿ <Ʋcp5p�) ��9�amt��6�Q��39��(�ɦ�[#9JΌ�.K���dV�n$�G-�Һ���T��m��7�@�p9�
�M�~no�M�ێ����f&G�fN)�bK_�N7�fd��3������UzG�jH��c��`?�ǚ�3�����c[�n��zh���u���9�^W��C��}�������QE!9=��M���r~{�	;���>����y��LU>��Xs��m��������.hbX͓���f
L@���_�W_>��]d���Nݖz�W��~C;*%dЕ9$ѩ�bu�]��v	1׻���i0:1@�c���G�uVI��`E���+��욹ڂ6V�;�a��C> ��	pv�����d�r �2�&�PO`��h��ɼ	WkUw�rd$�R4u�D�/��,��@���Z/[87�Ua��L���c�D���	!�\j�e.h��&��.>���1D�JkBA�����If��)�<9ؓ��t'���_��S��y*[3�7(ǢZ���y�[�+���k���S ���xk?�����>�Ɂ���Z�ќ-��%��ư�L|�<=F/{}�>j���Cj���������f�@'h�G�MH`dwsJ�ѹh
��ɑ�*ڸ��!����m�MT͵���S��]e�C"c;��+�1����0���l�5�1�M@�ɗGa�^/΍�ΐl���/_��d ����������cn�@��q+�IZ)H�ȸ.vw���k#�B��Ӷ
\���T���ˆ�=2���zB��/!wap�{4p�qpl:sR�߷�,[tM�v@;�S�lE�&��!�	 ���nr0(�]��r�A�C��Ō%��mĦDd ו: ~�g���&:���Gٕ3�p���ֲR�1����k�䎝�*��}̎X�rg�) ��V���c�Dˌ��wٓ�O���9e%���Z����r�%e6�#����u�.�"Ӽ��v�]����ѥ|ߛk�,�yq� ��ӛ�'m�C+�۰�������ߧĵ���q����0������h�}����O�3�B�0����i�T��#� K���>�^����/6�!�	�d��q�pM!��M���LjS��R��Ǭ�Zq?����$���A6�� �o�Zo�|
�_��:�_멚�{�4J��yO�Khq"8W�1W*tU!_�x��J��Є���_���C )���t!o��|�bD�$��l�`� ����@��M��<�M�gĆ'D�{e|�?��U ��	5eS�f�D�y Ə:E�$|������5���i����@&J��������d5�e��,-"��d�г3�������O-�!�XOZW�d��1�?�����������91������Z�J�F]O���1|���Q���p�i�e\V ���x�9U򥜘�6�NT���X<;�g	zgk�e��4QbҲvK��"��w�P�yԉ
��{��1Fd�M`�ݧ�ή���3Ӑ]�4B�0K2J�m:�d#ۻi=o��QB��Zk���?�^�6�hi�ɠG�rJvD�~���Fc6ۤ�>���c9<<ҙ��Y�e����j�e}9'��@{�-R=��Y�>�m�7f���c�7܂/m�V�	��nKt�9/(�^�K̝�0sJ���݃�^x�C˳.ڄ��o�O�"֜���u���K���u��ە��{��(#���\�D����Q5@��J�n/ӿ��Ð�&y�3Q5�]�nb�&`,f�#�d�7�Q�����~����&�~�������&_.��V�(0�K^���Eh��l��db�����֌�-t	ƣ��+iO����(�ɨpR����V>�{��nh/�C�����߯���}��W��>�s���q��������!���$��}�:�e/�����.�5[ݥ�Nv��|����z-'�1xL79���Z4T^8>9L��p���*��9�YnC�(� 4~��'�S(a�˙����_9����}�Z�(�ћ/������ �Q`
햵��t<�u� �a��P͝uy?6g�8_A�?=�AS��j��[ޑ�U��������,��k!���^�q�aʺiM�Q�+5�^�,L���w"D����@���M#��� j�����)o������������u|�������q}���F�
�9�8HG��� ���"��۟�0���?�|8�����@s�A�c�0w8���c�EA�rh��y�� %F�m>���F6 �(㛗�d����D���r�,3W���r����ʟ����{��Eh���w��/o���K��KF��8�"�0�:Id,F��\ty2'��mݺa��"˗1g�^2ȕd�^.5�<�md0pN�窂���K�������Ɯi`����*-�gɀ�� Lo�Q����eE���,�O�~ϔk�@}�>b�M1�c$�z���9'l����ڷN��ڕ�^�*_����$ �U��L<��ݽ ��@����Z��v����f��TT�*���L|�H�Y-����5h!�L8�+��0%�ݗ�&�K0mݎ���:_�b-Bf��&Go�S��ޫH��h���%[{'	�Tvŵ�Z[k%A�Z5�i	��&�c������?i$����J����W����|<�m������ZA��������ӿΒk��`}p�za�>���ogE������r�XA���1)
���lom��_�`���p�Y3�P]Q4xE�Z�=G�hcs[�Odcc[��IqY�#J��6�>K_q1��a��U�Xsag\�px�!��g��N�Z�E#*gh������8���M,em{�W2`$T�[����MM���K �,�D���w2
>%QT�rT�k��l��w"�/��(J���cV�+v���<���]���ZNI���Cj3�����}B���)Ժ=�vq�4&��(mwwS���uq@L����a0,J�.���4\�Czf�ֶB^���Y���M2p a(�����u�o����m^�H�^g�N_|B>>�'�w"�|~������7��Џ������yS�0_:ҥ�j��9<*<�1I��@��U
&�y�(�Tu�n���s1���������8yT������'��?q8���B��a�c��J�I:�N۴��D,��.�;�j������	�uym��2���Ɣ�uе\ ���#�?|�2di�!p{;c���;�T�VQ`(7�v��l�D#�_W
Y�2���H˺e�߻�p����#����B8Xg���s�}��Fk/.C/)���jV6���a�\\]r8:��㑭��V,yk'��4�\O�2�C��GÖڲ�Fv�}YW}�doG�x����1� @m����\pOA�t3w6� �Ã�my��$��@�<D�V��#�9�������C`P���Q��T�G0qy}�r�\���Y�h�ȭ����קl:K����Bu��S�s�������@>�X�c���ff=ff�ۭ��|�����?㩰��f����X������H�!��� #��1�V:�(�*�V5��9�ߔo~�F�x�b��.|�H �:��a�x�|4�Tës��`\�B���*O�P��j4e�J�N��6a�)��^�sW$� )SZ`X�(?��h<�Ó]6〾�%e/��%���N�Y��.�Ƈ���u`5��-	�:k.JA��"nQm'�N����8��@v�Q������F�D�Bf a���d���V�X\�
8�&م�����F2�"���ר`ܹ�D��	�%vz������~!7��B��4cg{-B�3z�W�U5Ϸt3����I_By����[3 vo���p���L���^�޸���7�c�4<�]{<�x�G׎��>'���:ML�,0�T�rn�N��f�AV�R䴸����K(��8�	����� e��.�U����UKɓ_ ú��*rXr��Q��83�wj��FV���[��l�gI�Z0�`m���=5:X�8p��}�N>]� S
�Nxũ�V_�A$q��J�Cm��8��*��׸<���J��`��m[����a�I�WߣE��a��f�{�����+|��sh**���2�juO ������{������=K�y'����4�}ڡ��f��~�-�/��^�x�A�Џ�����B�/����S���Ɂ챥���U�t,(�R�������g���Ѕ��|2�
����L6�v�.P�>�����Rݩ�.#��q"1��8�e�⥚���n����Iȳv��Ԅ �ױw����g�к��Ͻ,<z��x<eaŬ�Ъ=����6�3�Ǚ�a�r?�y��x���e���r@x_��W��Vjъ�/ tI�����SP�DP��6K��(F<��n4��������FB/�nƿ,u��S3暁Z.�c���*K�����v�y����m��C0I�p:���C��SV��s�v�z��|U}�j��Z~i;K횠`J���bƱv�D�pAy��0�M���f�y׊ �6�?AKr1��ۿMיx�n�����sd��#�Ѹ�`�2�~A��Z]���or�SAi�q�C��ev8Y�:�����:2��C��'��:*Bp�ք3��wg���q��r +��k��3a�m���!
�����ֺ ����{<��S�����S/��9��|ks�vrC��f�E\kF]XQ5~	::��s��U\�(�'�ʺ�w����"�@��z��G a�Ŝ��B9��&7�͖�}��5v����Mc@�?�W�J����kD��0A�=D[?}��C�f4*�	"s�Y~��q��<D���#���I^�zI�/d�5�&�0�C��D�%��j���WG^��=C�u}2{p���}1�x�O\G=u�Q �A��!�6����fX��~޹<*HY���l?�{�$\X�����A6�"} pU�UAه����ﾑׯ_��R2ȹ�~`T������Ⱦ�psڦ.f��2�?4I<;:��}�:B�V��?$���>���o�bV�$�QŬ��D�e�pȣƠ�����Q�	�|���3ClØ�E�2���R����v%g�K�� h�lݢ5��@��CZ͎��AxT a
�*$\�ST���c��ك"W]��CO�����p��c��uD���2>��z��%��_�����7��u=#8����=�+�<l�Q0F��9
��h'�ɿ��*7�����:���)�G�:Y��І4��*o^y������x3eƱq�=��0T��,�3�����1�SG�LA�8�0$���Dʇ��N4{��q�3�t��H|�j$�(O%�S[����sޘyH5amk�T,5H"�hf�'t~��@�:}d*ʼ\)2���Q�8)l|
A�uμ�������d膘�(�������ZpQ?܌H%�&�d�����1K�P	���5a�X�`ѕv�=[4����l�È/ZK��[߈��
����
��������r~a�ʆ��s��o=�7�ߌ���A�ܣW^���%�+�Z;K�,���dS�����79�(h&Y��XG�p��+�����{�����|ц*� %(I!{�5�Vz�M����u3�����`�)�c�`�G�XP�rz`Mw-�1�P}�-���V�aD4�^�����1b|ثWoR�y���M68�҆,�JA��������t$�Z���e�EK�����s�7a����WD���#��mv��Q�2�̥e��z�r���ϲ�[?����p��ǎ�9�y�r����s�SM�R�XQ�Mc���,9��cy��x�B��=�Y�5pqy#�7w��]RК�@�|T: oP#����gt�)�J:��6�	��i:�v~�5�������Б�΀t�����{�Oum��Qj|�����ZyX0��p��[V�3F7�Hkf�r:
���PT��&+t��B��O+�8m��ӻ�	��7=X�1F3����]Gp���Z37�e��
��/���=j	דrn�ڣx�^y��O��'�_2�����.>�9�wC�5|��+<$�
:��}��2= �#�6�1C۩$�rt���`90��h#�����~2[7��v�&b�����V�8Ǘ:cKi8�c;f��kf�C�?�0�V�&�Jgk����y���v����|��4g4a�������hf;�v� 7TY��$W�v�Q@��vL�M�DAY��w;�y�3`K"gtL�|��Q[���W��f�Z3��j��6t�5�c\s(�j�B3O�f�4�� Pk�tww[�m>nΜ��<��7��Mu���p�v�3xw�֛��'�������Z[a���3����6Q&����� r���}��|���׍�g��7|x	C$d�:x/��W\� ���X�e����LYps6ʊ�6̅D�LӪ����X�X�Ř�j
UG�s��"��|����zt=�Ѻ��:��ɦϧ�[��捎��ʫ4UTfN��\�m��f:��=�v�]t�((@�h�p<���K�1�>��jTP��b e�1�s	�������*�~���+���a�^�
��VVMߖ
v�� j�%ds�X�|�&�x�G�$8�/��:��u��э��l೏4����/U�egw�9u�|��X���?rn���yO� B����1?tN`�`F"��K69�0%���MfSʇ`�Գ����F���y;ݧ��� �h�����������Y�u`q 2����
�o�$Ǩ��=y���Q��v�p׽��\��\od���VMEm���d��B8�#�$�KX[�w���z ׳nE�u�!�^;��q�w����3��l�w�yg��C��ݜ�����Ap���#��{<.������+P���`V*���׊v���HE���9�k�h����>`�|YM��ٰ�,[(���?3<<�! ��ڑH:���g����J;�q�
�O]t�aocb�%FeR���d
2����Ad0�[��*�e�W�U���U@��AT���m<��:S�fE�+��Y2��t����͇��:͔)/�6��-��x�
OMkk:O�T����A�	�>�~�-5r�m�*-;�LJ8% �H�@t\ґ�J�n����~�p��ukOm���7�4�U�@f=�l� ��|-D���P�u�x������mV�`Xv߭&f5�Дy�o��ȏ ���Y�[����ӟ��آ�շR,��{S�-����Tm�筨�Z�at���ʝu����8<�'k;�2�RO�G�y��%BJ���J���;� ����5���0(B3g�(�&>���0{�q4)���Ĥ�zu4Xe��4Rߋ4WU/��CK*4�,#�/D�ѵ�ܙ��1�;�-��F�ryo8j�7T�qF�U5n�� �9Ȫ��o�5���e��×:y�V�p�+��^2M ���_�"�:99I���r/�n��w�����}�����=�W���+��ҸH0.�J�R��3YΗ������A����ƛ��EP�|���K����ʏ?�$���^nn���uaHU�QC#��N &{xuM��1/�	�����!��T:�p� Hu�6��V��k�˪�U4SD-.�';�Hv��k˅D���C�5X�g�y=��
�׬rmR|�ݧ\f�=s�m�e���C*m$���q�_��k�f��x��v�P�P_Q_�6l�tF��H�z���~�C�#�1� �fc�	."8��I:n��,EIkЍf��b>3����P��#ة���S����N�d��e֐+��$�S+��T_f�ߋ�3�	 �4IČ���?mh�TK�vPq����f ���tqr^Q�H�4�?;�����M!g��7�^�`ݸ�9Bw"[��H�^W�`
RLS���`�b��_|��>(8؆� ��[V��8��D��ZXQ�9<<d=�@%K/�m$E��'f|��I ��E�O��:�z
�t���z9�Zt����v:����X�3�Z�	e0+j(�*i����JK,��E_&���󍖵U�7qp������qE�G9��s�;A;k��Jf6qeU@Ry8���jwn� ��3;�zX�hA
����`��	���҈պ(f��{(!B��[��i-W��t\�!�I�bGЈF�ԑ��ã�̍�B��r/�*����5�ЮG�A �Xw7,?�완�D�Z(>wϳ�}��?�o~�B�ga�o�֓Y|i���@�^�Íu��*{�Q4����'מ~=�d'W��ut( �TٞNST���[ыRɷiuvN	��I>|<#M�%h̨�y2Έ5��`���5�R�	M'���eoik��ʴ)�f~�>�B���'���7���_���ȅ�:7c~����Zgw(_^���_~!ϟ�<����;9=��h+��ҕ����"T���[��˨�<Q�)�>�ъ�
�zC�����V��Y��i+����o���(�CP7����n?���J�@�7Z�g4:@��{a�2�/2[���l���q��ע%���!�}���:o�q����y��|ޞ��)琓GT�&��
2�Ʌ.Ix�d`<Ò�;#��8�LTY�ˍ�#ȗ婣~�J�_������Agus��1��=����9H.8�v����0�����$�'w�ڱ�Z��gC�K�5:�`$D����nD�_5:Ëc7lP��+��o�A!�U� =K'�h,ˈʑ�/µ�z�i�S��W'f�y'Ȱ8/rrH~�Aû���H�S�yY��io��`�D�6�goBȆ2Gk��?�����C���D�dݝ'�n����U�6}Z��ꆥ`��>Fy-�5� ,�KV@��*��p0���%;��C��f���vC��.C�a���v^0�u���}}.b��N���J{ډ�Y��F^7�!��>W����W�Ih�\��oUgdP���=< �U���%@}�R"���=Q(������ߨԬ�6Fjԛ��������)9?�K�u�Fjɵ_���)�3���Qm���,tTWTa��_����σ��o��Kc�&�ۦH;�`"@��ЇZ=|���ǘ�yj 7 �y�>8ޜA3���i�ϩNkj#ݯ��M������F���ا��[F�l�Xi��.�1�5 unb�z��jCf���t��q��m�a�Ɔ����_���~�5�O	�wY<�����}.6�S�OKY�F�a\�#��  �Y��0�K�FF�k��Y|��Ҳ�3��܄�+U9�����_o�<
}�c�u�� ���}0|�!��_?(#F��1��U�q��N��/1 �_����ЊK�&8 �g��ܲ�- .������F �*�Q[=�2����VZEj���N[�z���������}�[�6�d:Vi4�����qԲ��+�M�-��%1L�<<��}YCC×�5!���*��F
`URG{>��0�jPy�q/����R�% ��u��eV}�w�{�3</%�����a�y:!p9��9tqE���A�%%���ٮ~���|��|1l����r{�f��A�/_��V�s��#���"�	�Z�k8����;�r�1 �:^�o���N���y��|�£߲-W�E�x��\����&mr���|�n��s%w7���"����k����eM�9��l��J5��Sv�Lf����l&�+�Ƣ;Iwp�i�n���_��o�d�hi}��nѴ�_�5� ͛?��/��P$j� �EL�Ό���J�juK�I��Z�f[2Y�r�As����M)��ƤT8���ĩvpus�e�J�e�Q�T;"��\H���c��ؔ��zI�t�>}�(���S��7�L�Q����S����L��_�%��+r-�4�Q/P:LOdT+G�rӨ�\��i����>�ԋ^�%�J a����@�د�c�;���SX�=��)���L����%�=�I�dA��P�-fV����w��wܻ�U#��K��%Df\��{D$H��ٛEh�@ ��a�nnΨxh驭uZKm���鲨b�C��[�(jD,w�-�d������h��/���D�����܂*}�6k�qy��!X
�`�֣���wVq�B����;$�w�o׳�O\�H-4�����|Ǫ�<ب��#6���l����Z�1�i���+;���8�oX|e��m�����ZԵSЫ��BY
���v/b4����e 6,�C9Dw
:�+>��[O�~F���PR�9������}�6����T�S��^�M�U�[\[�����_��mS��
������J�i;�C�jn���͔0��&���m:=/��N[����� �dX|��.E�f�b��R�5�8�ЪZ�W����Q���2GS�Z�v�c`����	tm�vd��OD�"ڬv��������B��J�r\O�?��K}��$!�@�o�آ,��6����@�H�<�>��bچ�h�;����3*Ϋ�z���q��4�H���|16hP��ir�i0�;�Xy`�Q%�S���s���
��x��ε@+�(�G��-C��1� ��௡M�K	 ^�B�X����R��C(?���g0�m��Q��?����z�5�k�d�Y+l�||!:�� ���-u�4�����Z�p����sO�8��d1Sx/�b@��� >��	�A�Xt�8��ژ���Pޞ�����l�5{�v2�'��f͛��ksVoE�B{�끥��cگW92�K9`K�D��<��C�b��4���F����4�]�3*8��$�n'��t��h�"b��a�p�^v;�\X�ْyãt�o����a���LY�v��H��!����]z�~��V���I� Wח�H�@=7I/��c���׎Wz��UI
��{O�h�?m�l��3�������Q2f�0Yy���U���6>+�I��� 7s٬ԣEň�J�"r�l��٦$��4�{�gCZ�G�u�Xmͬ��q!� �k��p^+S�ױ� oT�a4.XרdS���*OB�l��Kd(�Sk4 ���/����i�h`:�k���w��iY������N��hվ!�3�M��4w��V��'�9p�;�HXX�� �s��% m��4�p�n#s�5���5�zz�͏L6�\8�ߙw��w���U���xYt�]4�֦_��ee��@R(i������9�6����� �Em�B�/����O��b��Hc?����d��3H��d�M{뎸�[�g}�L��,�.V�_�<jm@�
��.QCa*�=ܚ�\�q��yb�<�s�*٠�|�+.��!�xQY�uFY
���= L��DMi6�Z�%�OA�1��LF'cӒ�B'���It٨�y�����*Ȃ��z?EF�$�O�|��?~~�3�oo�p�EP���\x7�F7���c�q/2�!�%���=-�"��
GU�.S�)k)8��ző����%F#����Jn�/���J9:���X��`ͷZv�)z*�Q���n:��z��K��B�vY��Y3�u�<���i\��xu�JE�f:��J�N�1��3Ή���րL��gm�a]Q����,|��[��S�r�"��"���hZ�����?.T�k�>�����Ѿ�&�9�k�����ݜ'Cy-�����o��V���Q^��;�������?0MD�g�%d�ZX� U�T�o�����}u�h���<�������`�A��\�@���������w�O���f�]E�)ׅy�):���J�x�F���0=��|��H��[c�/?���߳����F��j��	�ײ%��Y����t��.#ؑ���ք�Ԉ;�U�S'K[��-L�tn�~�S{�ָ}�ƙ�԰V���l#g��w������Ȟ���%��5���49HUani����{�����UL����� �#j�@��F�h[�3]�	ro��3F@��A�X�U��6��0���1Zt�w�2��9C4}7�T�~��XN����F���_�� �q��=I]V��C��x�W*�ү8� G�  %�@��{��X�)����$ǌ�i��m@���m�^�<DWm_����@���E5*R���@�}���F��g����h�5��9SP���b!�Q��)K��H�yT�Z�x�5�ZtP��=���q���P7�}���<��D�پ��������R���Im����tͶ���'��~�7�?)A��Q��yԞ���) �/��y�YډңR> m9(Ҏ�C����U��-�G�������Mw�bC���] ����0~�h:Gs�(yE��/�tU�L�̢�N����j_ю�ц�{�wo��Q³p��,J�𺔻�s����Ǉ;N�����)���I��J:�Ǽ��G���<� �w�-��	fPÝ����K(��(��=V���ED�9}~Wo�*��ǧ̡���Xڰ��´f{e�t��{�@#���Ki ���K ^�h�(ٚ?i-r��\C�E�A��pw�<�Gy����Hp6��q|�����������?�;����wryy���\^`]J�ku*��{œ6�`.�O���p'mL{��H ���,��6�gk�t� e��	;��|���|����[6�s�m(�Sr��v�\�K�8 
����A���2�i휲y���/�������PG���7H�_�ƞUp>��ۊo��z��Ί)TR��0{�T�DB�6����M\p�3�>^��������,�n�8kH���4Y� =�nF�~ϊ�Ѷ.kΝ6*�cT��&���|E���>fk��S��ٲk�#q��m����`����08<Hmw]�%�����Q���=h�xȟ����oN�(�/	v�OUa7�>'^�sc�U[���.�����j�����r�t�R;]��]ڿՖhjiA�p�(c35�l�>�ԛg�k��z�<,���mo�+E�9tov��ǇG��]�l��&�p�rr����Vq�QN=�k�8�R��`�,4�X?�Bc!����l��h�;<D�p�x6M+��%xf�~�Lu�)�2 �+p�1a��`����\��Re�6�����C	1�JҗrvN�Ҋ8�(l�,��|�gF�^���*_<�Ϊ�&�b:�T$���ߤ�ׄq��>�|�)�������6է4��An%�[��	-3"n��c\�^��Q�ˍ̐��s�H��\Jl��F,s��J��V����0�+�v �uqv&W�_�F|J�5��NoT�
�mK��%��������}t|�9˛e!f��լ�8�1��R���b�v9��S�K9<:���Wl��v�25iMϭ�`���33�~�|Hōe(y����]wke��} �W��77o��yRjb�<:�V��;Mo̫[$����AnE����+� x�������_�Z�����q�y�V�Կ�|:���s k��
""���gۭ�z�J�'' >��e��	��e��M������kn�H7Cߍ��͛7{�Я��h��å�/d�i4�1�&Y �'�wL�]���[����>�P�q$�<��L�B���/�a�|\XJ��L�}A�W�@6m�Ih��њ�_�����aw�9�.�R�2�"]�����~膱?mr�5Ɔ�Mi$|��.��6P���iu���:J�G��t,\/�0G���3Dl�x��6��v�t�]�i�6)N��Yp�L3�+c�0�v��)�ۓ����y̫���x��Z
	@np�훱�.��Zd�9|�����u���=mh��`�Kȿ=?��\,�"nc�{B��Փ�{M{-��m�����m���s��^��J��!%xE\5�kU(,B>W��pX��G��������"o<�!F�..���*�ǹ����DU�L�V��11n�h,�*M$���|f7��|&��lȎ�멼�>mm� �@<N��;�R�9��ܼl�C� ⁌:=-������B#��+p���J�@�J���Fs^}���t,�h����	 {Y���hD=�l��&?�Uj�x!P2t�(�jBI�59G�-� ��uX����N�7������?Lzm�di@�L�
��~��?Ƭ��'����m��)�S�$�K$��oc��z�0ڏ�7	t�E��T�.�� @�����f���$�-Q�Sn,h4�  ��IDAT��|�,�ʹ��p�ޛ��	�M.J�ZL�%Ʋ ����fi��J�`���I�԰�����N���1H\Q5}�@��
Y��-���6�Hŗ�pa�����Pf��N��P���ô!j ����])7����?8:�O߄�H���R�M�7;3�wҘ���@H?'��wp����״�~����t�ư� �&�z) l�"[��{�T�:y�vY��;Ӕ����z��a���k�%p�����}RH0¢ykܣ���W�vDI�WX��5��h�)t~��T;���_e�*|�������ұ2iH�5!���zco��%+ڏR���9X�T��q�JX�Zv�짵)Y[t
�ӊFt<���<[M��������:L�K�Q�����^?��p�q< 0�㩥�q�+Kca����p��ۯ�2R�X�q Lr����i�u����G�o�1��WaM׼��Q0�Jڠ�����D�%n[J�X�׆9z���0��Ã}�ĵ�$��d{�[B�9��L�@�DU�n��j�\*�@�4B	n-�1:�e�̧Y:G�:�����7O���/�o]�S��DΆV ��n�\f��o��$9�ͭF� �a�H��>��{g����Na���C���64�[I��S�E������H�/`��zhG�&h�]�z�{�y2غшi[EH�5X�c,��`b��9�W@W���c��GW�ʃB��_��l��I���uTܖ.w�R�'�:z����{4ZϾ;C$��-?�F���LRe�#��b���h�����|!��'�ԝ��Ǟl���Ͷ!���Q`dC��yC>7���j
JΕ�1�
I�����X��(w�����;9??M��:�{������g(���ѤvW[�+�˰���K���6&Y�re�DeF��A��P�$ý�\3́� \�٣��x~������ۗ��oe��Dv�5*0h*EI��`��{g=Va�P�٦Hk]��C��u�,��A$`���9�Wo��C2d_�����I��a�D���s�|=x�hM����ps)���Ҧ�Q��8�/D�����k�Xhj��B4�eQ����Ac��"����7C�Vv����d!�ux ����)X�ô]F����׹��|�>���^�hT��ߩ`.J�n[I�J����2?�����sr����kR3����SuFLF�*��;miƔ����D�C�mV~�ꭟ�F+�"S���SC 3��oI��j��E��Q6dB�������,����F������`	`�:�l�{O!#�(Art犈~η��|�}�������i'�ο��{�M�����{�aH�EE�d._N�������\^^ѡh�������Q4P
�e�]� a�Ru	��!���nb �<N����w��^ЖF�\����������^5�<E�Y�!ϑ����[��W����{K9��G����uk>���#�El�kM��0+B������� ��ѫ&ُ�Q���mr��iJ`x�#���Є;�8c�r�����$�s�^��9�v��yd5.�P�#`�N��M�`l� �):�$U�l;h2�q�/�F7q�<�Sk�K�6t.�I� 6��z�����T?�����\�0VA��1޿��X���S�8���~�[Q���H+'%hՏ�d��I�_W��ʇ�ۑx���<n՟�?eWbn�`���J3�0lr qMȽ�r>�&]�Q��T��(1=WKq�76 �<����F�N?�gZ�>TDUvv�_0��V'�B���fs��E) Q�ܽ�魚G��Dc�(�^S����7��w�\���:���-������wHy���:&��;��e�g���-.��"�Q�2�07>��Gӡ�N��8Zw5Fb�1�b��}�W�+r�ZT+��3�p@@XxkKuW�!�XC��3�e�ctTGbs\,�:�*MK�xB��� � <���z���΢�u�ڴʴ���%Fo,J-,O�`��;EJZm��q�1/�\2���� �g�����Y���P|=�5vq�(@����|~9���U-���:G!����M{-UG��9��ŷ&�^+O��N$x^7���aPaݠ�8]lI�����D	� ]�y���GyD*s�dQ�����xd� �`79{����v�im ۆ�% ��0
-�]�,�O���s������Ś]�2[�ϥ4/nl�±Aۦ�/���_~_#�9*}�_���Nkٰ�}/ ~lyK�܁!���k��ibV�&'k�i��EY�����}�v*��I��5��O�M#��3W�����o6[�)	������U�����t����|�ɶ>Z\����T�zt<2U/�q���`�nb�_FK�cH'Q/��HcB�J�Țq~�eSc�kπ��K>�F���c�j�W�YL8zw���؃q6y6j�˙�Hm5<�h=g� �&���K��p�s^Ԉke���7/���tS&�i2���<ۂ:��k�&�O�ϲ��Ԡg�88 ���˱O��wx��R3
�4�?_R0h:Bܒt��߱p��zq�I޿�^��������Dɫ�����>�ot�KNJ��ǻ��k��,�	����i$1hA ":q���
ӹh��{����ϟ>�M� ���'�{x@YTϪ��m�����1�K;	�__�Ia��w�3�afE�8�����AY[*be�Y%$�Z*�7��cL`�Av��o��d�R��㒆g9[jE�tMc���l�UB^����a� p� ��&w��J������U�]4p=�AI�(�"mЁ?#�\�Z���iW�-C�8}k}�;iCq?�)�P��6���g?�c���.�r���BI�ե�/{�m(�R���l���j�d#�ٴ6P)�M!�Kr��r���[�����=X��)ӎDu�xq�}�0�noy����\��QYG�p�V{�<z҇��5�&L?�����ݝ�-�8??���V�{�GyHl�1��'��q6����� y?N�yN Fčk 0��\5��UT��f��1x���x�Nu���z,1fl��1���.ڂˣHR9�R �4�r��1L�|/p��W��3S�s�"��i�5N����rp'lWםA}����ٜ��z��@[v�1����2�
t�����MZ��Nkb�����k�	Z��Z�vl61;D~�ڳ� y����{�F�<sS�g��Ojk�%�4��Y�I���d3;D1��T{�3^��?�ើ��, �R�{zYΆ`����GPn�d~
x�ߺ������B�|�b6�������I�(� ��A�ڍ����={���/FN9"�R�L���yWM�'Hވ\֡q��ӎͳ�����kˠ�<�]���g9��I.�|�go�{ ����� e���F-h0ݡ�np	�S�'ϥ,2�ʱM�=	x�}"ɽK�Ǥ�ռ��Ŕ-k T8\$냻�ɴs���>8Ysk��<7���ѻ��<�PF/�9���F,��4v߶�R�;�DC2 �_#Ճ������J�ÆE)p 
pFV|>�?tAl�3������f�^���Z��A����Z*H�"��>��qǔ��n���s�XY!�XLcz���G�ֹ�Pm�]���H}o�����Q/v���[�Qǻc����[��}���}�ȿ�1s�m|�o�1�u�����_�:A�Z��e�xjM[0�2�l��q|���ZrY��y���#�Ţ@8DN���ye�nިXź�����}�+^�`mWuـ�.����L�k����G�P�&��1�Nh����9�D{�֌��
#p��:B{���K�N� � �¸���t���O2��(���`4C��D�F+
�BK�"� �b�g9V��Z���jN�l�˞�{
�n�W:������j���V�t&Qō��ʬ= R��T^#�a�WF�6np��C9�}��R��#�+�A��I���+n���z�8�NP�M�f����m�2T���WU����5�U5J'D�j�\���wMi��L��+[���a��sR$�.�?�Fe^��_�3|������Ww@��0�a`���9��V�)�~�����kt��㨏�'Re���s��7�r���/~�˯�3��k��,9
��o5/ P����G�H�3/J(��RG�~����@��%#���ݵ\^����?P�mVf�8�k��!�8�pᤳ�E�Rk]�����h<ep�e����?_����W�ظ���"��6�fp����/_�r/�?�gE+�փ���f�YU�U�X��<bQ&{����>�����k�dċ��`��%�H���1ڀ���3GZ�0
a��eN����.��t�Ua{{��x����	�.��V�:DǮ�n�D�<H.�F�'2���Ann�3��>Ru��o��-�]^\�Z�ãD��*���Bd�3����L�S�<g��Wʋ�yf��\�:0�
��mKu���s��<�ݠ�m�~�M�"X��F-X]۸�`���)����%��FK� �0���n#�(���'�@T'��Qr�,%��$x:X+(��8�^�\I],Y؁����tӜ���_(��ϛ��F ���mM�"[�1�3��9�	\*)qN f�<�������\ruy���er0y��1��#� �Ohz$߳rQ�}�=���\���b�k�؞�?��Y�"�u�K�u���5����o������Wξs��S	�+K;�߰.�����d@uj�N�7���v�&�ݬ"d>�<��q[=��`F��H3��d:ם䔣  ��ҫ�3���J�%3ֱZ�F&sU��6���F�#av��0�a��BY�8�>f0�E<J���33�L��A�X;z�E���N��˞RFo���������������ҡ��v����3/���~�KHj����k����|�7$�1��X�v��*G5��Je���	�y9����Ԙ�[�C^_q/��n�ע;/�FI�ݚ�3��c�<Fy�U���ԉ���򁑯˳��%y�g���  ��z	x��`�TPW��2?Jz� �r.��[T��ȻȂ.����H)3�b�]m�Ug����A*�x��;�l����ne?�	�[-���D��U�Y��2��7^�ٔ{߲�A�� G`���M�N���zM�||�S]U,|�@�?R5� GF)noo�2m0���4~��7���������K��@��&�dl����rH�������d���Znot���ݻ4?>3B�{�6el���@�%	�"LMb�U�,�u�� �	�NҳJ�p�4��@>Ј:���ࠎ������_r���k'��Z��I�,��W�FH��6Eyd�UY�ʎ��yS�᳂ ���2�WZw�ZE lH`��y,1�p�@��}B�c��E��������W�$�~}��v��r��5:���R�P�L�-�T�~�&Z���4���*����I����eMЂ���v]��^� �4��ۏ��s�}#.�;�����b�� ��`z��A�ǵ���)�P���fw}�w�z��� ��{7�T����Jc Ȱ ū\�4(p�[�P��Q6?!5���6D��G�#��Gh1���7[5�X5�r`�4�z�whKw�O�K?���l�������̙*�������D6"I���^)���9�F�U�VJ�K�/�⠕�^�8)S��E��BH?�QR�~���RJ������}�)�aWD��z�VX_��o@�
����܈��t�?�ؖ��LGQ�|�u��ч7�ּ��B4�O���kkmղ��"5u���((�pP�|S,Κ����u�%��7W����{9G���Ҫ޶���@^}���U���~��5 d��r�Fr*#�*���q�9<pӗ�i��7z=� ZMM������:;�F��$l����E���\���^NO?'��Guh��{��}�����S�b��k��Qu�]R�����XġZT��A�&�<�]S��d�A�:���Ǒ<,~Gô	�x�EK���c��)b�����c����Z~���	��܃V�1�tA�?�/hq<�\�	��ɻ�?�I� `�$��������==���>��W��GvM�4� ���Z����������K�E(�LP�`�h�]�D��kn�8�y�Q8���S�Vy4#h�q����Q0DM�B����چ����\�i�����vX_O��|7��B�,,Z�j1�C��>��	� ��,�3�[:�������IO�l�h5��"�֣l!�����T�/.Ҽ�~4�Ua��:|K�+����.([�Э5Z�D�Q�!E�;� �	�OhM�uy��D~.�N5�HHkz=h#�[!��f�&�R��ȶ��h C�r��A��-�	�V�>{�Dє<��A���>�/�Ӥ`ws��a�L;����#_=��93
YfE#F��ʅ0��Å6mm�+ �s7���ϻ�-��"�W@���z�nc.���Am�G���'�����P).�����E���*Q��5h�H����ґRMpq�Mo1�נ6ծ��U�7sj��v��Z��k��(��N5����areuLE n�c=����i�0�E��Wo����a�x\���Ni�xO<(Q�� y�������ϛԧ����Xh:o�t]���d����U�ih8X�?l�8xn(���3����^P�@�����^�$ש�$�T@K7��LϸAH~.W��������.������D����ձ�l��)4��\���_S&�ߡ|6ͳ��^T��ܨ6nD���P�͘�SΡ:�y�[i���f7��~v�6�d�|�����I�C���������	�5J���%nL�h:tM9]�����g�*�sSK���E�_��������2��˗FipM��Z���y@�1=��>WB�sZ��4}��#�,7�e���Jk�'9zMRw`$�ѕ�y���H�'�%�
��G�8�#%�U�-��ks�NV�<@xB `���L焧�2�^�[yğ�{y�]�8�Z���u�p'B�9�G��̓����z�
(��BY�(1���(� ��Jc=ee�Z��/h��F�Cv5�b�{�:�����HǺ���8#��6���;�2�&�U*p!R�>� g G8TK�~9�mj�1}g"\g
 �5��b�#�}�b�k����l��I�6��4'oXCW�!ZŬ[c]Ц�V���"�3�Y�KrAͩ��^X�Uن,	*��s��H��J~ƈ�V��[&����h��i7U��Q��;����{$#�
uĨNu��c�QNկx�:���|;�wA����MH��C�kagO�s�
��,��{���X�a����~PE�<���F�}�c�/���J�L5j�(nz�(����rq/��s?���>Д*�P�8ss���L���q��&��5 Wm@�w�`dǍ���T��~�C7�8�ߞ����E�w�VV�ݛdC}�G�VfA��R^c~���%?��\�LgU�s���r�1V@�Ȟq�3�z0��=�o����/�a��������͕�k��ە�ׯ�_KEyMEՔ��i0r�G�B��Q�6��@���MΧ���&��WӘ����ǈ1������O(L�>���Z�9!��H�lQJ��O~��?�����͍2��o�9�Q@M7����ɏZ�yVc��5�b���Iϵ��U"� h0o��1mN������#�K���H��-��ӈ��\��ѯɏ�Rg"��ȷm��[ !�u�6H�F�'p��xG�Γ�^ DG�)E0���)ثb�b�P�WNb�L��w -�"����<����޷9����lI5O,��$�I�Q)s�?T�N��R=@3���'���Q�c��e�"��JF���r�0s/��rz�M�	���Z������t�T �퍁_�n<�q���#m�� �1��v� �Y`h�N��t�{�{���_�׿�6�\yO�9^L�߽{O��wქ>{v�h��@ܧ����e���Ks���IW���r�4Z�@��9I�-��2:8f�A�ihd��&�;��(=��ٙ�����S$SL`o!9A����ɅE�k�a7�:ӈT��3i���ݘ�5*G\�U?V�&^�����IP�2��|G��z��B�(�:=�$��k�@Ӷ��Te����~gv���Y'��_�ͺ��΃�����lɑn���Kߨ=mڵE�/s�����������`��t�ԩ�ޚ����^Wz��+��L�&�tY3-o�yO��s���]�}��&nD9���3\̺*��K`kE�#c�����ަ���B7�V#e�`m,C��z���Pun*�ŀ���Bh:Z
R���3<�4���V�H���Dշ����y��mF(���׏L5^�N�4ثd�V�X�^���^'�u(��7h���l��rS��Pn��{X�_�@�����dfWޭ�D`�{4e]4� ���U:� G�iS�M�~&{�;��Y&К���]}�O�n|5z����\k9�-�l%,E����#�:���-�Ǯ��t�=��� E��%7d�(�]�!Z2%L�Y��Mu~k����ն��@�gP5th�M4��?�[����U��_�����ki���'ֻN�B�,څk�+G ��^�*o��VM}�� �f��z�����CԠ�~o(�^3Y�����s��>d�ѣ$�{��W�Xے��oo�ɓ����V��^\�����9�+7	,a^�i���5�c��\_�0B��G��s�H�W}0��I&�������v:@
����ݣ��"�s��~y~Ţ����O ��M���կ�|������p�]ؘ����L>�48x�#�9�c�>,��*m� �ﾾK�y���q�m���ą���i����4x�����@�>l�����t`P|���{����ת������ĪRv�U��"��N��<����3��ʑ��|]���o!/�V<��c��>9��h<:�4�z��^1��6P;s�]���
&����R�ZA�/��Yr�~�f*0T�'.YS�@ا4��%d��M����wl�%��yl�&jԶ�(����9K�0�j@\����i<Έ�*��,�Ѵd��Տ8�{��~hե��!�PI\gq�y�zЇ��$����o�5�{j�1�"|k)��ʧWhဦ���)�et�
�25)B���` b��."s���c��O�կ����/�E3tAj�keO� �����V�F����ͱ�
ݩ[V�8���m���'��r�����`����9���;�m���_��W�-��H���<�q���GKļ�q,����}e��쐾��[�=����}p�%��֡gٷ�t$�/W�qs���;nj�mMϰ��zK Uw�H��u�|���C�ǒ"��D��deEd����H�hJ���~������L�u�0��_΍�z�y��hB�W�7�?��/is\�7��U�=XHt�
��B􊕤�ZJ�d?�_��k9>�c۩�ل�h��h��QY�>0�Ҵ�g��5�����*c���7�Ƙ��BU����fYe����p�Y6�c����lz��,oQ����(Y��u�����3a�X�"#��4�''G����LI���\{�ܝ����/)C��Q́y����I<�,�5F�@¼Y�o���6E��U��3��o��
���`�_����g�ַ3ͷ4o���F&�w�[f'TBbIҹ?��9A(&���A�Q
F�`�Ҝ���]z.֑"�g��	|% �Rg��-Y��;� QEt +Bk�ZFCp�6_R#2p��8�rh�̛������m
�WŠW��δ�uR�����I�|^s7G�σ����Q6?Yg�F�N�Vp�� @p@��'Hwԧ��RU�rUQi����YQ�
��x�ސ��G�&M��h˥���.l�c)P��w?|��|*o�>��vO4�T�ST�7̈́�v���V v(�>Rv���z/��R>1��A�����A�G��%�*^��]o��贏Z�	��oi"���:2trОh�H{7�L�-S��U.��#׆H79���1uܢ�m�[x��C�Z�6k`8��~6����P6c&守ML|go���7q�>_-on�o��v>��P�#D�>�9L��%5'�J�!�x����J���>�F	��O(5AΗϨ6d���C�y���|�^Ɵ�9� 5�,Q��z�ζ����C F�5X��߼a�`[��]x9���SF��S����u�,�e��RDJ��HSȄܯ��zC�^�/�nMg����Pߘ@$ˮ�33�-�n �N��6�������.���p�D}=3;����wp ������W�e�ѯ�"�6zVM#l2р��w<��:�(����!�űmTr�<��E: ���c��O����R��lL��u���t�F/t�^���{�ߪ)��$����{�VO�v��N�@�#;�����_q����1P�j�j�{-�o{��ｍ?��QI��X���A�j��YS+�Hm^�_��l�#t�@b6�{oi��E�Ru8!_���g�_d;�c�g�t4����b���/�0������TS�!���F��)�%x�Qu��>k����`/���ڽ�VO�i��߭���v��\���s�s1�����kU`n�߳����g�n��c>e�8��#��z���#K/��~`��o,m%г��{����hε��ͥ��'�NZ3QBs��X���� �c.[]N�e\�c�XСi#H�|٣�\*����a�ނ:�%�C�ث1)5I��ϗj-��?� �U�� ��^۾����j�,>�}�� �FsH�sH�A;d��4�`ϧj�C��$*�n�w��2���ټV�RM��[�imr�4�?�N9\U'vbr�X��;�R���|b5�U���	���-������ɺ87ԗ���|��d�@.};ݱsh��	�z���h=�-M��v���oo.�iǛ�dT�輕Û��	��p���ϱ'?6�����l��?��r:6Y��ydm~�2����*.\�w�����\�O?�"i��N��R���`'R�>2D2��7+��K��f���z�=-�Az��0U���1�v^���$���l�D�փ�Q��0lں���.�m��ٓ���oi;�|���P�~D��=6���T���v�����+�̋����������=�T`#$>m�`�EE%�C�#Y�P���������.��-6�)�`�d�mlr	�g�����~�o?�a������جq<8�c[��zIF���M؞((����Y`��BJ} �l}���}�N&1�-��p���1"=k:�*a��[�c
�`��ܧ�|��T����-��i�=29���	������զ�����[s:�tZinO�I��,z�?��!;h�&��������4�ޘ]�9�]��Z�0�9�{�8������v�K�m�q�@�16"�v�`~�8��sE�S�/�0D竞K0#̶��Lfs9::&``J��@72������pf��^�Ԣڴ6fC��m�� _��M�K��v �k5(ZBD����rp�G��Ez|)�g�5�V�`W�3� C���ES]ױ�w?!REx�G^?�����e��֪l�����,ޔ�3�y.�5���!X�'��>9�i��l�VR��*`���Vz�1��6�ь��hF 4�f��-^11�r3�Q3`��T���	)W�t�HE"L���R"L~�bȣ�c�P��	T���֒�1ڒE+��@S�r课o�F��;G�j�v�*L��C�d �V���<#�	�/ld�9�K~��0m�{E�*�E4w����wϓ�K���lV?nUB����J��E��-��E�쮞đ�===�.���)7�Y2�Z=�V��8^�S}溪{#�rcY1/QO�S�nȇc�=I�=�n��KC�!M�,Tב��:�hO���Ui�}���r�������- �2��<-X̕{e��vf����wҼ�fJ����E
����F�֚Ηaz�L0�����k�2RB��5Z�=��{u��p���3�� ߌ'V� ��#��G��fzh󽵼L��ͮ)�T�E��-m���N�
h���Gz�Á��2��Lx��`YϤ�z�z�7� #��ER�o׺ƙ4������ �#+��>�^|�")=Z���&[���HA�nL�L�G�v��CZ ��M�$�_�9�b�fDJu��X�>�����ھ��a��mz�_���|�8  ���9��25'�2�2સ_�;ݮ���_Ρ��S������s�b,�qf�j��!D��KD���"	M���dke��u`��MI��=���]ʎ`c}c��ҝ�u�"�n��wH����7�����v��H-��b��*��]�J�`��x|#�{;:Vc��Z0=���F�"�:����5i��tDk6ʰO��>/��:,8 ��L��[$�kx���wn�m���|	���
є�Aj4 03�3^p8��[�����'i���ǀ�I�o(2�P�L��7�p0A-YM���%0��n�8�ix�J��V,��=����ap��@����O����V� i�����`i߲Pl��3�|��/<�|��}�ۻ���z|u"��:(��B�6�ya�v�?�
���_O�禷6~M]?w?6~M׌{������8]�1{С�ކ����C��z���a_���hDo�>�5���UpT�a~�" ��8��T����-����U��=�?��@'i��B�mrqw��dO�w�^m�2^82i�wH�`׵&��g;	��7���mٚw�ѠQ0b�[��W&6���#R�4�S��g��ގM �|j�M;-P@!�t��4b�ɡt��gss�T l3:�#2����ɔg>X�۟3��8��f���]�޺���t�dM(����P���s��Nl�u�hsT@���*+c{���V;�s�UU�LvT�
�M(��7��/l]��z�H'{��fM���%6��SL�[��R���c�S�Ϡr�|U��� �9�AS�l:�'�����j����)(�oC�c6c7�Uq�}h��=�\��R��߈Hhz�4�Cd�5
IE���b�e��g��3��/�0#�mac�we/��������'�`�����;���c��-�E�J��ƺ��(l���)�L;��O8�ا�o����㷴i�����Spl�$t���:�XU�&)�4X���xn��s�YhBՇu�,��Qg�p�G�)\TT��H�G��k�0X�MGD��eS��Ф��1ET�[�(2@�?]$���t�+f�|Ev�l�zr�  X� �M���9T�}�'!/ZR� b`�Y��b�&(uO�o��C�dӬ[b�"χʐ�K��x J����i�#��Q����@ ���₨���3��"J�@�#`�Y����N�����A�"�"�P����'�����1��NX�F�F/��ʯ����C�ӄP=�?�8�����ya���1C�F��S���}�����߽���3�M���^�$��G�ޱ�Ft���������/F�/�����ͼ�F��u��F���[:����	���0[6�ޡ�����+ݰ)�ȯQ��#�PО~mc��P������i�RPNB^�QAM�HG���h���V3�IV{���4�	�z:So�����3?c����/�Չ��(�.ӴX����M�X���z�<�\�W��5�A��-�2���q��ê��A�jk�ւ��$Zm��ZNm�9xe�V��}��Z����[˨w�V�H�T��D��|�M��U�N_��X"�2M��d�Lo��� �s��{�f���Ls�\���O�[F����+���
�B=Hs+0���}'׽��Z_�VI���6s�WUY��ㅗ�;`X>���Ǝ& v�y�PќNv`���D�cr>g�]T0o�)v2����J(�ų���X��U��%ߕّ�,�~���"�N�$�@ur�/�i'Zq�B�1�W�s[M����=G��JŶ�v41�M2��F���%.M��GM��(��ך�����ô�!�E&�Q�.Fz�(/��"��h��<j5���X�/��Z3�� 	He�_��x5�7������7�YȘ=	��ƞ�x[	���$4pf	��1�
�۲G�E��!Q������[9,�8;���0(@����ō����V����C�|��7_͙F��!kkA)#���6`P'e!��|��\������~�_�!Q��x�z�3�w�.����ke�/}��)��G� �n��E��6�k�`�Q���W_q�~���dg���o��`kۃ`��nr���O�t��!W�S�g�y�p5�6�y0�3-�	���2� �.�6J�1��4Pɉ��,]��������b�|��]КMF���a��Kt@�NƲ��z��;�k�6�`����od*��sD���{DE��Ž<˹JF�X3sO_>�j|:�O�>�fs$���Ǟ9v�Sq����%�U}�;3�&'�oh�ڊ-�)�����l�-F�<j��l@w��n�O�0(c�^.y:�#��p�3������q�(X��"=�$���� |mM��ԤӪ]-���]�M�3,��U��@}:q�R�V�6��';�
J\3^�Z�J7/�Y4���e��l�A?�����`Oi�4��qaWg/��[Y��s�U ��^V�b���F�st���/�O~�Ν�������2U�2�^	vmTG���S"��ftK@��G>��r{O��:�%&��B�K�������j��L�up;b�R'i]�:����C������O2{�ڤAҊ��0"�(��~�� "yw�����bw
�V�':�g���,ZZ����k>=c��X��cjBޢ�?����۔�#x�r��m\K���C�zx˴Ṱ�P�04��X/1��F��p�V>
ȿ���{me�UJa����×&�[N�iu�
���G��z�P56�"a>�^���aE������?�q�(m.l�|w/?��$����é<<��Yz9nr7�y����A���Z$���y�KV&\��c�ek�����V�"� ��s{���]2{�>h��}�?��zdz�my�uZ�vu��1a��3;::b�b�H"D~~v.�ݣ4.���қ���'gf�R�s��b�ʍ(��~~K�r陖S��
	"]��*�COi���
�ʜ�œ �ø���1��luis��Tt���I��ND{"�mm�������c����(��	�� 	��QJ���>��c�5Ut���_���-���Tȷ4���OU��	9��D�uY�/l\?�ȑ���Y��rdJ�dx�]��">Y&���⛣�UoK#��0�� �X-	�����q���p2&�FLEJ����w6���#�Jn��EN�?7�r�W������#�h]�!+ˋ�<݉��E)�����j	��_Y�J�@�=3KT`G�"�T�`�6ΕW"�k�	�&J��6@t������`v��T���3��n�UE[�ϳ�&)��K�
�c���431�E6>��j������#���������坦��oo�k��%'�#���P�t�[�aݧ�s$��ߤ!H: �cU�gH�ݢ�>|�<��٥Y<L��b���`jOwQN5+�Qոr�:��:�X��D�Ggu^��	��o;l��AqjC����$��ӱ9.�R=�d�p�w���)��&G�CI��iXsC��m�96��A�NNg��(�:��i�x�OPa�:(/�|-�=97ð�E���8*�(�T͛��k��x3ڊKa��VD��\��ޥj*u4h��-xV�q��_�o~�;���� >�������zӫQcX @��.��z�{IJ������^�K��%��P����kyu��t�Ts'|F���lp�\�wk��ss!n���Vl>���͏�fXc��K3>��LQrO?���Xt|�o��V�$���'D(�O����>������}���W|ᕘ=#O봱4�� I�=7�ζ���<���+��iYS�뢱qPw�{�Q���~AO���!�MiPz� @󿔡�F���)���-��m��..��ǫ�Y��
��i. "�Mb�����6�:��?K��l���V��њ4�̩ZY����<���)Ą�Jץ�7�7��oZ7�G����Ҫ��ɟ���k�k����Bn�4����.�$В�f�Fv�@�3'4dV�%� �b:U�K�$���a��~uq	��/-bP�i ��"�AM0^";xvF�<�=ҳ���ݥ���Mx.���n�;u����B�5�8Ɉ臞���T5*/��=[MbqÄ�e�RD��Ŧ��u֔S�|Pe���'�&��ޑ��9�@A����"DT0���t��9�"��)�9�6�ky_Mk��y�	�W���!�I��k��6�� O�l���������[���؜
���Xt-J���3�e�z�Ec ��1( �-�f��YI�g��/���<}����٥�����|���l�xߜs��Z�8�^��nÖ���4��U�z���vk�ݟ��8���d����։&��ch��W�;W����n�#Ah�He��K{^���Ń饄�1�(ߠ�
�v�^��y�X��W�d�5tL��hQ$�({F~4�VH���������R7]��!;?X_�>�Fx��oY�}�.+��j���"��ѿ���������"Ip�h���ڱ�䜘ڰ�!�`��T���^_1
 5��������r�r:�{���`��0�~���c�z
�6#_/q�<E�c��Wv����
Tc-�d��F,2�0/�����p� ��4���utY�w���WF3���b�ʸ^��PgFD@DK�=�'�����ե|B3�V5jD��>�ֶ�u�����4i��{��[(�/Lv�����L�sM��t�B��h�����,�y��$ �j	���Ed�:^���'X�������ImZ�M��hO��m�y��I���k��>�#]ߗ2K���an�#��x������=�P������WΪ��b�%
F��(8���"�,�J;�@�-%�c��{  �Y3t]���C�)��EO�M1�0�=�q��6Zv2�(`�3���d� 64Z'���w�~�`�Z*b{o�⑱,Ni�Hh�����F���[Q�4PRXm�~EOS�M�|�@�Xa<��	v����1�odiܼ�Q��QF��µ���i;��ټ�H\qݐՓף�qs��㳿������S4���S	��������=yؾO������-d>_1��JW�����M�\y�����P�v2< �+p%W�����2H=&;�6����F��?D?PR�����+p(;�H���ݩ�VLC��A qn[|������",MŚ�]��n�e���)�A�A @�H|=�;x"3��.$x�0�C҃��d>��o)9ꪬ�&��~J�ae���U���_��)�
IGF_H�DC`D}�����X(	Tw��Ua(��nM���"�Tx�P�M)\��ɿ��o�7��A�����`*׆�S��!�����±���|E9��щdT1��Eda���q̶wD`�;�-��������~i�^6�g�*��?y_��X
i�̓e�m=<<b��i�t��ig;��ZCu�B�-Nq�D7�f����J|ª�	\���"9өj���* ��������{���0�X��!"Mʹ�J{�yD��Uj���h�����U����+]�h����w?����"��h/�I�`�55�:|0P�GGLۣ��ָ0xmk����ܸ^��w�v��k��v�k�T��1��+�,�߳��ד�i��|B�cy֙��E7ia��6y�0�o(�T�n���5�d�� �.�Qm�4�F�ڼ|Q`ww/��k9�@ �"7�[c@`0�r��_]]SU\X��oQ]����T���=�" ���Z�GӨ�Q���D�d���@��:�#Ae�B��|v��w�+��d�&��\���E���{�y���UTd"���9Ȉ@_Zv���\Cd��m��qе�S�M޵�[��6f�(nB4A[մc�oFMK1�v7��ۖ�����ʁ����O���������}`���Qoui?��ٗ��#���7��y��!�:�y��C��	m��YD-�P}��b�&h������{>P���ŕ�%�۴��I���^���߲J~gwN� �M8�9��՟� ��QZ���`Lx�pt���$I��+��i,���S�[�i�YaB�|Ӌ�jS[�؞g�S�{�����߽c�������F��\_ʂ��5�`P��0���֬�q!�`%��M��/s��zo�ڰ<�J��plp/Fɔ����+�U�U��Ս�vE�p�1�AW�\<Ԥon������iP>%CwOÄ4&��_ ޺2��o6��=�ͻ@�m���=�_�#��l�Cc>�fp��s�qb�O��U���g9]?�����M9o~��jBrM�Ə�R#i��H��W	A�6��|�P��R����g���5��+T��0�}߻����./o�����r�6��d�P�C�`����OԊ�Ϊ˴x0Ϩ��R�=�Djm����$da*�c��;p͌w�h�e�yؚ�d���Ή�i>I`�h�Ql��W��,	�eʫ$���қһ��
��!Z�<�jJd)WeF�^�9ǩɜ@���׀���Nu�4ˀQ*o]�3�S�`2f��)�sB��V�K��-Ϗ��5���-m���(�988����_͞�;�s�M�����Y�6�nM���u�B�Ix�H���9��%�Q��*��w<��%�s|r��ζ� �ϭq�h���bI��t	T>���BS����㽬�~�x/g�m����/����[����F���q�����<����6��>�ֵ�c�6��Ȣ��r"x��P�����)�)����\�K,�s�����_b	��~�hֽ+���4�fr��(ٵU�����\�+�*Zģjk�хE�b)"�LN�4(%��uح�o=,s�.�TD�Au� ���lªIr�8�
m�Y����s�+VR`��N�	���ʹ�Ql2���f�3�k�6�β�w� }��M�6b��}H?!���6����>���6��j����$�p|t,���L�m��Q傁��3��k��>��rk�h[)j���ȯ[�`�#����HY��"�ؕ�ɨ��VC�ʴ��.V���g����H�=�ĠIih�ڙ��w��`s���}�F��E	�襬���"^\i��!�'0��{�p�m@^0�-�0R�t�oje��xEj��?mI�\sQ�l�=|S�b��x)�����يv|�^�.�n���}G]���
>Y�����|tU�5�MW�M�:(4�h�9}k�#�+|��fΝ\^\�?\8�IZ�f�j���(�
�޹ՠE*��`�ڐWuOnX��D-�˵f���ո���ʢg��7��6��e������3"���ZS�j� 9z�~2]������7��#U�M�����zH�E{���N����1�69��\jA�~�؉2i��و7��s������WF����-�A(�M�-�L����`���8���o~C�+���7x���� A�z �T`߿�w���2٪��=�J���gM�5���͛W��W����ɛW�C�T����|��Q�����d��N�������W"��UҲWC�� �d�->�%�t�#�L��>؝��o��o��[ve���L�����+���x�]hi��DP�W�/m�֣x�W� N
��7;[�༗����6�XA��Z�-G+3�p´
b��'�K�Q�+��Ge3B=W��眹jۘW�G}F����s��C,(t�a�@�� ��h�C�~�2w��,����Qm<�toُ����OA�>��Ê��� :@8���s��91�in��*������˩�� ]B���x��Ǜ7�Ӝܑ	x��%�E_����V��2G�
���*�ԋ�)��#j�����i���Z��N�kU9��ziɾ�k� ����r>vחi!\��F�Hp�fh�LH�]K����ⲍ��-#�Y�q��# �V	X��#N9��{uO��
�j�dȓ�6�*�K	L�~��_�k~>���}����{����Q����C�=�&�ps-��:�&y��bb���칗��}�.�!����8�]4LF���l�D�[b����g��c&��)�:��H�|�#�H�s� ڈ����~�$"���[�r�(aX�`���wc|�er�56"����₥Ö�yXh�xDM���(]��2n���|Y����ж��B5s*yE�Z?���Z��[@(�_'����<��m]�\��%?+�G����)1H 0-�+1|e
�MYS�H��mg�X����%ݧ��%�OY���Ab=���`	b޺^D�5�Q0}�W���ߍ�a֤�M�Uj�b>��s#(�Źca�=���O�9>�H�
�6�	 ��7�ț�o��i�+��v�f�5�����GeQ��aKs��I�s�;D��e�{��x�^QA���c�88y D �g�������hP���[��W���5{�e�"ͱ]F��vE�	>M繟���O�v��F�V���"���3����L��$����%��5�0�VX��d
���Ǡ�<|#tGױ�V晫��`���ך��[Y��1+�R6��h������g��_�qM���4�8�M��<|�kA8�~$x��S�a�9]�M�ǃ ₻M��Y�&�(�ժ%�@d(��Q����`�l]V�MP�V�Q8���#2������' ���˫����4]Ǵ��F��%sr�@4 &Y�@r˱h\mQ���ޮ��01�.�Aw�G��x J�O��т�����-i�j��z�Hq1U���t��)K�Ռ����,Ň	P6���猷4X��C�9�LR�Ps: �j?'��J��G���k5��HB���}:=���+����/�������R�b)!|-g�Ï�fpk&���I���*닥`��<^I��\�m���k�8B� L6��w��E�X5��lL�x�� ���G��QS�M!���4�/8�u;l� ��p NA�����NM���;?g���c��ńYUfl���b��>i���wiL��Q�㜞�Bn�_��@��&�Rh�Ԣ��ʟJ��*�J�9����X.��@Z@�vN�ݞ�����N����.AX�*�"�y�׵5��N��?� ��	$)!�B���)>�v$w�0iO@�N!��z�Nc^4��e:'jف3�&����Q�f]�J�pv$G�t~(Aڍ��0w�����
����V�s�'&yp]'^�Ɠ��r�T�c�(�@Q�5e7������a�*�u�_�祥�����&f_ lv�[���.���_P(�31hoND&�M���i�W<�^K̺�>;� ��_�ӈr�$7lW�e�����F�@��	O�n:��y`:�����\�}Iϳ��<H��B�t:F� ���vi}�ɑ�uu��&�X6�&�n�QK���u�ɪ�3��醿V�Z��߫&A�~|�p���x�^��_���S4YʯE��P��r�)�M����91-��R�{O�K� ��ҝVy�����I�s�^f4	+ p鳮]'�+��xHN P�l��:U^9�L�a[$�6ܡZ�BN�.������&N���g����t�A�e;'-��O�$-����/z4I�4�/P�L:�P���ƺv�<b1ϷƜd;���
q��D6�z�V�����<���Z�&@ȍHU��M���MOqp�00F�L��|>E��H�_[�Z\��ڷ��y	�tW��hm3zy\�H�����ϧ�ÇO	|]�P(
��9�� "��4Y��m�h#۴Y����	e��lxg��MrҨF��Le=��s� �no+��:������u��|�ά�̦�_�xn��|D�FM�H��9�V��X�w���vI�E���5kJK)��iv�l&F�Q�R�ȖE�F��f��!��N�׶εu�ݯ���L(x@D�a{�����eh���o
���6�hh岆�K_�f��������4��bD���T����#yu|Ȓ�I��f�6�=DŶ����__�=�{Ͼ|���f\�珹6�+_&�g	�`@�6�A�Z�ח9��۸`�f����Y ����$��V�G$��lө�W��Gy������v^�H�����3_q�\'n����S#���X>I�QG��������0� L�Y�gӉ	�*��{ў'{�7a��E؁��<�\��y6��C�E��<(����\]_�zrb�>��o�za���~ݦ���M5��`�|�S��	%uVv'Gi����~��i�n�Ö�%��5��H���l`�ZD�;?4��<?bw�hk�NT
�Z���m����5���Q��3��J����apsH��v�zN�/�0���AS�W�XM��}�s� �}K�$�2�������OhJ��0(X�t�X� �g(,ːhFL�V�8Q�է�!�X���#S�HhN�^t��*R�2�;F ���65{�m@��E�쓚���7g����h'���jHo$����I��$8��Q	T��%�Y.�'4��5!�\���Y�_&�j��T9I�q$h��x!�9��6��,�`zu֠x��~G� ��?Ҡ�/Tb`ݥN�z�������'���\�\���K�Sӆ������LH�Z�D֍�F�N#�]�2��[S�(>!�(�aȆ)�����,�/���r�-n~��ʛ'njS9�e��^恸^��������v������ǭ��<1����|��*��Ť������|�
̍Fb��Z�y���bɨ*�N��X�;�����B޿�6��8�\8k��7̿��ñƨ/~�M��᫻t��@�ف|�4ӷ_˯�yK"��ř����x�&{��D�z��i/ș ���`WN����}�����4u�>g	V
�H�;;��m+���n����@9!�פ��b�lQ��y�e�B���0X`�8+�g�r�4-� ���;���L9tdQ�3��3��b�-d��g�Q���z��������.�����sY	���0=e�k{k.}����\�hn��������'���a��=/� �шtLD���nX� ���hQ����WuA�V���C.�ױ�	� ���}�M�K�	�O 5��[��n��'r���хn!"T8绛k���#5�X��} j�PϿ����"�ɞ��J�uwJ 	�9D���̶ b+F�ǭ�	�G5��4��/����0!so�=��w��*�Y�A���l�����ص���!?=����6��l���{�TTc��:����|��%ZD0���(����<��������e�_���^�l����x�#��K�� ���Yz�`۲JBv�,��m�5�1E��'.S�?M�.�+��A��w�NT��F����z��
yE�!Ʈ����	�r�5jk?[-��9D�pj�� `&���@e8 $b��a�'�߽�k-��_}�>h���a�ĖꅭՓ�V��Π>�NȐ�L�d��Py�^j?`jc�f�4�4��F+`G��A�3!'p�ԍ <�{�h������0� 1 ݋�@І�Q	ɮ�S�B砗O�j�kpW�id�Խ���H�%h���wDfV��=+]���1���##�"�U�g�~_��`k頻��N���̪�A��I0ء��z
+�J�.��l<JD�eن�R`�E�A���K ��*x2������ &�>�:
�u���jP^�0#��f�0�$�[SP�8qš�_u=x�M�˴��W�'[�b;q�j� �~���J۰R�<�h�,��������,��y�p��oW*�������i���]�ʨ��؇*��iLO�w�����ﾎ@�dˡ|��E���e�˛��"��qӨ]�Da�ۈǼ�8c��--�G�th'�����J�Y�nF^,}�I��؛M[U�s����$�X!o�<J�0�0��h�+ܙNC�;q`t*mj�Qzx�٩���ק���ηd�:(#��iZѼl�XX:gw���H��a��k2�gX��Z�T�;j�"F��~zr�~�ղr�Y��=�Y�V2cX+0�6¬a,����Ժ�N�Г���%�p˲3��s���J&H���c	�N��E��$��2X�{��3�h��$,�T��,J]�\��������BBI�V�m��$��ZK��x�,
�ʗ�ߙP��-�,#/��J{��ޅBT��;�Ng}(?�p:���Ϡ��Wa���aͪt?�Ƀ8�|�|2��H�rgV�X����&��W��ĵW<�e����~ǉ;�
�R3T]���"�{�� ް�0��5.[]���nnM~S��}��}=)(�Ͳ�f!�\��~v�%~�Zß�8Q
k�K
f%S���p"Ta��(�� ��0�_͇��lʒ/X�<,(0��hX8���E��w���k�~A@y��I
���)p�j�f9	Eƕ���N���+0�v�R�� 1�5���v��ų#���m�3��H�k�|��J��6�,8yf	h�Iq1eC�.ⴖl���}K�}�9�p��r������)��o~���eK{�K|�Ĺ8-}"5�<�WB]^��Q$�]�V�����j���H�hjZ������7�c������=y|7���ߋsf��������^����p�����N������/���wv��WUV
�1�ο����?�_����ޞ2(����=}�'����`?���z�[� YD���'��"x;9=�`o�^aQ�x�U0�P��cR��kj@�� s�S%B�sL�V�`}�i��Ȩ2
U�(	d��aN���6ႅg���3'VuX��[jѼU%�!��
��{[R�3�U�%��VK�@S�e��E$V�[e�7M��X"����Q����=�o1 X]��72��l4�%	�0���Mk�Ɩ�*I����ɝ`�<y�~A����+>�s6��.l� �,�qMR�ͽ��"�G���q�q��.at	i�F�Q�IJ��Pp � .�i|-����X�J͘kI����Bad�u	��������D��-}n
z��1��>˒a�c�m��*K��1a�~�?�HM���栖)S�n?�❖q�ʓ��J�m��.)d���F�Z��i⌆<��5K�)$�P�������Yo����3&��S��D���(��[��7�2wV
�&�xu�%?�^�7Ӹ�ڧ�fV�I��gY��B䮚�y-�`%���֠@��mZ�V˨?>�B�V  ��|ş4)�%4
.�>�����<�s��K`#C���4M����+)��& 8���Ɵ.ܮ��3���:���_i���.5�BZ̪{�p��6o�I�:{��qN�QӉ�9�����X���*8��
^�A���#$�O[�Z�;�.Ċ�����Ԛ�Ak-`�u��u6�� ���
��ieBJ��33���]��~9��vIK�y^�M�}D� �]���MԶ|�����W���̶��޹��tIy�]��R�?�3�"���������g��N�}����qͶlo�I�p$](&�J���L1?9[I���K,DF�<�Pid�sZ��J��wt�� T �BVH��69��H0W-�w>Y��rP��u�lT�*u�Qp�Z��,;��	�DnBq�����*Ȅ��J��)��^op���`|%X]�7�t�z?�,qo����[��X�X��"dذvM�w�J~���ďD��N�X)8�_c��^ijV�s���c�èP`������,����$/U�X*�[`#�1ԯM��T6�e|o*1�tv�ć,�JW�CH}-��r�T�0yoځd˧��;w�g9hwD�lЃ,�O9�i� L���,2��}�kk���wo'��ȴ}}`,+(�0)�݉8Oe���xp�,Cl�5�ܯ��$��ߵYe0�ij�%v6hB�}�Żx��f�I�I�6�<GK��C�0����|����r]��vdO�P��b�2�ҫXVu��}�D3����*^u������K�sK�"0k��i��������N�l�� }�Įm ��WZXb9	k�c���O7O<?�7o��A|�r��H�/��gSG�1ގ�d���L��i�0�PnN���J�Q(,d�{!h�PǍYu���*��s����b�X�^�ַ� f��>&��x�Y��>K�K)��g�tb.Bf��fdE>|���)��2�?�p;bl|�V��ٙ��	�M�;S����n���X�d��s�C\؄�+c��3�f�R��ڵ=Af�X�T�6��kݐ�h����:܃5��:x(لk`��7a���آ @������#� `H؟�ENמRN�u�( ���aQ�bcC�Jx�$��:�Fu@	�@2kH|�uZɊ��i�p�v+	@��hR���9��@�8�f�I�!b� �H�c�Yǈ_:�p�泙D�' ��������dyG0���|ā{vvFVz�AW��| ��w�(3F��2lE����H���
�t�s�nP�Pc
	XΞ?{�?Fy����ymp	�bm�rV}ԖM��\W�D�]�z�Z�<C��"C�"@4sHn� ���Sƃ]D��V_ ����� K9��6&���Qv�Zr�¢S�4c���>+��]\�5װq
�	�qϥ�J���u#�j@�l캤-�)Y1�
�� ��@(��pmV�,�{�����ɤ'ٰS[U�JˑO�&ʛ��4&N�������\�7��(��B�
Q��"�o+Z�;�B(�r�e��+�2�X�]�0OVR
E1�,N��^GP�{sOf|Ǥ�L&��"�Bv�r7�B�A�?@�S\(���;._���%����1*�G ��%�j[)iq��$���okZb:t��UC� W�?��cy`3J��"g�^ X�N�5
�Iy��/&W����F!�o&��	���4�\�;�C]�)�b��º�"�c�����е�~J�링���5U��Y/T��YG��J�z��' ��ﶽ�Ŧ'�3��*
�E���.�0kYd��o��r/��u���Ȼ����ѣ=j��;�pM��O�*�Ui�x?���ۉn/yV��RN<]�ԢqTZ;�ې�~{����$��B��0[ְi�BB[yW%RZ�u֢� x��V��U���\YIiY�pA���n]F���C�J�����ҒBf3H�9��-AZ��:�5̈́(����ѱ;��ӓS�2n ��!�Yg��6�%�4i�4Oz��z���{_�� ���������N^����wwo���q�|�e����q~�r#!?�V�mĽ�}
��߹��Kj̤�I<��^��Ab���0��q���B��p�f�:u	�ʻ�b�B7tی{a�	�i� ����n�[��k���Ҁ+�:X6N9�J�d����r��-VwJ�(�o�����cx� k�D��֥�����y|LH�+�m?�HSا�*�M��@��b�M��ˁI�P6p��B����F�C�E-a���<�{]�$�+������J~Z(�:��2[;�&��
!*o38_����kU����0�$�	 �F_��H���Sz#F�+H�)f
�00s��hD���-�x��b���|\L�ҷq�n�F�X���*��@�4&Rg� f�f�H.�dQҁ-�V�ʳ2 3�yZ���]�b�^�`jeBn4�Y7J�>�H:(Da��VH ���L����6��2��!�?iZ��s�`�EqM�I����86[�~��g�ؤ�ɨ����af�Ė�F���S��̮n1w��C0���\~ba!O���N��R*.)��,n�F:�����b���!7OR/���ֈ�V��x9��!�2N�Z�%��k/~6S)e���,
�>�1 ��mʓ��n�ur*x;j�h���H����T�8��.7��D��4�ċC�����l]G vvz�NOOX�}�5���i
\t{�n��+2���'Ɣ�ȽF�g���N(ndp��_�_����[w��Hx��f-B���j����~xD����G������i=.ܟ�����oH���Ŷ��
n⪫�ǎ����a�|�⥖�h��G|�ԝ�����@oN+,X���2��c'��AS�>��Z��Z�-(j?������8��}�H�ȾKP~/VP�S|e��|V�t$3!P��lSX(0��{����(0�h���_���1h0 �YZF�FN�����7�rL���C�/E��ф�A}�;�����C�'�����>���֜ϗ݃=�k���� Q���f�ZY|���(�D�^K5b-1��1<��P�t5���6d4e���T��׽��BI(��~c}�\f-�.3�Wʘ���) teV�[�N�H+�]W��㿈?�(S��a��crQK��纫`�,��^|�nl{��_	�[(y���/"�YP��R@���2雺��� \9���`�6�E��%�UBzq��o�%s��#uc5���~�q-e�J3-4c��T�R"��3~m�-���ɢ�em�<����� ������y���p�ֳK�?���#m�x���;�����-�e;�A�tq�"�`�f�.�ȍ(2h�Q���۹���� �o���Ӯ�V\WR�Ä�ȾxY��Q��Ab��6�R,4���$&���A��m�v}E+D�6�����x��1�!��́*�q*{�1H3n,����A<H�"-ͣV�D��(�@���y^'�wC���9]M�9�z5�.���&�(sG��Cr��>��h2�^�-W���Œu����������w߻��c��B����%��Q�E��7p�	�k�Kl�P���$Ŷ��ZѤNk5��F#�,��G���Z[�W�+;������Y��'��&t��U�xt�?y��>z���S��kק�J���6���J����pk>~�D@p<��v}ǹ����}��Z	����q��/��w+w�<���E�%dnF���5\� L(�v�e�HZ�XQ�+�6d3��,��i}���+�k�Wm&���_˞-@�F��??*R�����Os�����m�D��}6�9m\O+��L�z�.�9���AI��! �8Z��MA��2eHv3g{X�ˠ�Qf"r��@h'�Nb���g����D��^�J]��'�M �*6���Q�	��eP,�A�~���Ҷ�A
:a�	t�1B�9�f)����[r !	-�}�e*���4vx��f����eS2�բ��M/ue�ڰ��Pm����;��^2*�j�� �Z/<L!d����v����x�kJ�+f�]
�]}�Yu��H����.E�l�w~�Qm��ez�ƻ$��ۑ���^��u�M��RHK���څ7��R }��*�0�������p_�˄xd!b�u$�]�+�\L�׼���T�j��A ��i|�sy}CІ�'�#q�Ȝ��׌ �&�� �<�#)�����G�xsv7�+w7�G�����W����	�-�����u�f��&|ta�fpw9?��8��QM6���J#n�7�3wrrL�+�0XN�>D���`�j/�+�Z���l�m��w�y��a}��N�iHj��i�K����ڸ��{�'c{,v?so߼u�F v�28
�=6}Z�i�B��kZ�P��c�:�E8"`P+j���_@tmJ��Kݨ�d<��*='�x�_��+wxx�/���0���nV콃����m�֡���K,��ZJ9Uj2�_��	ٔ����+ܡ ��vB	�Vq,�Lt �������}��ߘ��qÿ����r���˴�V�۸v⼸��u痳8��2~P���a�D�[��x>Z�Z��*�=7^д����^��=�'+����{A�<ÿm��3ܬ83)�a�����0���v����Wt�ɀ�t��$���}!�����ܹ!���83�EJ��Ī�H��w���`��Z~�)��n�R�:QO��%?�%;�Z?�@�06L��*=��{Z�3K�ƍ��1���PY�=�hɯ�MF�`��j=�n=VZ PX `AjQ���u�*�Qq��N������v�Aj���f>���U��5�:�D�)�"��ȗ���:FO��by[ڡ� ��b���>G6�&�4�U��i�a ֮���e��t���)ƥO8�{p����>�E�ک}��L9ȲyX%�uo����>]4�J3ۜOq(L�XJ�C����� ��q�iW2�Y�'n��4�l[�Z.�76t㥻AU��@��Jn(ٺf��׫$�NN�?�!�A�=� ~}�� %r�=�EA���ml��*3�����#�����17��-���� �Q�!7C���6N�ՈD��>�d���^��`� j�����#wA�U�ȶ�j�/,R��R�{�Zh��swv�bT��K
1Y��+M��ړ�������~�r���w���גqxU��)h5P�1�- ���]����u�v�_\0LCOEi3�x�׵OBF?'�XO@ŀxk�ٰ���z㲯Y)֨��ڽ����x�rQȠe�k%5�pm �Y�O ��o:Ƙ-�q��cp�-���h�Ï?) kh����{������^�{�����
y�څ[�Zh?�����ml
µ�@} cQ`PIb�%���2ċ$��^Z�m34�0U%s}~����������W���Z�6}o��l�
���2[��4�����g
�Z�۰w�@IlE	/���<������ ��ޡ����Jz���ُ�a�x�sZ���ܶ"�+���^d{�s�׀iȄ�����w1q�3��*�TJE՘��R�3�t'Ĥ��:���n H�Z5��=,"X��:�� Xi�sX�$�ς��l���W⸼��0����.��+ K�+P);ߪ����~�L��G�������@Y�����LV0o�Q��	��酪h:�K�6�����B���Q�	�����O�� ��ԭT@��@�I+���,s�H���1���2�����������Y@,;4+K9VxC�7ޕg�\av`�wQ��n���<��k�]]��&�J�����i��^�h].�n�O�ߺ���t�޿s[ V�<	}o����C�_�_���.����	����̽?�@��1�z��߇%�!q��R���oȺ��x�%����F��C�J�>���������ߘ����>�����]ӝ���[h=�����X/�[�6^޺�TR�%�%k(���j����*=ic$��k��| �B6;��D�,�=����慫#X��&0���űK@��~M��3���@y'�c��P �>?������� �.:ԈwrC3���]�XJ���o�3-�����	#zߋ���	�Ў���.�O�sb\������k�"���0������(�0�2afﻝ�-&�0g��FX?�X�Y�xv�cwI-1w��롯	ٍ�G��c��p�e����*2��J��DX"L $Y�>���������6�b�at��l]?���{ow�H�g}v\8Cdo\]N�S�I���=M�W".^��3D�V�����s�_t�9J0:�/�o�l8�#9kc�`N�.�䛓�X	�hk�%��Kn�4�Ѵi 0��ʈ=ʑ�KQn!�Dڨ�QK:d�V$�!����L�)rԼN�?oZ1|��0mw��6�[ ��7v�4�4H���
V��6O���M�F�%�2����u/��@�|����{�lyy���+"(����
땜���z��vP��������w�pR4_2�$.�#��`r\���V�f]�F�6>��/.���dX���F?�]%��Y�!��	K��W<���o�X��J�xd�B��'�r �$.ƃ�״�=}�B���w��w���M��6ϣZ)(�$q�k�	����4KR�C�Z-N�����~Ѐ����߰� @�����Pm�%I�'��;$`E��r�rap���s.T�TX��N�N�j���V ��wU��^��Z�Ρ�g���8�BH2'Ϟ��
�J���܌t�ip��8T� �-�@L�(�rE�)�Ǭn�ׯ��`��8?��3*��[�[҂���ZL��iO ߦ���q���-�ʈ��H��9t���
J�M+ގ��{��WKi $�0�d<!��OݓǏhy3��c6_D@y��x�`#�+*r-V�'��  ��&�j�5+�<y����)�'��㗁+�q��{�*���uG������q^�n���L5�R٪��<��`��[0s/�i�%��}���K.�d�0ޯ��ej ��4C��Ml����ǿ���uoS	�e�kU��A*��g`�S�Ss��3��7����p�妨)�82S����~�e�/Z���4�F�M�p�NLO�e��Rn��md�Yٵ���@ΪV�)`�7�Zc>]��B�*,Wz��DN4�EfQ�����M�fP�H��ap�/Ј�̽���C��u����\Λ����3\X��'l6z�a����q���_ 	z_0ū����΄�k,�|��>�J�[e�W��X�����?D�3�rFq]������V*H ^�8�F#�V�-���QpWn7n���Z�W�(lm�����������Ҋr��Hx�����"[�n&���젊4S/��,�ˑ +tş;;��|}3wWW3Z�zM�F?�5紒@G�  !k���z��F}��R7\i��`U�{Q��%�='��e�S�dld�5����B�F�+����癦�������K6_K`��%�f��N)@�a�' ��_�%�����.0��R��ruN�P[�11��D�R"��*Z�VK򰤑[l*�(a�a���dIC�4�w��3�2�\� ۖ���(�
�]Y�c*	 /_�p_~�ea��$O�/�t�͸`|�J�\(��<��d�q�ǌW���P<ޏϲ�K7g��̊"W��[�&YJ�,>(��J��9S�?E��{~�?��X��C�+~������z����F�^��z�-�+B�1D�+��8�!(J��!���_O9�k����C�m�!4�Te葃߭~����FC�J���d˓������v/��	8�n�Ul�xN�\�W�/�ol��9��TD���Y�} (Rb$fD����r���qK�jiǴAW���H�����^�;/#Q�^���'U�	���pi�.n��i�d��9�F��/&{�ĵ 7��ژLTp��l(��� ���6w纂����2�X{3���d�]�^�4lO�KZ�6/�f�X�;���/��#�N��hW�K%����4uNEгg��~���kK��^�U��Y 4\��l��@r�N��ѩB�*F�Ƙ4�I9��;�F.HF(k�!���-jn��O�F�p'������(Y�������81fY���$���hQIn�" ������׸PZ?{���R�=
D���T��K| �֜V�B+�䏚��!�d��~æ��{���Da旤t*���ܑ�B�ca C(A��2��������iҁ�Љe�I��������3kLb��E�88$U\^�0)ckYג� K����D�U�ILⰐI����k<]x$��`�-Ђ��k�}������A�%3Y�!��'O�rn��rlia��}������d�1� �`/�l۽��8���gڡ������o�3�l� H�%y�֗XZ{O��V);Ewe�
�Ϙt�af!J�K�r�G׼�I�+ ������)��0��?׿עb��FJ9�7��ZU�e)<$}�P�kX���>��*�RIG���!Ҳ��#�1[��2Xrv��� �����)�����ΰ+�M<��$`*�=a���b����w9����UK�8�ztZ�A�,%�$�X�x���E}UO Ac�P��YSq�%� �� ���
��`�I�MVcm\9arB�h$7T�ٗ����+I�R���N�L_t �,�+��&uZ'�=W���+b�SR�p���[J �&���Q��u|P��ᇿ~�%C��+;�'j�F{��=Ѕ	�y������s��FJ[`@���R	��Ұ`m��p��$��1HpKª�j�<�b�I̐�;�fڲ�"��k&�i�겓q�������&#�e�h5�]v�Hq��%{$��� l�܁� 6,�͢�A�@^O	&� ��;;�tǧ�nw��a;;��˯�v���oŲ��@qS���b�E�~=9=��]��;SZNП�� �����-f�aӽ��t׳r�<:�"�W�R{|g� ��q>��V���=
xd[�|XhH�����������;Er �]k�,33�Ia�, d�=���	`�V���{�߅+�X��<��͛w��F�6r[(����ix���V��+(*C�1��{��	�M H��_�q�'ǜ�O�<v�Ͽ��}�� m�s�ɓGt?x�8�V�ԃ܏c�O�����W3Zw�	�D������X�rb��v�� �8�@����%�K��ñ�����7���]|�z,�[�sf��ă5�k+�X��jɄ�Vk ����ѣ�Vq�g�EH���p��\�������?���VS
����==Rr��M)k���������Q��'�\Sb8W}�}���U䒆z���<��qNhIv�x�ƠD(�A�{+�$3��ɥw���@�}a��p&�]��3Xl���)Ɍe(ݾR�#�Wc&l|I(T�r�/�Y��b�V�2h�4k|����R׭6����z�@�=�:�_�"(��͆*O�d�
����j�[:>Xi���YO�%���ݝ��)�(*�/�;��bXmָ>&�T��a0��??��q�,�:�`l�2ESzq/q�AA�&7�F4��en*����������2�1�]���a��R�s'Aа�t�������v�'��,n�7��[���&apc	C������j��ػ��-���3��Ѿ����������_��Ȇ���f��m�X�!ۏ�CX� �����nC�e�6z����]�-&�%!(E�$2	��wi�A_��M���ZJ�/ ��hE�*-l�ۻ����4>'�
�#`�-)G ����k~��K��I���swy}ō�ի�  �V�Z@���`퀋ĩ�>!����#Z��6�2Q,����gO9O>��Ѫł�T8A֜��ӂg�V
��c ���s ���p�i���yuJ��dd��"�y��]��k���ߦy��"����+d��UcR2<�mC-���3Ho{Ώ��G��/�뒎�/.�	P�r��[�y��Qs��#��"�H���2D��a.7,��=�������d� �;�s������t{_ݠ�X��Z�տ ߧ�R(LX�2H�)N�
p\�{&����R�~1�hӦ_���DR��w_ZA8>&V�uf�_x|<���Y9/��?�:�-g��F�Z��k�����cs�Ouf�q?e���kk�>�Q�$f���Z���lo��[��9JJ�-�����O>D�/>�nqi�3���!���2a`� i�����[C�5��Y(����`i��f$9	��d�.�ESکh(��̒JZe�K�����	�6lu�zm�ؾ�1i'�Vѵ����W�6��\o����U�Đ[���q���m���<��k����(u�R������̯����B���m~w;ٔ�d�b���X�S&�|7)��s>�"�j8�cN�����bK�x12 w"0 S/V�%��[�l��	N0
:셫�d��> K�_���}���q�z��D`U�b �S5f���d 6Jh��Q�؛��O����%kI"��8�����u�`�\S�ᎻaO�*��й�q#𒘥	�0�[XK..n܏?�v?"~�\a����(�#�
�ۉ�>b��55f��.,���V\x����t���e6���*t���ZH ����೪F+��RG�c�F��l��J�V�� /l�mKk6��J�T�..	d �����h�_^�����){nA 6#T䘶K����:��V< ��w��=�$�Ep�r��;��QT?9=#xƗ��k�Z]�B��6\�{�������{����9�# f�!��c?#��������n؇�k*���S�Q�K�Z�k�k�������I������;��������ot?�;qGg7����X5]����E�3{��X�ǜ&_qd�^��k�>mV9~k(i2�ڠ��l�����t���C ��/��b|W��Зb�����`fqW��w���<}�\/�M�Ypy�7o�.\�E�SbP��\�YQTP�&��]���W�b�.�%�V �w�������<[�Ǘ��ޯa������!��Q�>h�z��d�� Yܵ┦��*ۜ�ĀGE.ҩ{ȕMCRN��r���ؠ%9�&��@����	���/�a焀t��#�g����:YSGK�4@[�̎J�2���ؗg�]��jH��y~|��B�0��r$�h�[�y�#v��v�y��z�R����`[YR�94Y����2��l�g`%bd�k��P W7F봦$� �� ��wr��w��{{|���2b+!:��9!B�w&ZyaŶ������={E��$��� .�H�
W#6H��	i-��`3����ٹ{��=��X�������?��l��|�,ؙ���2mhpK�@�� �k�	X#h;9>e��5)���<������&��G�X��֮��r�J.������%��n��׳�5��������|] �e���OO0~��kA���5\ld�{�N�)��H퀾��X۰��0�"���:�WC������!(�g�g�(2�	�yZ �u�k���D��Ņ��L�;����7ĝ��-��@{1c��,��q�g�����q `�+��g�����]\��6�[�j<n�,( �j�݉E�Ӧ�*���p<��!�	 ؇�S�.���z���?�� �9V5��4%,���%A�rϷX-���_�L���H�Vzy�����үy)�d_����293x{MC���������,_i����w?k���L�`�Z��T_�O�i{V�69��n�wZil-��%��,&|�>X�Ե�����1�e��:&ɠl=�َ<
#Jjk9�r|����Cg��0�9!t�h��/a��{�?,����y!)~� N�M9B��
"���B��tY��VN��N�Ԧ?�|�P:=O���{2�✳�`�yΪ�)�1�^��@�!:�C�F{�|�dhړJ�ߠ�SwR��ʹ3X/i����+���@(�·I��.}[�ܢ9�9F�g���#T|�8 �5���d�TS`�LU�䒅�k�<׻�;��s��@��"�R ��Ta@1ָN�ʛ��Mi�3��'�H�ǿ+7��튛$�����^��u:ZW޾=r>����B���ތ��J{��-y�޼�)n�[n<�ښ��@��e�Zh��$�n �����ܕ����HƠu\�ZH<�eq�Md�-������ �=�G�� <j�!���,�%�ooM-H~��\�V�����3C1�BH�R.J� )X��jɶ��V�7 �E�8'e��R*�,�)�F��p�ڃq	U����>�tu+��-��RKn������6�k�$���]���`e��j�u-������gu �N`�V3ԉh�j�����_�z��Gv~�$�&C�c˹/ֆ�������}���N���-3c8���s{~�D���.��j	T�D ¬��_U��myf03p%%̣tw�3��՞I_z@>��='�m��7�'ɻ�qW��9������d�*2�+��O��)`�$���[�{zˈD�Z"�&��2�ƤO[l1���܂{�`�PĘ�ߵn1�UVP�Oo�t�ڜ+�S�u�;Q�� �WóD�5M��6�g�,m��E[NhI��i�S�Z�N�&��"������@v$��}�w�>�sy���-wNF���4�ѝ�:�DK��������!�qګr�+oGF���sf��/7h''AQ*G�-ĵ�����]�����C\	SK߃ǯ��jb� �i��^�5�	�ڭ��	�de���Zs-��A�}*B�W�Y�%c��%������k�oQ��@J.���������76�&n�q:���Y��Q����6U��/tj�Z��iM���p9wrvI������;2����FwY�&�4�v����kRc\�~��t3��e]���$R�������D�k(�D1��x_T�`�5
�"��D��(-��r��Lb�=�7c� ���q��@ V@�l�j�q�E)�Jƫa,]Vp��|T=�BFj�ɱ..�	�/��1,��b::�^CX6$��L.�O�Z�im]XYq�nQ�-��	@�lF�c`}�"P��EM˫�Ki�[����RC/h�[	v�x��"��v���q�����$Q��k�bIV��(��p���p���;o]�X��
n&[n��2��J[֦Z�̪:)L6��l����s��� I���ҥ�Iv��{�W�����_Y�&K�����_y	�O��ޛ�F([��5��h'c�ؿ2����B2}E	ry�uJ�Q�;Z�\qv�G�Tפ�)���m��C�e��i�Se8���k��O�[���p����Zˆ5��z��5,Y�7�☾J�B2�p�A-e>h��$�� q8��4�Y��'�����5�S3d����\��Z$ ���)��e�ѦSH ,7����B#$ fЀn���%�J����r�P#�W;~	@�k?�?�$|~���.`�d�c��Sj�j{���c���,+������ M73��K����S+�L��R�]�v%>#ZmpXZT���#'����.o��:u׷��dgύ��P�̒����,������~p?���ٗ��͛7,����ʋH,D��+��Ѷ��m��Q��Y)WO�b�@��o�V�ǲP��/��f��8�[ݸ	lI�"� I��J��w3�v�-!YU7���	��
|b�pY�����8q٦��ڕR�H���񜰜zQ���x���rQ޺V
Ը4BX����U\��*��*�3��T�/�i�^�t/^>�X��x~q�
/^��%�?��O�u��>���rv9��!HV���+��g]=��,N�0��<ܜ�9C������#H� ����SK�`���u�Vj�ަ:����스�V;�Un7�{�E��b����o�p9n����UxL|y�A�Q���5qdѱ�ib��5������޿�qO; ��_��L7:UB\ѧ��&˱�7�JW�HSkI���	�-��2ր�* ޴�Բs8����%�m�q2�������w���	���z�JdE���-�|1��Vd^J9
>d_'�aA��I��
��
�.�7�V�7,nZo�Ng�-M�2'q������4�?����e�
���嚒�)B SCX�Z���0̵�.[(,�^&F�S�����[���E��A��q���3AX��	�{Glp���m���H��,`���ep�]��V]զ�Y�4�7TNK⬤�Nדw��ѱ��]�E(Y�r=nƽ C�Yw�Z�pJ� c��]���pG �y	VzǸ/�۲�/��i13�f<����<N���aҿa�EX��u�k�5�Nun��M�!58H�T".��uɍW4a��u�ੲ:fT̬͝3��b&Ev.e$i��JX K�MSqܚ P܎9d�L_����]U��j��4)kO9#J�v�O�&�:e&��'���'eC��$A�B�
 ,|f>=�F:c�G��cwx(�a������k��12�����sㄺ�������Ge�8� �f����[�֔l,+m�X�"�Z���f��mMF�;8�cܛ l��5Q2;�M�޶n�lY��� �a'�[Z��Z�1���(.�J�h �����2c5HALI��&�|�a\�P�59��S׏{O�{�?TJ�[�ܯ}躵�k�������|�Q%���� �%WX�2+�;̱L;K�tϔ�Zj��ie����;fV7WwL�|:�#�}9{H��!��ڪu�j%������I�Q�d��Q@�N�h�����hY�G��8��SʖH��졂ˮ�P�E8Yg���영�X�U���}�w�b������<�
 �ڭup0�%���9Ju+�۲�w��k�y���_U�or��&5K���ƪ�(�����{�6� ~MR�8��<I+-�Q��$[m��m����\D��m$ɬ߄�����h�Q�b�A6Cb��;�,�r�DH���^�nQmb���,3+Z�p=�n\����X�:e��0�i*�A�����c�^	g%6�f�����5��נsq��~$mT+n�Fh�%���z��U��>!S�[t�aXѼ*Uz�Ţc�3�xAV�����h�m��
��I�Q����ͻrզ%�C\ V���
�-�Vdh)p]��g�IQ��yPW4���[�.W^�yvv~�g@.�o�7��N,��5��%�7�rߋet _��<v/^<c2�b�����$�}z���בkɳ���s�jT�7��r�M�D���%��g��6_���á���fz���k%���Zʒ{ Xʍ������$C	��ۭ8lbe�g��b�����v�tm�ms���˶8[W�������G��O|<���2EK-��/ ��#.U�9�nv$ut�ZP�İ�+j��8[1���`� �pL��6��w�[�G����|��bx�R܁7�}���^�S����Q��;S%����3Dc�#o�c_et�6M�:´IS1���t� hHi�^��>�����[i�2X$1�G|W�ͱ��S���R{Ҁ>7 ���f��iA�����U2�f��+���n�����=8�=��b4��~|���;���gEDc�,˶���bs�4I'����Y���L�*ae7AW�-#�5%\d�*��l�N
OǟcNV�[Y�l����:ՍL���\0�>��V���������6,��t'�P�t%�͘��2E��W����j/~�e]W���{#����t'~>r�El��Q�ڳ�JP����� ��?a]jX�:��z
�����[}Y��Xwr2�e��e����V�TdAk�O��1U���j���K֡K6-i.(Ȩ�b)d��Z�X�������j���"a�Ӈd7�$)��yN�uP� `V�ɸv{{[L~ ��b��������u��87�.˾�>@x˾��IX��v��P��;�t/�,f�����\�T�dmOt˚��$�4a���UŁ��3���-�C6�^�NIg�ڤ�m²�J�f��:&J�+�������oM@+_���,������%���a�2�3��������ß����3ֹR��r~;��RA�C�󂌻�r朏ټ}�B��5�{{Q�f0����5��Fzn0$���!�x�{�C9gR�\K���K��W�����x�e\�-�Y�h߶�y[� 0)�mG3�`���#���j�����._�R��b�SP9�ʧM$hb{�)�a�u�=hr�Ej�q�=�[�����@X��0�R���+�D��Bs�TڷUўr6�����E�|�I	>g�)�>�,J�;�B�O��K��*�)�<�n�����à��� W_R�4���%��V`%�#��o4�Zb���o��*�3�?Ω�OU_��(㷔 �G/H 7S�+q�	xr�OB��e[�΋-�� ���uDm J��:e^�,OK���&�ߤ͐����x��V,j�8I坨�������ۥ��:>1,:`���^��U`< 
�����g kG+%@������&�lv���@D�����nwg/
�5)���
2C�pQ4����d?���
��(p~}uM@��d�(�l<������}S�+2La�Y2�����s{�p oZ�<"pB6"�Ad{�_\���ߓ?%� @��ʵ �1\������_�?��"{��V宧�6���ͥ��<u��uƷ��B,��Ȱ���vO��kc�q9�n�Niֲ�KIɢ}����y�����@O�xM\���6ɠ�^!$�W�MJ�ܴ����*�>�&$L`�$7����G�x���$��
�	�����{��?�X���~��?�>>�贿��l\d��!YȜ�^+c=,�$������xf�WU��~{ǔ+��Tp���1ǰ�w�Or#��k{�M�!��|mZ���T����Ib귶-�j��L�fdT2@�-��f�Y̅�IIXY��/� �f�������D��j.�H�VU�	�oepdv�y=J�ȴ���@M�ɲy��h�i��)͎�����������T��LX�4��W���L�h��YJ�e�.�2��1 ��p�;�����?�z�e2c�2 ��;�B+$�m���r�X� �03�A�9X8�Z_�BZ�!4�6��t��n���-Q�l���H��4x��ۈ�%�J���� A��ChW��^�`��#��:4َ@E��C�Ȳ&�`����)���4Xa�����V���K�c�PW�s�>��N�D,K{�`��~���j/�C�d�MX�Ɩ�r΂�2��+�� �+ Xt@: �|�^_�)�A��L8����llOk,X� �FZ�=ޮ�u"�5)�F{%Htn����"��5&G����s�@�茰Z,��� <}���������f6!�܎|�jY��hu�6�Ș|�����s����$�ë�]��zv}���N�E�c�0��ƨ+�E+]SK�Yp��{�Wg��T�\�VH���[#��-�6k��U��>(�Ql7���ʳSKB�Ö ���ؗ=��.�����hS�Ӟ��{����d{� �I`���%V�9d�����o��'��>���6��ÑI���EK�S���uU�E9PuG+�q�G�q���\�7A߫�J
Y�SEcz������.?-+2z�`��yT<U�g�o�J�Qh8��a��Ţq����m~'F�V䧤Lb���})��~���Qu�����T���ு�ܯ��Tʋ�v�>�D��:�,���Q0�n��H>�c��i�U*�PF��Y}zN]{ijF�M���ks�N�KCU,��b}�C����L�d!���kg��~���>�v|��XO���A��Bg���mw�è�h�$��Jؤ*�hUq�:��v�@�$A�J��  �e��Uv��o ��7�b��8i40��=�yW�K�<`A�n�"�f���i ��eϩz��8`-�=~����?�޽x�� �G�.��H4#X9;��_�G�K�m�T%�;ɆÆ�ŗ�	^����Ϡ,R����R�X��	�?�@�7�j�C�C��\��u}}�\O�u]H���J��~����-	�b�`������V�--��<�(\��k���s�/���"�y"r��r= q=::"�-�>��݉�C���tB�PF<�� �����;=]1���S�I��p}-�<j�o����~A�A,{( � ` y��2�R��0���{(�pK*4����;;��E��t��/���{��1�@=8�DV�J���h;�\������f��ŵ{��=�)$п�K��)��u�k��Ŋ��w�Vyґ�noG��C��-|��V��	x6�B��cp��B4���幟�ݿ߱�>���WR�T�j\��4�n����h�I�S"^G��>��;e)��/�,�9[a�Ù������r�mr ˼O4/vN��Ce������j%�d��A�G��`]D�Թ�݊�`U%9x.���d��k���f �����*n>�b�WXŅ�V�ǩ���'�Q�f2wOH�Œ����;f�I,��A�Y�h:�d-�r0-eM$��ق�b��DMg M� ��nf��k�W���feb�W%13�L��Z�}l���v��o���_*~���3���t�(�R���5Q(�E�����i���9��mdI�d\�|c�g?�vWϊ�r��Wk ,�P�iP�y����!���������die��teZ�rJuE�
S�n7�f�v�dbD�t3����<��Gq�Ś�@�w�)Q�ѓ�!�Z���ވI 8܍���_~�?�X2��_�Ķ�uG�	8 d��2����Z�x��=AǁX���`�?==� �2��;?���JZ�e<�V���ՇB�_}�2�gKb�h�������X�c�-����� -������O�X]ƶ������ij�+�$q������^|�$��xM�"���OxH��w�H4�b��=ڏ�h�`K���Zl`��-J�B�P	��*�\���TZ�H�h�� ��{;üXh!��im�����˗��I��[鶼 ����,�u����P�U��W���:'�����&JI�(��i݅�,�E_�:,�X�|���u�3)b2��[�N�%&�\)~5 �QԄ;?m�~��1eo�6�y������P�����خ�h�]1z���ǔ8�ap�ϗא�e��U��M��f��Rů0�8�y�r� ��B��%2�����kֻl��^�����n0����͓�A	IJ��ͨV���2f��{�-�T$�sѓ6��Cƀ���H<H�R�8Z�5��`	��m|�Dm|FM�G��Jx��1���NK�8g\-L��1��ai�{'�j�J X��i�R�-U_�kv��]5��aY�:0���`1a./�4ՂY�xn��he�U�%\�gj��DKA�.�Xq��s���jm�n��p�����u����Ђ���?�	$��aM�9�R!H��� ��]3�c�Ҭ����0�rW9G���"����@,K��:�;әu�?��JkF�5�ݳ����������q' ��<ަ͉KT�0PLkI8h-c�b�@!�8n# �9u��򻸐�n��7Sw}y�no"�:܍��w�q����f0�%�_�̑̢���%­5�4nwo�����'�l!�Nb�����NYxh��������k�h�+�ѣG$������'܄��ҋe��y��B�_ǾPs<J��vqq�>�ci����"��x�K�cdF�+�Z�M 0�,a��3��;����~��ߺ'Oi��X�:�5�c{nܟ��\�J�������L\F��V� �"�u� 6ZE�ZcGU�krE]X�	v��kf�z'�[���=y�ޗ��/�L��t-��]�ޣr�;���2����<ltP��n'AX2\�K)�J*�u:����$�BA��8PN�͋�{���]�ƗM�j��� !-ƌ�ӵ�\�����9=���J�@:���R��e�s��p[���ϺŃ_�����A���`�x�ĕo%z�<��/M���nI� �f�^AC����ɶ��5�x�ԕ��2�U<b����k]�|Y�njC�HJ��fz{�¨���x"$�,Fj#T�p���r^���Ȍ�b�~���� ��4Z�k)��j�5s�1�����K�oEm�ʟx5���7����.t�>�`(�{॔���­��X��*2�����
p� =>ޯ�y_�89��P13�|ȋF�$$X��/�_�zӜ��ip��/��y��1�2	kڼ�вI�O 1<��O�6mҩ�I9��o����u��CM� �9
f�`v�k�ȗW�j��u3�Se��}⧢�5�^0̯��$fE֝d�u

5x�V-�r�+��W�0nj_�z����/��=��-��<��U*�����&�B�i6.-��É�k:�sȯ�\�/��b��j�[��0 J�*$܄K)���S���^X�Ro�}��zhb#�%  �!kj҅F.��%US3�>,K-[p��5�$l̚�[өl�L͓x���@&��1�`��+��x�5�@^�bV_k�U�Nb�F�Z��(���=���貖mb�GW!��# ݚ�9� �=\��*֠�%��<b�[�k�be��NǼ' D�Idx����䏜�5���B�p��|���;�/mw}�a���sgk�g犱*�p#|�8$�n����A=V��Ǹ��aQx�QE!o�\O�O��2�9�Jvh2肌si,s2�}Z�Y��t.]��q����Ȉԓe�Y��I�Ja,C�����A�\Lv��s�5Yu����q[ب�~�0SHb�,PX9���:pIj|��5�C�sO���]���}v9��t���b����l����v�EU�� ���axR1|Ƚ��i�-�`LÖ��"$�#�@<qE��ܙ/�&���D����5-��I��8�Q�s4L�t TKW�ŧ�Q!�)���A1ݫk�D��Ƞ�ₕ�q���xaя��͎��.�Ы�	נ�Q75jj+!l��J� �6M�^���!~�b(�aҏ���#�lfZ̎Ƽy%���W��x��!�ɐTQu��8�s)i"Ŝ-,�6�శ����r�������u���O�f�ơ8���m))M�Vd3� /��%[_��DgRj���8��s�"�*�)�CHM@��(!�Gt1-���(4� ��z��c\V\Q�;S���孖��eM6"hNmۥk�I�ba�G�"��n�������ş8c ��^�!��c��-}*d��-����Vx����^݇����[I����Y̙I��f�Q�-��Jp-Xk����؛"kr<J�l\��O^�9�5�[ɝZ 6h��,6Bz:"����mE9��Y=����Ge�:9���o�//����u ����K�^e��2FhC'֫�K�������F�����be�����,��l&�ׯ���kwt|�z��B/A_qL��9�s������؟�,o�����w�}���;_�}l3x��v}u����#���SR4���+/�R�`N���'�;���Y�wIa�)%��;��L� j�b��.}
ʌ�@���P�dW�%�P�W 0_��$�P�� �\{ʻp�w_�J��sQ�����������OÝ\���hf�J2�bJ�"�-^�!�Zu%M��2\���\��k�X�̢��Wv� �(r���K�.�_��I=�FP�`������V	E������a"�yl�ꚡ$�@��A��r��O)X�G�o���p�X|��F�&��z��-�Y�\o0
3rɃ�- ؒ��/����(.6)%�u�s��Pn�Z'�m.uo&{a��X<�!L�|6Rٳ@8Z<���~:�r���G�`��V{6ݦ��	�B�D��H�qg�JQ6���6� OX��@s�*�v�3�V��lR�ʃDy�5!0y���Rg����׿�j�l��V�T3�XI�B��9N[��6q�xV�����"˰�l�]�q��.bb���ȼ��q4ԴL����
"T�ħ�k���E0� ������dZ�m�`����G6A�*`f@��x�nBMʷ��F v���')i���-t-�f������Շ�8?��`�4n�W{�)rw
�Z�V}x7�oپ��]-h����	)�q �֢ ă��a����A`h�۷�| R�4�Ӊ�X����>�ׇ�,.�yP��6~���cj��Qh�����������6A|�~����ױ�N	���y��=�x}����{�s�
f�kwrrD
���"+��p�}��~�ߣ��5�2����;X��I@��ߦy��g�r�^��#-P���� F۾��{����G�6��y~~��������i��򌴖�*a	N��"��S���)�����*I��t.�"t.Ke
Y�l�^܏f���R `�2�ﳷ@�T���\1Uk(?�6��SiR� �l�ț~!7l���>��51�L�4y>_�����e����a��,/S/�æ}�\�����j}J]�������k�Y����3�!���k��D��i�hJ���0� s�%zØ�+V[�C-֯
J<T:)V�Zes?K� �);�>i
��D_�č�U��
h�0Z
��n$��U	�#``���
Jq�ѻ�0+Z�l_Ǉ�Z�دH��x� @�W��AW=i��K:�1��)�}�|�]�@����n����+��Hy�\����b�T�v`��kP~/�R��;���9.|��=�!�����c�ؑ�;iS֨4�C�5L:��F��Ϡ�����=e�-�@^&Y�Kh;i]�_R�
�w�ؼ`�8m����ֿ_L��)z
 Y|?X����M���L��.o�H^}�:ы�����8	�B(Z�|pVC���,�����~$��Z���W��f�u�{)�Q�8>�I�ї�=
�z��5�u��3��
�h�x]���?��D�"���C��We�M�����g���Z���!E�yķ߽;r��:;���a�=�+d/~����8��I��:� �\<y�Ľx��]���/�.�D����`�[HN�������p?���po!�)>��>�8��R9��А ���"X@[2�Շ����������u�p��f���u��Yl�����V�h/! r����b_��:��^A���������={F���%�.8��3��K�\���v=�ݷ��]]\�7��PN 1�lxH��P0����1[�?�9>�;�@�F``�b��T)�QrO�g��?�]Ku)$BjY*)���^hS�.F�����O�ًW�y���S$1��qō�ѳ0��5�_�8�2�O����*�z�ʹf��M�1�7ZPc@�'Ŝm����7~��q����ְ���N�ם���G9����P�h��N������G����C�����u�������}�Q��8IFq��>������_ڿ�%��I�@�tk�mE��}�<²u�$�f�$���B%�Z���nA �6�Ҭ���@��.b�ʊzP��H��Ȫ23�D-��]�[d��.>S���|J��`&��{I�!K<$�^�JA*�'�lEqe�(�F�������*������ş~�Y���(>���F���V�fsjj��j?ŋ����x�҄?�̌6��v �R"�``�E�Y�@˛���)L�Yc�3��H���	PS�E�'^�& f�*ɂ5<m�g�Rߵ
_C�!�k��]?-D��h//���w�+��`˗/�QX�LSL_+�חW-h����Ӹ*�%��t�r��� Ұ3ĕml�w�f�v�f�H�V#��R���u�$�yX��r���Z�!��x�9��n����n��N\����)n�o޾�1� k���{�VJ �ֵ��`}Q�b�66�L n���x��l\�_ -H!�f���-L�_'����>��a�1�t��R+�v
P��#P:f�����OON�~�ҥ�#t4�pÊp���)��@`�wdў͵&�ϑ��g���"p���ry��z.�kT#AlV�L���G��V�7d<�9PX{Id'�V���8ՌK�	����}�dU���l���t��hI;b�)X�F(%����t���p5����\�l��ᦡ��VK:-R^J%ᚇ��^���s�x����\�a�uil�����ԊOG۩��eBݘ� ^��7��`�D���B����r��x�|������
u�]1��BQs�"��c�ά�I�Q��۠쥋�r�#�l  ?vް�~-.'+#�$k�$dcV%�ƪ3:&)�$=f��^Y��\��z�R	���$��c�,Zǵ�K��\�X[�N^��cI��j�>k(b�2�=hn���5YBm,�I�b@*��l�49o���끒$eh��Z�
����O���$����%�]�3U��,|&��NX0�e\�nk5�-�v&c2pc�"j����)�(���t�<��G����KB!( Z/��͝՟�,������N�v%�U�FI��v����-�YfM**΃sq"3������{���1;���ZNE����zqs�y�R�M#��pn��a��4��x�i���u�
T(��.$�f���D�6-�͋9�d���w�)�����ߧ\�w���N'"�V�A8���^�-�aI<`A Z�|��l`����` _IY��b�%0��x�I����>�lE����*��:*.���k��-}��n�ؐ��Z��+�bE��-�W ���,6�z���j�>H��l�sw��,�p�eN��p-1;g%�(ߑM�; T��H��NH�F�~]��]��b���3��4�x*hU�>�sI�-1`b�\�.e�2�>Y�d\{�6�Nkٖ���48����5X�ҍH �&.x��r��c�Y��+��
�^c[��ꒀ��� ���p��������H٨\x6�R��b�:]R�:���CMő�ދ��H�Y���~d;?}�v� ƶ$�3��3�]�댙�jL��4��t-�P���\����7:�6B�5ܺ��Χ���h�'e��>�J��so��:��rc(�� ���Qy��?��6�E��N�׀���,�zz��>�f:��&7��ـ�]GW���0��i�ʊ,G�|�s1���A� �_% ^�	8���X�Gr��OF�ۙ6�Ԥ���#�ME��GS2��^j�!wm���<[���� �a\��I�'���_�Y<uۻ�L�8�/o����%� 㦦u{C#�J�q@t�&��&��$++���l�5�zXp`۫ ﵈��ҋEL \��� ɲA�&-_����d:����xo$v�op7US6�o�\�,����P�T0��a)���TlGW@`-_�E�sI��'n9ͽK�H1���H�\6��ˮ���_?��K��M���l�L����Qj��:�-_�ӫZ��X9�!�g˴���x��Ok�I=�%�f1���AI\��d6u%R��k��J1S�QL"��B�P9HL��� laC����$ �d���aI���>�<kK�������ܑQ��5����Y88�E:	�d-���d�ʼ���\��׺�ƾO]D�"��!���\{�W�?+,^���.a�/��� n����bs���`C1kn�x6O+,��Z%�qZ�t��l�d ��������ˋ~�\G�Z�ޡl�QI�P_YhI��l�q�^������.p^�
 T��i�����	�k������h�I�Gh�3r%�&����fj�K6C�Pq_��pI!��e�dc㭵�{�^J }�>(iq���a�x$Y�Q��Tu�&�v���S6���I@���	�&yk߳�4�(�TI'7dp"�d`"(ڔ�ۖ^R�ղua�bv7�(kG��5r��Q�6��z)&�t(ǣ�va�*N#��B���q,jx�s����[��Z�$�R�Y�n�g���� �`HRAv4Bp �>�àv��;�� ;:>%��,�6X��
fp�17����0��͠��/l�rN���J0��(�*�V�;��F�p����1
)�	���4W�vr)�2ņ"�(k��%3�+�Y{�ѐ�#䞋�/��#-n�5���Щ��Pkv�׺~xi�&����g�Xh���q��(�����c����"����c#p.����gf�.ϭ|:�i閐���M�6��U�R�s��D�|�B��Y4;ՒDy �ͭ�C�c�R���Fk���<�sX�p݇�j	����o��t�y������w�XT�܇!���k$sx��K��^7L%�T�s����� N�0x�,+%H2���P_c��]��hM��a-s��E�	H�����u.�jBt��X�m¦yo�d[���)�3���%2MdQ���:0�c�	���:�*�a�x�?�z��3\H��Z��3ߗ1�j5���j�q#�MQ)3�� �A+I4�	Cl$��Ӥ�n��N;M��4,]�����?��Cɑ$�Ts@���U�]C��W�dD���d�v��Lwɬ$���Δ<55"�zw[֫�8�͍�=eO�3Yob��jfi���}�VH<:`��d���p�y#2 g_��^�D�f��Y9=t|M����d�?M�裱��=!\���L�*\���C��M�H�)���5U�Vb����'\.]�_���-}���yqZ�{�6o����Wخ1�V�f���^-x����<^��am��%��%�{��s**�]��e.����1��ޣ��꥛�_~����
5�Ta�DL��V7D�����
B=;���?܋[H6����΄W6_�� Gl*A{ɮ٘`��GN���$�b���� ÛL̀��� M�fFꧧ� ��N�[��9���c�|�x+1?���%��8�a!�r�pΰ�~�fmֵ&��V�FL�f*�'#�8��ӣ�z��u�U����ơ67�~qF���s��=�^t͎��>��kV3H۠Sr��k��b*C��u;��H����B�BF��;C9�=�F�]oesZ?�)y�֦���3������ŏ��B��|Q��9���LQ!%�=�8�D ����9 }:*��D�n�� �ٵq��� JTbjm�M9���Ol����X���~ނ�xm})�P���k?t�n|��Z�F���hm�������q�{��&��v�W�u��uYT-u��ڜ��6�?[�X�+ J�ugM�3YY+_��f�6w9�:�V�����/��ӆ�F��':�~l���"c+�TZ{��2�>x��q�k������xn���3W�6�����}tQ$(1#��ɓA��=N��&o� H��Rw�LdrL�J�ˆ��昨n�Ų���+�y�����G߽{E�g+:�d�d���)g�05��,~��v#�'X�|���3Yי�k1�^�:[֤)2���t�����u��u����]�<�z!V�]c��Xuv�(��\G��n���j��ll߬尦���k�����ru,e/�* �B>�[NW��Y�P����Z���7�y��$��^�jG"�4�H�A/�.�L����0?�@?��sA�?���)��aMm�t�f+K}%!tF~f>y#�W$N�)[{�g����H�|�9{���T��~j+d�4���!\���c�3@��Tst�̤?�7Q��@&��õd�m<�����80X���ƥ A�-���Q���( ƬY@�^��ZG��W6fyg�?�)<M���5}��==��QW��,�O�)@L�J��+���(Uw���+��eȮ�`<G6ٙ}� z�{���@@9��d�'��7f����J�n�n�,��|�M�_h��Ϟ p��C׊ m
�F�W�3}��ωv��2̮7��`ݮy�`e#
���S�Xu!릦�]���|5V>B�C
]v�]�pG3���%�x#��=׋�k��q' l��H-@�j�.[��mT6_�KY�j������o����S��*8]�K������V�xYu��4yQ������;a�)����ĦXfЖ�r�0Ģ�NO�C�GPk��&W@�[� |�\Ac�y��pͲ�//N����w�{Go__���L���� 8.|�:4����1c蚵#�}�@|��-`rf�y�����M�%����#�x��6%qb�t.:��ׯ^�sb�1�%�1`Q ��Y�si�����}R6&0�³5���>�?Vu�dj��'�*p�^�3gW���
q`\A�w �5��ʔ��F����zyN/��U��~aN��o��ӗ;	P��L�4r@6��)1c<97�_S-�Ţ�2`T� ���~g�X)L3�J��n��d�lo�㏜QM��cOƄ�������KӍ�����1h@�D&�2�*ń�j��N��w׶}��e���Ĩ����Q����$-��R,_�y�Ϣ���Q(n
�g����'�uuq)��`�*���Ī �@�ʻܴ�~#̽���o��^c+�& �9������A�(����n��(�L�����z%l�e[^9Ǿ��}�dI�Z�9<s״+�r�{D��N�/�`:V�Qs�p����ZtK���#�fSRyՙ�AX7D�`�5�S�Rh�0%ɕ�K|K��2I���u��D塖���T�;����&��@S9�q������Aj�8M~�
:]k)���
H;����ߜJ9����6�a� lPV�$I�v2!c_ XW�s�{��������@oJ�q��&��=�ڵ/�zK߾{E�E���<Ú�V���/�5$�/[m���S
a��VT@���T_�	��2�g�̻���'amhX��gMP�ڲV����W4?Z�c����F��>��/.� ���L��N�T��-t�q�`����twh���,�>\N��F8z�^�K�S���e�����Z���;$��i�s��+�/�����_>~��������J?��I\�Z�lN� ԣ~U&�����A��3"�P �y�d3�Xy5}���O!���lr�ř�O�V��F�ϻ �r���_�(K�E�k�IMkL@={��|�9���`�0~9:LJ��F���|3-����4����Ղ��cО�D�P����J:'�4����E�{IPY���p/��,x9)�D/Űo�\�$ě�(u��"���� �"��s��
l��7�,���rm��63�ڏ���1�	�Xž�?q�)pܳ��MA�n��������c�p^��=G�om�2����}�[@�d�ܭ�cO�_ӟ ��[rY5z��	"��	X��c�����ƍ&q,V�@��Խ��TC�B�����3���$�LC���_�Z���2�Z2�
'H�w69�}W�Yꁱ�sA3�c)�VE�^�9 ���Y��+ܺ~��v���4�!
�}A��>�^��&(+�R��x7p�l��������}��$�!i,�oִ}*��tI�}S����Ы�3Idw���X�
!�P4��%��Y�67"'�HU��.�7��k7_,$~��2��-���ϫ�}��/�W
}��%s�HLXya��l����ܐtZ^O��p�q���y���h��m�d���9]��t�YT���t�(�}�U�j�\d�J���ө���)ŷe�o�
!��kl�,XČPMS�5 ��L�2нg�p��j9���i��zMo^�[*Ύ�B���k.����ayW��B�"]@���c�壹�<Ƿ18d�t��h��3���}!�abEj�z� ]����ߨ�:򁿣�x���2s��ęH��q�v}3 �fMLc1z*n�h�a�����rU��P�u���`��@���:�ѓůx�Mo��2I�[X�RN)����E���JϦ��&�����73�g�=\��O� ��?Zg���K5l�<<���.�2�����XOϙ���#��k������mH��߁E�5�=�h
����6�l�oc�i"���[������.�@[�U�F�`J��@���%D��&#�0Y�WҾ��yo.L�p&�d�H
����+�]6_ӭ�m�L~-��� L�sA��@R���=q�0��\~ڍ��-��+yc���0 T���U��w�]zR+T�%rF��-�M�8�*���Ȇ�6��0(��p�6-��JjGg�}�楼�O8��̉�Z��Wm"����T�$ː�96��d?�m��wke��Fbw�6��օUE��v�mŀwW�3�z��w����PW��nҍ����Q��⨣��#)���q�R�;em�M����fZXmO���ū7�\�$.l#�L����H	YhP;Sj�� M��F�Jƚ��2������ 齳��3��8���~��N���~I������o�?��/��/��Ki͛l��Ril�i�p\��3d�d�زr�$˂`2�v���w����"LItP0�9m���o4n�cMX;R7�!�v3n���K✞�i��d��{c<x9t��Rx�Mg&uWe�/55~��e.d՛��y�t�Rl[�TR�(�Z2�8�ر�]��h\\�E�� ��^4�\���<���p�~T��8(v�Ym�QH�LCX{S��=m��I��DK��y�םZ�bP���O�	��xL�����9�U���Z����[����C�|�iB�E�N�5�X��N��O ���d�`�.;#ԅ��:��VJ2I�Lsѳ�˪7[�Ă�� �������k�Z�fA0*��z����S���X������Q�B�K��j���:^��P�4)l�qO:$;��'K��+��;ܯ8 �#X��%T�f] ����7j6�f_H)�x�`�b䊇�v�0o�;!��ˋ�I�z|yyJ�^_��חtuq\��`��-�L�匧q49�{;�D�?�%�N�{aN��\��]�h����N	��A�/p{���]�<����2�j���Z݌	{K�#�m�	w�zDx�1����C��T1����r��tVr+�au�gg�Wtz���e��=b�EsZor&�_�mld���ҟa2��D��F�!F���J2	�B��J̈́DV��G�贔�b1��x�WmՈ���ߴ���i��/�b�\�	�����蛑?�?���� �jJ/����yw'j�dڳ����N@��RO���
��iOܷ����c�8)��Z�����!�h����$5�rM�\�O����P�wz�f█��`� 7i�#������kv����)��_��BRr��{\֦�Dޘ��Z6�2�ΎW��ŋ"$����mwf-�tn��W�1��@�f��z���Qj7n|z�L��kO�� (`-:��!��^�8����O��\{둼��y��T��mC����UkW��r%�} �4Z��h�� ������q@��h�E����E�J�h�!���֣�z���a�����宂�N�^N��mI��r���֋��:��º��d�۹XAQ�9����Qk�&����X��[t�����Ӕ���#�N?d�����Ϯ�Elm��w�t��Y���6�yz0 ��;R�� �Pk�0��P��*���Rq6�kӼ���\���^����3��A���'��A2k��jt9�;�Ǐ��pL'��nt�i̚�Rm����?t�2�:%\g��f��H{�[W�������㔽g�� �G�~1��a��[���~��q~$�J���U�y���T���L��v-d$�}Y[��n]���j�R���0�~SF�wm0�0���>x�Hl�)�"� y�<g�q��P�c�v��γl`�99d`�ߗ;�cƆ�����������e�yvrL����;���)H���^
�4e���cG�BTGW��≽�Z�?���k�D;Ʃn���YTE������S2má?U�e_�yf��
"y\o�o�x��Ó�qW�t$/J&HX-�I4�^t�b��Se+��V��FH!����Κ�1�H�Ta

�\�^�ָ� �<�����Wtʟ�Q\��b���Y7r������e�6���9��h�9��|������4�*��y�l�Դ�'$�8 ��L-e8���\�b�N��L]�SK�!�[�uW��s�-e�Sc�T���Z�^!(1�����+�h�>�T�|���o\B�{h���]���򇫛E�C����ZrY��1+��|�{�n����$ل�T�mjY��1��I�fNh,��d�(�,˞��<�1�պݼd�h�sd��'U�jY��h�[�<�~��o�C�/J���$W��q@6���l�jk��KD���o�1v�E�b��$(��n�7�
���� X�~���o�0�mo�ۑ��g�x�'0������GE��8;�3NҐ���\b�Y	~|z��!le]��y�.�/�	o�̳�&��}N5T���s=[�S%�����@�X��~��ی�����&q_�	[ڸ�z^�zM��td�3��	��Ii&)�Ŀ���,�v]7i�պm�h� R3�d���_5�!�0Ysa�`@�H��)�b�����l$Ў$>kF�-X�����Jb�e6�l-���y��,"��V\*������M�d��)B��idA�x "/�3���w��2��֠4	Vo��$��D4�"������I[ǿB*�q�Ӂ��
U]P�	��Z굲���.��ق�����Th�]�s�l-E���P���l���U���y�(M�P�z'���q6�+�ǓՊ�/.D���K��I�IJ��Y�p/�p���ڠ�:#��յغ%�.?� .��P:��i��}b߷��ڰ�kN�]ߟ��?6�95� �4�-�J ���<:wZ
S�,�D�?�-dm�B��R���j?��~f}��G.k��S�hj�b�3h����<g�sh��͵��p������u������v���|�>�(~1{��>{�c(��puaǐ1wY;y� ��%�pU��c*��Z��چ�4
�ղS%n8/;�V��E��Ș��W��{6� �ڇ�"^+�6�U.��u9��t`J&�m���=] `s�4F��[�0�0��d�Z�Օ=
�cݙ�l�b�M'��A���'��R]����|^����.�Y~q�R#Jb�]��5�{�>�s'�%\���(�
 �RX%�	������@�X��`񾣀���.^���/h�\	6|1*y�(xna�x���,.6�q���z	~�P��fk�eb�� �ߌr��4��SD�6�����w�������N���b T`J{.N/�l��2�dk��f��^|�R4w7<
�_���n�g�!y�7п��{y��+�=it�X�� P�DX��2x�H�7{��xr-�#�����R�S�����T�����|���������Å��~�_U,�
����cu7��ȋkY�g�p2�lq$وR�z�97�+
��R�Z�����Ա�͂)&�1#q!�NR@u0"Jބ�t�y*@눎ˋ�1MK'�|0KA/��LS���Z�X��/�#-�љ5� tt�����@c��3X���-Ma�e�vG|�hY��\��H抸�$ ^�Φ��>�=��s�PjU�
�����JsA��&�'W�/�����5��]>�|Z,�6�,��Vn�:]�=ާ����s<W�>2Q	��E��@�d��P?�y���Q^�����l^L5����t��VM2S��N�R9�D���e�5�MJu�����-��U���L�9)eB��d<tC�ކ���d` ˞P-bUqIAR5�^��?tYwh꓁Ō��A,_�vZP�IL|1@���ue�����1�U�0A�������%�a,��$q�ٖ��ʋ��$�ˑ-,�e�n+�l���xA��S:?���Y�����4UR��2㹰Ȳ��������\c�t/.X	���ɖځ�)�ըT&cRW�F���6;q7�~��Y�b}�~D�����?�6�|i#?/�~Р4++�ПI��0�L},��Q�\���䬍��k���d��p2��s���L�3������ �Λ/�����DxȎ�d��F!0dC�I�D������?ܓ��ɏI���Q]�Vb=X!pyqN�|������1�����ZcK��ʬ�ɷ�h��,2�o��̣V�9��� ��&���r���T!���@cY��uL�'�I��!����*�z�/ 7��)�[�/.�@����3�,��{�9,J�	��:|u��(��H�*��V�5���&M�ފ�1s\��RڊN�b��5��m���F�%7�7���%P�fH|2,�a_M� �X�l|�({Œ�8�v��ϩk�k@�!KTuc����r������v�տ'�v�F{��A���:�n�`a9��($�5���ˮCl��W�`�e�}�'�k�z h��`��{�&�w�_��"�
�xS�	5*���O3�x��ƽ�O��Q�_��RX�p�U �����Q��Zcϴ���������A� s(�����l�̹D� ��=�U���g1�	}i��y��>��,k�i����<�~�M�+i�]̡�J�h-F����x���Q�^;���1�\���j�i��Z't�l��x�~؇2�T�H��V�'|S�$�G�nm�p:-����W���Gc�j:h��
�:s��F�"!@�־d9�J6g�ZC��5�K�O��G��9[���+:;;��oºNf�uk��ĳ�+:.���t�'���2���@wtl<I�\m.qL�l%3,����k����P+��F}q-n���>���F8OO/Ō�A��6Sn���u�UH�#)�yrv.]��;-� ��d��);�-xX�����?�y��5+��?&$�̅3wA�@@�on3��9���O��$�j0*�H����d�M�pc0m��6�b4��AZm�ފ�@P�L������u�Q»D4�G�����`��\!-��2����|)LZ�_�99�l��@P��1�m�ɺɈK¬��%g̤>ݬSm��n�;���5�h�E��ű�<+8�`�y������
�&J�#M2	ϐm!�[>*��nY���t_U�X��|X������I�z���n;��;.�hɉםZv�抛Z�b;�� 0�h�ڟ�c�@/��^w��n�ܛ��0���bl-���뼇�Ly�*�{�;��P���������e��s��k��Ȳ���h�p�,�Z#�SQ�0n�3=@V�S��b�8fs�s�q��,���|!�7�yY?}21��%kmk.�lrn�=b.�+	gEZ�%@�XR��d���oT�#~���x��%�v|����Y�S
{[�c��ٺ�9+Y��Dak���������.f���lf0M�
�� �˓_��G� �|)���>B�<rپ���ޗy��1g��	ǧ���w��C9�� �>P&A0�O�|��R�5n��b2�{\JZk��ɷ�җ�9Z�Xv���n
�!~U�	B]�n%nM�#�4<�]�]Q�UN�E�0�tJ<'${G/���hN�#`�ӓ�I�����mˡ�l�����
{��9k-pY��Q�������2�k����οbqZr�\7D`I�7(=�E���OZ�N�������5y�³�W�0~�+C��X���..GǱ�P��z/° �W�^�P���3-�'$W'y�Ç#2��L�^̑\�[�i�"���U� ���M���y�s0|�y'�-��?n�_����!�[2�$%�F�����q�=K�fY�bؒ�[�����..�a�U�{}>`���t��s����*`�}�����w6��=��uD��f����O���7�A�^��1�݊	��Jd@��po��y�:7[��xL-Jp9�U�g8�%�R�6f�?-x��5_�`M�fP4 ���T���}��s�<���Y~sk��;�����d�V7��<�`	�k��s��
Tjb�����,�?��ЋU��F�>���<�#ȴjy��p0EE�u"�,��UVK
W�fQ��Ļ��74c}�E��*�L���FA��vU2�dWЬk�3ʐZ�ހ���
��d���l.>h_�2ęʪ�覜�և1g�r��	dq�s�� ��9*��������=�aJب\��CTu�}���$�n#_��8��-ǀ� Yɽ�vq�j�H�����`{�RGRa��I�2Me�)	�J 1Yv���� Z�x��(Onz ?ןb�@Q���ͩ}w/�H<�6�r���j &s�p<z�]����ޕx�h~��ιn��ެ5�i��jm}.}ÿHY�Yi�B3�A��(���?l���q4�����O�D~2?:���7ᬛ��{1y/��鬀/q=����C&36�a���
�L^�����v��|6�I���$�E��t�S����1�;_\���H��9�J�	�eo-&�| ��9�[\�VvM�V۩v)�f�n�D��񜽺;jM�+G�����j2`�wVj	U�YK�;�f���=���q~we����,�,֯�/^`=N�;T��!��iM�|�XdH-+���(���\FL�K��P�O:r���1`���� G028��H,��:��ڑA�����b�{�j �l�y���ѽx(�(Z� �Pj�a0����p�}�c��ϵ���5Z)��_|����	�@}3� �[79T��J	EN1���驌=���ZR�����9MR �^�<:g����3e�3�ղT�B���Y���`����`�`��wu+��lBy�d"I.�D\E$[���T������[�n�K��W��y�X� ^]�����]����fc�Q*�"�%T@�BV�6���ip.��x%�xsH�ݵ�#����3=�������W%L�Mf�2�(Y\�����^�S����M�sOϨ�yf��U��d�F�jmO�bMڦ����C�P�
~F�[(�������CO22@��~��08�����K9�i�XJV��4��'�T�4⟝0��i�ޙ#�K��RP����x0%����ԜqN���t���Y��=�S�gY4���,��	�V�5x`7�|a�"��pvB��Z����f���Z��}��9���K�4�Z��W�Mʹ���d��+�/E�3�h�4(���K��`M��"��q�d�l!�M�S����)A�3�)��F9Ȑ�����
�UCc������� ���9�͈�~L]A�F�@�e,Y�Ə(��7���hB˞k�|_���f�	h�̑��t�c�ژY?9�/��.j_�4F.1Ç `��I7�M��GXm�Q��	B�AU��!���ZgV�}h��L�,aE�GNuc����.�����V�1� ,Z���:$S�ʉ���O-\���Xh��з1�)����]x�L�>!�z�F��^����f��K뾜Z�Ϟ-���ې��B��Z�����M�z�=b��L�)`V�@��k\^�l�`�Cٝ��Y�,}��QS׈����*O�H����֥�EQV���lb���/Ǎ18�&WU!�>��"�Y��H�Z��H��	��Q0 ��	��������d�]Bk�wzzBr���]k�S�.,'}�u3�=�V��>���l���_<��F��>�������)j��?=���A�9ޚ��e���SIvZ*�
\� <޿���" �֯�������[���],�� 0.;�^�~����Iz�}�?=�_�&mOur,��q�oi{��[���+�&/rPc	�U�f��T�M��p)4��\@j:oT���aB�c�.�7W�ؓ�J�X�(���z��oإ���e�D��oHM�r�5�L*v�*�=Z��䈎�Ex�;���l�T���mBX_�Y�qi�L�.曑�?q�u�b��67̵h�v#4\��-o���l}1_�0���Lа�<��흟_�㚮�ot.O�鈟ň�\0$�W�Ko/��1�	���WY�����M�h�q�z_25:�|%sA�����Q�_�}E�����g`��I	�+:g$3�@7�T�~C[�uY��7(}w�O��7V|���@Fʬ$�+%�4�ר5Rk�{�aݕ�g�21����U��1j�ղ�t|P���M�pY�
��V*��JBj�hW�#�<V�W̲L�i|�/k� x�Z����`�Oiʲ��)h��2�j�B���~B�1�.��f\g�J���pc|,Mlݖ��r�O�����=���΍ָ;�r,������H�!����ov�F S)5�:���ٺ��:Y�^��2�5Z:+�Sy���I�[L�r��J6���{zz\��3���/ZlL��K�<0��X[<b3{�X�q�8ޓ�9K�ūI\�J�77��WG���մ$3hR�*��P��As�`�ο񘊫��y��wG?�kn��?�� 2���_*�h�~�������y'_�tq���٥��*M�c+rU��]�F�D�>A��xV ��Yx���-/CB;*Y}d���~ϓ���n}�.�KK����K6�r�d�p& l!��
��!&Z�� ,�������5�0��kof;b4��R�R4(�y0A���uJ@�����%�l�Nk)6YW�QA��Cj7�N<g�ԫV�VK9q��L�����X��QbC��'�r�#˶<ԁ�#T���9L0�Ƹ����|�$�5�.s����8�v��փ?�t��c<~#�jc�~�;��G�P� ���w:��k���t�@��\�C��V���I�._�Q�,���5@�����ld��l�2+�0.ow�BMD�\�B�^ޞqxE�@�<��  ��IDAT��[`��X7A @�(�AQ;��%�̭ŷ=�@�=��3^A� _�
�E�G�תւ
��R j��ȧAp�=n[���>}J�N���-�6��&C4���Vݺ�X�N]i/0�����|�Y�&�vmD��=q;ڳm���l���Ꜩ�u7�^�$�T�ީq�ά�P]/�:	g������:/���� �~�Ϥőu�#�V��W�����<�AQ�ʽɁ��XϓNk\KK�)r����S*��.0�tH�3��Ý��尅h�8�]���eg���ϧ��'��u.Q����Q	���$9�f[���#� z��>;�ts�4�:�N.$�J �|�O�ﻱI�>���>�HzS~����Ř�dq�=@����0y��0d��g��Ж��e�778
v�'�?ҭ-��:���V�_A���!<)�Å�j{ִ}���v[��+�x�����Ah$Y��%3�<�tI]~�<�B�2��Y�����	�J�������e�n�ڝ��j�0����p'�B�Uڲ�>I�-[�?�k@̰�z����W9�A|���Z�c�x��=��Ӓ�v3�0�d��@���A���ފ2:ئ4�pݧ���<~`kV���J
��S�]6K��3 %Y�wb������&o߼���|G�T����Jې�"�9��ܧM�<,t-?�++�=��(����J��4�i�5 Kc��s�rO��<<<ێ�"�k�	�K�	�O�u�qX� 7��vM��Z�\�<4�{��4lj��5��xm �}���-�������=Ԟ�����Ek����B����~�ңŭ��}b�E���)2�	'x���3���~��h�~�L{}� ��d�q5�s'��k�'ǰ��i��Q�a�^���/����n�~��-���ӬS�$lwIc߸�.9��.f��e�s٠�~7;�� w2�+�j�uU��f� ��v�Dw׷Z�����eM10a�[����L��-c�l'�Jnݰ�����A���(�ɿS-F�S�_F�:��i���������첸�gF�T����)�G���1ρ��=>�^`�צ!5*ն����e<`���-����y�%��ZU�Q�0��=��n�W�cna+!�.�X��)s)���%/ޔr���x�I6foW4�>���4Ha���.Vr2D�V��P:{mq>;E����ͯ͋��w�j4�~&��!`�,D-;#�D��>3�w;��T7*� i����'�TW��ɯU�{�k� ���<�\
sj�.��>�?3i�E ����g�U-�pA���x.���w������_�+�h��'�{��� ^"�d��5f�f��ӧ�����|\�V�� �Wo���� �}u� p����,<ާ�X���h�|�qH�hG�|.��Ak��p�_'˦�ᦦr��B�q%˨|E9�ْ:P0`�jU�nL�ܞ�=n�PD��rn���CM�O���nlGlK�s%����x��3^g��0���O�#6(������Y���-Ʀ�g��3�ԌSt��vo���h-�ƪ���ذ莔��cv�/�V�z�,]=|� $uL9L���o�����N����)�0H�,��\�m^�[&�d��c\c����q�ڳ��K��v-�/Ys�9����z{���"�j9� xc����uB'`<����r�@߭�g	K��.���H���U��{F����������c=��u��T��o�f�sV[u��.�5�����|����%�]�ly*��<S�߮���I���lx�(�!�O�Y�/�%l7����Ќn��k���ɼ��p��)��-�������kg�zPa�P7�ɽa����q���Y�9�*��[^��������'p"��v�(�q^9�1���p1�Pw۲��C��`黂�9�MG��mv�N��:o�D�h~�b�`�Q��xM-yĖ	�!9WF`,n�t���-77�5Ygϔw����[���Dן?Ѯhf\��7n7�6��$ F3\zu�B��Y������{ט�g �A����@%JR�D����2�|���~~O�
 ������]�yG/_J���`K�n�?{Zr��s�щ�; dR���ҲB�e�q<#�v���,�A\4��U�̞��ʂ���3�}wqyA������/_詌/ߗ)H�������d����F��,���E� �Ckm�=�^�s�@����^t3�6��C���r4m���L�v�C>��5l��H�0i�i��h�� ����#~g�U�a,G�>��S8������?fh"�+�	i��S6��ƫviZZ��z�|�s�7�?�x�:*��5��?���2���/0�FF�dɟ�o�/?�L?�����y>g��W׭�K���S��Kao^G۶P�͹�[��xd��L�Y涉*p�G�O�h,V�t��d_~���TIY��s9��f������A�.029볥&>X�Hr7�3G�� Z�WNl���q*s��&1_��6�1b�҂����E�eO'"p|�$���*cuvvEg�J߯��`���65�9���bY�e�ϡ�e�:�G���^�I���K����5G�^���'��%-�R���m1~hc��$��Ww�5�uX���??@����3���54Hj��h+���2����Y+$QΥ�`l���Ԗcg��6ɻ��
![��lSIe�j��1r%s��N �l|;��P��<"0����rv��Ņl�7e�^�����%0�߻���\g���8�a����Cj���}��7��w7�i�.`�t/�Wbv�FU˽ư��r'�?s���X�8����wS¬��y�PdU��~s�gl�#3�-��~gZC��9v0�L@���<?./���Hk�2�b���wo��:>9.�y+EeY�gK��ǟ��W:6�����2QkR7����r~�DP���Z������#j��_w�?�E'~Ǉ�0�� ,|wڞ:���~�]7�~?-؊�}��o@^ �p��g�����Mi1ಌ|`����t횹#�f�.���B���x�l[ۥ�}��޽{G�}��Zu�D�L]�k)�|C?����g�����D=>>�� L�խ�V2�.p�}?׭F�p1ǅ�kt�Xoqg�,̡`i��_���e�W͊BϤ��L�tZ���F�N�Y�B*[����awz�@qj7XW�[�v�ş!��5�x��o �jqE?X�ϝt�n9�����#=��4?��z��|���ruA'��\��_���5w��2�>Qģ+��j1�V+���7���d�K(��z�:L@]5�Ð��%ٞkV?�s�N�c�ά ��V���X�=zLǉL���YuΡ3C�6À��'�+�6ͮ�Ŋ��V*���z�f��f�- ���D9�T�
p���FdMuf*v����l]ه��L���e��<A$��dH����"Y�D;�mY�		�EK *��>Զb����k�)B���˗/J[V�|��n�e���E�5���f���
n"$4׃ 4�C����` ���9fe�f���O���/�����ɩ�<��������h�B1�?!��y��-��'����g:��^_6�đ�]��H�g�����<�����V�}��AR���_�H����b=8-`����c?п���?�(�.K�[�Z�Dg&M�8+ϗ�ِ�����nh@�f�N??D�0�K�#2�����nz����M�?E8�٫�{M�ۇ����s���H��	p}a�V����+��h���r/Vl-�@M�L�J����U-�M�(8�7�*������W\�������"��П���o������(�l5����s��r8�(�LT�]+����!����k!E�k��W��������c�Rqz�B�-�N����qS�t�tl�񝕬+��\�r��nb�������l�6n��kgd�'��{��F��4,�L�2��<=�񺗠���ۢ�mDn������� ����)-��v��Dϋ�{"n�� �Q��?][S6���N�>2p&w����q��V<w���t%Sq��q���qu��qH>�|Zg�1�C[�Q9A�C�V��~.�ő:Bڪ�S}X\�7�Yc��@��739��̿)@���pUdo�uRTf����}�X`���}_ a����Yeе��"KTM�
>Y��Rl.���,��O��R����n�@�e|,�NM���9��C'�$�+���gBO��������	H�ge�����f����ýf$}��QHWŊ���|��.^�f�cJBC�{�n
<Wnޭ�]cw��Mg�^3�Rg�����Φ�v2~�L�rѩ�䅜�\��Ynd<��u|�R�i&�Jt��L�v�͕�[���I���#B�"�5K�C�}��d-�s��m�;ټ�fn>�9�ύ��N�}
آu���Z�ة�r�V����-y�8E� �	 |M_��ٔ����i%�,��U+�&�F�[�Yǣ�Yn������5��/?���t,%�z���R��_�������?�D777B����Fa���5��-_��{{ؕvIA��Or��)?|��P��>�?�@�W�DX��kaSQ�-��U/�}7t{���noi�ZP.}��Js�hQ��;�j,���a����2�̓�*���{��s�&W fʙMT��IM�_��6%�U��q_����_�'.�Gw|r^d�k`G��e�^Y>v�T�l}r���3�3&*����S}N<��6Q��:֙%)U9�����XA����q���S��!$"�b-�^0�����No3��ۯ�2�]0Um f����f�`�T&��̉���c"����t��R��;����Dm��l,�]�fI�@^b]�u���]/�/�L%a!m$i���l4>Ok��\;�{�2�X�%j�˙D����;��`s1�h�A�R��Ġm��,J ��"4uO���G@u`��z=�u1Q��:�@���dfI�GsmI��'������y�{��5���;:g����s�r�����"e�ɉ������nJ�U ���8 ���~�����D3�8	�g���Γ`���ap�b9{����O
��{��ݖMꚾ��Sy�����=$]�v��s;Q-�3>�d�"ZJ�ق���Z�"��׀�^���@�y?|��E�X]�Gd��x�S���>�އ@� �W�����<birOX%<�k+4����;��My�p=P4 �����9Z�9�\" ,x?���Zzn��R�]�"F$q@c�qS��#���:-
g.�R���cʘ�~z/��fU�t�>���V�՞:/�%�;� 6OR�r)���~�"�����wh�7Q��EW�Y�*�&.~y�����{zx��������ݻoh�\j�1[i1M8�lyI
@�[h�?J��0��A���RȚ}��q��>7�
Ʋ�C$�Y�;�C\no�~����#��q����YT��3:�|I����WE���~,�02��n$Ӡ�: �s����� ���X���+��yu��T�����=�@��Q��`Qt�Jj�F��F b��Ҿܚ*���ͼ>�9b���E5#}0���)�x&;Kt7�'��ݏ���Z@��!�y����NW-|�Ԯ�~>��%�`��ƈ |��1વ���C�/��48�K,�s?�ވK���ǻc`G�"v��*R{�y�}Q��
[�����'n$��3��R��
M+�;X�`�l�N\�ys��>|�H�7wjN�/��7����o���c߄��uK7�ڤ=�����g�� PJ .VAʁ�|�S(��b	�*f} �kf!����Ef<n,��g�~:=9�2F�?�us{��e��Ȗ�(��a��E�<FK�=0�4�g*j����i���/��OL�����?�0:�Y������"���j}�i�R�vNAY�/ܾBb�|�	�������!�8}�)P�7wN�a-H
B<�H�D{�غy����0 �����2_9��cR9�d!5vI�x������V�W��hk;:��`�b�~�)�x�J�Dx���u���hn�d.�����2��/y�䚻��x��t~)�����\�+�7�;<�l�3qM����Z��zC��oF�L��^�ͅo�r85| ֜��c���%Ŵwr�n���/��Z?���Z�Z�X��Wtrv)�_�4?B���T�W������5u����T���6�(�_��x}�=�{Uc���������hO(V���`���踺��A��?X{T�)� � �F�!{aI�Ŭ��}>�jZ�����%;�2��a�l���JA�������=��R��`~~f�\J�`?�Kɐ���k٥��',pȔ��+��:�mӊE3M��˓����t]6�?�H�E ���ۙ	B�q��)�*l#�'��~��Сж�~V5M{b]Y\Z�Ae�v�O�X�l��|x����������|�{z󻿣�WZ��y�f*��,,�h�a�㏘� 5Ϫ �� ��s[�>y�Dg4!�7�ҧ"��ڤ�:����N�xN�^�{���u��Sk���������+)7QG5�Y�DL�BL��y,2� ������C�?��fj�I���M���q���5���Z�TY9|T!APH n��.!}�=�e)����Bc��=�R�.��1^1�����`E�A:x��}�%.��������pr�N���C������yvf6�<X����sP2ǀq&�%[�%�l��DB>�vB�ݫKQ�W�2�Y�1���{>�^j�MX�����
pCKd���@�1`[��<.�����e����Ï?
�?ן==��D ^��keJf�V��a!I*����l��vtO5Y����e�^\��:Z�m��#�>;������
����f���\���<ۋ��'�/���{,syO��(�ch�l?��i<n�@���o��}R�3�"W��#PQe�F;�;`�������X.�!���kۣ�ff)�.�*��ۑC�9 _;��)����k �nl���,�$�c�?��qk�f�:��T���$j&����O}��*]�ˋS93F\�aS��V���.i�g@����O�lө��m0�	ћ�۲(��q����,��}���%��4(7�Sh?�s �ge5!��{8��? ,�8�[-:3�Yؖ�7[������/7w���z��w����|��Qnbӻ`�c�]A�Dp�V�*��!$���׹���I���KـT����_�Q(6�eC�b���?t��(���b|� Ѯ�t�T&�@A^D�\�+؄U�����*�V�{ h�G "q~탯�̺�{[�-{(N�����1T[N��S���r�{p�@A��j
ھf}C�Bs��Cֽ�� e��ѽ	��p��F��Vp}&��+p6�Ws�����.��m����-{��}ʽ��<朱<l�H�б촔�����;67��حO��6~ZO����ٲ�eɌ8�������Ky����sG��^�,�����Y��[==m�u-��,.���Q�����ڐ�V~��M��h
��ϰ�;�!r�Jo��us1�}f4�5�y�x/VE�T &��O���5�c1���N.^H���啐\'㜬�J"8'LO�>i-��P�kvV�Y�xb����>(ֵʠQc ��ǽ��=�����v�>Ρ�7KW�,�����^���P�8��aZ�y�Ȏ
�W,`��F�"G1ǥq���2Ӷ��EAa�PO�lu��ng�\M؈�Oڞ��7��1����Ó�!��lVk�\�3x�j66JbYP^>].8�f�p�9xB�9������z<��%~C5׬\��L7_N���_�h3�9��E���\\`�P��R}� ��ds�@B�F�y�]����@v��Ŷm^�����In�$������yp������7��������i.��LyUd�����	W���>e��  �<''��X���ƽ�����;&������������X���bq�PF�2��*`sT�-!Һr��>�T�)��1����s9�o�Ĭ��k�n�����5��$��x�R�y��hׯ�G��-D]�+Ǝa���iA�n�m���H��v���/U@'�B� 
����:�C�Jy)��1�*Z��X�0& ���)��(�eY�,Y��Y�a��$`���PQ 
�V9J�������L��w;%+�:�k��ӢٝX�s[�#'�����8Y�[��xXY������dRJfgO��}��V��-��w%���h�+Zl9[����t��!�RW�ƅ�b�����A�@>La��$.��39@�6�����RH����˜9�~����?	o�X������Ǒ�
�S���;͒ո��m������_9�:�T0��4e���3	�N�ĖJ���p[-+�����q=΋��fs�g����$bO��@q�n|Й�R�u��b��q�7�e_����Y'��U�/L����WG�[3�����ܫ���/���|�I� +;�ҡQ��6�a���@ /��j 0S�_,��;- �����U�b�,��M�:��me�[�^��F�M`�M�:����C:&+Ze�O�̔�K9�f�^�!�����]�&��ϢE�#��Q�����M�ёb�Lt��cez�鉳�n��g�	᧥tKOga�	��� X��\�C%s�"|�!�%;��4���+k�� XrYhE����_n������⪧�/���~O���]_o�&vJ:�V{̳JHGm�>���Ӷ�9�}*�k��y�H�b���쬁I�HA�����Q�.V��[�<�
��9e�F���`ZWK���|i���[��G�'������ܘ�s��쁃�פ�#B�Y�4��.��ς�(�C.J��٣:�rMʮ�R�#j�.Q��N��U��z���k����>b�rc%���
�PGׂ�nCp}�����Z�"A+o�(97�Z�BP��;ps9�fks.J�gS5�C3��1@�~S`��<s�	H����kԹ�����T5:����;�ϸ_��Ǽf6[Y�,gh�V����GX0q!��<�*(���)�<�LN��z�����8��d����� ~�	 ��[�Ebƪ��Z�TB�{��ֵ���/�,�P�,�|g��\���(?5�{T�')����ʧ�/���N/^��z, [��� ���iw��S߬� Jr
����ds����k`�77�Y�� ��(�~G=��Lu.M�=�`�LuJ�i��ߦ��9���b��N�٘%���0�QCP���^e;/�ԛx�G��oĿ���n�뭽,t0��8
+h���_��F!�V#�QO���;��X5���ߘ(I���y!��5�D
�Fj��Ԉ �6���&����hF���v�LV;N-5ٟ#A�b����'��f�-�nV�������|�ӓ}��x�,�0K�8���d]Pj�Q�1-��� aɹ���խ�5V�Z��n��ǟދ���ቖE�|��^�~O��~'a��B���kTN������(��l�ٲ�{.[T��f����eb:��bA�@Z4ޫ>$��8О�s֫`@6��������g��T���X���
�B�X�:	���e�b�\`�YIP~�L�gLA�<����D��!��(幼-"�E7��p��c���i���2s�/P��c*���!@��O��2se#5�M���Bmq	�B�1 ��o�0)fY�h��Z����v#2x���ub�#�>�-yC݊p;����;����5+�TT A��-��eㄷ�L�47~?Sm��]³��Q����1��������Y����3�����N���K&'j���y��#����/����V�s��� ���T^���t4�D�v��1/Tj^�9L T01CN������	Ml�boQw:����ɹ,���(�\YD���V����\�iŕ%p]�>�]�x�sR��hnz�u�a��/����˫+: ��l�(���k����'Z���:F�6���4����86"��j	蚔*���c��lIRɧWk\Ù�s�M�w
��M����9��\;Uk[@�^)^�Y7t
_�u���e���>��f��s%c~v��)�V��Z��j��;K������	mM8��|lX��Fa��v��&o�-��%��)w;�S`ޝ�����ґ�a�C����09ExV��v�}�ᅴ�jn3��h�f�vbcE|������=s}-�IN.����5����ћw�����/��0�gs�l>x_a~y�5#�{B�>QDY7w7�M���V�/�Q!�Y2R���9D��$�w� B]�V� ����\���D�;7mi��f�֙����Ū��Ϟ̶�8��Okf�����f;A=�Օ��<o΍l ���r��\�~����㈹�w��j�~t�NK"E+����s���|�}`!���,k|�F$n�)�^;`58�@M�
���U�Zh\����X&n�P"�0wj�b�C��<��J:7I0�Ô�q���q4e�W� 8�N�A��\�6�����7��>H�q=K(P~q���E��Y�*o�?-ǈ	�V��X��R6N�i�Z��#>Pb�l��
��'{m6w�AJAS����q��
�3gT��,�IH�L�깰6W9�z)�_˓3!ʕ�c1ej���^q
�a�����i�����ogc�vUV�b���5}�tM��� }=���a<(�6����Ӏk�Z;SH�:7����'&��;C�4_jL��ԍZ�����]��5V���$8$ካ|�nw3�c�>��{]\ X��&�d/��L��e��
�M�s43O�2�(�1j��4�P ĨMD�Մ�s�J�{Bj~�P�`��iB�G���
�?,[�i���k�.�%,)3QH5N�o��bP1�����LP6�G�~��-������|��hf���tR^3��1
�$��,�n@Q���� ���@�s�b�ö+��i3З����,�ϒQzv~Io�+����/_�i��V��H���W6�>Y��=̦�[�B����ھD:Ȱ��]o�j�?2x���=��`q)�`��9�%9g���EP�엲	����n�5&E�����{a-TM+l6x�����/�����אn����R�������&O�nBD~�њT�'��i�'�*�}ؐMP�Y'/�V������ԥ�
��K��=�����ಋ������ݜтq�{�N�=�7c;bF#��sx�O�\o�f��4yBc� $k����e���t<�p��A�9���Fq?vҕ "�`�A7�aDܬ����-T�7O�g2z�8o��ImLHj6��̏2��k��<I���NN�������/����>]�d���U�������h��Ĳ?Ɍ
֫D��+}�v���=iu�O�~ۙkV�]�L���גeI��y�8�x!�/�x<.�K�I��d|�9�d�ɲsh��l)�K�� 8��d�r٧���2PᤀO�n�_>�#gh �>�֧��I���AwXF�"�$�\��ֽHw9�<bOK(���rP���h$�d����n� L�Wè��<��-4_����y�n�ԕF�pF��㤗M�Yg�c�p���p��0�U�q6Z
��{�K�yg���_���h����N[��๱N"��Tܽ+�&�� Q�588n0�irAk��,�bT�o9i���.�"����zG���z8��vE�KP�
�Y,��VgM�p��cZ܏A@UW�>�`�����z�L��HOE�~xZ�-�[��`Y�1�z����7�r��K����
�V�4�Mh��M��%�3(�ڃMo��p�"(�3QM��kr4�G�{k������,C�wީj6�\����R#]8������'Ԝ_��|��[�pXMLN�/ Z6�mz�$6� �5�6��J��F�EG�� ������!����� ��),�1�+R= >k
����;��EK�vg��UK��3��7`�{�c��<G�
�`#!�_?CLYo\ZC�G\��2x rN��,����ֲ�wX�dp�ese#i�m�*ZF�V��,q�w�(��}d1��C.w�x� 0�]s�БA�5U(8�c��sh�#gǿ�*%w7��D��X����cÎfK聅����9=�Р �ب�)�p��B���n��N2w�Fm��~�����Y�'Vp	���Z�]h���[�-�\����ޚ݇_����BaM�0�y�����{���}�|G_���c-sW�┪"V��/�s��j��	h��vAw X�GoY��j��V� C̰����i����]�w!�j���B�@A�I<�V��
��������ӱ�����#�?�@�
l�n��`[ S.�����Kfe��.N�.���M-�f���3h{|���M�1�?��k8�<�NP�������*�q���,�dz����Y��^l���0a+kfw7���������BL��/��ha��F�3�Y�\�UW��d�f�R�Y���p�s\=0���Z�������Y�gW����^J�����Ӳ_i��^=�+׻����	��c�����@AbiJ��K-`�m�te�Z��4��TP7����:q3�]���t�5i��(�	(�Qm��̉�O##d�J;�h� ��Dz��u�7��F}�C�Y-�.�'V>,��@Kk��*M34�~�Zj�֩���W{ع9��kf��L-��׾�kO�[�g���FȤ��[������ɪV���2$�ðk�ْ�~$d���z5�l��� {r�j��`Q�z����ݦ�����^;��;+��X��]dx?��Eni60"��tZhF�Ν�.���d$0�F�G;����ڼ�~�*�?���Aס$/���(�EW</oH����
���ϟ~���t{}M_�$C����e-g�&囓W�*�{.XS>�r�:�l�'el��<�KV��y�=�����9�uR@[��%����$i�Qa�e�Ȍuw���o��hzd�ϻɵ�=�Ӛ3[G��.	�������Kz�����J�h��\Aso�ӭHma�8��t��T���zԩ3�Y�X�I�^�u���SE�%� �;�֥?�������0-�r�0T#^^��f� !� ���{>jp�b*=��3���I/q�x*�Ҷ�Mr��I��dopu���pP�j[){'V�ET;$K[�!vޞ��Kz��J	4��O1���kU#�v��s�&�\����e����/��*�l��2y�L���KNȤ��F?�1[�9�������Xj���7���f���pW���v�)2�z�����GW/_KOH��r�e,o��Ԍc���>��:�ا�0qm#%K��f��Kȸ��ͨ��o�X�sM�"X8�X�Ac�X8�6�%��|��L@�*l��nEǶ�'6��'��Ǎ�C��*���r�Q7���N-,eS �~w@�K
C�L��*�DE��������U,`�yNA�L*
r#H��-a���Z��g��U����ش���q��ێS��UZ�M��%V�ypAg��b�J�.Օ�Kb 3೵�-�GBĺ���sm����#q��zg�_yCDi��``��y�n��*�f�L]G��V>T���D���I1|��t5M�=F��if�	z�,���i5���(w�q(���(��y�6��ã�w5#�{�g
:a̓y������|�?�)EV�17���M��RQ�y$|u�#s�i��/�$�=�.	�:1��������0��?�8	m�n�p��ġ��6��>�����T,�����l(X`����H�yɞ�d�^�`�<���
$o�W��5�q�Ry��� �`�F^3[��h9S�v�!��;��Z�MNa��X��<�S�%ָ�@l�sV�c�"���wA�u	��\A��۵XF �ق�/w&kkm�rƆ-sKe�׳uRf�0q�m���ff�'��A����ʚN�m�����r2dF�Q��Y�v�D��7|͢D\�U9����@xH�w���5ȊP(}ԯN�Xo��������R������d���{0f�e�J��el$[�2����f�ՠύ����=�l&�#������\^	��j��.bѳ*��l.���FS�W�0�G*4zI�
�&n�K�3v(v������䛘f��h٩�����n	�,�gy4��E=9�rZ�8�ɔ�+��Zfj�&e�d�sU7T�=�A���8��LF�t OA���t`�m�V:\t���@���־�L�5 ?m�
���X�c L��L�z�!T���K�s���)/*o�$�/����g/F:�i�=b�⫺%�-]��bZ�v��%V���U]U;X����V����e�ʣ�I�ON����.�l�ٹp�1 ce�闏�/���M�磀/.˕�E���")��҆N�ue4�D׌~���M���]�U�T�f#���%5O~K �&}Ρͪhq�ꋫ9�NυO����n�|��������3�sA�h�t�K��]��*U��I �S�ʐV����k�56ONhU���^��J�(��q��u�n�V��w�������m���ɧQ��� R�%���3��Q�SF�Ͽ�,nӫ�/��������=��lHi�`��>�ߋ�j�Τ��c�%B0o�}�#���\��Gb]&1�Шq_n���?ֳ�����x�Ї-WF�\l��yLx}u�=�B�lޚ�kj��@��;�S T�keK�e��l쒑׸5ӟ��8�eթُ��C�ڣB^Y<�{�.o[����P�E�a�{�o>����"���9qɄ� �yQKPF�гg\ ���@�W���2ʌ��ؗ���~A+������Ni�xAw�_h~s;@ʳ�ҏ����`��n��n������qz1Oy�s�����䥬sJ3�L;�xI��p!��E8��pp���5R��� db;p�u��/�b�;�ࣙK�q�9d͑p�,;��q$�<K]Jms��4ӑ]�ge�z��J
�UQ �L��Ge1�f��ǹ����S��@(7��֩�\�Ʉ���*a!�+�5ֿ�^?�{�;)��h�Q!<��6�pz�u�\54��:�� H��X�Z&H��ngE�'@&Z���V��6�}� �Mf������a�xU�n��p_3߶���<K�����&�dU�H�Q���q��Kݏ3_���o����`�X��������?�������H_��Ǖ;�e�J� ki�.�WkU���>�,e{���
V �b+@�=�W��b�l:�mѸ]2�k�.�Dˢ�����Z��s���B��m�ܥ���(��&kмdƛ�(�5�B6!�s)�!(��לk92���߉<�`�
�#����8O]'R�]�3i�N׹�����u^+��k� ۖ7>~����z#@lQ��y���^4�LY��s/k�Klu�V�>]�fe����LjX{��S�$�syzT�Di�����d���`:�g��3K����n)6^��]��}^y�OW����T	�%}�w3�*�h��kDY_�R9�,��P�hEL��<Q��qV`3L6�ɣ�H�9��8�޷,��yRM�3���Ӧ�`�_4�i\��h&G&�Dc��=R�fZ:(��M\Yx,l��&���4a��s�
%���S%d/e1b�F=��_K�̊�s2����]�]���M����&ɋ-Y�#�Ϸ<HZ3bf*AdA�����º���qpgW  ���0h�f�$b&M�WY���u.ֹ�Rj����͎�Tb!0����];��r��	_]����}����}}I/.���xi�ic�+z��]^�ͫ�����~*��{����n����[��9���
��Q(|��������T-K�Bk=O^|T�U��P�Ri����G����vѽ�C_�F��`���@��I����ž��`m?O�Ej�� �px���;s�������*�v�!��Rr�hVW\�b�;�}����~�Zһw���#}������G���o��������?�@��/�^~�H�|�B��k�d�{Vtp�a���	�$mkg�Õn�rğ�5�3��!SY�j�����z���� @������c�Ҫ[�P��+���<���J�ƣ�~�l���ҵT���3�4�I��r��.r�]�l%b�[`U�L]]z]�����XJn��=31<���=~H&�U�w�Tx�e�"�k ΎDYx�<��2g�����pU�?��U�K׏��J<b�2��	�){֗�s�C\�o�G�Gank�����7�9�� �WFfVfU�I�gzf��������>H�*�8�`k"�jf@Du��7^F�p�`�&�**z�}@V����H�
R�Kzt��]I�6{r�Ÿ���":_���f㣶�:= K�/u k�-�9b�'�}��z��=G{Y�h(1S����<"�x>j�������zH�o$�J.�u��c�:D\�Z����ҳ�+�����@�E�'����8��4��(�g<�Y���X�YxN�x�b�1�e�����ץ���|W�*��X�l%�don�Q�����1��
�AJ�׿�h��s�(r�ōɼ^��_S�fm�/�B8-$]�Zn�|���^���]͵'�az��Q��i
.Z�_[�J�l|7.d�u랣�Gi���>��MD�ݻ����{��)7���훴Q�����v����������k��M<�c)�{��f[L��/�Oy���u��7����x5pQӐ!S�����c�`�p��00K9J���xyl����,j�U�ḶV5@�s���W��Fs@=}�G�R����;k��k�\8[%�V ��I�wn�D�jY�2�.ƪ��*��mn����m#@�G�����(�����v��pO�ގ&��](B4ӯEi-��UM�l�ɀF�mx��� ���BM?�@�[/�q��6Ӎ��J��ytjO��x ��P*$��H���S�X-���ޥ��d�#Z��}��TV0ު�-�V{�s[��1�����33�6��)�a,c�v��,VXf�Wa@AS� �I���O*�߿�e-�~�hC��=\�0���5�l���a���k�]`>����m���s�-�t�U�z5-n�z������~�6���1�6`Og}i��gboi�3ϣe!Ί���r�v	�w��?
��f2�>�ѭ���e�s���77(m*��^���A<���X�|L5����P	��ʣ�+�$�>�` Q���m�=��F�K(�$z� ���+@fd��F@N ��Ji���4!�Xy���5.�4f�){Q'~1����^�4ʏ��
�r���t��5���!�t:���Yu��X_�2]����Ղ�=J�?7�M�����z�+P�Q��B,�u����*��߉z�g�����6�l�:,��^w&J3����AI�b?���R��M��n������{������f�!���0}�N<�8M1�~g�C�V��J��X��;	����E��M�����虈�:G��0�+b������ɓkkl��u�uSG��T�6��</U��z���rݵ.G{��i�li���\W=���u�$�*�'e|<�\�5��n������U���C�R�5�s��u�hYNUz%w�����-=���mڴ0�hD�h�r���9���
m�ǧ��Z�9�ax?A[<[HϹ�\�VEB+q�L��UE����V$����(s���j����\�?Q���<�肎p��!W�E�1P��kZ��^���\�ͼZ��&3��E��1���SkM��6�B+�p�����Q��v~�wZ�,z�͜�Lį�[����v��[q�r5.�Z��!�p�!���c�C���������������U:��ޙο�NVQ�˞�r�vV}
�� ^T�zs��Ev�����W1�}��!�&��G��Y����Y)��L����%�����4�5�)͑�,���λ[�	�D�֭t@�6�l3��i��R�c|�V��4���	�9a�c�Ѵcc$xm\l�ÅW���1 �4C�˞`x���'��
aX��Ff�n��5��P�D�)�2f~OoU;h����$�2��=E:�Hk�2�¡D�tF7�b��y	:uouƹɟ.E�B�����}s�g8e!*��C�!�b��7����k� �K��g�3Q(�$L�C�(�=�N+c���
�NS�.?�������<2�"�ڞ��̻���P1��`��rp�V�����y��"��y�����ӣ|��M��m ��\�x~9=d2'���{��y�p�f���|$� �q�����s��|浨�L�����U��L��ud���[5]Sz2z��ys��������ꈩ�악�<����g����u�"� �>�ߏY���(m��!�:65���[,���S�}o�%���>��#�Ln ޴|/@�n�3%	�9��1�B:Z�ͦ7%�Ʊ��3m�H7�?̖Dy�D\�XրTV������k�,�L���G}��/D�̱�2[�X���n�6k�@T�q�,�*_��ޯ����U��Tvy��\Pe+ѯ��;˟ِ�������$NG�qK5�Y��Жa ك��kC��q/�ן8o6�!Ǐru��������j�&Z�ў�*�nՠ{`��.�c��5mL[����T#�umO��kb\I�o�S95f�������H��3e+F�~$����7���??i��C香Q�A>ģ�8�v5͗�/  %�i�hT��c4�R��C�6�U 3�b%c�q�J�>����WN��b�z������Y12GT��b�3NSN�?�f�� ��Y?g�1�TO*h�ˆu��Wgל7M�*Pr�b�\�ɧmA߃W[���m#�^�j�;�g��[e���F�bvH�*G�*���j�|D2��Fi%}P}���	�}���Y���+����W�EQ�/i!��)��fR�Z�0�[���)HU=憗A��������p�H���[�o�9������}#� CZap��w�=�@�[�n>dS0T�y�5`��Rg�{�=�����gǮ?�Ꝁ��L�E�}/�N���#Q��=O����U��s���3	���G-��ǚ�G8��V@��4�F.�}�G��T���?/U��~�LǪN�:���H �p�T�;�k�����o=+\=��=���D��_77�U�m��&d����@�����*�vA�x"��;�E�!0��ѵ̩�%4ENs 9_���lI|Ŝ�t窷��w��0s��!�_y�b4�Cn6��f�Xcv^�B�X��aF�*ɧN��<V�IuM:X2�ffYᘭ3��|}��o��z1Z�Q�Z�"�h�n)��i!ը��H�qTm��<�g�v�M�������{�o��_��[��9z�B��.//y>N����]�摊�][<���~fY���/w6_��(�e�%��I����%q�ɍ�}��f:�=�����\\ݰmT��>��	�z��kI�N����@ Rj��I2��:U$M�;�k�%��bh���*����Х`�J��)���\4��ے4֒GA�0��6��4|K��G~��dy��KP�L4��ԯ�Lr-7慳'}��SL1�7"� 5L�h�J�0�(^F��5F.�}b�#z�e�����:��C��.�g� 8��p�
$��K�|k(ǝz�*�<��ٸJ��M��0;�"z夏��)���I�L9��7�6h��qWHط�v��j D{w/�� D�Ҧ����_~�ǇrA����\�&/��F�c�*�.)#������2�<"�NJ��e//��c>v9�z��~��>��1��y�x�Z&��|k��y�����:5W�3O��@L��X�W�y8К���s���ծ����ÿ���5 ���4�Zx�u�;�r�����qX.;ާ�n/"c�y����)c���8jqDk�jwO ��B�䅁��!�����Μ)��[��i�.�l�9Dќ�ހe�v�8nJlv��>_���~�
0d�[�P���eN�g�"���(�j�wv��d�����V;�b�_s4�J��� ^(v[�|�}(�q�~��z��W�Y�N ��>֛�eg�"�|��Y,$�P$u����ߘ��W"~{s%��ܘh��sp.�\r��\��蕠nbu\�������ׯήQ���q4!虝����
��~w� �O[v�M�Ǵ����Q�� T���r:�do`^&�;T0�2�i3j���0C�e�h�$�a�Z=��E
O<���_����`5������3ꬠ�1y���&�E"U�J(�m���5���\��J*X�0h�,���������9����}ͼ��IM�2Y��C���W�ʺ�!5a�4s�#Zї�< ��#TL]
f��k!+8��7���Ҹ��~�=�w�ş7CG\��*��6 �8��֟(�
Zt3V�DN�c���x���'�OOr��6�]/�\`�B_�р[c�ª�\�·��G��v=*�*9�Y$C�}Ѽ-�mh�����v���-�'\7j��Ƞ�/���؏����>�v��/�\q=����L�I�w�t�1O: Aħ���H�� �t$�E�#Hx�8�5������=x�Vܞ2qݫ���y]��"�ZSk �� ���6�EF������sL����XIr�8��s@Ǳh�����}\y�\���дmh��M�Z��.,�o��
��9�5�c�{9����D|1�`�93�0scc1/>7y-Mm�C�yee�;w |A����4��p@��)JQ�#:{����U;����Y�u�(�(/l�x��2Yl6;��)Ų�'�W
���;?���&����,�  ٜ�^q���-Ó���Z�x����ӿ�$ߒc�������� ���G�������$��R,6�LW*�uT!ۋ2���mL����s�^&�ɩD1�#����H���{��.��Q︀�H�n����?����rT�wh�p���w�O`�YBM���B+sc�v f�H�!1a���*%��eJ�8z3L؜@�g�����]��9_�\����J���`�ME�u�Eۆ��}Ǵ)�=�6y���+�z�A�qh�:�/���d����7u����sd��u(��nT�aڞ�4KjM%�q�_6��:j���2��+���X|��ab�&�h�3S21f��c�vf��+/�q[yg}e���8����o_p�U'�Ҹ/L�PE���|x��5�b$WnpQr�F�Vq�b>!M�j�݁�J��~{���該�Jc���fQ�7�ʣ�k:ʠ��_ޣ��h�,�{����Q'�� g���dc7���TYQ@U�1}��%�,R����ѡ���eHL�4R��*ڟ��U��:��E?���4%�G��T!uu�߼7��O�d}�A��s4��ő��)�
�<�#��Y;���[��-H�c���<\ثN��ƺ^%]��0qL�<-&b����\��Z܊H��G�*�y��c�&{�乖相���gs� �|��e&��e�<?�/���������������\��r��e�78�g 쥕�:C�R�$-pPq�E�e-�Q`�{�R1��������B�O��<����R&��]�>���N��^�A����Sl���r5��k�ն6l�12z�\�s�҇���:ѡ8��_$_�[FF�����Y��6��|��<?��q���d��;r}u#�����m) p hy$h@O'����,Oۨz�OJ���S�t`N���F�7CI��1BARt�JG h�ԅ���B�S{��#�>��J�b����Y�0��{�o�r����;y��o��@O�"�W����C�U\_�=ݠ���'~���Ѱ��M�GVq`\�V���[��Ek�
 ��ӷ�eU� �zrM��za�Ӱ��kf,�q���W� ���<�^�����[�����M&E�f=�ߐ7�ƆR�bߍs�9���V��xR��Y�m������H�K�͂�6AT����~83��'�N�8^x|~�0R��Z��0��R^n|ӟ�5������1NH5|��y��� �$��Rէ�=�ҕcO�����5�﹜����T�L�{s~^�����*TZu����Ǳ��y�d�����?[_c}_�Ƞ�=��A���_���&��q�k� �u�<�7?'���3��r��R��j� ��h���Z���9bJ�C4G�aN_ё/�汐2}|zN��%��zWM�ϭ���88rP-�2�8��^����ņ���f���-ǚڹ��kz����g�#ϟ��������s�_e�'�TR>x���8ZļD$���q�y�,wδon��d[����b�5�H���E{,�C���X����1ʟ��Y>}�?��_���Rnn����޿{'7W��I�e�
� Z��*娵�De )�ς�ن�*@�8�q�Τ8F�9�gM�6j�
O6���Q�3�_At�9�G䁼��-[�!��ց�i�v��|��[+��^	����$\���6�ju���Ϭ���o��֣���r`�h`�#/�曤�-`).�S�?��U"�|�tR0 Vy�=Cv`�{>�Xy���,�|���Iv��|�6��YUu�H�尩�$�hzb���S��[ɪ�u�/�����m�,?�sz�I��@�	�UX&�Ƴ�x]jp_B����'QeO^{��iRSf��������,����l;_y�x:T���^�2�DK�Y�d_�[�h�����6y�'ٝ.�54���k���^f�"!5a�}k� �bK����t���1/�b���w<Z��l���|v����@���
���z*���E^Aն�XZn�,�,cB"x�|ڍq�P��͔X΢\�s5߫\s��h?M(Ͷ=2�.`N֯#Y�c�Q)?��89�U;>�b��5�)�:��������WB:�DQɲ6<�Z ��52'O�c�j���<ߢe�}�W>�^�A��Q���6�L�p�mNOv���	r2����6$a�SG�����Z6�?w']_�Ղ��(�3�����0��������r�}n�T���3�9(�wޙ�l�q�W�����D/�/�r�A���Wv�?��s>OPQ.����:P��&��*F#X#��4oi/���0D/��,��o?���j���y��A�}{�H ă��9�Q�	 �9���(>]��3���Ӣ��b�=�-b��2��
f�,K�׌�p`[��{�jD����Ϩm�4 Zn���$��>y&O��=����l0��E#�K��~�'��;sepS�s�<���H�����Br�d�4�p�{Bf�{� ^��YުE��N���k�X��3�h<&��[py}-�~�k�65UϏ�vD�1�q�A��5���a�j(��u�x�1V�
 wi�W�-y$__koĉ�m��^]�B�Lɘ9?��ʯ�ߜf_���W>��{�����A�2��8P��}���d��ӿ%���z�.Y�&���)��a�������at_Z]�y0h?;�V*)@l�����!{�`���M�S6���ԑ��x����8��4�{���96"�"�$t�D�Ʒ70�7#G��>��l�X �_G6u���9Nv��ȯ��1�Ѕ�"m}��Ov��:N.w~V�
ȣbt<��#S2W�¸_%+=�z�_G�'�k�4�����ùk"��i[g��6Z���������:×h�(���<r`�y�P�n��}�n:`b������a�s�NQr�����-���>�2�d`hq)���'ӹ%2��������4E��'wk��[�$;N��a��S�XFS����H��>��#�|0w�b����U��f ,'�|������<v�Y�,�� `ph�	Cva)+���#��Y"�ɦ�N�=Z��
����3ґ����x��1B�P4�w�zB���*�l�u��&vʷ~�ot�>4F���!bvA��]D8��K����k~��@�4ʕĄ� 2`SP<��ɘ9pw�~�����Ŧ�Rxd���f�K���?�6�<�\��*z:�B���|�"�
��)'�Q��
�%@s8�5��ݝ|�� �/������ ���ay����U��qS��8#��-���Z�uP`?�Ӱ!���
��&��U�vQ�c���97'�:���+���߯k�\�ȫ��?>���:4��K7;��$�.U�kU#��Rr�o��H3~���ҧ9��#��{��C�D5y��ɖ��������+$�"� &�dM'Zwm;��rO��k��`�ۯ(��䱰��=���V6+m����֬��CI���J�K��泥f��9�V9>ql��P���_����W=�Qb����{^����Kz�&�ב�Z^�ǹ�
xR05А�5������{5?�:E\�e�y_�)��6�+9ujd{\z��|�����ȉ�R�Q���T�s-`�z#����d�К_e���V�d���$\����5���߿��'gz��M�W��b�9����Q�3?�L�2���;�8;�����3>��'�s�W�����W�?]A�b('����8?;�wVq�;|ww�s���z��~w82���p���ٜU���u�p�ҲȮѽ-��ߦ4;����Q�������t��t��Ѡ�%��)���MMp��v�6��P��mN��}Iy��6Qm�p$6�3�d�g�(�A0�Q�Z�;d��	 �J��- Ɠ���ث�$H�lf4�:�Λ	���]�U<�>N�B�p������za\����e�ϣL>����t��z�D����j��ait����B��Dln�c����.Le�u�����c�0���ȯS*#)�g�9���'\���+NLy�ڻt>LY:�D����z��y����yd Y?�WT�����/H6��dxu����쟽�%s Z?z��#��\�EG�n`��W ϻ��X?P|R6C��cZ2z���a�O����G'�Z]�㳓��Q�b>���EK��+�9�R�+1��jS�S�uZ�>�(��;K�l�_+��Yj����W�A%!��И�NA�HU	�;���&��le�Uuo��:��r�_u��� �F�Y���N�Hy�*�Ƶh-w�VDu$����װ�]?WWO�Ǩ���կk��?�T?�����j�el�Q�S�n��S��E���t�Xsy��� {�)��������9l�w�h��ŨE��S����3��7���aā�G����bM�=�� �2�-x�z~�נP,D���S�=~�8Dԏ�d���B�~��䐝*�*�_Gb�(��nc����zQZi�Ύ6��(/��c�Q��)ݱ�h�߿���FA�������n�;[ˤ1(�"Y$���{hM�^�;0Ta�r��D��1����ұ��4���.~��3}�z���V�F�ap]����.WP�Xj��Ф��|}`��|(�D�����἗��z$0�=>���#*$s��O�Bv��7SD4.��T��\�ֺ���e=����J�u��h]�lf�h�L�
b��k�a��f�R�<)�CV�g���Hm3�v�I��ix�!���b3��3C䎅r�M�׆�Z�q�y�iҡ�b�TD���!��
��]'kp�X�iI�>:���������+�U8�B� �fvm6K[�������n�P�wd���T�g /�)r7����!9y#G�~U�G����(w`��(u0z�+s�	`���FZ��K֪k�L�����Ʀ@��H�u�o���3�Befת4<04
_.���l��֢�Z����a6�����"���l���U�e![�Wv��,������+��`�D��?�@#Ld\.����5�k�j�	M3��Tl�G��Q�:�U��l~��ϼV`�G�Bi�*)Fo+T�v:�q���^
У8~�sw�6ZV*#��K~�������0��M��l�"���/dk��{�Zԑ\ɞTD&�Й0Z��Q���*첳m��� �	@�O�)��Ϧ:�U9Q��)��� �_<p�i��U�{�Vs��e��D�&���vKB�v�]lS���:N���S�$<m��v���!�k:L���׭\r{�Q� H�xB��z� P�?&GPH��H:ڢql5��r`Z2�
D9�VM!Z� ?�ªqw�$ح#�G1=@�j �"�pm����	bcO�.=F�b.c#H�B�Y�e�.���0Я:D�q�Rr���*\���,'�^�l��z�\�J�!ku-=����+2�6��D��9 ��f��֍\��+�Fy�kAxs52B��9�[�8�kY���tlpڱ��G4�=93�8�0�*�&cq�+5$z��F�*��m&m��fd�-Ej�j���K�yD�/̼k"9+�:E0���M�^]ԯ=�/4��T,��9��c��)�YE�\>�p{^~���{\��ÿ��W��F�ν/�7��B�����O�`�%'�G禱6 ����wsY��G-��!Y-r� �bi�l��F�}�A;��3H��>L�����W��F=��QQ�3�("n ~�po�H��<�~(B8�֤>�Kk��c}����Y�����q:��#��uE)��tf檥�XD���lԼz��fU�$R��Ȋ�)�~(�����Y-��Z��E-��M��Yۯ�b�k�������#b�<"�~�%�q����o��sp�m#n�d@����~l]^m���=M���x�1�l(�-�����`U������H�O�!$sr�e���؂���p��e���`�-S�)RR��U{u�Q��Ve`_��b툖���H���=�l���ȣں��0�ա�9������ZfG��ֿTd�^d�;f@|_Ҧ��������Ŏ�9�\�d0��6��?e�F�d@@w���E�"a�ȹ�\�C����t��/�zO˽�=OM����TbS���cZ��h@���g٦���Y�����:�}�y܁E�tV-M����gt�� ���\$�uA}I����c�TV���OD� cX0���@'	����A��6 �^#W�|(�����3F'}Ɯ^qC�{�hX';Z��W�P��o\=����E�*��Í��˒ 
Zg��wG������O�β�唍��^������fe%f$hu���F0xٺE�M?��ua걷��>(zԴdh��f�!�XQ��֍G�̛�ι49tꞳ|������Y�I,ϗCNf}��-�#����L��Gu��r��DBYb��0�#_��r��9��u�!�� ���(��v�j�Ki����ۘ#5�g����4���"Z�r��r�T��M����ao�F<B�N�4�_�?nk��8��u��)&��N�٬(�)OT�z��f��,��Ϩ�H��
@Za��~.y�:*S�ni��|�F+��>G7j{�D�&��kFX��c)^m��Kʜ6���b�ύ�T��Sy���O�"��$
U�yZr�����N����z-�׏�#T��V�Vx8p!x�y�"�i�d(��S9?���E_�������;y��-�
�E	�o�b�����N�PU|�����s@),9p��NB�S �F ��l��A�u�v\/p�I�E �)��kf����]����XN�57ux��A�VA����HR�����Η�iz���lp���v�컸s��)��~����[㜗�>��"<��+Wr�@�M7�̥�W!�ۊ5۲M�����Q�C�:�^<ƓP�w���j
x��?*Y�0�c4���n���k�Mё�Q#�u,�ejs��S����`�ȉg5�5��"��RJs��q!��g�a2!#@�,�J?cGXF�5j�/�o�6�3ى"i9��!0��\2xjT����	\t�I���kD�{�58��<���4z�A=T�щ����ߨؕ�L`o��|� ?�"�|�*7o.��j-k�5�F�2Qc�n H�,��ҷ�ǆ���ݼ�2�UWznk��8蝑�LƧD�:��U���ǡ�\.����T+�Yxip��@b��tAY�h(O��-_���Ҕ�e����à��~�y1R�C����� ��ԡ�K���* �D�\#�@a�˗/�)�kl0�l���L^@Ҙ5�|1c!��TJ6N��r�M����F޽����pϘ��\�U��=������C>�߾�wdʉ�\�]��2��-�a������L�(bldo�{Og �ϢC'�#�|�C�2��gkՆ�Z�K���L�⺺(�dh�F+85�{d�fD�{Aߊ.L��WUϋ���9׆�9F�ش9]'R����iW�"U� ����,�"m1?Ǭ]B�����4�\c�S�~z�9V��p�;�����$*��H]�tv=7�it���&���?�A�������`X{@rv���Q���_�����ϟ���{��j�.��Z�v�c
gR+20�JnW�^�Ѐ
�U�-�d���{�n��Ҥ5D�쾢�T ��-1؆ٴ@�s�s9cU��W���HL���Z�[��q)�
�ٲ�� ���Z��uP�u.��U9 �G�[g�qb!�~Fk�ǧ¶�*��øb$���p2�>�)>����P�Ȯn�A�h7�:�C� 2g�s��q�������u�8*�,�UF��,��I�{�9��y���Ë�x�bc#]����xz7���P,�~�lR���U�����NK��ι����4�p>;ǖ@u�|��u@�a�ްT��eg�Z :r` �r���"�Ht�7j:r����6Ci�<I7�E��U�ft�� ,N�	��= ��FM��ڦ�G�Q%�ҿw'a������[ys��E3R��U�~�7f�tӈQSV� y��"+A��|�0�E�N��<��B��7&�s2n��ʁSpT����� ���$70����ϹD��Mܘj!m���pS�O*^Qm�"�iy������A���-c�?ߘ6�䅅�T�P9�aZQU*�>�':^�`�������JX6Ⱦ�4��@�aA~R���@���(-
Q�6�QV#ߌh���W��J�g�`�	т��knd��}C`��O�?����/���`!`]<��(��%�)��	�qS�גD��I��jt��	`��W#^�R����*�z���K��6')#�P5��d}C(�ȼ4�u����tʃ�	3L�;�1�ظ�ZG�^�P�Z�W&��j;���Ԥ��V�S�����눹x��Wk�:uY�2�]���J����y��x\dN��5�i$���c�8��Q���~��0?�;m��k�����_�֔�Qa�46�$f&D+#�����B�m�
�-d�ਙ�����Bgr0��Oi--����\^������u&�ɞ�ve�x��x����ˌ�T�MK� s�(6[�'3���*���Z�/((B�Nd�����lӡ}8p e��q��W^So�y��� أ� h�t9t�,��K�ӹ�} `6МeDT�`��uo�=�u�<RjM�[�ޟ��do��
��J�䱲51�G^jK��0�� >*{Ei!|G4�����"pL���@i2�q���q�r{�}��cW�^`XVE�}.DK=v��.N)#]�aDZ)H R�>�OP�x��.f��[Q�e[z��q�.��V@����$G}�r����ӟS �[d�i$�=�F�w*��[?���N��u�ۼJguP�K73������X/�_2P����Y��������o����ʏn�j���"�&Rn)AlR%f��x��B*��'Q��*C��{bjk���[f� /��!2J�Q�9QY�ڙ�z��7��^w��,�o��5
�c�5jx��J�ί���@�	��?>���}N����6�FR�P�r����.P1e��Os��N���Se��X���.�X�1d�x��?"_�w��O?��o���>���;Y]�����."r��F��[�\��Z��.����+����e�3��_ ��w����&m\?��#zC�^�{���B�}��6����|��y�a�e�֜��{E��|)��7m)^q�4��������Q��&� _P*�Q|0=�:��wi4)���Ȯ��Tc�">p(%m�e=D&���1f���^%-+�Kd��+#kN�^V!��kL���	}~���ѯ���Wi�Y���j�KN��
��9�h��Cدs�i轿�����XzBj4��a�EOƇ�{�ӫ��_���M�w�}{K"�h�ݥk6i���"J�R�O��jU9ČU.��������?��Ԡ���_(K�$V�.d�Z2���Ⱥ���5�����ٞ�c�Z��Ta��|\:!*� ۰X��xn�� ���W9ȷ*���"6Ж]��sQ���f:`d�yA˨������(��ڐ�������r}u�q�������Cl~GO�y�4_�w`�mO�ud�[sDe#�T�~�21 0Y2�v�<� ��(O�	'�5Cfl<����-�h;�4�FӚ��7�-"tg�Z���������w�3}��w�(��2�	��;�x�B��9�v����q	aS�T��F���@����_�O]-�D�ū�0��O.d@zU	͙Z@(������G�6Y�d�c�2L�(�GZ���=����N�~�����%ۙ�52`h�����Aw5U�G��t�Y�����eC���3�[�^Ӂ�4���/	��Vӑ2Z��š 0'O�(�w f����ּQc^c��w�da��0��&�jĠ���UhJ�;,���v%�m�V9�S�g�|żert\�����6z����a
�T%��i �2�bm����t~���@$H�ca��3�k�u^���fDOr�Z=� �k���A>}�*�|�Ĵ��nǟCp�f}�� �aa͘��5�\��Z�ˉ�:��{��}Z�YwL�}���|��A޽{�+�ކ�����	R�Jy�r��N�/���jm�ͥ�qg�+=d�{��p:���i�$�j,�ҙN�o<�M��;��W�:	ڀ_��� F�4�R��*���-�AScQ�!7�cc��D�܁�#n5�J�Ǣ��ʬ�j<�XG�j��׸Z��b���S�u4�轅���bt � �7,֜J/F8�'W��5�ȬLl�4(R��?���"e�E%k���i�a�߳o߉�ƢJ��mP�Jc�{�qgMA�v�/�S;:f�n��	m��҆~�X����K�'H�鈞�vDQ9��m�^45r��1�W+>�� 5�h��,ЦZ$0�Xlԑm5D[ՙ�-G/ci�̥:�0�Ǳr�D�8@��~��5 F����G�>o���`@3���u4PT:�i����g��~!�B3�8*V�d�XҶ����*Z��E���7 !.��]�.�qڟ"ES��a,�&��9��^���<�I5f'��-�Q�<�l�H��n+}��̩�����Ų���1V�� l� N0P�� ""��6jdX�W��>�*C�ZD�����|�����4�;%�!ڂ��\ڤ#���Dn��*�$=���T��r�K�I�v'��Vb��$q���;s�mqT#$��r|ъYXȘe�����
�ҏр��Iv)��?�����||w-�4�O���Dg��6){��V�0z����o4~w�̍P�]x�C:��O�A��<ӐA+�u�:k�[mH*���	ahM�ǍN�;��M�g]6�F+F�'�b ɍw�.w0�tG�6U�&�]C
�7��oq#&�Rpa�.߷дW�a'*΁��1�A0���1yx��y �r8�r�Ϸ�Vl�"�6�n��G��*�
�� ����l,}��K=O�}�UkIڤ.���q#���;�^���1�� _>�}:�
( <��(�Z�9WEO�:������V$���`ʰ��r�*cof<�t��ŝm3�H,����Ѧ-z6s9��VN��Rx/���@l?��	 #79��IJ����A%�
8�ﺺя���_�x_�#B <\�����G#\�Տ��z�˕��}޾�����rP�2���["���j������ U�7�>7n3�z��4���h��n{� pJ �_����b*s��#��=���Y>�����N�GDFML�m<����@>�RZjF)K���E���F��C�0D�QP�����\]]q}�;����O����}O��ޢ��D�-�Gy�:fZ��BV�#�*i�Cz @��֢?^��-���U���ګ������I�4g��E�/u�ȝ��S��� Ο��4W����0:ed�9��WX����}}���:��V7]Ɲ='0�-Y=锪��a�ļ@3�_Ҹ{|N��gƘ XH`u��I�bC����r��ޝO�JF�>�P3Xq�f@ZNخ��݇��c�F���`0�|�R��A��\�=*]E�-ؾ���x就�[�h*��@��-#���POh���ɵk��=栟�*��v����M�6��g|�HҘ�F�M�X��x@Y"AS\�(".����Րc��E���gX��m�ўN:�����[ؘ�6�M̏�4*t�4�Mv��߾� >�F�^��8$	@p8X�UD{��MTނ�)Y ��XnH=ot��dt��p��l�95i��Ȱ`���&�!J�Mo��6)����;�3I�������ij�OV[ �FO?����q��xe���qc���Z��<7!�\����&q@�҈���lt��@���w���&���
�^���Ö�Ǉd,�	����p�|<[bлUÅ��H�ba��#<:gX4����o�G���_�߿I�"$�}'�	���?==�/?����ݩ4#g���F�k<GeW�L騣fZ���׊���*����d�'����|������z6�a(Q-),	�y��_㨍�H�Ѫ��]l��ԛ��>��<x��`�Ү�գ�>p�(֔/�B4s�Xo�SM�k*c�XJ��\���?"E7�#]��-a
����_��P�0_p�Z�܄�Z_�C�ά����I�|\�97�n0�0�iD��R8jV��q'�?}Kk�9�Q}m8ٯS�h߭@K����,����
���ֈZ��2�˴Y��;�DҮ�Һ~�����FJs@�;;�Ƒ
b����-L^FnDuϑ���5�(5-�\�h�T�N%�-�ZM�e��N��}���*�* ��l5O����@5ױE�P����m�Lw��B���� �����P�^a,�-�v'K��[ӯ��c	���*a?�=�����d��-/eu9�b}N�[�qX���-Z�[qBQcF�"��,����#���
¢F����r��A��;�]e^�b����x�>��<�/4cT
�5�FV�O�ѴM��b8��T��5�C�ܹ��4!\:��l�J�C�6�"s@P\��&;�ڴ���m�W��D3���*��כ��7��y5�P"%~ў2R��m4�G Ҵq-�d�������4&�a�����ΌF` ZuH�`��
�&���Z��Σ����/N���/4q|����4��z��di@1^^�J�޿��I4�D��*;F͝�z9��
o�0��� [�7z�-f�r�Z���������<&ck�#k)!��f]�7<�ބli�{+O���(>��H�<�ХϜ:�DM��cQ�e������s`H!0�NU�R)�x��,�8�P$��L1'�C��N
��W���l���B���}�x������}�*���o���h*�`���'���w�Y�qF�w�#����xZhM�	.��2y��������e눁rz������w;U8p[/s�f�Z�4l�Ѭ�y	z�0��h��M���Z!u�K�_����<K�^m�4�m;4J�Dc�[v�t~蘘<��J_�V[S�}�}k`T���Ú<Y�����͝�U�A�=霳ќ4��Rx�¼
 4:5����������tag@�^. ����_��x6J@,�M�_�y(P�	�p� �o����E%��pϗ˵\]�P���G�7|��bF�X�n�E�MhT�0�QM=��8��}�c K�r��u�`�e�l�S/�"J��,.���`A�a_�=�|�	�m��+���;��p��@�Hv*0dI���ؠy�	_>W�b/��.e�,@dӺ(�q#�9V��'�Q�㴪&O�g�0��m?�
A:���|{x�`���Ն�A��7oe��`�����BU��������ܩB�qvX[u�E�xBD|�O?i�<"s48rJ��*h�X�2�����Z�(�4���N�A��UG*'tAۥ�`�9��"��<B��������cl��J�{v�Z0Jn!����"��q]OO�tr*�-&�$X�mm[�E��"�]�Mc�+Z�
�c�`KQ~Un��C����^������^�Xv��k��Q��~�
����j7PӔ�+{6��!�̟�a�Y�0��Cu���V��������vqa�	и��R�]�i{����jL��7��7�Vu�C�tp�1��5��XnĆz��8joN�i��(k��]'�b�b���5��SH�xK�NF�i��%4�R$�I��XXT
�]�0t#"A��^�nq��~���3y~�M�ŀYO�mNΊ� Zmˠ�k�s�:3��y��^Kd��x���|������]���乡CB���
b>�h�S���Ϊ1�z6(:����� ���
1�i���Hz�V����/c\�t^y�c�:��C�9s���$!�:\_�1/My�ۼ ��L�K��F3ߋd{��+03X6c�d{��s*M�G4�mKJ�(C�A�SEbx�px��3L�K��H����T�Ъ��Λ�$_G�r��=_ҫ9H.��c��+Buu�\�ˣ�����</�h�	�[!�i\�ڠT�ҳ�{WZtn��Kp�T�� �W�����z���s��������h��Q7DK�Xݤ��i��4�`Q#�Cl]�`�$�����F�}���+��%2*wbZ�FD�J�U�FQ!�.��Č���B����v97m3T�M"+u����h:ysqiѯ�\���ĠXs�r-��>�&�e�{$�c�I
?̫/��ع�.�m���$�d����%�5��ĵ.舢���..��߶N���Y���#��H'�k�R�����УW&Ȏ{>��9 �י 4�V��L��8R�7y��
vN��u��}��@ ��6f!���9����G9?gߕ�Eh�|�&����G�^��ف1l�4k(Q��"��>5���1�nbҰD%�1�>	���z�>{t}�s��XGS�#F� _V��U���Y�^q��I�0@��V�yy��`���vԱzM�H����O�J~�z�j�7鞟��͠5���	e{!������*N�����*�9h�d@(��͸&xE�
9��[똴�)Lث�a�.��7H��|@���Qɦ�]�q����F߽qn,,�~�uh4-�� %SP���HɆ��EK*���4�F�!��H�il��H�q��p俱.Q�Pt�/g:$��)�J|2v+]gFeʟ��A��͂R�Г�Q?/��Wwqu-��=An�HhGqr+#���h��٨�F����t����=�U:���\�"A�J�L��>�8d��`iMq��q��l1D#�����59��\�1 ]� ��J;���s;׏��K�Ś���D�Z��0�H-A��lťrJS�<F����MӒ|��4�M���t��j���x��ZKLe��+m�
��k��G�ӎ1sM��E1�>��A?�
�N�����޺Ր���A�֩S�^o���8�f�ƍ~���+0]����:�6�"IK������#%lM1��߯��v�z�~�HFu�t�-#ٽѴ����� ��j������)4�����5�2#l����r� ��:Gk���F����Z|6���P�Jõ\A��Gys���+���WƵh-�-0����4�.5��@B�k�������0�yB'�.=�����Xm��t� �*f�/�D��͵r�@]��ڌ-% ���Q�S�M���>�8;�8���̒{jh���?F�󮞣�.��D����+S�`�s��"���1z���%�Ls���[���`�X���9�7Z��@,G�2Tţ�Q\Q��w�>�-mTHl	|J�=���R^�1*=� �K(x�z�����Ee#��j������P�*�;���J�û��$����+A���SFr�j���K�Xw*�)�|���J�;0��$�dU�B	�����h5z�s�(G��W��(��Ơ���2��Y��ڏ\'-�����q�6���\�̹y[K��R��^.�;���g�<���(���7(�� ���w
C�@Uf��]��ճL�j���b$5UH�#��+����Z�������₢�kx��5�8R�в[��v`qpP/.W����X:��r|�7=8_�.�h��4}�?j{ �~첣Q6��xU!/��ي�p���=|�vUg����v��#�b��ȗ��E&�g��gHd�grp�\>�ќ�"k]i2�P��T�|M6���j��L�����m�g��v1S�Ss��d�	�.�㕆�7�AX�c�m�\֡���y�sޘ��F�$����F���������e:+ �4��fԖ8�)G}0����:X� �]��������p,�1ܬ�s���BS��g!2���¢ΐ�Y]\8hd�z�F^4��*ϭAzp#77�V���(�kE�Ѩe�$i�$�P��t�H��d�@c��GSr�X�ț�����
Զx��{�b�+&@�����2�m�}�nfOBk��Qv�z ���m[ m��d1_܃�R��FQ58���-������y����wy�Q �S��8o�3ǶRM���h:�ʑk�B�	�ςhЅ�X#�:��3�)�-m�*��i��H���o#�S��x���<C�2Tى��P��#nN�����8�7��*�)u��0Kp5�0z,O�L>��Ơ�E��EZ�˗�b+��@>r����#�qg	a��Ɇ��6y�_�5�w��U�ɰ����.�g�0���ʔ�V�`�N� ����g��M�Aל�û��������n�i��ë�l�6��.mr0��r#�o��a�ލ�\9AR��� �"����H�Zth4A����rQ�m$i�eM�5���!����L �����!�U�U�ԛ��4~�� ����$+���_[G�c�bVþ�>08+��yn𢡋rV������:�S+V!�FE xB�a�_%�us�����:��w,��V���XY������� �n���	6��4�\ˉe�QE^�˺�;���h�~S"�O
�V웸��0��b��J�Ǧ,jK�aAK�5��Y1����=���Vޱ��^LA{���/Ogy�l�ޮ�����`l��д���x�r�7�1T����6��o)�%�ޖ+oB�4��%�綡<H�"~�Yos��`�� "WM�����W��~�=���jͰ\�` Gu���>�H���
 ����>zu��:Y���pZ�\J����Xҝ�}�+I Mw�5�ٚ*F7�U��l����Ҕ���LoCAl�����q�	f�NO����ڿ�����urn�s\��� r�շ�!Z5����;�r>��E>�mH��޾O -9����ڑb�m���m���&�k��=�,>~w��l�_�pV����M�7�������ڒ3��wk`���Z�g5��>2cB�9���tm4FҮ�
κu�Ud�X�m!7sA�ߐ��ٲ3x �B�9 �.�o��@�>#� O��I���8ǁ]Y�m��WZV���<<���?����`7�F.]�6�F�^�%_���g�iB(L�1g&ڬm���c�b�t��J�.W��q����I%��W4@��!v���Xr��� �G�b�sM�?���]9��܈Ao�3xO�x�9^�_y�����[��hћ�:��7T�Z_>��R�PUHI	wS\��MKׁ	~��`���*i#��a����%�D�F�ߩ��p�
<����8(J�[˙P��_=g��������*H��w��7E�I�_P|��{���s�F��Z��7��"��U�`��d̛�h�B�X��D%ֳ�������6���W�R'�� �Ϛ�!@-^�ak]#��|G�$����g��Ũf���b�I�fs�F~��Gy��r����Ӎٟ�!n9��o-]�� �������}I�^)u!����r��xȿa������I'R��<�dռ��9���M�ejՄy�ji7*��}�tOCA΀R
��Fx�raª��^WlՒH������9�Tm�8ӼHD$�b��CT���@X�Ō�<�tZ�^70W�+S;2���@���[�~-����������9��N���X�����=#�H�Ԥb�����Y9�ȁ����1c�MO�����\�^?=>% &F�W;�dCb��A��R	�LNT�WbN!�/�^P\␋Rjki�!�i�� ��s$#��pGg�D3t�P�uu}����M;�'X�����v^��9�H˜Ӽۢ`'�O�#ϥK�E<m������>���z�z����R�M��{�R5����9��cت�k��3��s��Љ��h����JM�g'�?vAU��Rtyy%;Q��>.x�&���p�5'��
P����ݝ��ݳ�?�X1���V�;ޚ�/T	:���"1�� 8���MM�H{:6en{�[y6�m�l�Vĳ�mlV�?V�Om�ϳPE��2D�B�B�����F�E��9Ds���^.TE�������֠��%��fŐ�YSU� ��Ȇ$�|�~�� ���
�7~��A���!_~ 5���z1�>ZѤ�aL�Ң�r/W�%-��������m�^����X�f�f���8*Qs��`iĉdt���]!�1U�Y`�.�ْ@��E6z�I�aۨ`�_� T5]Bt��6�4~�@������	z�a4���M��0�
��Մ�=�E�,����z��dp��`��˫wܨчlI ��] ������I�#Y��Ʒ�#fD�#d�~V�	��dD��L��l��1��f:=�%G5"��
��M��е�d^p�n<lO1X.��NLKl�<YVm\͎�n����\�1��)���t��Lp�P��F���Si��5N��p�]c�`�k0�|�x��PE�2��b3���5�i9��mgDr�ʥ
��|�2������ZJ5pzi"���@�����x��8֟��k�X]�5��CM��_�jT��Ttf{l�QW���G�6멘=wB��é3��UDv �K���Q�Bӽ��Ee�5!(:�,��<�G#����d}�ɳq��C�n���
������m��-v�hts'(A$
��F~���H� ���@Κ:tu
U���=NW؇-~���垺f��I�7r�p�iX��񠶣UB
��¤q�f'z�T�����Ӟ��R2�3y8�{Wl-eE&�e��R7�9�T�E�l��B0ՠ�H{L Q�]���� M'P��`٭���-���ϟؚU�����a�s;����h:l s��e��;�A���|�trm���ڗyT ����k�,%����۲]�T�����Qi/���~o�
�+߬Zo�'�E�܁z�������>S�zu���=��2e*�NP����+�(��+�/ځ�L���~�p�Gm��d������s-9�r՟R���&���/��y�3��Ioh6%��S()M-���1G�ZF)O���S���(��Y�/���.�������!�k9p�`]�R�����2�&>�Yko.MW����@��
7#,w"����}6E�.�!(c���~l��εx�3��,����W0t�2@@{V3ᣕ*[��!�7ԏ�g��h�{�Fb��ld�Vzm���2�&�^�ų�Sԋ��L�(1A9���T.�il1N�����ꚜV/U��7�.h׌&! ���[�/X�Ir�Ƅ��Uo���@�91�C���E�K�F��lܪ<5�՚�-ؼ8��>�%�Dwbm�DӐA��&�Bz���BL!۹J�5Ϯ�]�&t�3ɝ�zF�'�3B�wZX[�q-��LI�q���O;w�F���D�w0���Q�a,<��ᩊ�+�g�e�&t���:mX�߫�Ȓ�ԉs8�X�k��E#C�X_�7�a/�p"�#58m9����ű}-+��3N�8г�O�?r��l����y*�HSY�e�Ja?x�8�@�W?j���5���(�إ9I:9S�9ڟ�K���47v���?�?��Y�����ajK\7M�\nr?O� v�vN@g�UB�u� _���qT6b.����ן~��?}���I[�[9�;���j�U�:a��S$S��sc�z?�ՓG��ZP���<w�V�h,eר��Rh�L[/�9�gr�NJ1@���-�R��vʇi�S'�q]?o���{ޱ9��d�T|��~ �0jJ}�J n����&��Y��$̵�6������xO4�9�G�c��lO�Е����XTɧ�:5>��L	��p��
n�ݾv�����g���5�p�G���k|��%�ڠm�췼u� ��؂�i��on�����Ǜ�9��Y�9VyᾔL�I,f?��b�*��>~���t�!�P����1S���z<ǓQwd�
�: X��l��K��>?�������|���ۛ+�n�@ֱS9n=K��{�6 ���w���7�rq}#W���d�}���(NJm��R�dV��Oq�j�'�����zw{èB˪-$����a�"�
�%�EJ��u�8w[����\��W�'�IXD��ȇ�a�'������Q�M૱{rLv�)W�<���F��Xt;$��|I�2y�Pž�ژ��뮤�fu�B �ܤq����d ��FS���\jԪ��q{_��i,�)�`�mJ�FR�Ʋ��,	kG��,�7߿��o.y��tM�ӟ����4u���C��/�F�Y�������me��\���!��G%ݻd���{�gޜ��O��(:K,X%�&+^hOs����GN�0��7�K�2΍w�ȍj����ʋ.�=�m���E�vr���*7��:�q��q9�q�堌�)��0j�1��G�Q{��:5XR�V�T�8��/�Z�Q"|�I~,Uu�5,20*�<���t���`1��Y[J7z��&�`W�,Og�e���E�"5E��V�2��E*�ot�Ϻ�o� �Y!�Az������VP�ST�]\b�]��u�Ay@�r��F�N{��v��B
����\@�Q޿�N>�𽴫K��?�$	�Pk���=����gM:O/D�0/-R��W�#�&�W��J��ӧ_(`�1�c	ΛvxK.��'yzު�4"��2��b	���#&Xg:=Z�W����kN�l5�N��(���r����@��J����k��Ï�����^��O�>�����K(5e<H��Yv$��+p3�B��$!��G�,��M�\�������%��1��F���Կ=�ndqr�V�����y��=uj�� m�6�Vv�ޙ�3d)�ӷMw��	Ina�����S06�� ���RЩ��!G�����Th��������2�70��^�8�{�x\}�x)�}���Oi2�,�O'y�暲	�yg�F�X�-u`�X��,�8���^�r%��H��3O5�B�e��~�����ɋFTHR үd��? l L +-��=���aZ���{���k�*��ՠ3Adj޵:fܘϪ}�냁y���&���@{ 4�zj�:�����!G� 4q�߾|b 0�|�J`k�^p0N���t��t�ɻ]/t��M�܍4��Dy����soQ#�_D*�S�c�v"�:-" g*���yR����s6��eb�o�w�ㇷ�����M�ᴸ(*ck0�'�������0J��>�y4DLI���+�-�h�˵��?���EnBd���ϻg��������׎�<������(�s�A�UO��֒�S�G������*	���U7j5�غ,���d������j�{EuԬx���|���=���h�i筽|�7O��ڏ�?��X{��|�1��HOTт��d��#�AJ�7�P��^�����R�-�,r���n�a��{�Ӈ�'ꮼ� �V/�f�.���]�^r�r�P�Ҫ*[��.��4�1���wC��;9t�΂O�RZq	!WlY����2��䴽��{�횑�3�A?��{@�?�7λ�N������a]��|����M�.��(x��VpB�6ޥ�uh\A�g�l���������ı��qL�f�隀�r�� qt�Y���Et��_�A/G����[@p���l���ƛ��������?������~8ȧo;	����F��[�t����B�"��2|N�z��Eb��1�<GsOM)����J�ڿ@�~�K�y=�%.1!ˢ�d���B���W,k��E��-�k,ZjG2ax��R��e�x0*�f���[b@,������
EG�V(2�2(��g�	��W�>�d�u���u/;uca�һPD%)�RP��0 i]ֵ�-�>�D¾=��'OkP�mV��بXy��K�Ӑ�D*�r��Dd(��l5Q "m��L�l!���=� �<!tD2���GQ���ӱg�<��=w����0��ń�l��G���F����FC��T�����Y��"H~�v�V5�kj؎�  螽�"�L
��|�VQ�B��T9A�Lf]֋��/A�gD���3��^���\�T����0��zލg����1���Y������8O���N�A��k�X�uŜhsD������|��V��g~�۷oY)Ɣ�B�����; $��֖D���Y��6d�O�!�dh��ۦ��gJ���Y�
o�S�=e�4.;��+z�]���%����QRq%=W�f�Ϸ&�m"I�t���wt����݊�W�#�V���4Ku�������c���ﭥ�����L�Y�vҹ�z��U���{�29�߯yZRA�2�Ϊ��G���=ɕ�Y��-�4�:=�����Mr���1B��gk�'��ׯr�l���m��N����u#�(��r
�8�27&����@�&�IQ��l<�鼠=�9>��BqPl̃n�h^�e�'p:�2�Ni�]�t�noߥu��ܾ� ��[�!]��=�����U6e��8P4� �F���o�Ez`��=�|�Q%V=��wu���F�GW7o��xC�&�<4�ܡ���J=��dEB^@ƿ��������+�����(��޼����!�	Zu��\�����\���3;w��q��\�DMZ� �}�]�K���=�k���t-�O�=&�?tTEhL�Qy�l��ӂDj"�X$��RU0�urLl�V���j�5���v2����*�����{��̞�?����a���k$��0��|�l�]([5W�yK7/#Z;k�7',v�*�rGV�L�rwn���-D����g���V���k���}�����C��V��&F���lFŰ��O�sQ�t8�l׫H���!|�.�[%P�I�g�	��4pSeR�h���X4�h������^�w�D\$��fI����1�<��4�� l/�۞^�`$Ox�+F���OF�ƭ��g��ӭ8Z 
J�3�ξ`H�.T@��G��DMI���p.�-EƘ��ݤ%����|�����$ct!����2�~(6C�
B� `C�2�s��� �^��h��	�������{Vݘ���<M��:	��-U���4�$�"�}�ء_ &��`�>=>�С)7Z��x���GN���vu]e�|��=B䢄=��Ɉ�*���iIƮs�W ))��ϩGO�1Z
Q��ܻJ�V¦&<��"/�^��a�UQO�*���8c�q ��T�c�&��HKN���StM��R�ܯE��q��9���
�s.^S� *pWn�|�`��P����}a�Y/F��42=Z��ܓZ��'sqq�L����J�_��>$�����o����p��>����ow����I���_ɛ��&�P+���T���$��^���"�{�ȉEJhἽ³�~���>fпB�u:��ye�_A���t����ț$ Լ~�%@q-�>�	"�Y�KM�v$G�5�
���𜓨�\����(����KF��1i�v�R,<^Dp�i�ά�$�=���=��u�����/�w��֨{˂���x"� .�M�H!�f��[�t�ו9��c�@DN���Y�[����dK �b(�/����=�j�qng�e!���bnu��9�x�E�!d1o�\����RPli�ת���M5C2�@Cj$Q�t�猽�m\�$_=��[%��4�pi�4}p���F�B�{�����d�]��P��wRi��n����FYW:j�����_��U������j�#I���#"y��*i��}����=ޏ��{�۝[6��YuP�$�,�������z�;@�'�j�����]����˹��Ҍ�]����_M9D�ީH���!׶R]0ͨ�yc��/vpŗX��%D��{�A��ddw
�~����_tS�3�a{���'�<�GO���O�ڇ����_��^�l�S����x��)�����t��%(�6F��vM�����{i��ֳS	<���a�k 0�]wKs��Y�^Kƈ��-MU7�.���~������g�]_������do��8,�������|���-�r��Qp�u{�
������^�ަ�Lc��e��MN�`x$��e#����X��������������v�ׯ_�S������������\��<ij��><\��(�Y
��`��9�X!/�yd_r�Ⱪ6��-7���F�1X�~�NewHX���t�����̹��C�0��� �Q;�S}�(ua,VSn��z���3��*�	P�3i��ޗ`�}����S��w}���[mX�k0�ת��0�|��]��'g{7��������9M�2�/�m2p�����������ﾷ�O�jNb��)���p�y�����g�K���/��ǋ�'��8	$I���2y��6� ��'�}@%K=w7zhB�P,�!�^�ܖSBFg�|B+ʶ�b��bq@������d	�������3�yy�S'"�l#�6��{r�k�)G�sZ����1��p���r�^�}o�>~�ɓُ�?psG6�#��%�@󸣏┢���qa>UJ�7��ѕ9���c<4����$35ʄK����D��AZA����3�<�>��iCI����Q�N2a���ɟ�Xz�$����wr���܁��1#���6�،�������f;�H����d�k� ��0N��Ԟ��Y���&�t�dr��@k����)<3��ȅ�����O�.+�,�)�QJs�����y��"��	�s�����ݷ��D�h���z��~V��;vr�}�q��geYe�T��!�+�����F�`
��y��y�Ú�����;l�a����n��lM�ɱ�U6s	���8����_��g���o���%����;z��0��g�aӺ�jb�vJ���#��EI�T���%�U����خ�LC'g���J�v=��2���;��3���.8Ͷ��Ʃy>����n��ի�ږB��#�W�)�)��xH���L�1o�-��yl�A_Y�1ו�t�sg�_u �߬dr�3��C�_���ާ�3�=����)�`����G��Eb����B�>�w�ƺ�5q��00N9�O�S9�0�M>�Ds�	�W
t��� ^���A[0�0;��^0�?/�L9(���(�3:�[)po.�0�oBm��(��H���p�R��'�c�2do �� e}i������
pz=Y��~��^��Iu��:�����}���	��x�~�e��!�m=/�Iq���h,�B����׿����9�r_�|��ڻ�.�1a0=�h�:�A!��NS:!�Bk;��w�䌮��GM1=�}G��hm�����Ѓ霡D�̬�1�qv�A��$��=
A�l ���Y�~������ߺ'���
C�KXBj����8(s�f�D?�n���^��]�V�=�۾�u�������6��U$�� �zR�'�_N�<�eg��a46�:���|��b
��n����0�/t����ku�p���'�@XD�$0��=Xj=2~���Z@���b�D��ƅ��?_6>#Θ��T�(^�!G���ݬ����6�*pLxi�>�l��iW�_�
��Y���;��C�=$�Ѿ1Z�x����Z	�@+n�߂$�9Щ?4�]����Jaz��u���%?ǚr�[�Us�ʻI��}YR�u��d�}>,�pZP3���h��Q������e�{�n]�r(�0سC{�pi��00S[����dN�]�jC��Q�s��F��	��\�w~��$��&��]@i� $Y{�&��\��S�k���P���P=m= /�! +=8��-��s��o~S2�G�kdɎ@`Ki  C�{��h��>i���4-h�q���v��b�5���:���5��1�排̫Õ�|�ڞ<z`_=yĵ�Q] ��X f���wO�Hn\��(���X3�을�,�,�� �6���FX�a�� �� \�Q��WF�itPF	���\c(=�0����VEw3vV<Om|P�0iL�'�v|��Kz����6�1u����{\����(�߳^��kߥ�:j< X_�����Žş ¡�������8���ƺ�a�fm�n�����;j�޾}O@���/�<���ݷ��P��b�~o��
�����
����� x �X�(5sr����RH^+�m�莝�j��|Y\�X�J���;�k:/y=�k]���b��Wp���xkݬ7�;�M1$Q�-�y1��$dfb��kX�hvA������:��=��\aS�� ��ܫ�c?�L�j���X��y�;�M�h=b0g�3�%�����)�MW�Ƶf=�DlFv�W���2X�1�r���z 	NEzk���8��Mr���I��U%!5{6�F,�$���^�K��҈E��&���u�t�LV@\�͝��ZR��H�o�k��_�m`D�ȿs�A.:�Yـ�g"�5d��T��_��L�����l����?'��5��Cj%����$�t�js��"�z���y�u�@/9��O]���߆���!A~k�W�c��c�8{���LOc��_�(�$_hꀐ�ODԸ�l�P����&'�i{��z��!��N�&~l	]�����ͼzA9(`f�Ȫ4E1�y\S,j�nbRh.��+l@*�{5��3�i��a|���� ��4-5�3��e���~R����|��m��d�00������۬u�(��Z�0��	����-��[R�y����4H#��׃k C؁\|����?���S/��vc�>}�wo�ڧ�n]\kMS��eT�8:�3x�i0/�+X,��R�����	�+��C�M���A�'����gk�vl�s��-u�\m���s�+(���g�Hw*�T��0y؈�TL�Xz�@_b�Kqq�������u�?�����e�Z��:*��Y�^<���e>ۻ昙Mx� `�����j���Ĺ�9fƚ��u�6���>�'4�p����cZ%@��rt�,���r��~ �K0�`���1��ks�Nq�����7_��|�7�5�m;�
iv6�RӾE��5S>x�TL�N�3u�f#��]�akD����`ٷF��X�K�w���K��,.�d��c�( ج���0]1��b�v;M�[�������P7W%>"�z;`�l�,`�}Ge;�F���N�e-�1iD=z�I�<�:���V��c�z�([t��5����_)~��gy�V:F��@��.�$�E�7�{��T_[���ds�C�V���0}l"��l�����#'��h![�+�u�C�� _��,=�ONh`�#��^t�N� YS%@nJ`E;��[��P�����j�D��˿h�jo�������3=2��R;�����\\�$ve�)2Q�'��<m�}�_8���h!$��x�b��dJ����v� C��PceHg���48z��xJBi�V��98���fX(1���7�	�� �m M�������y�|��I c������؂�2	x)���?PM���H=��f1��|͚9�1���`Z�q�ܦ�@>������{��y�M2W�\ @�ũ�C��� G�Cf���,���c���H���p��X��6�=s�b�����%�E9��ť��/�y�����~|������{:L_~�l�WW�L��D��@�.6kw��}� ��muw�.����Cv����5�6�����9C��1��w,X�n������%�ʧz�ܞshѠa�'K�a�"���~+�g����*��>�k�_�-B�1�׹��zWo�zW���`�/�E�a?������">Ã-��ЀU[�Γ�~ne�����	������X�(BH�N�M_�8��.G���g�M%��3
F�Tem����h/��
ރ0���*��׶�N�K��af���Q�D�w)�G����If��}�='�����:��{�������w͢�1"�LA�*��(��~!�l]�)P%�+��zr�2ͭR2t�eٴr�$����9���$�x�� Zi'�N�@�5[��l��ܐ�����k<�$�'w��`~�`�b������1��VC��;����~�`�A����pe	ڵw(��Y��Mh���e������4�������J�X+GV@>Ismn.�kr{6ɗ�������1ݖ�ٰIj��E��"����`�����6���ث�B��:x���9`�ۊ}2:&L45�5�r��ۻ���� ]Ʃ�\�#�A��,�5	��B�;�/lpe�!(I�e����ݧI_
��/le�.��8B�W�P�x�Tg�MC.�C5�k��B9�h��I�t����ue���j�z&W����z;3@��Wb9trه7���y���林d�H��-�ōKcmL�ZI5�WЛD��0�t�����\�%DI�5��Rd����f�������<��M���-O����. �J���R1" V�MZs����$���5����&vp�g' ۀR6�-���Ĩ��eK���?_�6�ʛuO�f�5~��g�9������s���;m"c�����8��>U6��-����	+Iз4�� 
|t���� s���#��c3������g��E5�0��������C�/�������Iq����,7F�"�κ�o5�'t�8�s �^���ˈ_�(�u�gc�:�����7L`��Z&tp�y����7����9�n�Hvr��q����se���,p~��(G�����}��8r���gvj��͚q�j�F�:�)�DZ�`})F,}]��>UV$�cܿ�j��a�3t~�u:��\�k1�c��{�Ϫqf<_!5��Q�5�]��I���e (����rl�]���D���J ̽�uĵ�q���qH׷k2�)ع�%Gw�?�Hؼ��	��꽜�f�$ :S0�mz�d g�YW�l�`uCJ���^D&l�.�g�������.���"~,��
�����5!i�;	�NHʾd��.W.5K�9�
�:\4Hь��5>�{�n/1%CH��>�hHA��%�JRD[�&\`���Ŏ�!���F�0އ�5h��2�_po��R�+�p�ɱ�����-�m�<1�"vZ���K��*}�UBW�A�-u�o���e��M��h�h	Ye�V����,T�eq-����'�l-��kK��d�Fc�}5[0^s���"��[ci�91(a�����Ζ�I��x�jb����,�(��`\���ye�:��|e��"��4[�C�9�L�'�56�-�6C+�Y�{9"�um�D�KS+`~O+�BO�9>��b�AY!���%ڼ���o��Ǚ�Ĉ��!1	����`����F�Ġd�p-��]c5-2�
9�5��LF�{�(|����/(�ų /0��W|�����D� �;��9�BW��P������b�^D�Bp�q�
��bl >�3�w1\x��Sh���C���1�Nh�7�Pd�Q�k lY}�L�On�\�k�"۶Ժ�|�c��[���G��g�* 4��V�n�T� ,@�ތK��:%%���a�9��z@�e�(�Ǘ �h��7P�n��it36ͻz��:��p�./y�q��]i�|2���A�r��ݾ���j��@�F�	 h�'�1g9)8XҖƼ���Gy�38d:� a��Fȃ�s�9�K�=:��L�e���|�rH�vV����DM+Y�)�_j6�,��v�U� Ɍ���%|(��Z���F��N���Da��ٍ[��꾑hk�g�Y�[;Xj�wv�c��ǬR��}�Z�M0�3�&XP���V�+)5ۚ�4�斄�>�����]��n�&#�p"����*�*Cb1��3ѭ��)�g�ޔ=���O�Q�1O�l*�,	ħ���\�
�*1�%t��Qj(�^	
R�Gg����W�:ל�^���6NH�p�H�ט���P�S-8���擕�IPn��H	��?'�f `3��m�<|�) �ڶe�d �4����	���*.��͵�;r���ϥhE;����L�9��.6��Pi ��]	l�J�	�����?�����ձ� 6[[i���5��ŗ��93��y�����v�N����c��*����_	�s�����44 ��������i�䁅 ,�,��{8��5������o�D��U������8	N�Nfn���o0����Ǯ*��3|K5p�1��sd�D��z�֊�C�s-��fόor�Gh@j?���^�O����kתe���k�8h���جq�� L3��	o1�M�A�9�X�SƎMj�'�7�3U44'�|�f���Z���k\�݄�����	��в�C�K�2\V�v�@9����o5��`�]����	�vB�d�r /)u,Y/l�˒{�|;�\��3����6���h�li�g��}�c�%������%Z��P��ȝ	&���%�Qe,]��Q����/�nY�����u	�G?@�	�3|X�E� ���>;Z'J��FwÎ���Eh�L�lt���M��Hk ���"���L~mV��z,�H��|V;������`�U��<>���h�q�M�kEA@�%�E��N�F7K�r��-�ö���fG�E��ۍJ��L�_Gk��%G��u��(���'Z��K���!�ax�Y3M%f��c:�&��3Ԙ��D��)#�n��5'�u.
�Ş�碛��]��K��^ڲ\����'�&���(���d��uI��/��%i]�*G�u]��̥p�O�:�Gh��څ�ä-=��z�V���,��Iq���v4pP��E���:|�˛����x'���,���]\�K&T�U9�4($��4y7JKƉ$�H,8�1��z���'�P����Al��g
$Vs,�*�LUx�	��Jv`�pFu���f��ϬRc���r�0�P���T�g����+6*��0Sc���(}�üg~�D�!�� ���&)|rR\M�~G� �s�P��ʜf�Z�>2)���C���i��0]׈�~�\�l_)�u�9F��?���:�G6,e�O0��k,����v@+c���wY��'Ҽ-G_C� ��e�{��ǠuS7d�(�;�A���:�v�yoP�AZ@m��|������N� !:�h��،���;ַv��.� 4x�dJV�J?z��I{�{�ڥЍ��� ��,@u�i��|��3�֕�9�#�)Yƚ����gu��r�{�*N8�*d�g��b�f[�*�X��Z���٬�r�����u虰^���/?zQ��͓Ð������ �H���� ��]�����7�!RTފη�v�+��+�j���"��O��p�X�9�xkC`�O���*%ˬ1�Ȼ9G����fo��R@�]O��A��X7s&�ى���g�Z��D�xr��Xe���&I��Y�� ��j'#k%1s�6��3u������C��n%VT�Ȼ��*�^a�����
�J��I�>��d�*i�L�@��	!�����i�,�=߬뙃Asm��)�!����ea���+�MG);r���q���AW]��֏/���Rf������
p�#i�@��n���'�����׿zF�����g;;�������m}���آ� �4����,|*�?sa$�e� ;��#��
`� ����\%-w`��l7Ǩ��-���6�_ӺH����^�T�X*l��<��G&1��=OB�ѲǱZt��Le�=���]l��a��7l��V]��՛I����00�Hրf��� D�i�Q���1�Ȯb��sJΠ��#��6㖽�b,U\�1>h�c������u ���ۏ�>��� <�IR����D^���Iʘ�uwF����wK���� k���}��hd���}���oDm�_%�v��1�N���C<G����6$���+3�6|a0�&��␁f
�jV�U����>f�Ӕ�JN2)luv����^�^�ڮh$��5�9�����^��}Ԑ6�V�{!S�\;������8��*��V%�h� ,�[? �>#q�9w����0{�$/�� ��N��Կ~ӤY�� DQ�[���w?� �2q])�n��޿�;�_�u��d�ɲ����=`�8��9�}�]cSIƼ\��+���f&���֤g�Chqs}�kL�{���
 ����C�9�Nz�4缩���i�3�q`p�"Cz�Mvv�|/K�Cp'�S�4��E�/UY�|%N�#��i�A��e�rRv�D��Ϩ�(�L��W݃؃R��E�*��D.�i�Y��c�X����X��s� Ru{�4b�,�R\��&/�n�)�9%k�#��^v��&<��ѯFA��d��Y�(M������#j��>���F�^���z� v��E��	4���|[�S �l��W���q�2�==2�x\�Lv0�(�RB�S�<�ً���aY}.�����=1�ǭ;���	F���8ט��ǎ���q���NM���j	cڔ�m	��a0���u9�f�A���,)@��C-�چ�u��N�U8[�䋖]ҫ�O�{(`ͽ��{��]7s�̃	S����19�0�OL����5�|�@�c�<� �4��'�'"�{jY!bsL��d27;)�Ҩ ���D�-����./�l}�,�S�R�~�Ď�'ў�i�@6WXF̱������w�b�1�F����OK��^�#�;����mՖ��p�SA�9s�n����A���FL��Nz�p�n>�Ti�Ę,����r-�ٟ��|p0������pa�A�x@�%�j� ,{d��:V#��*���Ս��l"7���u�p|�YS�/u?�Ο=�TF��Iwi���Gz�-���=�<7�+JH�D8S�<u��龂�
���`� t{&�/�M1O�����Cr�D�z�a��y�Q�'I]a�hQ�\�!�W}L{��]�F���8�8��8
��� ��
k�k:��;��x�i��5 W4H���p�ξ�Y6��J�����|s=�������(��{sǍ.��������,��70��-68����^I{K��_04j����b��i'��Z�t�sg�i뺡K:{�Puib���BHnx�,U���B#�;�5�·�T�v�&����8��~09e4;g�m�S���9*7�����"-U~EL�΂��5����vsk�|�|ލ�}�qQ��Z��/1���������)u���!�l0�[<��.��0օ���5��y0�Z�C�ެn��[���FM�[4�����}��h�󜷒-@2Un��KQ��Lҝ?c�|�uP^�ĄJ�x}\�� }7M�-{C��3u볮aE"Vc��#̱y}�X�Jl=�M��Ҧ�����|Lt@k!a���nT	�L�jQNrY��jgG�7H�U���;��'��.;�1:���1���*��1��乢g�`5S�ί%\T�|Q����e��կ�Z����r#ǘd�� K�J-����8>iZ� 3���U_-bi���(QV���]�U�4�C��'������,�3�ɍ �ּ�лy����Z��'A:�Ǭ��בg�Ņ��/FĥUg� �^�ӳf����g�j�� ��y��H�_-������K	w����z���Ah��jf��iǵ��M1��K�7�6ЍZ��M�,�(!�~�����,@�>+��u�Ԗ�+鋦ru�Ƅ��QL�֫�X�!�IF����<�v�DcH/C��1f��>Vj��/	N��z��v�b 3"5���57V�9��Sn��i<?�ݝյ���g_/:�hhB+���z+@۷��G��u�����j��B��>a������ķ�x��#�-�XS�nuV�.�B�2d{��������z#�����+K�O��*��(�ZZ�ʴD���ӨF,�ˌ�|k�_�I^M*�X��� @�$��
�%�ɘ���D��$P/^������|�^�Fn6�)����-���Ɲ�뵽}��~z�3G+��l���0�y�4}Vb�����E��--tmݶd;����.Cl��qǨ�x�(�0�{\� $9�B�N��[�ܮw�>�˗��ݻOv|t*��YRi)͟�F�5�}�<AX��/'�eK�O0��3O��ʆz�X�p�XW�w�X��q��N
0��L��A�� _%N��qr���c���};^�g2��s94p`��7OZ�޺���E|�����'�~��!t�k|�� �J��cK�H�g�����d�Z������	�b���V�f�����3R��Y�	�Y���Q��}��,��qhv�Xe��
��#�m��e9�E	FK�G��I�Qю�-���58՜��h���"<��sٔ��3��Ƭ�Ţ�s�RI���t�NQ溗�m�І�"�r���9�����:��7$��A��4ל�@�E�7UR�)ܘ=����w�~f:(� ����L�������O�+�w˴+�o�>է���!*��A���Yft��U�T�x@�6ٝĞKY���k�r���L���͂!4�Y�u�P�'�xm��-Ӝ�ĶY�"_G����I�5���
b�J���l�������b��{4�+�L� .Ӊ��;M�%�:̕���H����g�����Q�Z�Q��>T�Z5�4-[�Gc����9q�ee6��&m�@�$����o�[�ǂn��8w*/Ž��m)m0�)L����ח)|���_�;�a�>l���+/����lOD�fܩj�f�]c����(��g��6,�N�vW���z���$�˥�v�����Q�7�qh�G��J4�ɶ��\u��d��>�6U$[��Y}�H�$�"4j��HdVԴ�8gYҋY{�b�:�u�������v��`���I��Fn�p���;��F̗��7|���<�������������ޞ�x�=,�C�4�ź�*�*�رs�$ށqt-���Pcy�J��U��!��ӡ������ì��a�	��k����͐оy��$H/�'/�5>�G��с���Н��7tw�����}c� y�A,�q��w����[��l`��M��o?�y�ݹ��@}�C�4:�oY�6Щ!����pa��s��/�睳S:0YXh}?�������=}�Ȯ.5����HR�v�C�S����G��:`����p����*k�G�4 �����W%��Ja��40�{x�!f��˱��v�%f:ے!�^m9H٭��Y� E���E.,� �"�D��b��U��Ȭ��,[��j�y��H-ӫk�KJ�=8+2�;q�쎴�X�h�rS
 |�\4��Z�-���{�zgg��8E-�	&Nw�����.�nx0F��Y*b۱w���V�|�l�P0�����.>_Ӹ��#��~�Ka����Ŧ���c�\��@/�����į�y^�����`��k�z9�\�?����Å}(�7O�S{�l���n!�Zj%a�b��ޜ����ϸ���������\'�� �H.8{-�����f�u���s!�'׬h��',�ϛ�+셏�i�����qv�FǨ85X�y���R5T�*2�`'�T8�����]���F�dXVD�������RK5��8�؀Ȫ��I�85�����Ed��?�u���X�Z.�"{�X���(3������{��0�^܃`�u��˺��l/���j+���/5c1KO�������n��P�� ����~;��sZ��S���驗�[����\�iX�N^OQ�����믆�&L����ϵ�+�f�*&K,<����^(���=|������v~z���8�;iO��Dop[��qM9�ʆ���>�?��G��%N��g"X��5���{�%�9lV���f1�E9��[RG]C-�@v{/���&��N�-=��QnvQ|h���&�|��Xts�����R���{��
���&�;)��-��P��������ŕ]��+ObA����\l�?�:ⶲY�z�C�Yj���׶(�xt�I)''�vZ>�O�y���z�Ў�]��!"f'�<{���=;�6�g�G��q2���m�Z��>K�%����z1Лl���+����	�#�gw�P����K�]������u&g�'���8������L�.�k�%:UV/m�X�Г������+@k������ƥؙLd���m��M���$��p�[u�]f��M��g�w�ޓ&����6n��ېC)缥X�,��p�	à�/+"ܧ��,!�����<��Ƒ�`���f�7MTd�/r~�,?��5݃V��(�ùH����w����xqE �<�m@b�А0W����5��f_@^��Cs_�_���9ڞ�y'�2�h�`�ܔ�A�F\hn�1���~��;9>�o�>*��N�hKV�cZp<�H����F��-]71�ލ�`7��(~z����_�`�����ׂ�?�GY\���M*`Oc�<\����@�n^��>;=)��,�`V$Ə0L�K%q�\�Ur��� 1r41���Jys�� MI ����,Ldrf8�h\Ph�²�]�ay��!���/���ݡgr˱Laa���gyߙ<����M�V '�^!�R=7tbz�P��{�\�^g@��� 'f[����iøt�M{��Vjl3.�G,@^���,��`�[>ԃ������r̕{�9�g�-)O��??z/$�Q~�SxX6���Sc���0V���7���g��&�_3{73KG�\���Ț�l�`(���v�����*���!��ȳ�����o�h�%����?���Wvz��.&$�'4�F��k�]���~��?ٛ�mM�b���K� 0_�E! ��O*�t�x&s�C�zO?���h�j�&��ʷ��Ǹx��R���*����@�s}����?�M9_L�~��G(ו��Œ�h����h�A����7e�z��k���W���;�9`� ��9�ڰ<�v߱~�`�u�`��36���f�����f#�J����޹=~tϾz�� y����$	'�%\���mZ�)p�-v�|�y��QW���J�\��u,f�QW��i��1�dx_Tp�xߒ��{6��

�"�$7�G�B1U`"Z{s� �{�p8��i`�N�c��h����U�U���M7w�d�4:@�8�� ��#۬�����@�	gf��/>}�oJ�V���Ks��G�1V�������T̆�k3�kPsޮKvVP�jc�|̍zX,k���ॶ�A����a�g#+S�7o?ؽӃ�yD���]�l�_�z�5�����O/^����s�&��T��b�|�5����g���'�{�4�ׁ-�}��ʏi<Dg�k���KGL�. 4'c����)��6`f��{�x�_������6"Բp�x杨��$�L���j��?p,X08�O6Z��L���*��֬�2Q_���Zo�\��8><�{w��Ǐ˟w���}sj�/>�IڊM������T��o��� ����D�N����3tM�VQ$}��g�C���F���w��hǬ����(Ճ���sfYk��h"90cD)�i��������F%�"�|�y�Rkc����� T��E0 e�ͦi������������_���w`h/ӛݮ��U%>>�)f�U��Do��S�P�1��yt` f�`��ݻ�F ���<��� Ø�;w�ګ����\6h�����'J��w�뜂9�sM;�I��q��U�e�b��cv�q��+�|Y����k��ay�f�KL=Xy��ksk}�!j��e9����ۏ?�(	ۥ���l5&S��� �gS�o0È!�9���i˪U�?�dު�H]!�6_w�gj��8��Ki��)�a���v+MQ��N���ve���޿�`|��̶$6��������Q�]�` �+�c|���v��.�e�������/�^���5�4@+U��Ϫ/vf/�2�[IC����v�J��~V��ûg����=}|ߞ ���y��W�JZ��8����_�WȪ�h8�u��s8�/f�����=�Ƃ�c�漹n�(lZ�]����(�au��%���;�ʾ0S
�1�<��Y�܉^ j��C�{�=��7偼k��r�7��#�׼9��N�m��:G
�k�w@R.�AɮV�$�P:�'���F�z��^^�*����ˏ�wo�3�Hߤ�l3tPl�lPli�����\Y�<�M����v���m��\��%��3��7�O�P}X_���\ ±T���k�~B�BLZ��g�uc�H�/tS������_������s��BeC+e�~h궩E�ݗ���������Å�Q7�s�ͅn9�B{�r!2�jj�%���L�݆,؄Y���_���9;���n�M�YAw�3Ձ�f�Ο�/����_���� �/8��Ʃ�Ns���@���J°ٹ�[Z�6+.LD"@��0nȚ��s�}�Ⱦ���ꗿ(��]���Օ�~u�ø?~xO�|8��7��&����=#���!�B
m�~gNP�����2=(����=ﻳC���~QdV�q[�J�w�Q.�"��f[Q��o3�SJζA�T6ϡl�rݰ4g�������e�m�s�V N�(/(���K����Z�j=��۰����\ ��������6�Y`�R�J������1�w0����%	���|�UWj%o��s ����W��W_�ӯ�" #�P6������?���~��~��?��&}}�U��A�W���1f�1nJn"��VeW��!�QV�^ ��e��%�5 0���������o����w�jg'��Y�Q6����cn��w�)	A|���-���r��l�ϨȀͅ�h%崐^��`��hk�1�|����F��"o�e�/a��u�O��r��q�E��> �u9@VVI_�ò�"��O?ڛׯJrxf�>{j�����=��<W�ѝ]�w7��P����&�o�^��*�p�r0��&=s�#'��3�%��ΜK�w����־{�ؾ����_>�o�~b���uH_8zP�z��#��Js}*K��U�wQb�:k2��o�k�I��O�<�pе�6m�Շ�<s�zagdy��N���P���et��#j��m]xq����l�Q�q���g�QyѭJx!5 �,�A��Bs'c	������3����d�*	\U����"y����ٽ�MC��ӹ��p����T!)���$��3p��>4%�
 ��<�[teb�n�2��f�+^�N�{�(��f�ǿ�lH�@�o���@���.������xV+Q��,�g{����/��Q�����7٭'�L�fɏя%�zj&� ��<�`Q���hʴ�i�XLw�`��6!T�z�U�,��ӣIUs5:��|�tU ����w������帞���|��`.��]�.Y�?��d���2&M����UL�C#�@��g��1�zd�1TF���㒡��_=�_~��}�������ٝ�3�!����8/�����s�6刽�4��u�9O��+�*��Kd�����()�U�S ���g������v>�%���^)5����b��_�Ko�6ekN���Ɇ�q.*8
͍����g��z0�'�����`���Y���/�w �b8u�T�zV���R{ƭ�d�k��;�fF , �.�/ٴ� �a�2O{��S� (1�_}�Gw��ɩF�8 ;;;#�p�<\w��+�>c
�zs��͟>���,9]ˈz�ƫ��2E+Rh�tg��J��2֜��:��x����������ȱd���ڭ�UC��h3I��9;u%�=-�e�mQR����sv�����h�\�a�3,,C�F���(���j�$��r9�s��Ȏ�W�;O�P�������1�$$�H.p~,�Sr1I+˒�@���%���>r���ܿﹳ��(�Ӻh�����g{�ᓽ}���h�b��7��经W�b�T?yR�_f������~��~�Α�⻯KL��~��3���=;-��p5к�H����S
��a��m�M��Ε�>B�8&�s}~�̵��������N(��Hw�f��b�y�к{�A�;�;>=����=�r�7��ӻe�O7ܙB|0`���Z�ҍ�B�6�4���ЄԸ	� r\�up"-I��l�a�����!��.(ՙ�M�n
yv��.�J^Ki�y]�`8����-7h��-���s[~ �*Sy�w��5ʑ�Rr���Xo�9�������:��=6r��~����o��y{V�=���,�[����I��?9��S�d"������C�x�oA�{�cv��8�юu�a�� ��� Dw>�ppެ5��"S�����<�?�����-8S�z�3�p�ET���f�v��������$�t���f�2����Ah�daq]���?���_��,���k�ba������B[��)ཏ�=e����34��j�ѕ�i��������_��-�%D��,�,pq�1��q^��XKG�kS��΃i1~�d2W������ *ƄѼ�ڻ4�[-Ta���;	 ��a�S��*�ZT9�	����:�b�9|a����	�a�H��) �X���W0��e�/AX���_j���zQ�F0q����B����F������(����{��~�\}�it�N~�b�3ׇOI���M�t� �ǲ�B��|�޻C�����F݆��`�3��NlyxZ�e�^�5c�.���A¨�A��Q'�t��$���|�u��$�C݋ۛɇs�������FV�E*=��:h�1�d�%�b�����g��� �6w�.��n]˧�K�8.��senl�-�?�]��j� ,*�=�d5�qaE���;�4ƈ9���C@?����1~<��+�s�,}a"������+�65���h~��]>�x�#Qz�G��F�˄D���D-ȝMYO(e��[�����L K�4�X0D�ox�z�e5��8
��m9�۫�����Gw�W?<����������OJ�L�/��@���>_]��@yG���L�<ԐT�Z��vQ�
�%�̥?����'{m��`l�12-�&Ь%�옝�Y�*I�ݻX�g%�9��_��ztr�|�̼������A�Qg�2��7��R��ѧQ́͝O�<\f�|�"YP�~Ȗc
�-��_�stj��MuV6�v��3;??%낓ƃ�uo ��4�}]���˂ܯ��"���q]��<=w��`�VV�.m&`W��-�_y����&S�jI�~���ᘈ�?_������^��f�Cr ����f�ׂ���»�����d$��,�	�{��k�,�]'L��#k�z���v�[����
��ŒR���?��hpɃ��H���95�"~q�Ep�Q��ߗ����g{����~� 0,wt�>��$(@F�����-[����d/_��x|h=��Z�]�h��\)X�^{�Rl�{`+�B[�H;;9=�Ǐ���o�|Ax�,k��`C��c�.��Ff����\��Y����D
):�\wt��g&Ӻ��)��w{v�~?ӗ�Q���Y���ʱRplP���X�a�FM�=w����M��Su��=���[�c�Y�F#ta��Ρ��{� Gc���.��^��b����{�E��݀\ �a��Z}&���_�|}��~f�J�N��D�����åc���Q
p>��+Zע15��v�5�}�x�����w��8���?.�	�b.pt:v��$���rtWzy����˻�Y�ڒ��$i��B/-��!�4uv���*��Q� ����;��Ai\$*�\�5����%���'�U۔����k��v2�ɷ�Sa��8rvz$�����]~�`�^�,��=c����;c��!�]3<!7��I�:&��ׅ.�n�����K^'�y  �b�g5_H��3���9iXy�#���v������6��<ٸ.�Ji���_�*m�^9�_<{l��g��o���w{a�q��[i��LA�p}}Ko8Ȟ�ɏ7��-a�ґ����MY��ǻ���٨�]�`����-~���l-��9^q2��#��rAn��c�긜52����N�}��J�w�?���Ѧ����0.Ey�݂@�Sv������%�������T�0HG����0/=���b}�13Y9����G�-��׏�}�0Pc�)�\p#��/ ����c�,��������7,���AN�/�<�2S��9�m�%���<D���d��'�f(ޗG�Cwl{6ww6�ت�7	h�%��\��������ŧ��uӕ�p[[f��1�\.<0`9�O��0�9�-�ځd��$f�2 �݇J�(ʎ��onJQ>׷�<1Keju�OuT�9���ߍ��(y�j�n���ð�:����	<l�{�>����/l�ӫ�\K���x��p�-�Z��v�]2���h���r]�@]�tsW�n$�O�<3�\?��s�e>�*��^Y��>Њِ�����?��޾yC!����J2p��Ya�12��G��� {���q��4�Gf�2;��ѝ��(}�f#:͒w��z�Ɣ�6WZ��f��
����0mS���yyǧ���c����-7�'BxŃ�Cn(�50�j��&����g׉�85���#��Uư���h�ճd=�J�������kӗ#S}���k��unF����d���@�d�և�7}=��kʤ|��P��{���z|����#�\]]��x]��{݋�#{Tb/b%���p��^`Tޖ���k������KlC�ɸ����;\�a��:Z7���m�ph�=���-�@F�%c]��Q	��%�ML�9��[g�ǺN���U%_2�#Fӵ|�F4裶dZ6���1�⣗TC���Ý��%���d���~�����<7G���P�T���܏7/��5P����UO�<��ŉ��}���&�������&v���H>Ky(ק /�1-�X"������/%o k;�;�����٣�N�kl�Y���8+�;	|��Kr��\��;?[�_?���w?د~��N��$'���Q5B2�X�R'T jN���&e�1�2��A�Ɖ�F�*��ܳ�r�V�'1�T��;C
۬y��,h�䤃X�L����$����r���E�- � } ��yQ����r�X��;��@e2xid1r:z��ql�jb�A�f���w���(��w��V�Ƚ�1X�X����Օ<�w��A-^�rZ<2e�BԀ<�g'GgB� �����# �E�F���G[���Y	\4�Th�|�`��ۍ��(ABM�J�D�x"1�Iu��"h:�)Sr� G�
�d��Q����b^Rϵ��8�<9`�!�L2'��r�2,�Q�m�jx�F�ΞqN
�ʘ�~�J;Q� �[_��w�qrq�}\C�c<c�2273��;S���p��a=��������[�2���,���[gD�"�x��K��V�4i�Hv�Ϻ?��V�f����^O�?���>�
����S�,��2l}����_�,�{koN4W����l���� �x�\_qMo�!��b�r��FF|	5  ��IDAT��fd�"4F�������������3{*�C�#"�˹z�Nȹ� �? �u�NV�eS$Y��K1���N �|j�SҰ2����� �>#�M)5��)FӄF-�>�dg�\����S\�Ơ��c\n�]i�g���v�ڲ��y�_������=J��+� ~�f�N	b�|���vq��(7�0�;j��z� �����a	�l��xf��&�$77[�fܖg����>���7#!� ��3	lN��,4�C�'V �ٵ��Z�h���k��jF�PA�9�w�I���ͭg��܌:�
B6��`� K$�ۍ�PИ��<O�p7y~Tנ�0�1J�K�<Vk=���Or=�&/H��(���4�;�so	8Y�._�����(ѡr��5������r�NH$UTzv�lV�4�.��Įʞ7�J�=]JJ}�'h�7�9�c���2LǴ��|���<�ӣ�~x���ݯ��_<���?����x!�B��-�B�K�s�^�T��;;?Wy����kg��%�ؕ���")�<x�Ò�«w�ĭ?��wj���#�w$�Y��<�����xtLBI�'l�X���u`�[�٠��+SN :��|L:'� �.F��P�g[�W��&��LQ���@����޽{o��G���K���=���dbO�<����v��qI� ;:��}�;iqkSi��..>ٲ����3�������.�x�wo�ٟ��g��t�k�YY�ao�F��XB�Ndˑ�Kv�@?���Bfn���av��fd�8Y~��@�!9M,,J�,U�E0>������h�g<�ԫ��#};x&	T��x�UV�����QgˠCÑ��2a�����g�%i��4DV琬�xP����f@�|�d6�جA���7Fm(3�v�9�=h�Q�7���O�Q+�Ңܣ����J��7t&(GFT}�f��vb���y�夰�}^�����dE�(��ѱ��J�ؒ}�h��a�r��n�p�$�<G����Fɶ��=1^>����U��:RY>�bt0:I�b�gw���hI��0�����N��ņ��K<�J�@Ҁ��@� /��5�+(}����ٺ�*tg�e>/��)���������k(p��Ȃ!�%{�{��؝S?�;�.�9���}���ʝ��P�9�s6���� �\w�ّ��ɨ�����i ��S����V�n�#����x��5�2��J�(k}���$�i���ZҰsGv���1�%����sa���2�*�u�=�<'!�[Cd��m0�L�sl�>�V�:��'��4/^R3�VIk4�3��H6C,F��	�[M�S����e�`��Y�k�����:�u�=g1$�6�M��`ҡE.kq� �4<��x�������\�zP�� �r$��F|q~�,cuj�xٓL�灂�)X~�u�K^�ƍaT+V�{���Z-��Ӗ��I"+u��h�s������o����v�^9�af���T
�^�t�޽;vt|��	�NL�<5Qs��
��Ņ]�k Fb�W�хʄ����&���pgk4�s#��8�u'�}��x�|��X���z�Ł��X���f�f�ʌ;ߘ����h�ԎY�\�1�r f���rt�V����-�x:"ږ@�֊5����L|qY?߼yg/�?���?ڦ<t�].�6��<��Ǽ?�K�k������ѱ�� �\�O�>��@����׼y/~z^��SY�>�;������l̧�)�])�x��̃JU;x@��K�b��B� 11)��`�T~ZE{�NY�X#�����3>�|1ZD]&�Q�
��A�f~���%+-iP&�F��6~ϨMc`V�G�0���X���ݠ�:˄`|�u7ʎ�R�	�X��d*j�q�aw3^��l%<M(c�!1	G��D'�~S?���)�������`&�t��e����ԑ��8$yra�C{S�ɫ�K���V�|�,���غD֭�@`�S���9_��rn�+X��j�m�k�ā��H$P.y�`"w��ה�X�Eg��<ɿf�4ܚ9^��q����p��H�R,@[�0�i	��lȈ��Z�E]�1<|�s���E�Q�~f9��74�� w=�j%šv�5}�U{�h6����T���G�l�C�㚚	tH"�҂q����<� t��>�P�Aˈ�d�M7L��KC�VnFǅ{�ڬ�1i���L��k��Ό˴�]�S�ԒW	F�Ȇ��u`����-�׋��.��!5 ��sRą�|le3�a��ㅴ����L\�Zz���S�k�b����	2�Yc�� p:�jf�r�'��H�^s��ڑ>;Pq�!�g��	`������S�X7�{��7��A3��u���u��4��f[��K��^�4w*�ީ:�+ѴL:<�=����xr㋸~�(�q��*$���ĵݭ��;w��g_��Ky��� [&� ^F�xpp\@�I`��=��ZS
"�DGplE���7�ԯ�eW�a辷��i�iɛ"�of�΀_�1M0� ��DQ�^�#����[��"�p���Zv��bG�fG_	�G�g����q6ir��BI�Z��Ã�\,*�'>���f�g(a.�b�]_|�����1��Kjz�i7�_��{���=?+��vv~����n󎷍�ц�A%Kd��`#�f���~eBz^~�ww�����ӛ��By�����$>�e�E� ����C�l�ߟ�u5ʜ�.�vCZtM`AF	z
κ�I����@��Y+7��|��r19�0K�8js?>ĸ}.x� \��&>#Ԕ ����J�CK��(�:N��� �*�tto�N�YIJ:�\�pG��rXQʙE��.��P�'��í� �3�ݬ����%E���|��:�l.g����ַkQ�%5^��o���M�YĬ2��Z��N�I,�wߠ�An��v�n��5�\�a�W���y��1!m�l̘�e����+�J.�[�������#������ \�u�8f}jƙ�U!���'��U
)?{�a���h9l�K���F(a�I�5��G��Lu���D�u�J�i��X�X� +^���r���\� Cҗ�n�\���뙶����>�`�0�;%�����?~f������a��N�W��Ȭ�<KZǩvD��X�9`�{"q|v�|{oݗ�ɳ��n'I
�$��^`��G��4�P�:��$m}��u�!M50���=�*Fs��f`REvl�,�8�{�ޱH|����
��C3���2|�Y�q��zk�չ�d�X�������Ov�*�F#g���cӬi	�,v@ݱ�1�`�b`��Gs���"�]o(�CBsprdc��7y��w�ޱ��;��k��$ɍEh ��ġ/\S���PWޒՇa�R$����/��9����I�|1fp رD�y%g%�Ȑx(��쑿�����|gw���=��hB1������g�'��n<��%��N��kH, En������|^_.����,� �~�8�a�������9d��]D� A�H?;45�4k	,�=L��)���{}��?�d��=�j%�,���"_ҔE��2�oM#���PR{��n//m�6�H��$�������?�~�v���{��7��낌���<z�3�eZ���͡i͊�Mw�rR����k)�
n �<�)�;^��������b�ޫ���~b���ݨ%$P�\� j��jӞܻcg���؃Q��a*�g���H���C�77b��� �:��Z� 5a�,��O�#�������N����u|��؋�%��#��'Yf��4'm���-}9���6�Z��+>R�	
?ү�+�!�^&M�4E��+��Y��'��->�����vt�JǠ�FY����U�.�����<�\�;ϵ^�t4i�HӘqZTN��U#D���G��n'M_  ���30؊�w�n�UF�9t�q�v�,��9��y�D����!�DtcV������L��PdCn�VW���̓�ˆ�1�%��`C�?+@���y�[Y�w�X�@*KLδ�.�����إl�G��ٳO}i���m����vnQf�g8�#X�/}�t��o_��� U�3�Er��E?������s�.���ĐJ[��MbA�Mx5z.�ԤO_=*�-h�@F|�<W�')�&A�'|��b�fs�X�E�s��ɶ�H�fk��������,��*VA���3�:���o^��Z�A4���q1jͩkY�"M���&ߔ�l8�D�{� =���\mZ��<��5i��L4���.� �5��^uv���[߈�)�r��;�w�q��'$�ٵG�\�NB0�e�*T��d���,  A��̮�����8ı�7d��Q�����-��E7�����B��w�ڷ�>���A%I�&�
x:/ �.%�w���%>Ck��Ƽ:8�1��Ě���5��X�)d19�k��~B�����h�_�I�/�.h�����~�qV�[�sO��w���8Sȼ�,�Je`ƍ���6z7]\13������D�(��b�}����|��]Tz��{��3������ٳoi��!�ٝm���v���d�p8E����f1r��:G��&;-����s��x�����Jw�C��Y�c>)ٛ:u���|������?؝r��z������^ۺd!�做A�6���<Fo�	�<9�5/���M�wa������e��p��C��P���lO�>�g�ܱǏ�5zD�Q��U��±&�G����u�wx�����|���/����wM�����H_;�ܼ5 X)�΀%�|����v��A�a�N*���VG8es=���MS,�n\����*A|1�� ��bR� ���5�u�%Ƽ C���M4��Om� C��CX�+u���{���J�%7��C�[?b!����k�+X|LSlF�L��;����+7��CR?�G%�^�$��������Bz-78�gnX.& �a�υ�b`�d���.[g!L�����X؜�kwB�� ]��5��m�g��l��k���(3JGX�#�?���r�Q�֎�5b�ky\�g��n;FP�,��BiTI�';&�`9�9Z#����[s៶���ݞ��6�4�n��!�Z�ԁt�ZU*�>����~*�s@&��e1���t^��e� ����Y'��OE�Ai쨩b�����9h�͌��Ce�g�>�0+S&���)o��ȟa�M�v�n�Yluv��<5&)y7:�2��9��ؼ���4��futb_}������)A�(�\���L�J�s��!�(��c5���P͂�1���Pf ���
l�{�<F�"�g �yۭ��1e:�:�bя,�*��޽s���S{T�*4�]�M��r,3�N)^?,X�<1�xT�C}���w�[��r��I���/�+'&Ni�Z����6����1�0�z���eRMs�$���$�ai�K�J��̰u�#碏Y�$N��V>����^g��� R�9��0/�M�+QN����D�p�������_��~��_�ciE���P8�l��n�-�}uC{�B�5iZ=��3|#:ʔh������z��=Fr�I�lQ^�ک����q�5��9)7����ݵ� �K��|kן����Cy*.�s�N����*���e���K���mB���G���i����Z�\Ї{xo�'w{|���1X����=���cP�+�T��ؘ7��p����.6v�hg�N�{0��H���=H�͙���<��NA�g*9�E��3N�ٙ�ӊ4:Gw�C��D�M�/j2�>k��i\�Mx��t�5���k�k
�P'�Sf�C��6�
���k����=mHe+�jlP�Cՙ����,�M�ˮ8��Z����g ���a�"ZiR	��.f�)tm����Z�d���G���6z(J�,�Rl�e"6�;g�48x���J�)3�sئ3j��]�j�v$�X>X�^;�3L��LQ���P���,����k���+J��g�� ]�K��4��o��/����+�p�ޢ�a��=�D���Y�}�C��}Gg�V�#{�� &Gs���WsP23#!�� ����y]���AeP(ϲ�C�k�fy�=��:�8y��r}��k�[�7�C��C)ܮ1c��Ts�s�-Ě�B�@-�C�hP�����X���3g�kx���ޔ3�$�v�-	ʆ�����sz��'�Hxf#;�n�i���F�o\�L� �R���2���Dt����w�Ǩ�Z�d�7x~_C�<��~i>�Q��1�5Y)�e�<(�� ���r~.�./6괥t	�W������OJ&I���[ͬE�rk��N�%���+5Ќ�sž.��:dA���17�"��d�X�Tbi��� _��Z��7����94�ƈ��owY����3���F8l$uy|r�@{s�k���V~n	�����϶�|a�����ㅝأ�����o��_���߿KO��#j�=ԍ��C�xk�}�����CF���l���W1�o�)�T���޼���4&�o�]]���Տ�P��;?�������/���??���~&�¾��À[���'����af �����˗�����ƃ�F��j�HtN��gW�J��,�kg�2_�n_���?]�|)ڕM�T�|��q{@���	�o],μQ٨O�7���C{x���\�B{_�/so��Xsn��~���^7r��H�
�D*��lU ު�o�7����Q'P"BñF'","*�o
�9ޣi�`3x����7�1�C}(��&-�qV7�3��O���������M�����a-����aMPl��F�r�Qڍ`��E�q
���'��߼�1GCM��Rj�����Iӳ�ɋ�fn}^$�'6�Df>}����-?<ce��;p�D(2a|�	zB�jZSίT�ς�A���?�v�/����^������-�X�>;�KS�8cgx����l\��ó�I���?���������1JT��*1��Ϡ,�㛧V��g�,7@�Y�.�O�T5?22>]�^�1S_��	�%��PH��"�#C>P��nh�I��	~_Kű�;bC�8x�ʁ���fo�ٹUϮVkB��-��bs�����T_�j�a�DW˥�h�����k�/7~	�.vx0v��{��òŷ��7�!���FM4�`��n�-���H�/P�g�����ڔ�Ø{�CS�e�f�uC��B����֚٬n��o�C��3z>?�zF�R��H�a�	��ɻ��vऽC�|�,xp�\F��螋��O���r4����r"�[���L���Y�n!���ɻ���2���H��X���E�&�Oc؜�by�]퉄Ԃ�T��}P�y�)�3jID��Ⱥ���+{��u�P��3Ϥ�ۗo���	�=j�(%�{<���sv9�5�'�	�F����k���\���X1�6#�V�^^��q�YC G	�￳��{������0.��ݥ3������ڬ��J9?=�������Ջ������O����dɺ��\+T>xpV �]���C.�;'��;]���]_�X,F  Mzv̱6+9��q, iU��V�;D���� �L|8�ѝy�^�D'ӈ�iI�����p=�	N.���j��=2�{r,��1h�-�(�&��eV�.�ih�b��I{�G�$Y�#��jݣw���{G~���|$�V�L���
�3w��D�ܻ����Q@"32�����<�=#����J���������Znn�2�� ���VwiX��&��[%�(�B�	�H'F@�q�j�K��2w-J
��	��0ڦ�H���h��Ea�� � �u�)P~d�N��eag��n�*T���6�Q���j�ٮ�vZ��D�|�U)�D8`$:�N!e� �1	�7�P�]7�٠�6m/i��s��k�+� �(=+��ԋ9���5-�C5�/�>-���c9 �z���4��
�h��"~���F�ãiMW�Ϋ�_W���~���M����s@
���{J���u�Т�m�P��Oig~��սT����6�Di���e��1-��{�	DK��FZuND�9�s������R��@wJ��4���o�X���6;�ج�b����Bɥ�ӊ��	�6y�{�8���^��ЁN���^{+��@� 0
�כ#�i,��>�i����:(�L��A�E&���r�'~ǔ]?,�[�A�	EU�r&�a�|Z!�L�.hcq�!nJ� 1e���ٸ�Բ)�Ѯ�Y��U��n�A�dG�Yks�א�I���@�Aq
��L�N��0�����] ��9T
���=��Kr4�
ly�Y�P��}6�jG�M�m�}���N����Y�ףˑF��F&��`��F�MD
���q/��H���Q� :�gR��͋�Q!�`yO�ɩ�)@��Mh�+�An����29�ڕ����ɅP֧����]���_7�Q��LGȍy|8f3D���z3���e�o߾% ��傀�������[-P��kj��^���2N���	w�)M��p&8l@J�P���wX�2y;cTP�����:lH�,����pÇ��L��*��Uh��Tz���t�͆�@��e����Z�
�~�鑎�r<p� ���:g�H�����[hJt�K�}3!�-��mY�y�����������>��HW�=y\@����K�~�L�	L�Z��d LMo)�hF��"^���-:P��͂��m}b�P����0~(�X�*ϿW�d�
JJ��G$V�%kӀ*i>�p�����]"#�(�&oQ@��W��n�X
x���j6�M����RQ��K��5qcH m6gsV�F[�����h�05��$v�\���mU�yT�);����I^ݨ�d��E�N��mF�z/Ba5�+�����{�|���t�GK:Y+G'ʯ��(<zU���X�G�C�c�O�����6
#Hn����.@��R6I��xx�8��X�3�>��S6�nU�
�{a�°�(�GY�o�/�fWSm>Z����+H.t�-�[���2R�	�%,:\���R�?;V�}�5SUi�2O�@N��Tuqߖ� ��޶��jK>6�fU5޵6�?�u�(�2��t\s`�H�X�Ks� u�}�"��&�N�{�Sݪ7��RnoG�~�G�H��˰W��Y��.q	�H��#Y�x)]�fC�5�&sp)/%��"�u�#�T�U&sc9�R���G��;���L���Ч}��h� ,;C!��?!�Xyw*��x�C):�f�4��64fp���|�:�V�@��1��m�j�����ŵ1Q��Y��}o����Ρ��K97!W/��X�����q��TS�(��'P,6�t�<F�{Ed"-ܭ�9:>����@�5]	��[k�l����X1��{m��*j�#w��J��!{{K���"�M�����<��ՆX�ГZ��vz��e�P�o�J���������h�" 4�Զkv�_/f��
�<H��i��GE�������4��2@��VwJ�].�S�7�F���
�b|�1i#\Ѵ����(ٌC� �1.���Q�w��ɞm�{�օ~�-p`����8�\R��S��� ���"���B�Y<�m���¬��jM�0���7k'� 覅H+�R��
����O���ӂ��q��b��<�4�&�� �$�{B�4�����Kk�h���ށ�Fb�Y'7g��##_EĪ�K� .����Z��$x�q��0G����j���ѱ��HDO�?�W1Oa8��TR,8����-��{*������"d50)�nrN���C���WE�wX�X>��VW<�2/&���/��L�m�䜻TC_guQ�G�&Y)tp@�[�/?��{�u���Z%�e�&`4R�
����Ux_9�*�!��_�wF�&�
�5�}
TƟ={F���}N� ��a�g�97W�4]������h&���!i2�Y�Vz-#P<�l��W#E�b�*��Z[ʨ���~R)�������[���Ƕ�;/N�1][�>�ߑ��ML?P7}�q��\A�qLm<pIA��N���P��Ո��]��#�U$,����<"��i� 5L��#1���/P
kK�����L\��_�naT���^%!��6*���W$:��Z��6r�c���xi�m6Z�'H�y3#��;���� ��*tmQ::�r�Mn֙�������<��-��O�'��FU<~�5��V.��]-�H�6-䛨$
�[O����C��9�
�������A�$��hW)Y.��|y3ETi���z>blW��r��p'�2�/��钪�kd8���1�0�k���j����U�F�bw{�z/��,��Ao��j�0��{y|����C���֘-�(�y�w Ǉ�i�����M���H c%�U\��,H�'Ѕ��܎h����h�������J�t,��i-ݛ<��O�;b����V��oU*��.Ѫ�D=m�����x�\��Vfά�>���z�6r;<�h�T�泧W���:a�oN�$���6�#�Zc�&�8�&i9:��z��?ȼ�$sH����gЖ
�.=v��&��Ȅ\8��8nV�I@F�h-��H.la�QQ�ݻ�I��C�:4���j�#5\�p�n��{`+���C�NG趰%�G��:���8�,���bK�ˋ��=K�hZ�q�#�6����C�s1�ѡ�S �;��9"Acr������8�Q�R�+��b���vmM�D��i$uj�-��c���m��-�9���!6���|�4�*W��r������ '݌�Iu�	�>?�o���Ә��8_8�<w��i��LX�~�Xr���HzK�W�����k$L�ym�:�X�۠}`��.tb��e�/�,�~\,հM��U���t�!���N^�����ɏE׀����}Z'������L!�L���E6N��:�] �Q��2]��$}b3�&�� H��{�3��Uy��re�^�qҗJR�����ɉ������m�}8�Lt�!���H߹�l��v��-�G���C�����Y ��gG������-����Q[�E��T������=���O�wqy->}"��&R�:UW�#�Ժ�\�;S6H��Uc�U��h�~����,�����1ݟ� �-���an.m.��XD���V�_��j�E��͞X�! �u��Y��`�)��R�z�����]RD�y��M�3���T���jU*�@QI�s��� �5��N��Y�`���XT�%�,R��=S��M�C��l�
�˶L��J\n}m��6_���F\��[*�"B��GGY�!�c�QIQ�4��s��F��s�E���=���W<gZI���&6	 o:�ZgT���N	�b��	�C�t3Z��cU��(τ�������J�[ V�# �(��6t�P�'�K����%&����2 ��	W[��an>8�kT<\��B�4��y�0��Ss�x,����MH��T���sB�@�6�&e�g�¤lu��m�@���q�SJ{;���*��3 DA��{�͖�8���Q<J`�ĄwY�0U�5e����O���FK` ��͒����\����-%S��kհ��6GB j@�=�?�ý-�J�k�u�3�H�Y���޿�fK���N�uQ�g�?ݛ�H�U�@C��hUb
�����T�X҉���Z�="a��]�xeo���ϻP���Y�����z���kk�NI�59ꬽ#��˰�t���:K���Du��ˎ�&xr�
�9`~�:];%��9���Z��t������ѯѲ(LU<1������K
����1��^��i]��>�(�H]�*Ȍ���4�!� ���K������^ۊ����.��kڧ���8>#rjq��v�)#��c�
�:V/�5uLʆ��6�FK������L��uW���O1r��D�N�p���I!M A p���<�dL��7�{�t���p���dv�����'������|�����a�]��4ԃbT��s�/���0�n���{�iJ�����/�`�V��2�؂�~L�
jUpV��,��u*��(��2�SB6v�n�l$C�(�����^|Y��R��Ս{腾�C�w�S� ��:� �q�z�þ7��3�}{�n-
fr,f1��jq����}D
��Z}� ^kL��$�ذ�-tW��]�x��"� ڷ#���}w��=}ھ��Օ��t��^�~��^�h��K�y˖#%K31f�Q�]���h��;�]ݾ-�Յ��l�ޅ���w�"��I�r�NQ(���������P��ȓ�jޟ��z���c���~|n�"`¹?���,0H�,-���x�,7Ftdw�O�݈(�T�y�Z��sZ����Y��#�R�hQ�^�F�z��w�h���Z=+�	V�Fn�J�#5�^�
��6�{l,�_T��8�Y��oZk֞~B���'lJKz[��a>�^���=2ztx�Ǵ��/��ų�4����6P ��B��WL����o޼���N~����ٳ�Lc_N�k��l��b��j��XI�H٠����^>�~��y/��%�����E$is�u:I���I^>?`$�o_�"�c�����/NOO?��幥�:3�o�j��e���3�q}������4�L�ʅD	�����c���"� �'t9v�_�n�ݨ=�����*���"|ϣ�f��կ�E���%2���_uJ�(����bgQ�!誁�{���G�>�?�`�+�gb/���<}L=�V_#�؀{&������ք�:uYҼ:_T�Ģ�!f~t�b4�c�h[97H�����u���� 1��ԗF% �N(�U]��������J��������r�2�*�kk��M`�k��6"JɆ��/���|�x�H)ljN��R�" v+��/O�_��w��7��wOI�@K0�a���`3S`@�a�xB:j|�����s�Lv�G�`Kv�a{"}Z�/ C����Ǭlal �R���is�@i���M���5Ӑ�s�g���9���lMZy����_�E^�~�(<"{�?(�M���A^�i'Q܀=��=���\Nϯ�����m��<��52V����T����gG�"-T��u����Tև�n:�ؿ�9�춹�RVbvJTrʩ�P�bɼ)����B�ڊ��/�1�G�p��%����z->�}S/R j\kU:C,�T ����l����.�-,o��u ��pZ��z����>���X�j�4_�x��g4���bWB璣!�p$�*�'_*f~uf���������bF�}��!�Q��9 ��d��
:j�nV֡b�i����O�vmTK��^9?{{�[[iC^û0�O,��]凍Y���T���c��b��ڄP�.jy74'�Xˁc�~����c_6L�P�����Y=�����E|z�lPI�>j4�d�O�}ʢ�d�l�X�8R�0v`���H)��\"5ʶ�7>�����D��n�'$��kM��%��ųg���ɏ?���?��ɑ=���b�Hk�D㛎q׌7D!Ш��ww2��E돻��b�t�Uo~5��Y�@���	t=K�fF�޷�~���#Fpg����ѩ���hr�ם�*���k�p��j �*��y���S���ȴx����k3��8��#�c�Pz��G��&��)�0 �+��t�����9��h]֍�6T��Ч}%���Ћ�#eC����������������"�eU�rt X����+E�G
��I����\��{�҂���&4T���=1�hk����^�}GN��dp0�kC!�I�����;���_ț7/���Wrr|L���P*����X�+B�s�{Nm��%���3]����D��]c 'R��� 9c߼��������K9<����d�zEG�e\����V�Ŕ=%Tl����ե�\����T��zMq��n�}@����]�� �f�( �,���?'��z�G��'��̇ǹ�Q��� �:� ����.�:
�k����;�a�/TH8ȴA���ǳK������̖�B�1e:��ڄjT{mݕ�������'���
ě�J�<cfc��,�3�~����ң�e:����ۇ?2p�~b����C1�ڧ=�LE і[��k��ѵC-O����Oۻ�K���ٸD����zD2�8�ފ��%F�D	�U��\�'�Pˤ��a�k����*�d�c�ź�����<��22��!��G�������VXa⧍g�jõ��}�1r�@E���}u�J���b��ū�r��Y2j3�1r�"�0PƸ���鍶*<KWq1i
 �Z�Co�.ݢF6Xl%hk�H]�.�W6!%ۣ��C��diʼP��0>����`MeM�?j�o��D�h�u�r��*s@%[�[%0;of����M^���X���Kٙj�ph����w��& ��o������`�����[j��n�RJ�W�1���ʨ5�owo[^&O���w,�@q ��+��JJ��esrr� �u��c��T��/6��d�/.�����6`�=!;����W���}��C��3��+ �򫔜��ɴ��T2���U.��Go:��o�T�Q� Bk�)�QxEFٖV-E>���sȎ1H��5��s)6V��`fd}!���#������U�[G��q�h��{#�HM�ה�~�&�����5�H��u�����5D}�pt�z�\u���#]oQ&�<�t�(�0
�Y:�i��}hs�(
�NO?3���ky��yz��� ��*�~�+���K:�x��M&ON�r	�Ӝ�쀈�ehe�� X���!Cdub�1$j�8N�mM�7o���߿�Wo��pJB?b���F���D��d�M���f:
h���x��t�.��{to��H��|8��q�G����*���W�@!���h�B]G� ��:�XM�6*��=�"����aU;�3��Z��ʱ��*Ͳ�E[��F�=Cvx|~�\���,���;�G-l��"�<�Kݮ��3�UJ���dL|��׹�X���I#E�Ŋ6$�7=��b��T�μ��)����d��O;ˑ*�7��wBN����Y/�Ʊ�x���6�B�6pT�����Ci�I�0�0D�F/Y��g��p��y�4�b�Ѽ6�Ȃ���,RF-��|��21��<�6V�'\�_����a��g��5�?���Qř�o��m�g�%��E��V4""���E��RAԔ!|���v��4���p���^k��&5v	�d�C��/HǑ-}l�W�6>��J�u77��TH>�J4@�Z֊ �My��W �[Ӏl�N^�a{�tu�{�V�,NXC*!��)�{ZB�l��+�t��=N����w��e�NN�x�ܢ��<y�7w�r~y.���a�^�2�{f��)�y��w��Bb+c�34l��8<8�~u}�6��d��IDEQ�����9�4-g�'p[�[�?���u�g����g���S�a?��ģ�>�JH�_/��z�+Y-U��9%ɳ��������hTRZ]וI$���S-B�:$; 2l2�*�鸧�P%W~>��A�~�0m�9[G�<� ��M���Q��rz�/�X�R]�w���f��ϻ��9h�+0�թd��B�͌��άr�9�E���r��\ �/fsV�ȁ�uxxhN���⃃�f�\]��>�(>y��N����erz�̤M��.�v$�� �P�qil�5+��A[J���Y�J$�^�<�He5�H;�)���*?������O9{
Y7T�I�?9<��ݡ|I���Vm8
Z,������}�[&�I�׺�U��x�cd"�
�z�!��Կ�����u���@��vw�"X�E���\m�E�6����q��<�_ڛ��v�{m�[�����\^�k�O6�Ɲ��V���wǣ�ḬR2Bȸ��Ȑdv$6�3�T�K���uzSʴ�Ѻ��7y�Q�o9���*���
���&8��`p饲��C���������@>��"���J~��%���K�G;J�,Vq `�ĵ�Ԃݼ���1����"
������SZXK�SK����׸ms3rLz�!�ad�?a4�8y���H�x'a�(� @�G�ɃJ�[Դ���,>^�\ ���G�މ��zjH�X�5��wm��2	 � �X��8Lf����ʓ�۩��p��ue�l=L�ѓ�A��� ���1E��ň � `#𺠄��e#�Z+Y��)ǌ�����������T~�)�W����A�_;����;M���O������_���=I�lH�x똖s�#�4^�~��o���R? ��+��>~�$w7W��?$���HS���<��dL�u�_?�Xy��|��I��n���j��25���
y�WS���f�f�تHg��޵+�(�u��*$��)����P%���Gr�J�l��ĹM~}~��k���P��r���������<����7��S=6Sj6:H��w�s��R��~�Gs"wU��=U��2�J�N�U�=���q��EPW�õ�
@�Ys#�ٞ+V��3���UB�����kf$Pi��ç�N�ᇹ����MrtίhOY���%;iM�8_ճZ�� e	�u:�d NaY��]��y�����]Z;�i��p-5�-ɘ&<��`ha��l�-����d������_�_��}u���3G�ªͱF����@�<N�-�~<L�]<�����Ң#����1����Z[e{g��F4��nQ�w���A>~�"�>����\�u�QM3��GJ���VN?�����/��G���t�ymYd�Z�&��żg�~���a[���/^���K�}������C�o+-������Ɂ�&d������E��@�p��f��,������`�z@B��|�<�����J��ng��W�����
^�au���Y�B_��9`����B`�K�I� V���S#b���._���J����6)�-��	8��[���~Z����G.r�����갤�P=1�bF��H:�S�3�ygka�w�|�t���V�e%C�h5�zu�Y����i_�X�I����u�*�1(G��m�?���sr�+`���au�XE���+^���"$�����J 5��	�M.W�*JC�k#�#MGC��W/N������OZ���o���R���/���G����
Y7΀/�i��N����>�G����^3��Ro��ߞ�v�(O������A+-�hL~@2�(�@cvTA�\��|��n)�D`zO�Q�╅�ސ�J^
y����¤Y[�H�m�+)ݘ�\�)T�x���p�V�*�AV� �L�) ��_����V}ޛ�g4��Щ�B���e)j:r�i�͈��d-Q��<������5{
���m�:���G-���@�*�󜪀�]#}#���j�}>C;OS?����&� ����ɜT���X<&@��` %j=���ݢR�������:�����\'�t{sǹ2F�k��Z �	�FQ�'��j̭��������^��}rviǥ0� '��̵�3�Whk3Kv�!�A���A�QX��S{��� ]���[�,Bx��M�#vi#�?�������4�G�4$k \ѯpo�:��A�i�	����=�����w39O6@�\]��Z.�R;�� ޏ�0ju��ͼW�}�b˵��#�7P�����+M�?>y&{��ܦN�DF�j�L~������/���}�`��:D
>���T��`�!�J[��s��9��l#b��s"E��k+�N�<�k�v��A�@���װ��"���#z��z]�����r�����o=2
��g
.�,o�d6}����#��<���[�^s�Dyg���}�MZTwrq~ƨ	��sp�v���@�������gh�y�M��
���!;z?�M��>W�=�cB�
m���i��� �����^����N��u�FYd:��Zj�=��O�'͕�2m��k��=�`�d��wb�A��R����F�$z���f��$��b���]h�=J`l�˥����06��� �$`��lb��N������˻�����/	�A�s��"A��<�S�9��9;���ە|z.?\���ܖ���`0^���I�t(ȹ��?H�h����R>�B�2�K5Ȧ�\P����T%�R���E:6��|=�k��^��6�-W���M�kU̒�{xZ4"1�e�jч��zJ$�%:�M��8]=r_��Sj�� �_�/�M����Go�i-��9zT�ݫ;K4ik �j����0�v b���d��{j�KY�
�~,���u���V��<���(Ҝ�)?v0���|M����0�%��౱�����-��vR �:?��B#�C�{�8�찗'��T��#��.x��u��/��	�����c`���UC���/���� �b��0)Z��� ݪ%l�|��z����c���t)�{����d�)J�ڹZ�Vt���U���9{��|�1T~�˿�������'W�w	����˯���:�d#Ќ�� 'h+�Y6%��x�Uz@w��5Bc�g����!�o-�Up� P���J�|n�߳�to��b����|b�¢� `o�y+������?�~�Fܷ�������~[�p?3&�~�9AE��m�W�p���֕G�<�-����' �g�9e�F��@LS���x���뛶�������q��Q��Ye�!������8�w�����U
�	��_���B!:w�\�T��J�:�'�b7�j���@}P7��	o ܞ��N��T��O���s��(8_W�3Y�K.�$�}:kp�4��c2XaE��$M��5
�� ��htA�"2�FT�@�Q=
�F��F��Jqb�����"Z�O���˞�h��z����t~N��ʙ�J�N����w��ai���z�D�k��0բ*�XZ�� 6�X㘑&V1�U�Q�O���_�ɻ�����3�5����j:ML6À�%�[�Du���O�,�W	PA�̀*�_��ƕ�A�I��!�	�7a���ٽ�W�gL,��)3�:��/�jYT�L�Ͱ�;���]��j0��m���7��ΏHYټ��u/<�c�2~=�D�tg�m�z^�bk>Ư�s��}<�Y<�R9�`ȁT!���>O��U�sC޼ij����.���YG�~례��Ez��%_�_i�}���P�ԟ=��گ#u6��`���tA�f���"����[�C������p�F�Q���t���3
�*F��5��k� ����5�}}��l}�8��m ����Qg��J�֣tɵ���L�L�9V���Z�hVށ|��)/�)����o�}#{b��4Z%��t��~��l͹|A˺�+��m���:u�JI0ʣ.���
���1�wU��+��������@��B��1ʷT��Fh0Ɛ��)6� ��5 Cd��ۗ�{p��,
�n��ewkʮ�4��>�5�k���>��u�����u���1�SDVQԴ�Fʢ�h!`����X���lcꎚ�� �"�	���;*��?�";�����#��.��Ѻδ!=J'y�1n������O{x9��G�~:8��m�)�Kn �	��N����"�	����(~�V���K
��Ԁ�����)y;�[[LO�1k��.�˞9qhiE�	�tab#|ws��p��oo�`��������8o��Z���T�G ��q��76&�=�����az��l�T�7�F'��o��*��I�i�/V�����J����S�D/"Π.�S�ӥ��@ݒ�E�p�}W*S�J�NL�SK���9OF�o�Y>|�,�7�?>.y|��qF�����Ek����YPZ�Mfv/�%t0�;5�l��M2�x�Kre��+�-b����:��jDc�9��!�jW��ܐ2���󛛵G�6͏ϣ͟��"P����騆�k3 ���S�u��Vp��k،�T0�~�{s�NJ9�G�
8,�u���x��$�ݣc~�Z����)����z��S�O��6�� �n�h����Y5��J�4��GU~��F�8{c�~_�9�wCMsv���VVn<c�R;�4!���!�?X�k�F��竛;9�r���ӊ,�7Z��IܞlK7�Vm��rHKP�@D�q�k��́}V��\(U]�}�)��TRlM�Y�&��a��V�*��w_\\���ό��R�A��X���Ćx��݃��>P��og80
�]˝oܾwy�/�5��P���wEKysr�$�ɅU��[o�iq�c�b�r��/�f�8���AF	�k��xYU�rȶБ =�v��
�iM4��k��ږxv%�w�n�M�׉����'���ۚ}�0�|���(d\P.�&�!�9z�&&�M��+w���*[��9�ǜ��N��aL��z{>B��:s�4P��_�k�XNP�kg��6vP�I�с�5֌��h��h6�C9=����1��̐X�$��
 ����I�9��Q|����P��a�|�-�k�.���l4V�m�X�j��)�v8�j˳��3�<es�Bݘj�CXB�0.ₒ"*)�7�	3\��1�^zj�=�
����[��t!=̃C�/�u^���R<��<��Š3����habB��玖ڢ���)���|��҇��z���G��1
ˮ-�����q��x3lD�I�ST�z���z�Fr=����{��������/QQ����F/�_Ȫ��F��O,s�A��X@I�'|v^���Wr�jb���1(kMϥ���z.|U%���ae�$J-�6�_�������m���.�k�1���uV���-�+/0����c)�
�=���\�	FުT���#q~l��aI��lg��z�L�v�>����;붣׎Z�c��(��ͽ�i
�)���Q�,�BF'd���Ǆw"���fK��ը��lն�'{;ی�!� �{�����-�n�<c��^AJ���G7T=�>�?��/Q�H����69�H�ˈ|��8Mgg_��p���܅��U���*�{�͢.TТ$ޏ�u1ݿH��_��~�7�ӥ4�"�|�|�2�0[����#���ɽ6�>�^/Y9��$q����4'.��z��o׷"g�g���G��ݒ��c��v � ��{�B�j�u��E��f��[qXo� ޶SF� ����x��$}�D9��>X6:�{~�^��W����|NC�Q�7��䚁�����s��uic��X��Q�l=m����8�F�|�0�s�4�ü|dٯ�W�7�	�֯�$DJoM@Q%�83�Æm�9������)_�;�I�M��.���_�����b���錇 �B�l���2]������/�?�qX�uX�Τ�N���Yk�8*�GTG�S��e��]����c����S��o�:��op�V@\US�E�E&�����F����x�����y�'�d*�]KU�̩�sVM�h�*��iz۴�GG��n��ޛ�y�l�,�j��fZmc��E4���][�d�f�#j�E���Oic\��-x3�K@<<�U2�)
T>�ԐxCn�p-��X4fmN�S�y.W��FY�xv��5�C\o���բ�7�` ���U���}	�o���ܲ����m"uo��ီ.,�cd�p������n��ܪ�(��k�X����߇5L��7h�rn�Ś`_<�~�9:�d3�V_�s�4�1p�� H;����4�5O��w��5yI�qi�xq}MU3m�x�Vz��-
`���"��r)�wC�],�����^�K:,���h�5��?����M��� �j��^&@����M~���|��9��y��b�hK/"��9��Ѽ�>}�i�
��V��
�2z�u�1�#~���&�-��a�-���drDnWNI�4��ήL��+Z��'t�4MlO��O��/���^%۵E �����=Θ��V��k���`�ПE�L.WK�弾�"�y:y������R�6��~�5��{��9�&����/��)��N��_�U����&���nR���P��g����r����{)� �79w��,-C#�����̓\^�0 ��^u����s�t�0Ӓ�_�P�l_�Ŀ�>�Y�*��SP�^R?��;8�F�kb��h!�j�
ը���e�V�]~��0z*��_zԶ3'}�����a��in��K�!��.v�rdr�$�_U�N�����*@f�(�4;���ٚ*����0��
q��r-�O�I�uo��
l���XF4V�{2i��ؖ)K��J��Yy�F �IԪnK4�'*�tR�b�u�_3��ח��(�\W�f$${2���T�ᢓ�9:�7S���ʑ9�x���d��`��i}�z���4`�<K�KS����(R��«T�7AU5=�" �1&Y�a�_3�����zkF�q�iɝ����[[�MA�>��5��觶Λx���W(��������̎6�R�nNA�3:���^��~)s�ap�1`ĸ���~;�Gԋ�$���37���kh֏�k	O���! ��x`]�w�Q+�YZ�?�j�P���(���C�}�����N�׺�����>�x�V��������iUo�����W߱־>&.l�=�#���ڑ�y{�����Y�'}縳=��P��������;�O��&_ 7r�Z�7���o����'*��|�tl:^�� `5�]Z�EG��к1��SCb�lc���v�֟Eߐ��ճeZ��x�����#�TCo%w�'�i��nSAo (��ȸ=%����D%^ @�����￑���E`�i�Q�������A;P�����S������� ���͠5x���4�f]v�۴�M��=��-V�n�l���T������lɷ߽���]��t:J{�3?7��'Z:44�'���(��XJ>�#���d��l��{��|� �yY���(@Ph�5�v�?��AMd3X[�P��m��͐'|Ѱ�V���ϴ#�6�C3t�	'����nYi&F���(#]Q�S�������C���󥇍n@����$#>/� ���($g�M�',�op��䎋���;Հ�9�������䝠����D�ί�nnn��F�!��j�=������-�:��	��k�ЄU���
����k$��(g��s�6���Ə�q6�%4D�fI�8?%��c��e�B�0y!:������!+q7�;�'M�%�PRY��ط�9�m�ak��A����
9��S"%H�h����j@�Y�������j�
oE#
O�U�#���mT-!]����V��9$�=��g�C��7pԆ������5�,��Ӏ_(h���gY�e��7��
�\_��?�*2htUD���;�Y��\5 ��6������_�@� �u�R���d�.%Q�������k��Ӌ\T�n�S������m���>V�ju~U�_���f���C�����`��s��i�E��^b��X�W�U��=��*��� :�6�֪�Vc�U�I{o��Z����9%'�=7	P@�6f�Erj��������C������"��L���9}�2�3Y�g��5�1����?S���3-�Y��W�=c�ׅ�f*�\/�4m����B#{l[�k�u��=���;Fd4E��2#�m0���
]4`K4��3�Z����oS=2�R�4����������Jߞ졎)וE���M���ӱT>"�����v�iL�m�|����X�Y�:&�fk{��C[V$�C��C"�?����Vk�0^���������YD4���J��s8��
��vh���
���� ̨2��C/��#����ߧ%�W�ӱ_(}�Vm�&�}� �&u5��|�HZ̄33u�~���Jɶ2�V�G#��-Q�1�u��FxO�/�kL���HG1��Q�5�@5:��u4z��G�9O�ސ5r��,�w핒�Q��2�
N����$���/�T(�֯���(�|?J�bxi�� �]��U���a��:¿�#��e<U��L�q���9z&^Z�C1��D�
`�>���D����xxt��a�#�v�(�����AA�KbxJ0������5�þ3���9Y�9y������v���ă��\�/����R���5 f�?�Zm�SUXP3�-*X߾}˔���0�4�՘�3�(p� r�#5��+6��-de�eZ��d�Q%EI��	�m�)��i�������S��g4�^�Eʲ��e���)ᑦ�ԍ9Z�C�7�G7�Q�'�3!��A����^Gv�;
�n��$���;~����'�򨁄~��x���:J��B����o^c͗��36����8���__G���~��9�+|�b��G*9���m���+�����˼����6IFOG��i�u��1ޡ)\��b�=�����VH՞� /�n>.���6+�'�|�����'�����`���M�R�������1�)W��_�V�,�X[��5��Gl�|����v�5h?_<�JSԌd�������,�'�\�lv�߃���wC�{�j�س�`��RE�x` x�Y����־��U�"� 8LGf�����j�r>"i����-<����?蜭�zL�%��kd��}�?�L�'-"uH���>7��B��m�?+�����
����+*�s��=(�C�(Z�d�`eb5��ϣy�i�<�cߥ9���K�Ѡ��~]���K�MS�]QP(�@��U���פTP��/�W�.�~�~�G�����/߳�Ѻ�5M�%2����Q,�'D<��]��)�����SHӀ��qF���:L��U0�kF���X�kl
&�/e^re�so��<���A�k��6~6I��j�V�aq�o����� P���0w����E�ǃ��x����*���l��!wh払��oKP�]gh��n��h3%zD)��R���h��PR~�F�����A�O�^�ko�x,)"W@W%�B��fKb|_MP���!/м�7�X�fV�@�m�iZ�>�ѯ�`�⩍Ѕ�aec��>P 2���W�@"b�����?�QN�O����Da"c BlE��6��y����O���	����h}�<ͻ�n�r�5��Y�f��?99�&@Q^z�����͵|��?�E��E�7�>�f�;�Sl.4`��9���C���ҟ�rc@�A�N�D�����?��WU)�EG��r��ߊo�9��7�N! ������CNcK�YE�ks��fOL'��S���[� y̏��Q�߫.�p�G�]8ց6���0l
�"R�Y P��
�{�hl��P�'6�s�A�^���5�]��B������[�t)�: � �x{��SY���n�z�-��Z���B[сה�(H�-�
�n����^~�9L�J(��'Gi]�6C����6l�K�Sa2b�)Bȿh;�ƺ�l1�jt��+�M\#"��ǰ�6��?~���>�bNEa�	��1�Ħ�9��NQ��8����O�y }��x�v�C볝�=y��B������^Z� R͕��`}д#�"���[i�Vv�hu��*?>�yuw�QV\/[��q���+�Y��+��pl��4p�1�Kcu�����4�,�F(>�f�xR뫋�s��im͎�:U� ͈5�H�<Bc�\�v����a:��N/
J�	9J�2�>�9��Z�*��S�B�����$	�,��RG���Vt<�Ҧ���
�2%�6����+��'�І�F��0����1�(_�oy��͛��Ѣ+*9a�󜸓{��}�5���aO�G.����W��N���˅w�L��3ϻ�U`2]�$P�)(��szz���q΅�q�Qj��	�cm��,C�隡ƚ�&�R�AIm���V��gJ����4m�)��b�S4v��4�e�^�_i=���vedF� �}��m顔h�#G���Z=�Eb���>�ύ��qB�[��y��68��:�k���-��(a�%�������Ǝ�Rl���l�b�#q�Ϩ>@�8�op��<M�~��R�W��H������Gc�����#y���|��[�5��$�K����4�u��7���Uu�8�F�D�[Ш�/�A���6/����W��tW�O��xĨ�/"���ޯx^>�cy�N�?em~ۤJ6fbQ?r8�C2}[Iz
�ɼ$IK���:�W?6#a��ysQBu�%E[�^�|r���u|�n �y��b��8���qC�k��ő���E�;�u�q��ш���q�駟���gLy�Q�� `���	x�1u���L.�o�s��c��^�t�bU��n��dKo..�� �W�rw})��ѽ��&8] ���C�y��=����e�-���
��ۢ2MM��n7����ۡ#4����o���m� F�
�c��^���/mI����%	�v��յ�^35e��8��`sK���N����]:���Æ�� [��I��n��{k��_���p͔�,x�����Hũ��"F.�ހ�H�U[vv�d�ޢ�����!(Gv{2��>$wh�=R.��=փy�)��S��V �ݍf>}>�ݭQ�]6S���ۑ4�G+�7�q���D(���� ���	��̛��h:hP�#�(�:���ٙK���K��1c�����]0��W����7R�_�����`��	��_D�+M�D#�E[��C�+6^Vo٦|hr(��,��s!ˠ0#�K5<j�ܒ��.�yT/:���)M݌��TVP �|������X@T�x�@��i��/���#O3e�U�\�i��e���g��w �א��͐2�Cf K�k]�h��Ҕxd��Z������=bO*�K���1g�Ta�ϕ��DD��-!j���ͣc8?-Z��_�>t#F�Ab"���3/�?1ϖ+#qb5H�h|��������fDrm4-�Z�����������_�|I5jL�M���j<&ɓ<<>�
>�	�q�j�C�w��Q��T�*9(��{Ƶ�j	7�T��;�>��D�
����b5��US��c��S l@������?��D��8`F`l��J�O��S�`-�Pw�r:���;�3f�6���>7!���\F���#�nm9�`�u�6Ǣ�0�56����u`�״�%sy��?�ډ6��7A��m���l9�z��	_�I ��cgb�XzEi�b�{�'x���������C����{:�|�����C����>��d&���b���WN/R]����e����7��yH�9g���P���k��ɳ��;wh;���$��=y��OF����� ��Hk���`�Ѓ���&9�wr}uE���`k����-k����7o^3	 ���i|W�N����T��Aŵb��ӹ�y�R�����Er�V��Y�U�ˢ:ʈ�J�^�� KW濭+�KH��F����uAq���@��RшB��QG�`:ڝۥ�y�j�T�`�|��R(�N��c��*�^�VTF�c����(��8E�	��x+m����b-�>��q�����	>нO��d��	,���m�~�F���+� u�Iy[�'���4�슠�b��@ܲ���� �o�+���+Ri�� [o<�&sc˾hU�U!�([�*�T�XF6#�bB_lx�Pd�Z�V�&+�m�e��"|~�޷NW"�d�mi��ْ�f����H�-^]}�y+���а���X� ���~$_�jA�<-��/�rqu� X��d�1�g<�a�q\�%�Ϟ��$-ʛn�MtM�&�x�O��h��r2���EkzOj2��}k�"e�ſ������H�5�����H�`ʟ�͜5m7��Xe5�0�9��;B�࣏���;�Z�-2��C5*�y.���$��˛�ҳ����!�^��s�e����eeӭgӜG�>�wx�8-VL"�4ʀ��*�t�Q����K^&R��{��|.��n�"4��a���f9J�>/��ZK��I=T�$��x}!���7���m�/˳&�(�b��2�p�V�9� ��r
L4Z���K�!�4���P��:��E��g7�Fե���&`��x�{j�T!�Ʊ��e���k����h�O�^p���@����~�6��ij)�QNbk S� ���Av0�W:���9`��DC8%�;{\'� �f_h�c(����g'��z�q���am����H��IZ�,�B�fw_��Y-��gc)^ �yZǏ��zS��'�B����cy�*��=ޮ��� �$x�����V��p���i��5�Mδ 
�b�ށ�����P׈z&;�����g��t�i�ONX�nD�9�Qr�,�X�;�v�{��`E��YF��3�FH��������p{�y�$p薔��=��tXC�Z�tl�d�{4�;�A�!�=�R��,�ި*N�g��7@�p�9�(�)�s5�����|:�"�=؛2u��t}�Yi�������*S��v*'J�^l�O��L߹�k��ɨ����m�<R�����xͤ�(�ݳA�tI�H��5(l̂0aZg���f����4b�P�{1}�����w�7���3!fp�H�(.�w�X��xx�L�Ң�E04��=��J�G���b�	�e��r�5o�J�(T�ņ���~s'��5���~�ҏ��^ڠw� �X�|v��l�r����Z�@P���W��%�&�ڦ�G�����)�h�h�r�*�:[d����Z�r�ɵ$�[� ���5h��+=+f�}���y��NRw��}���
�Q$��#LO,1�,�lQ6��~ �Л����v�P����>� �ɋ�#b���?�,�1 :���D
���|����r}{�mD&S6�=<Q���CC��;1��2R7f�d�Ff �d��)R"��1���x�pp*�Ye�kQ%�h9���Q�|P~�a�'Ȑ>:��b45�$�Wsij�QZ.?�{��>k��ע��5r�l�7��eQNr3|�9	y�L�ѹj��_k��@ʣHA��s�j���4��(��I_RwE��5A�̫����4�O�+��|�Zt�1<\�߫����%=2�H�e-�E�=�6R����P,��k(1��x*q ��x!
����B���(N�������������SL�����+����@�û_���-+���-�:r<a��f��9z"�U?��U���¨�a��qe�u�`�#R��V�ۻr�~�lmS3�|�H��s	 �����c�@>b4�zZ���m͢*���[1�Ϙ��8.���,�zkMw��AB�ޡL���� E�7u����!�S��p�7��(P�
=��[ ��}������tI�/������kyX�d�c��7c5�"�u�X�"�� #i��hH-�߉����
�	�X��V�������(��հg�Z�t��w�����t��ۙ�ʵ�����f� ��!��B+�d/�5���l<e�X��RޤJ���,��� \j�Ϟ�7mF*����[*�.�v��-��{�V)�If��ִ7t����p�4b}�Q�_s�|��tn;A�1��G�I	�'<$��qA˹���j�o�R�U@J�ӌv��p�`P�UIv8��U�H�6������>1,z�6���MZn-ɐm�0�5�l�*�HT�4,'#��^���$hH�ú�*̃RP�^p���Ѐo�u��&G9����xT*�aM���P��Y�߭/�(J��Y$�+]T}\t��o����+�[4�e&���A���[hب���'��ߓ4��@�Ԡ!8��a�xm퉬1�I ���QFVC���v� ���%����6�-9yԶ R}_ξ�� ��C���%P�%u���e��w3*���*:�c�*�����������+�d���2�Q��=���[j�#�Qyt��Dq�;�ё:�UG�Ꟶ��s�l�u4�+o�`e~J1���*u�R�_�n�T�:�N��Z�|��W�����#\��?V#'�%k�}Z��`ˁ�_k}ݛ��ڲ���vʸ�N�k�eG�֮��ޜ�U^���i]���BhJ���s:C7�36�h�5P�����kV_^N���S% �i����j�dA�k<2�.2�
�! +Nc/��D�78���f%�R�#��mF��z��&a	����]�O��H����t���&���݌k��ܤm�c+�Q���<}�B~}�+O�=�;���ɖ�e�4ٱ��GF�q�β Od^�7Ftʃx4��e�f��bA[�@R#�����}�j�@�h2cO��d/w!���"���l���F�Z��k�?D��\$�|vu�� �  ���N���B� �
�h�Ć��N�c��[3�ٲ���., x�k#�{ ֭h�U0�<3"H��3j����b��5����cm���$�]�E1��,}�γ=��,��\�z�74��kXP�t����N�J��IKN|Ǔ*��^]�`�j;�#���=���m�F$&Κ��U�'�V�2��2V���8�oQ�]7O����o�M15'	M��tHl�wg|3�$>���15ʌ�U=2��(]OԌ���gr~~!���^�}<K�Z�s�x����bn�5w����ࠠ����*�$��1�.�q�:�C�:疼��Q"��=0���3pse��"��|�h����Y!�����-gݖ�t�u_z���j�u��]�;�N��}ǜzm�8���QA����Z��e�Xl��ݑ�{x|"?��'y��~�k���%j�G�_����bᡃ�q��T���/���?b��m�+�;�����a������iZ��s���8��
�H���u�@ݗϟ��������Ü|��^�:#���ܾG��d��`���{ۉ���ѕ��Sq�|�8��^m�9aQS�B�� e � �#O������ٿ�&G�
X�����1�ކUTI׍~�u����|�*���uy[����S���C�ڣq 9�S�o �1�pb>���a��ϱ�4��mF�r$S�~��'fz��f�����^��7oy��	� � ��'��iM�������e��c�p"����d����mc��msK6����%�����ͅka�C���x\ek�Xǝ;:L����'
Q"�	$|܋�ӳ�V���������Fd�`�0;�ynK�~0�5-�D��/��|گ���Lcy~vFG����<4����Qo{&;z8�a�@�ܡ��d��o�� ��r�>��u� j�5�u^���}T`&�{�K�Ţu~��ś����39�����}�(���(��f-P͊ԶO������s�5��s��x����;	<���\�=�����#��Ջ#9:ڑq�)W�o�-����g|q�m}�4TY�ŋ
�3FS�
�T�YU	�s0��L��vl�h�N�M�ֺ��,������`�=p�XS�z@i=><��>h3V~]VD��Y�W�� � ��w��kt3��;M���D]�d��F*��Ȑ(â���cT����@��DTa�0"�8i��B�c�F����^qo���#�b��?����H���|���w�?˗�k��L�r"}��e�E*i�� %�k�\ۨ�� Y-��3Da(:F�X�f�r4���
dj�-�	7��-{AU�3j
���Y�>܈�a!;ɍo���aoZ���g��t
g@p��7"�_\�apzu̓��YW+�+��[sV�^__'c3�W�f�~�k7@�9"c ޽E������=$0���҃�& m#x�0H�7"b����:+Fy���d��VJ��i�V�'�k��E����p���*��nV4����`@${h�Ջ�4=�6Z�����W@*G��M��5�h}>��ڔ~ȳ�{u���;_˞n7�q��G�k�/Ѵ��k�=*��k��`ɫ��q`\7Ϝ���U�I��p'+��m&�VE����+���s��ː�&l� ��v����#���#��*�z��ԳZ����8��=!�]7|�^F�l���Ԇ��=�% ��̺fb�i��jAS�,3�:�q��I6��{H��ޱ�l���:����ڑ_~�U~��/�����[n��	|��nۑ	q*�R�ҋ���D���ca��A��6٪�d�({bcS��:����ӹ>��l�v��_���)�)��*]�\�#�W_�?�% w�&������������d:R�~��h㶽��ƈ��5��H�E�WW�JS^�p?�J�R�09��!�"� @�na�R����&a�
t�~�5����ʯ�HGx��P�Z���i������Z{��2��=�zhǚ���HoT�3cKI����+)�;��g��R����O���Eq��d���!�98>����%�I(�bMs��o���	�fT7D�f��iD�$X���\�ik��	iy���ĘN4m�|4��-�g.x@DŘ�l�И��nz���x�)�9{1݌Ɉ� _	t������t.�0�fJqA���$����ѳtN{�34�}�"�yn�S�Δ��E��*Y�+��f��g�e�&���9�1
Y��|��Mk��y�~�	�|?�f�2��d{V�Bj�5�_��v��d<��<�^��F���>���FD�(�x����2MhmWT���%1�Ol�B�4ߌ���,m,�L������y2FM��	�ݧ{��t#_/��b&��|��ƍJ�yC�%K����س�&��(!�S*��
o+�]�j���^�e�`��=�>���}�=������j���n������4OFy|ï�RK
��[k:G�)?'�; e��Tz
ҁ�����$�2nOE�r�����7M��KNd��Y�Κ�V�V���:�#|z�@�7e-�`j����W�qw��ϩ���9�ۃ�|Dd(�{n�2ww�i�f����C��zy�+��>������N0�ƨVTm%�TK-^WZO�Eǔ&$! ���vL�^m;��HӉ�؈�!+�q��k[�t�>|������w�k����B������/�kV�����Ȣ�֪�E�LQ;e�΄��k�j���R�������^�v5�w����t�_�(�/����ޝ\\\�gZ��O�\ự�nM�Z͸�+�u�^]���5���ZĖ��(�ȯ�wڞ)���-2Jk������K��o��W����gt	�GTK��ˈ�3^V=T9w=%i�p:�,Y_���((��������~jȋE����E�����0C�1�M ��X,&xf�������J�ުL%Eyedo�v̭�2��}�}Qm�����Y)i��W�7�,�(k��i�K���u�����J�� ���4��I�B	X*Y�����S1=/(�MA����\F�7��\!��,ѯ������K��d�fŞ| %W�%DŐ��@����_:dM�wc�<�h�^N��OrX�ӟN���_����>��խ� _(7R;Z_4 �M��E�d(I����$ѱxӒ=�2澩5&C!���gVH�C�QJ�#(����׆5�6�v�b���'/C�N=������������f�����/A��SZ�6[LHrڙ�wH�\ȗ�ό�q���GB!Q��{�+A5t��<�.*1�����	R�ggWr��K 2V�.{�2{����$'f���V��jD,Z�����s��\�\��o�p���PE��>ћ!kj�FY�9�^[x�su4�粨.]�[3O��$����ܞ�_�x��Je�J3�U�]c*�s��S�d��fd�#Z���<o��e��6T�����5��y�R��O��T!��Ħ�>_��J��{\ۀ�����e�~oV�jT��Y�֗+��R�U¡�P��M]�w++$
dw�b'rs}LP2���G�d����HN�uZo?|�������ś�J��?��_�1媣���'�B��.����l�H������������("*������D�J��'��EIj�A����	+-5}�N!6v��,������р�l�@�l� o�|�����5tN@Rn�]i��ֳ5�'*6������R�*M�BD``��� �Jq ;XfHO̩<����dF@������׺V%��)C�L�D�L��hu���`�xB��J�B6��p�-y➂tePD�"*P�1	������G�~��Nd� ��.0f�Ǌ���*�W�L�b��E���>�5�s�}����ކ��*���X��'��0:��ˏ�E�m��ߦ�r���"ͫ��x�RF�I5#�	�J!0�����@�� p�u��4��s�'и�7�lf}��tU��*C�Y�hP0�O����n~�Z�Z;QT�l����U�M���L���n:B���>|�,�ϟ�"��t�%m��Jf�I�͊G /L�E�H�|�l�'�`�aŝV'a+N����p���P�E
��-yA���.d�,�_~O_k�X�HWYǷ�Y�~�J��j�W��z!zǁaw��@�曔�k�̼�6M{
�W���5y�f��f�i��(b�2޳�I��/��<#c����77n\chx��({'���R�8�ǅz�����2�����#S� ��\"=����1�&����A,�e@0_{I�:��I3.�������o�*��4�eY�=5��m����{57���kW�{���1�!4Rlt�s���uڲ��*=�}�{�5��v�Yr�`��J}�:2��]���������)K�|9h�y����1{6z_,r�c�] �����\��IiB��+��=��u[9#���)6���͕6�II�͐����`gl�m灖;?�s�����ո�P��ގ#V�@{N��O��d����1U����׈B���!�Զ���*.Ԁ��3� �`��.�@���J7���q�>�M�'����~� �O���˛���ӭ)+���b0n��`
w�� �N*l���`����S��M�¯#?�`�q �@�DJ�F�����#v @J8�o�*&ު�"���z����������	���ճtm��?���&o��V��v�+�,8'���{��ujcq�\^�W��4+U�k���R���9v��<?��X�%Q ��dl&i���	[��I����3�wo_����ҽ�t�bŨ��h8K�]�Xx�&ςP�O����jg��1�V�m�_�ppi%�5��[��7��Hr�+�s�@���9����'�0�O޻�E���(�Y3�	����P'�H�&JLO,f���Atޏm
|���~m֪�G����b{���ϯ���bӭL��a�daE��0n�
i�#g����'��/����U���oՊ�5��B�(�M���@80,	�B�o1��N��(������%���Y5nn�{��WCy������؛vGn,ע� ���ԳԒ�ѱ��]���}����k[SO��Lk�����(��]Z�d��!bǴÑ��s9��^���,m-�ͅ:88S�������I�׺���{�������oQ��`p�e!�seP��׮�,�a�.�ϪGļc����bF�6��D�u�#H�e l��a���&��b�h�Z�¹]>$�#Y�4��L��P2T�<AZҭb8�����g�����Qo����<[[�H?;�5�͟���>������[�=�E��Y �<Cς��^P�ߧ�z�~={}�G|}a��d��:���"�ڰ�������� 5�6����?��u��A�cY�X{+�d��s����,g�Ρ�gLa����&f�����'*_뇇��ҳ���Ȼwo4_r�$[<R> w�{9!�SK rw7�®�� \(�A�1"�Dҿ�������)���k��suxx�i!6�?��g�󬚓|fA� ��g��O?�۷�����(��{+�\E����7x�IP;�re��P�����Ng�4�1W�6��.x�
'[��;&��-����X�ك�O�=hЍGi,תa���\��p�h��Z��䧟�_����G99;�Uz�G�g\�X����h�9S~N��n5J�ei�"¨�Z=���.��N�8������OcJ}��.T�.W䉻����!ԅܜ��8�Žݎ΢ o{GKAP��|��1)ft0BFz�4�^��rٛ>�u��^�&����$à�/���f�_��J?2Ag�� �]P^����/�?$t|�6���|CºG����k9M_��3�����,���çB7�\��k�fk^m��߀��\W,\�a0�c�( ��m��&@�N�4Ṹ��O��W���\>|>��®nQf�r�� 7h�Io��.������mo������X� \NU�L����~�ز`�N�2t��r�xΓ�!M���j�JQ��	^h�\���R���hq{1F��PP���"+M^����WIr�PU���c���jJr�����'J_h�kƫN���=�0f��A6]�j}9����( -���a .���}��W��XJ���|?I{e	�s�R�����F4�$��# �t�\��}�>��D�A�����T���8C3���N�S��ߒ��?}�x=��?π��I�������կ�}�;� �B`�핪����j�tMR������*�m{�j���[�߭�X6yJ��)�����^,��:������Ľ{�9-a֘y�8�ƀ^���<y�̽+�ͮ��	;X����7Q9�h���Z����96�7a������r{�m��`ca$AA3e���	j�g�B���ZV0�Ty#"ه.$��PMJz6��k�����h�P�����`�<��^+�;Ðә���y��02�ؑ��ac�nx���} @���ruqAY��Fڍ �s�y��_��<���o��_2���)��S�&��  ��ᡜ�8���}`���J<JU�ϥ����0Z7���Lks����7�7�)�>~�\Ĝ�W����{%A�n`�mp9��DM��Ku�`.�
p4�ޜ)K�����'t m�n=��{����Q����y89ڗ�/O����!Ȱ'�0�U�!�u`�X��G� �z`�G��^��ڰѺd=���br�N{,y�<G����O�m�A<�,+#?|�e�ʥ�g$�p��U����ײZޥ.�T���5�dC�����]�5&���YqP5����t�b
�Ds�r��2"j9�ǔ۠��\)�{�Ak�Y?L���M��x�+lER����\^ަ�~�6׹|:����n����nҭi�'��<�zəN�߄,�H�_�z�y��e1��{T�|�����o�ib�`�g,ؘ��m�מ)�E�~�xig��� W�#�\a�@�L��m�fРU���
!)I�eC�y���_��}��WH�ֆ�\r���&LL�z�����Ҥ�=�bks+#�o��{�02�B�Tu��]���m݇$aE2oLV�
!�e>���)���X�A��=��_�q���I���:oǬ9-;5"���T{;�������G�=;y���;�.�5���������W�{��޾���5J~J5`�>'�{<?�@͕imH���f���lO��z��B����I�/SO��M4�O���ږ���E�����-y�n�m_<,N�أ1e\����z��F��"!����j`z���y¿��s'��}���ٿ2��4.�F%I[A�Qc�ã�޾��o�0�^�D}�3�P� A�:ue �3�����f�z**!�b��AAWq� ͋�)�<��H&�쁗��7�.��?���|[P���hpW���k7�Ҙ��	��ƌƿ�e�X�&'2�Q!� F�E��=�Ցi��Zsqs+��Q>|�� ���K"ΐo�v&�\O2��1@�Y��L���e�T�k���槏&��Kے��_�KÞB���t���;r+�\���*=���O�ٺD��ٔ<k=�D	�7y�2_1�����yJ���_m:N��!�s��_��qCg @��J��C2�'�ք��\�kxXM���Á{N�Re�.�9�md�U7$]र�^IM־�ů��676,;lL���Ԭl�:�YKaeX��?SK����]Dt�~�7I�h� �fx7>��/�0XR`]����l�D ��M�d��G=O�����ņ	�88���y[2�Q>��e5����{��Oev�c1&k���^�ӎߋuj�-�[a^-,k%W~nl^�=E��"F	�b:���]�u�`i0*	W�/`˅���������D�{�i�%�\���8�P�D�ig�/U���\�8�����:���C������`L�\9e���fgToE��y�B�`:zFn$C�P�j�	ys,��|�&+��سCE"<�/���E�D�ޞ�ٗ���@_c $"2V��敏O�����^?��W?;T��L��y:���?�T��WT��?S����)p��p����yu���9�Ǵ�t￯Cb۞��z�������yN����cfoj�\ḑ�j��-�gc��ޚ�{�E�
H%��A�5����
����q��Qs�����������W*�~��(au�C�V%�����tm ��iD#|���&aü��m����W����_��6��!���}�8�F�H�su�0���HZ��<R(k�pEn4ܸx@Z�z�^��@�W�	%O��/_����]����C�܅w(8��������_����vrt$΃�N�]�SA��4q�5ه��t�YZ��5:�HB������e	���O�oB��k%Į|�U���zYcT
�M�Tʷ٠Q�F�5��/+s������<<eeX���bMz�.������\�>�������b:t3 ����0���g~�=Վ����*Q$/:Ԩ��[�� g|͵!��f�{���B�A�q��O!�=�;մt��Z���.m ���Dh�H��Xǔ��P�ȷ�_��+`��ݎ 	��fUB��S]�i�26ZoH����O��zmܙ�������v�C���&m2��x[0�t�r�mw���MV��7�2.�<���xĘ-� Z
0����A��si�����Nߡ��$NTZ��ث;��P񀅐�M��L�I��G����gKί�"��\���"�fȞ�����Y��d!ϭ=<��˧��Ȟ9�M+�q����Ҫ��o�T @�{�tNEkz��9��[��h2��։��7�P8��J8ڕ���,��
���"Y9�GY���J���Ëe����99!�[Ys�|��\���1`�;a��	�+�=���������|��ρ�<�^t�«�Ί�d��u�i͘غO}���;�j�ISY�m҃
��z��(����U[�ո=��[�~�t'�X�w4��_�=?gF�(MN����'u����G
�*F1ē�գ��;77wr��B�>�� E;���15l	�9��r��N</n!n�+
�)��{�z=��'dGgz���^&��u��up|��1�Y�P%=a�� �\�*f��y� �����l��nl�hv/���l��3���7p^����3�d��0s G-�$G��	0a�wɹ��O�c�.@(�yx��Hc�yx`��ݫW�w�b(O����d�����Kh'ܟz�1&M�q:%�&����F�^����*�����t����D��Q|1�ŝ���Ӝ)�^'ؤ�����;�U:T����0z~cõ��z
q	�oʆ�Y��a�_Q�Z�������ҵ�UЪaє5�ƪ(m|�=5�����d�(�[�������$�k=��/�m���t��A���>o�?�Mu��,��u������q`vl^$J�"�`H�/.OT�V<`�:o%����V �0�/��?h�Rf���a�4��H�'�������O�� �l��՘q�$d�GaC3՞\<T� �.��]�ju5����!!�]4����e3�����{�ez�R�uoM-��{�Q��ufB�D]���S��ʝ��q����U!8��E��)Pl
�y(�_%`�;C^Q��)`��8��I�LYv��?z|~�.�������{�1��	���M�׷2I{��(	�i`GX�әz��5ۛ���_���L����\�2��NA����6�mY�>��x;�*0�z�IV� ���T�qa����d���p�4yG�w#��J=mς��{]>.��RK����k���߷=`5�XV��	 �Î����8��۶��X]��n� |\؟>���,c����/]/ pﴂ;_$Fө�T)jhMC?���-n`D���1���6�.�R����:\�r ��o�wp��_���ߢ�k���s��a�k��>���;��*�Ne�
��;�����hCk(B퓷�5w��x���Z>������X2�6�jӖ ��]��F)3G���V
s���!�#�5�}aa��s��\������?���+�;�l�����X޾|M�yV���ʊ��f�d���̿L_��U�~8g��7]�9`J��^�\�Z
a�ъU�?��^���5�*`�g��X�m��m�� m��P/��An��Ǉol���&ާN�{+>"4hr���#{��φs��{�~ƍ�_�ҿ��^�A06�'�D8:0&Ɥr���$���3�f�F�s�}�.�.ڎj�P�΢���w*
z��Vƞ�qnEt��1��F�׉V���gL�"�_;y�}�~m������X���hJ�V�h=����e��|!�wجm�P0k�46��*^Tѻ�K�ø����C���H���ƒe�Հl��:���|L�6:�l�${ _ٔ!E�J����U!�&��$�����v�N��J�{n>-
��x�ʃ錩���G�_ҼK���5��)�G�N-+/G�k�]?��e;���-��=��y��;׫
�d\�h��<w�U��@bf}sO~fw��9(�>.�,H[��|���]!7��Ф��|o�K�3i5_�Ϟ�F=aHu�6�_v ӵ�s�*�w�Nӄ���z'�o^����1��I(�G�bA����b���JӋ�u�J6>)Oh�g���<z.{�#��Jk��,�ۀ��,�}�ۺ��z���;���ly���w�#��(<P�ٕ�?w���ǟ�U������|��ն�����~�lyׂ���i+Z����0,�]s�4����P������ܨ��k?)t 7�8�~aH�� C����-+�ၿ'�0�YIW|�(�,��&�R����*Bk̏C�	z�&y���0p��j���ϟ��i �����5�mx�����Q6_���o�Nn�Yf�''�$1Źm��r�Z�e���i5^pΠ������.��>ȷ��0���BQAg{�2�(��d1�gLW	���1�)�d*=�~���nn^�F��	=�"B�Lm����2
}lQ}9�P)Y���� �ML{@:�T��������n���+��N�iإ�L�;L�Tz���/��:l5�'2YE��������"*�����J�$�s�����;3:��h�Z�j�F���#7�l[�/��/��7Y����8�ڏaM���h�uV%+�}���!Ʀ1o�;�2���R�S���Ү	d�K�&��5%�HČ9.̋���$�U�2��?���V	���>o��Xf�� ,�S�8���1ګ�\`�+�B���ӿ� ��~i�B�%��F��>�t G(`���a�X��� � ��%��L,���5�a+̒ȹ�E���ry�;S����KL�|�*�mъ�ױ$rS��Xa㥤�ţ5��?�y��3��]�R��缾g`g7�+.�'%���W�;Q���E�o������\5hm�j�8ԹS����NΪ`g
�_8�m��Zm��K�ݺo�ܶ%�A.7
�vfrzz"o߾&w����n֛�� u����?�o���6(
.[5HDrN�{����	_�F{khɼ�U�nt���6�K�¦�eՀ�쓸���C۞�z�{�|�kUZ�@�9~/���߿4�W��8�]�l�������v������ ���*���v�e-!�1���z�fLè��}��k-����[o4�\#��Y���V�:侩����i����ū���?��db�v Vy����Oٮ�� �aK�qu3����\\�3���J�+����&x���i H�гo�M |(���˷$�%��(}�� WW_��?�J_�%P��������{>S��BASFy�M�3h$���Y7ԃí��#{"��h��붐ˋ+��?'��B�ͷ���º�d�̉Kנ�B|���7DG��p8��I�r��� ���@�NA�� �ӧ�4���{�W�r?���qPJ���1������k�����Q�-QÍl��i����q?����t�dh0�N�M絈Dz^�wgbFtG�.� �ך���ѻ&�h�U`�7t��<=�^����S�b�c*
��Y�W���,5E|$ؤ��9�n���C�0��̔WO��͒�]���tz�#X��c��1Ļ c�a��C���~a	,H>�wx��})Q��4�6�v�5�+{��d��q%��-A�`���%͔��ī4��Jp��,q1�����x�f�����Jo �5'chm�F���2r�Q+V>���R-�9@)N��P�>�'�e_�:�d�ZA�{�d�?����h�]K̼h�=!J3Q�<+���$g�w�ǥ��a����|�Am��$_� �5^/
�.'M�c)`�a�@SJ��T*
�s�k�/=��(�F�F���8�L������I
!)+x�z=��vI�	��Z1$��An��y��ռC���<�@�*.����
1Z����
��]�pW��e�l�隔=V�3W^��I�q��ρ��J�}(^;�?��Y��g���M;���Ό��g��g�o5�W�>��T���%޳����_��g���=q^A��R��~yKS��%��@�K �T^�~M������B_)g���1�!H�F1~̨A6	�,��֚> *��)i#��c׼�`-�:��0@�Q���� .�h�1Og������0��A6_7	�!Q�V`%��M���!�9��;m	��KX��p)�X/�a{��l,��*l쳩h���I���ǖ�TX~����<9���S�Vg�6�5u��,Cq���k��ْ�b�H�z�Hy��$d��B� �Ms���p����W��|���;��������DR.�= �O܄Γ͠�6�ߡ1ǈ��z���ծ�T�&��y�>yAa@Z�j�R�VD�:��ް��@�2YeK�5h �|h�f0�5�Xr�7�C1�TՕ�����`�˦ǥ�xD������C~1S���'gLJi� ֦�(6A��T�x/͌�� `� w��o���1ܧ��(Zb_	)�{t�1q�U�W>��Z�:.\������hg��W�Y��7��$n0�M�3ǐ<J@} �>����ChA�ٰ�F�Ʊ���b �N���t��)x82в�gŢԜ?�@��8!�K	M�	��·%�76z��y)-]��UR��&ŷ�����	4�����U���PX���
Z�������wOl˥s&�ZyF��/��Q�P�!�Vs83x�}Q������dP��J��j�h�eP^ZS��G����IX�����3��ν��D���e�ڝ���;vy-�t�����d�_*����ش����N�B�=�9m(�vw���K����3+����h�� �*T�[����ڨ��s��/�����,#Oj�� �{�Y�z��';���
�G����읡�]y�^�d�m�Ba�k�TS،���V�}�>�p��"�z �b�.��u?I/:�wa�u����nx2���-�c�N�Tcw���R��H.0�(��`����L�w���CU��͎U��X5��%���b~�}a���9�Ll�f@-�#/0�����kwJO4Ș��*S}g}$�Ypn]�\Qijr{�������M_ `���bp*�W��ĺ-LH���X�iK�݀\�A�:ÄQ�����X ��o�ͭ����7x����d��#z!w�3M ,��e��3�{�N/�i}��\���p)!ȟC�s�h�|T�NӜIv���D��/� ��aI7�u��c�,�U+5+jj�Q�]�I~0�PR����y]��~�y3)EK�3Cog����[��Mo��s�3)��b[?<7�zt�}�$����T;�>��/Xs�(v]	��0�������"7�9̴���܋������/���[SR|`
��:�؇���41[ �5���%�)eë4�rl�\�8��'�<`M���3/5��EFեԞ"��&?���®O��U
��qe��uwsv�	�ˬ�|��4y�s��"�a�x,l�+x�]T�]Z�4�Ai����)*E��h{����s���	���Bt��A]�}?�,q�8�U�z�:��B~y>y�u����N�����%�m��~�h��Q5?���I�3� aX��I��G2�R����Q�����C1����H��G�C� ܳ�C����C�to��D;x��=C��'�hU,l������j�`K(L(:$񦣣��l���%�<�+�8��r�A1��qRQ��;�g��ÿj�6����!��|O�����{�����=m%g�y`7>CO��\�3?������B��{���Ʒ�A��W&��ë���y� 9�3�7�=�>��85'�ck8����$b��58�B�8@��K��=Mg�5�~/���^�e��A����1��X�k�L��4^�B_��.��� �ɯH��L�Z�� 𶡯�Z�b��f�+$$�V�6(����>���"�G <+�'C3 �6\��aZ���b͞|(@�Y��;]TJ<�h��o7@�Iw�,�	�3�0�A�9��|5�H��SF�4� yِ�&�("K2TOh\ޡ8h?=�n/�2m��O;�j���д��R�r�Fb�A���A�s����#���N1�y�f�g����_�F��?��Е^
�vg�C�1r�<u�69����uļ��G;��hq�1����U�95Eχʱmm\��zN����RI�]|Lvf�Zc��a�z�4֥�c><, ���`1O5��ze�&��0��-�*KY����e�
w���Hb����c�%5-�~kE�A�z'�AX&��7E�mIb�d���lx��:_�zt؎�4��%�m�q7U\Yߡ�N<ܐ�,����:%�s0�X������>�Il�����#w(��QL�*�!k���{�i~�\��Jn(�3 �Yě�������V;7a�OS�H��\�吟�:���{���9��=�	�sx������*����]^��1Ǥ�G��V��\*�H0?��EZ�����{����F�YϹ�O�|��L~z�C��~��|��I�9���C"���$��<��|�Tf�Ї����(��י���Eɽk�d���'ī��ɽa����=<�#���+x_�R �g�tk�{��/Uy�D���oϽ�UkՓ��_��H[�H���m��߻^_����Ӷ�Gx=���^J�sN���8�!w�7�9x)p)��63ܓo���{o_s1�!虅�;M�X�R7�\~f0hJ����h��� M��O��?�/�(���7oH���AV��|Y��"2�2��W7�S��NS<���6od�����Jgf�^2|�t	ج��$�{Ғ&(���D��zyzD���b���)\?�i���D��p�WJ��9�4<i�y��q
ɶΙ�����5i��a<e�Ga͇��ގȅ�x���Vr+��+cR������-�{ȡ�})A�LA��M�9M �����Ok����r��)mN�)��Z� ���I���u6Aס�~��ws�(Pܨ6���l�sP�1���CX�	�g_�E�F��g+hω����T�D��P�~�su�Y�I����ʾ//ߞmu�g��J���	uEF��?k4,�E�)P(D�t�G�ZC����"ND. g��x������I����TO��+y���b��������aG#k>�aKѻ'�c�
Fz�`i_�&���/���*����?��g'��ʢ��$(�����%_��Z�����C�UB^�
���V�)fW���-�e(#f���Ɗ�7[q�YecՖv'�V݄:��
�A�����x��ޮ�?�x�6`���B�+�:T
$�4���y��e�z�<����\�~PTU`��V�<&a��2NL�G��yg��J���?8f����[&�S!L��h�PIsv�9�����;z�non�˧�����0$/�?�Q1�k_��R�N��]�|8X(VK�]����\�;���
D���
��j�;1^�1�r �}p5�f���F�����20ʀ,�> ���^1L��]�O [�+����I��סr��u��q��A����P��ߴ�g9Vm���<��d����|{�m�>nC�z�{�������j%	��5�ǋt���
��
���<./T6NvX��2d�����e!�W�1[�|��&�[��ƴ��� �����y���&$���L�l_m�� Ds�� ���G�t��]O:����B�S��WO/6 �~2��NO��o��˗�����T�&Ո0�z���l�<�B=K�Kc��(b:!zS��jj����~x����r���s���x/��ᙧCAs�@ҽA�y�ܴ��kָ�<]�d��*���î��qc�x��Ȓ�S�M��N�|u5��=/ W3��q��l��#�I�g?*|4ߚ�c� �o�<��(V�r�=��Pz�@����Ds����쪌�h���He{�鐣�tS"tǪ@ � �W:@q���Q��'�n`Q"���"��F5�����qҿ»R��:�`�O^v�>OA\��p�3V��2i��Z�y��:�7�`U�ނy=��[���s�F��%�= ��K������@�bu�s�TgP�*��wS��z&o��\����y���۶6k��)�]A�Z��D�aT�Hu��F�a���G�Tݱ1"#;#X��}ُm����:*��Zek]��-�az��?�,E�����=�KK��J��
�Q�xx�/��a�`�롅��w���i��I@����K ������u�����yek2X�$��Un�⺿���~\��{̟ͭ�"|�YRn53�� Ƒ��C׈�s� �P�)��m
H)`�0��b���ptF� ��=Ͻ�A�s��[
�t�nW�U�ec#�@���.��k���>��P�T9�޽fue�s���|��l�No�$�n�={ل�tT�*i�D�h@ݻ]���F�P�׫�k�~}��$�;���N��7̉��]T��BQ����?HgpGs]`�[zJ���UBnV�@��|����1��&􌾰��+
O^'����O�_����'��F��c'��5��#:S����'��G��1�V�����T��E�'N_��C�{�SX�������y���*��~)��'�pj�yB0����q}d�F#6��[�I2
䗟�_}��e�W�W	��1�댊U 0����-�ʳ�g�%����L�N�4��؍ �����A�a��m&^%�=�����c�<T�<f�]�^��Z�JVX��Vr��p�l��& l2ɺ�%�~+N��d�v��H�YEd��t(�,�\1�hƭ�%Ön*�r��;���ƀ��F���H����._��:u�6� ?e�j�����	�گ躝E�M���`�y��r�j�Et�n���uUf�,A�)�z�8�N
���=</롻&���.ͫL�y�g��8l-f�j뜑��
��M�ZWx�����zHe�am�����Ѕ2m���Un�!V��Ayl�ޓU�9-�+y*�S%���h�+�!o1�ec=��s[�geN�-��z�⛰L����KJ6Y�(Ç@R��ŷK���?X��$�C�n$O��+Bp�O�qj��zVQ�د�<�۱�|q��2W�z�`?)��=�,����:?���9%����|�(w�7�+
���[�,�u���6���<�q(a�1)��^ZS�������x�F�k,\7�V��aeߏM�|�_�ާc\#O�*Ͻ�1�}�p�����sT����G�Gr|n���]�E�q�=Y��!^B���	�5hۦ���On��:Uz�(R�*̘+�bɏ�hM�ap:a<��2��;���A9Nwfrv�����F���MD��'�vSe�G����&�\�6����J���K�u*3�j��t�`� �iN�R����:=9��t��f�v���g	��K��^&�ܦs�����1��+x}��!��,4��֜>��+�L��	�+�����!�P`��)� @�� ��ى�{�Z~��'>�{k�φ��jB�0�ގ����"��[w�;=="�C-���Մ)G� ��w���=R4�3�M��k=��j�6��EA\>g���E'�����9|��=gt�C�u�U6��xD#,�b/I��`������-�4WW񗍣�2=+崺9�e��;pj}^�۞��w�=�B;����g�.bѵ�+*GZ��-��;���$%LI�v�i6��%�t	��X%����j�5���`8��Sf��S$�Y/vٌ>�^K	A`I%`C�&y9J�]'%	��B���]_-�H�4G���%�����V:����{d�Uy6����)��]����$���}o����o(�W��z M�C`�3�j�Wo
ïA?]�3�ಷg!�{V�ڼ������skT�U;a��r�k^���P6�&Y�����zuCA�M��kG 4�����!_I��!��0�Y�ɧO L��}��6m�*􆡙�٦5'���D�rE�2�Ͽ|Nc�g�@$��J낭ړ΁6� �b��PXo�W��3(EG�9�%	9�e����0ƴ��z�)�K�O]������� ����_Te�6���[{��Y�o�V��\�7�M\����g��g�~ey���j�����3������?���{���Ɠn4����R,ˁ�� W��x�lz���� 3@�	�W�?<ʗ�o�:VܱW*�x4�#�NшM��{�1�U�y`�����8�����"���i �r$��%�����ҹ�����-��������z�B>�as�9��0�h'=���IxO���f�:��Aj����^�=>��3{	P�swyy���P&z �{�� �"�#��c���c���v��t6��Lk��h�:!8Qq���k�%a�Yĳ^iL��������L�����EEZ[�/�xcY����)s��� m�W��xd+��)��|�����M��H J2�G�o�f.�����Z܄�$��]�4���Ґ��4�0���{�
��aE=S�ӝ�oZ�?�D�d,b���.�W�1�
5&|F���VӋ]ܭ/J0ja�][����\�g��@�?��g	�К��Kt+Jj���ա��7fT�`�yB5�t�V��2!u5e>Ɇ��o�
�W`/�o[������p��s ֭>ŋ�u%傒3�5`�\�Ds�x��<QŃ�sB9(������G�(��/�/��=g�֍�� �C��*�OZ��oG�­��V 1#�t)rTo��z�d����@�d�C�\�@�h�a	N�/�	�G��T!1�__X/<Y�wXZQ�)l١�#0��
���*��yXЂG������2L0������pf��}M2��G'�KU~mse�Ɓ�y]��L�眀W��r�/�x��P�e_�z�����ʶ�[߇����)>����j��j�mV���QJ�u����=���c��m�)}��Y��S����<��n7/�<��@���V�33���v���G�l�+���{ϗ%Γ�;��M#�� �&�L����A84�EżlQJ���A��z�W,�b�z0���	�P����鱼8;�<z�>�j�dNӌc���%��#��w��W��';rpqE ʅ���H=@o�U2�6��'H�͎����ׯ^&��+�&��(��1Ɋ oT�L����{3�g�O��(�s��[���t�G-&�H�7'@�JJ�N`Ŷ��lH��HOf^t�>���t���]7�b��c�{wB�D�֪�j���R�S�1�HI0ߊ�Tp?E/@�b�
&��~QUn��F\���	�Ux��}��<m�f��i��qNU8#�cTG�B�NK���Q��( ��`��������W��l�刘�ite`�zY6�ݕj�
�{�A��2��ǭ�T=`�GOŕ���j	����$*oG��~H#Ik��`��֛!lo�Pͥo�0��8���;����Xw�GkHJ�m�:'��pA���/^+��3��������3�)�+�y��T��>��6'<��66D�����r[�FBB(��s��Wo@�f���fqy�w�(J߁�Z~��?��Ã�$�v����aǎ%�=�#ջw�$6�I��	�������@�m:>ܫ��yu������+��esJ�;�0A��&�PY��ƪR[+�p��5��=,�"��+k�Yz�\�ѹ��h�]���8u�5ĸ���*|��魚UJ��6&�%��>�nhT�? ���=��b�4��￶��s��9��6@��]��L��:�2N���d���׭�S}���9_���ޚ?���=�S/����A�J[��6D��kee7RyaaK�g{o���z���nn��I��]k�Z�\n���F�cN憴E��c���h�<:��^<Ȱ~L�v�	�Xϰ��t�I��;�A������M���Aq�"�z�L����O�J�Wrys�Έ�{~���1}�Wس
&:\ڼ�c��i�;iL	t��� ��9�D$�',�N �W	��t�g����w���Z������r���ڗP�5X���R�9�A��/i@�#2����/$c��� `>#P���ce����k�∛d��ʢGað!|�#��"I6K/D���V�5��c�XQ�S�x#��sV}����D��T���>@��^9>�ʻ+&�bgՑ����
!Z4�}����ňt<����X�W?W�o49���Ob5Ѳ�ݸ	ռz�"��c���G+/�
��"�eg�,V�_a��������<G���ccop���E1�׈�{4��R�P�2䍐'*���u��]�I�����D��
�
+�'Ⱥ@��
�*�����ms��b��<=�#$�.T���ś�	܅��(k�X�'�7�T��)Wm�}��_���-w�V��K��[��r� D�\�V�ʆ�����(�~q�Bک��<�t}���#��� &���+�^L�jgT6b��"�AY��Z��Z�?͏aȔ%G�n������?==d�����<�.���):�(��A�XA���{X��=�c�4TFE�{1�O'*����V�b�������o�=�g�-Og=�����Y5����Ws��=Sa����{~�O�k5Z)k��:۞��ð�_��={��>	e�3^M�c�d�����k���}6�Fb7*��0��2\2���U���C���;��*9hhO������$�^3�,< ]Spx�����`�����]�I��KL�P��x�q.� X&`r����4}�����к��K !��Hm ��c��Q�����8P����X;8%WU$A'��V��(�a>����;l��7L��	��c0c`��:Cf@����������r>n]e�Eh�-}������W���gY�57��3$^�_�:6C�	f����XI�b�,]�����񼟍��*�>���5C�AJ�?�Xk�y]���PAY�{ΕH)�h����3�D�j챜��C���΅`�����V�#U.�F`yun��J�Ƭ)� |��BQ=��/�T+�v+�G��K�s�AB�I3@"�Pz��ɿ+(� <]���6~g��������ߞ*f`�v�R�^ �83$��l#�kK[^��Pࡖ���jh.VYe�>�{�rY�)S�ָ����$n�Ȣ�Л<�M��R����<A9�D"����Uk��t���j�FJ��c�����kY?�������)����cg�؝sf���{��#c�&�wN�jՠ��N�u���c�w�}�4�=	��kϩK���Ga�a����������:� 	pQ�}=�,��;�"����xVj�5�2�bj�V�WE��gáV��CTwk(gf��Vv�wW4�18+`m˸x��۟+�������{L~���=����dR⦱���̼�k<1������j��ݓ�׳���ss��w����ak]��_�r��r�1�Xȱ��޾{'/_����������/_���5A�.R���6�H��g45VT��L���(�zǆ�$� x�� �b� ߼<�#�z�3��c�����oO�����<���{���
��Ym�����#��q�c�O��ۧ=�2�(��{���=n�jz={��*$-�"�$غ��������_������Ԩx��2�k�1^��&�膊q�Ө#L�wL��As[;�c���h������������y��k>X��&�)�4gXcJ�qE�� �<l�ЭD��jE�rn��tt^tp˓�LS;B���^���rGD�����B�n�U�Lñ�H�����
@UN�9����]޸���+V���M1SLd��-��r���p�g�]?����V�%�>��Cƣ���u߲z���H�3g�w��`�TV���T�����R�ߐ����*h�h��_�DO1�-��U�]�t�4�:ǋ��p�W�Ur������x��S �%�^�V�&�h��x������T�j�������Ge���x�B�p�8?<,{G�Ҡ!
ψ��(��m^����(*Q�:�����ᒮa���f�����JR�¦�i�h����'NR�U������R��#`�|:���vQ�>��P��֏��N�_�!���_d6kXR}}���v����	pY,����k}�����(�J�wC���@^ߌ�G���G���{��b�5y��������?{�8��Ûρ�2�m�5���<I��5��$3u����=��r���&����4d/��j��3�J-/�wy<n�͗R��]Q
��U&K]�1꟦���`��������\>~�&�H,��PZ7�Г��@4秵
�����YgyI�n^0�x1 j�]�l'���~y���{�!7La���y���(�͚����Wc_`��z)W�7$`E�áoyn����{��L��!�����) ;�PG�!Z�F6}�X�a��7�����N��n���]=�4渇{�\��QӾ ��YE�2t@���]?o�W��a�����\�_���hN�hU������m��A�y��>����.�[=D�y��r���3�P�SD����2:^+��Z��`�ѰPǢ�]���ݱ#����{}�L�s��|�2�Q=��i
�pP�aΕ�����Qu~:*v�xn,�GDs��d��L�}b�L�����.��e�n���I}�|�*ԥ��J�r�0xr�N��h��ZI2���ƽ�H��eP�¦?�ӭ�*Q�HY�r�\��+%�E�RQ�MoOd����o$�����B|��)�M��XU��[e\����_c��������w�����큒���&�2�P<sYq�u~���hΔ�+���u�A�ﻻ{	���/�kڟ�B��m��Wh��@KUG����*�>��^?��[E�Y7KND[N�:=D����ih\`������%�`�2�R�E���$��p�7>'���=�ź��Fg��	�d:�g��Y����?U/����������j���թ�Զ�����J_��Q�T�Y���]m��4�6�/@���<]��d!�c�2N��X���#��U7f��8
f<{�2o�H�+5]�(݌/��&�E��{g�K970T��V=+���^���t�J����"#���i�n���N�3މD+��
�N�3$xq���iG鼾}�V��� ��<Z.�G#l�%��r�l�wȟ��M�������d�\�r���d�nG�&�=n���v<wx߿��^~~�C�y�,��a�A�,��� (!�i�+po�4um�B!a��}E��%�ꃹ��O2�ŉ�{�Z~�����ö�2���3�ZQٍ�Fv'��|�����˗km�4h���|0Ӂl�<_f��?���*����q�6������Ұe_4�g������5�b
����{�1:X�#;���~�G�O۷�e�t1c
?P��k����S���*#x"n��t�	��;͜��B���̨��C*���v8ɇ����ؘ�q��\�,���\H�)a
��/��I��2��B�N~�=������
<�P3�&�h.��f6��tmeܥ��d`)���&
e!�ߧ�n��t`��!�^٦5ǂ�L�MR��-@MQ�Vz.�w:p��#+!�_���m���^�ɹ��Y���]����fu &R7H>�J�<U-վp��D�7�w�Ha;��$F�X�����m$�(1.��������%���w?���	C��_�2���Ǐ.˳���N�'��e��ʜ����)C�h7f���]�F��銴<����~��g-*R�m0�է-�$��4�R�>�
�*�*��WJ6L�7V��W�sυ���c�\�ƕ�ޙ�-�H܋X���Aa����KN�S������2�G�תa����{������󺗮�;E>z���4<2��J��Y�I�x�@ �w�0[���=�t�A�8F���P�NmT�Y�V��!,t+R�����)Ð�=E%w��%;�e��A���J.�� �����۟���s�����D6ٰt.����ՎH�?;9N��*^6��:)�j��C0Ȁ$�5CoJ���>�r����>r���h����O����y�����j��t$����p��)N���zD�(����6V��av(@Jc�a�����k�|�R���KmA2�5;�p���;(Q7��{�P�ch؁���,RЪ�З�/���;5��O��+�|��=�>��X�Y�E����x<�wx*A��d�jO2���T1�Uo��s��u� �mX,z	��[16���M����UT��T��Э�J�8
�
��`@��P�[9`��m����=^�=u����*��-�B7��`�	���筏<�}{�7��.��uS�I)�K+Fc.3��H4X�ٸked���!R�J�r�zE{Br8}��o)D�>�T�.�����������աj�q�k��m� �5j�
�v�B�s��[�^�% ��NO�����~�iAt��ZM`vpp"�ۿț��e>`����D揲����ĭV`1��&�v&�ɢ~����ߙE3PP���h	v�$(������ ���ʻF��%���3J�����M���<!�X�Q�I��X�����>S�W�W�9�4��p;�؈�����`�G��U��!�g��+���(��d�� !�䠆�˛���Z Z=GꙓѸ5�Cå�~���k��I�����C�.�
in��!��`v6-�`z)��iL�{%o�jzCc�&X	����6�BDr�z�!����+�͸ǹh:P�\��k�^����=�����T�/|�]��n�sT�8^�h����/>|����V޳Q�>�mr=���ET��P�������w�p�@Y������҉m~��F��M���gޒ�?�C���F��<v�B�ުJ�D^̑ D�)7�\('C��F����� �\�L��'@t�@@���.����)�ސ�s�yrys'_..�a�.���SBJ�ʌ~��eN�`�s�d�ie#��S��P�Q���D�j;��-���~�ߺ�:K)^���:�>��'�����-�h@Q���8li�uV�Z%z��,1�H�|��*C,��@�d,�����2N�b�>1O���}�$v�V��6cȳ��t]@pU@�Ye�k�%
M�)�5RM�tF~�(�1����=,^D7�P�ﭢV�@Z���4��<^œ/��#%�ڽݚ�5n���7@���hI�y������o���Åt���r�Q�p�BX�k�9}�����Mcd�Vͤi�VѴ�)�ku���54F�i˦��V��Ą�P������d��xi��3K lg� }�zX���Ra����r7���uXӢĲw]IB��Nw/V����P�%�{k��Л�C�&�*��z�r�n��k��&��J���"�c�5)�N2 p� �=i�T���\�2��jkj�1���*Py��{�艖��kxh.0?P��+Ʀ<����q�x8We`!>�~����Y�{�|6�M.=���7Me�pl#n����EG4D�A$C���Y��
&��f���?�e�ͦ,���'Ŭ�,?_As�l�Pd��5��z�+��Bv�[�ٍ�șg�c�-����I�
�����%2��=��X�߰p��No}e	�M�}i����F��Q��W���`�V�$o����k埕z.1]F��ͻ�s�<�0�qM�<kIϡ�C�yC)�����Ez�N����婼89���=~�
<�$�E�㊼j���ie�|`!�`�P��Zb���!�51��9?�k�x@�m�<��m�\~��QT�\�{���K�6G��|)�I�ZP�I������B���m�a!&C�~t���E�,���8�:*���Ib쏊����^�2�XXKQYi��0}[Vu��~�AX�W��'L�U%��a��`��@8�ٍ�j�4�ᐘm�E�����r,b��ƺ[��l��ak�M?a{&�s���G-�`I�z�4'I��Ѽ�������py�� i�Ϗ�ϓ[����UgR=\�!z��Y��b�MX~�Fߜw� FGh�c�Ѳr��+�S�����nN�@O�r�`%�����Z�MY�I�y�m��s ��!�2q��Gr��BVm�������s������+���B�O�p����V�sbv	�@<�LĢ^ԜI-�I�k�P�H�X�$D�Ǹ�zM�0�4f5+0�y6@ ���!5�F�§��VV�5���yؔ�� <hK#���J:09��j!s�"o�=��~�c�{���r!�r���P��*�>�5C�Z�Xr��̽�����=]��V^��\0q�����uV�[~d�m"%Ͱ#���Y�4&ơT�>�>iv1�#�W����'G��)]�)�Lc���h��y�^%��I[�3݀�KL�t�錡��b��M.�WԒo�S��c�i`z�)�(Z��M ����fU���/��\/�;�m�U����6�;Y���Yb���l��,j��6ކ.C^�nz�u�6^��Z>�p0��8�&���s�]��54W�h���_R2��0�9`��gTo��G�^L%�M$d٨��Ak�y꥟�[���A�ʄ��d�8��D�\�{#�m����pW���?�(~ 
&]޳X���T��;��g���+٬�.E�M����P��1�fWpb������T@I.�olq�V��s�}�c� �(�1�)���^7>��Md�v�${kC�5n�(�}=�>s��|2���Ɣ{Y�u/�0s��Xܡ�Ij�(�a�vY\�*���5�3�
I��^�&�2�]�%',�h�&�^�Ȳ����6�P�*1�QU��{��7�VȐ�}N��y@֣�8p�YZ��,1�y���5Z���E�}i�)#�D]��"��\���[�T��r�'u�$ؓ�Ԟ�"���0��*C� �*q3�&.�;�<�&[��#��� ذ�E�i�Lɧ���j�|�j�蘄�Kj�ɣ�a陯�>i��@`а��������M�$��$���z�ꕼy�ZNO�)����_�@0�I���>���������,T�����$<[�=(~�$`���0ѥm��+�����r��t�6����rn�	q�N,��A����;%�$)��k�dp���ϗb�ګ&�y�$��`	�qL$f.���@��t@�}m�;1q��y�치H>d��6�V�����U�7��ek���8����.}p�GЖLTT[����Q$�P��+~s�s�RGA_���Y���:���M4�F�֔�1� �����a�|�t��?>2%`�8Wn����\�f�ëI[�b� ��(S������wv��y^e��!�"�
�VFN�4c̃˶�o��}3lH���~��U�QN��LєGH����{r_!�t7k��z�=����ߍ������8_��T�(�v���8?=ؓ�g���Չ�{q�-�xe�y��m���7C^+��^s_��&Q�L��[Wc�5�wf�������h*�`!L�חq���Ɉ�)N���ۼ=�|w���i)���+`�J&�-G��'�8��Ve6��y,�h��9d0��g��B�{0�\U�U�g������b]�!͊'OY0>� %?�]���8�u�y��\�P�q�r-0�yf�ߕ���KE�^��!G-���sV8��	�b����pBM���r�ɮ~^�+��N�ɏ���JNMFV˼�+����ry��qd���,q֒Gs�RTX���%{ot&�h �ah���!�F���1PJA��i4���I��`P�3��.�7�F�X���g��L���^n��X�aL������ƿڐw�������S��������ݏ?Ȼwo����{j���k��Ġ�@t� O�X%"����i�9^'��KT�Ů�o�Sqn�s�rU�*i^�-�@��j3�!�cߣ�%9���B*��܄�J�8�B�'@��TLvF�K#"
>��Ri�s������\���:G5|JN�QD�c�+[�@J���)Ʉ�XfQ���Aif8.+�)���5��
ـPS2�~
&��[�j��9(�aT0��e��c0�9<����k9-@>��\G�O�Ǥ���Uo�H�fd4.w�5n S����;j쨛�D99��kϊV��a0� �\^I��nV�E��{�M�jH�1qqp�^�MzrL^�L������oߴ�u:��ֻ|��g��#��Oq����h*�c�w�{K���
���&�c}����1�:���@�ٮ���nJa�
�V��|����kAe =+Ea�V��T��m{������5e��	��p��ڟ�W�# :�\_]���u���$��,���5��d�1��х`�@޽~)�߽�ÝV�� ��i�Y��	+�y��Z���i��?�N�"�eԾ���g�J*�������[�j�3x7���h<�pL�=J��y7�\lk�F�:V�}�%�Ԍ�+s�6���y`�k�K<4��5}�F�-TƓ}u��9���Q��������lѹ�/�XLzL:G)��6T��Y��'��ddn��Q�k�?��*K�d�����P�nd�fL2���g�4���;4/�B�6��Ѳi�&�ޣK�9�.�'�V��9=%V��M����"]�a�M���6�?��Kx"F���o���	��Ğ_���kĲ���Y�G��lm%��4���jXw��h,)���Kځe�p-O[mrMbDsRxՕz�Txn ���!y�d*'gQ~�?���!��eB_//� ��G���2�k������ʦe���T^�~%?��.})���g/�Xa�Nc���'�3Gsճ��~�W�8��z��vX�$�;X��p�;�vt����WO��연�wzS�*sM��0X~�����[]9�G\o��}�A�nR�C'*�},O"v�ۛI9_�Ϋ�g���q�HYH)�9�nU�t6�D��4������b);����Z) �K���dP��f��p�q���=����YNg��i]6�--�<����q��旄M� (��S�&@�V+��x��.A|P�p(D�e��x�����V4���$��D���:�����a���F�E�) QVɈ]<���{x��ŷo�� �Ջ���#s�H[F���f������u2ή�6�f���}�!U�Z=S��2s���+A�@&���_>'�5�p�<�Hys}u��w!˃��'f���s��%��Ț�-��
 ,�̜?h�cn��zm;�����U�{/O�>hQ!��|�'�1����L[yyz̾������B�T��zű"��*�Nʘ!(����2����\��P�8�� T`'�{�d`�URݼW��)>&)�V}�P%A��-]�`F�;/�h&��[H��0���qvpe�i�;1����4��y���<oœ�g9o�0�P��ṔDN#�����1��.K�ʩ�]��=|�����0]p�)SX�P&(j᩸���*D���ZBnK��H����+�@	����jU�M;a�COK~l��������}�=�\��������QF������T?T8�ѵih����j��k38�Z�t�{�zK�A����5-n�̬e�		���Ps24�ؙ���)�b5�b���t�n<KBc�`O����9w�I�_^ȧ/��ׇ�r�����k%2�f�)|N��o��M������~L����D�%*� �}�I�]]��y�{�?a�)+�����I���dQv���v��
ógX�i$��F�g!�\�#������"�*Bg��J�jv�ɢ	�ҵ������$W��赵�x[�'��AK��Y��Z�?3�Z�9fm�g(4��ܛ�S=�����d(_��>s�S�恅�bi�m�_�F��"�3�w4aȾ�R�,x�+��HV��{�TB��Q�L��MmW�8+o��K�{˳�yh�yJ��2��T�K<��Ӕ��E��'���x�K�<��s�A)��8����̀א`�T��;Sz$<G�x�u���9P Ž�3m!�v��Ū�'*����]>\�EV�S�C���OS �4nn[.�2�߱@���EN�ښlhH�
���8�����R�6�1h�����~���h�9>��G�s���S&���G��kK��dMm�	 -pƓ�����!175��3^;�P'�)� ��������MQp �EHm^T�>@�]\&��*�9����͞={�� ������[y����G��l�|�k��W�(S�&�(G�Qlf�m�@� /+��^`�w�@�+��3�����C�y��R�z��H���8 �Ғ�=���zJAot&%�l�S��ט�L�p�z�U^kx�ɞq^���Ļs�j��E߁^ ���9�0�:hJylK$F�5�6m�0'�rSjt+�Ale e�w%���=��r/ƌ�j@�=r�G��y臲��$���K.�l���������汁���͗��{�Y���T��j�;A٬�IА��0��3C�t_�'�[D��8�-�=H����6H9ɻX0ި������<�,U��n�X3�M�ɉ�jBn�a�����9x�����ق �Y3E*D�n����%�	��=��q4�]���͗r}7���G�?L�xo�����=
1�o�Z�����T���G���L���SZ���S����&������k
�������������鳜���˅��T>�j�i�`�<�t�P��������B0_�%�GS��w��[7]Z?��j$%
�&4-���s��Vc$HI�7a(!4���ڃ��ޔ�m�� U��l��yj�n(�<]A?7�UiB�=Xjd��ˮA@���ks����h�TLL��
]F�Ћ��L��90�3O��Y�X�D�W߬�7v�P�'�½	N�m��)b��7��kēxk��z�ۋ;T�ڬ.A��Cm���A�5N%���/&ֶK�h"�Z��˫;u��
Q�je�s��5�J�k�	�@���OF���9�VD��	xO右��0�M`g��vyu�<P�#=s�TV7�?�ۤk�ޯ-�Jv
����F.w�I�/8�f�S��\� �A. ��^���%ǽb�S&"J-0(�A��w�;K�$��q�p⥀���nG��h2��@=��ZiMI.���i,����n�+�
��ӓy��$��Y����5��h����.ɸ�܌Ð�Oh+'J��������k4N��t{l��h��w��N��R8����X�zky,�Az% o4�X�W͜'���,E���H�!���
I��Ï^q���F�p��$�EԱs����eԐ$��X",�"B\��Zk%A������ ���4��^)(��c��1�ͩ+~�xCY����Zt�/�;��e����a�His$�D��EN��W�xHr��<M��}+w{����� ��ĕ,�|�ך+=(kqwC~|\�� ����\B��ki^�W���ş����6s�m��<�C�t��2�:	_�2Q%ɜ�^[K0G����Wj�l* �^"�a#��3y����`����X�Zq���|�6�ͽL���{��s�ӻW���5�/ �ݗ/����?�:G�p�K9u �w���}$ǧ'܏d/FNG�ߒ@��O�;���"��	�E�t5{���h9��֖��k)؝(�O ��<"����I�B|���}{U���b�����coC2tg�`ʓ��=@�R��8���q_�n���5��[<�~u�$6��| R�tY�{h�T��!�܆��5��q�!̴)��/��^�H�N�=1	1	 ��dF����ߌ�`�[��x���* �3�}����z��"fc��)��U����\��G�9@���
@V�C~���VO5�`�qc=��,/XOG^�l���|l��^�N�s��f��� �;��5���on������2&ϲ��;�B����TL��Wӓ����R`]�)�o B�(��j[4�+�:PPdzS= ����k��kcF��/�
WΒ+@[����� �{�'虰�����x�=�	!��;�za_���W��)���+�=����I�q��{��]z��{��L���u�͔|:��Z�OR�0�<Q�_V�n(���cQ�M]ogОЭ�C��t�k�i�"�Twv�r|r(GWI>>�˰\���W�
�h@��1��ֆ�愷AF�ϟQ����M�q�5!G��ў2���G=��Ωv6D��R^n�6Ve_�ju���� ֍���a	�\��Z&L�� �XM@���Z��
%�n��cR���߫y��G	�*�:ugz?&?fZJ��?����@��ٚ%�2�'K�/	�i
���q���G�5;hS�ߵ:J-i��ѭN�⋫ ��t���$I���$X���U�{v��������;�w�ⰻ3�ӤXr���TDUͣjqٓ�UY�N�MEEEE�߼<�.;VP�p��M�V���Z�D��M�;jd�� l�ʽ�r�Z�mW�E�v���ʑII�o�<�:�,�2Ec��Ec�dXh-��_��}SB��Kfo_9.��ɰ_��V�O���9L��e���7hk�-2���m+^K ���{�t~+w�O
�:��Y*�KN��M\�Y2�Jt��e7���"���7c?<�-�����O<�G�Pa2�ǧs�����p݋�{��p�gd̻�k�g["0�A|��V��y,t�^�)�\�5I��Y��]c�R�6���f�a��������ܡ�:�k�d:���Bȋ2�#��V��й��ݙ�;�ks#�s��y�͚�����n+ �^
s� ��i��63m�ob8o��ã�!���+`?:�E/S98������<:B �l	�;cL�Q����{65}���	x�����G2�������˰�O?����!�@1#L0$k�|�u��Y�������}E���inڶfW��da�w�5yt.�1��9Fʹ2���X���x��~Wz.k|8��8�Y����c�8�R+��nK\�h��!�� L�YJr�]JmCm�{!�.ɲ'���%���pz�Y:��ϣw�R��x��t4b�] yQ����9�U�鯶�7�b�B�2���h��mO�R-�V�f�?^��R�F ���;&a;A�-?MJ�Dv��Rz��Ľ���@a�;����-`�{��y��[:՝�>ޘ� K�[�/MՃ�z/�6ƁgZ�ß���#(�/�<b���AU�B3�4�N(L��H�$+��I�e7�צ��	ɳ<��1� ��y!q�M�^��l�A�|�X`6-����gdVb�K^��(�ɂ�N�@�*��
�uB��ӎ&�|�+���I������P9;qBK�<��l��dM�lD���|�	=���֐�찋��4�W*���n��U.�k��k�����{eg���'��(����'g��ڬ ����
�Qov��x��	���Sl���C�<5>�  ��IDAT��̓�5�Mr<����������87����՚/5����u&�//2�j��J����U�j�7��z�k�v��տ�Ŭ.�͸i�ō�5�� @�Qr�T�U�S�X�n�dG*��nͮA�[����<oit���Leo��&�tb|�
z>}��ϗ��P�M�Vo6��{�w�B�!�vL�f�� 5������&LPMkƌK���4�Xb��Hr˵f����Q��|!.��) H�;��E���VVڰ�yc�D@�ǎ�����H�������`_Ξ��tˀ�kg�i;%�J��M��t�]ҟ���5D�����iY��f3L8���������r}s-��M��ښ����ܑIH�7��P�������8�����W�7d?��X�X.��_{;5��>
���&Ԓ�)���K��noo�/�E.ί�E
�4%6;d�ɞ�9�ƂC�����8��󹜟��Bz�/ ���K]'(;���[7�Dy�c>�t��O@з`#^��<��&���G��ּ��������;���?�!����uy/O�,5�7ȝދպ+�Xf /_�c�{����A� u�`��R�@�R�t�n}.�=��7L3����X޾}�ǱW�i�\_^���h�����P2 *u��� f����������<N���]�	��ĲE �;�����0�k���G��7�/S�Gx>[�i���`|Xx�U\��S����|$�����z/���v@�����b�W��X,Z$�O����_�c�W$�`��b�$m��(<��(R���!M��-a����rx0��lޑ�X�A
��W˺��k�fو0�+ �~H�yr�k��	��	��^�����H��1倌+n��<��(/z�aRF��A�L�c�Іb!go�d�ݴ�G�X��-wd��V�ܮtM�rv���$�S�jH�no���lW�׭lN0��'�Du'�R�d쬹V��5�%�d'nh�J�����-O���+ӝ����_�]��q�����'��0���f�	�<��C��AJ7����U�	|�%���T�q��y!��\���.6����f;�{�
�z�/D��KC)��	������FL��e��S���H'DR�-�ҫ����&�`M@w+]�+8��0Q��	j�P�C1s�� ��eS�:$����;DC�&�F3R�h���l�Κ��6�G2]��x�a(��vK�7T;�~6�5H~�x����b{i��,� \����eC�^��ʦ���_�=��y�(���S��kj���`����v�`�Z�f���(t+�C��jmX���K�`Q� �

�k�Lx�b��{_��o��aI�*_�~0�v�6=�D	+���Xe �j&
����Y�����߾{K�����脌J]oe[h�Sp���ݜW��rO��`���K�&�g
�޼z#�޾�I�z|LL�r)}�~k�F�Y�Km�'��?��ى|��@���eɲ���ug�g̼��+O���[j� �&���Vuyy#w���:3���H3�����υ��>S���)�kh�a�I09 o}�{��s1��=��F� �l�[+��5�<(W� HR+��&0�"Vtp.ϟ��o��V�4��\�絞õ�����`��ѻ�#�qK��f�u@�z��^�~G��%�cclg��2%+�Nt#o�* {����X
�[��4�k�]�gz������LHZ�q�.����m��9*����~�^����850h0ۺ�LW�w�e�%��"!� �je���a��lt~�>	?���^|�O�=��5<S]�e�-�L'�1��յ�q�,W����bE1 �*�A@��B^������K�V.M�U�e+����^tw��cA)�$�Cʴ}����ұ��l�'� �xa��%�Y�T�d�Nk������X�fsԳa ��X$L吭Y��`״n77s�~��7�gq��*�UW���8c�,��;�*�]���SB���}=��s���S�� �1M�~7llʘ<B/ŎR}2 �L�y�|O^�|.�������>$��������,�ƸUב�a�+;��\Ia�Tr��rQ��� ���D�VDɪP��8۠�z?�4a[鳥�j�sk���ʿ�I�o��<.�<>�ƍ �;�	���Q�-A7:�:��=ndO��F��mHQa��\��.�-�P\�rr* ����Pm�SK�2���8`V�Z�|`j��j��y�O){&'���0 �S��`׵�k����B���k��e�6{�2� �V1��D3��l�� Jf�#s<\����KnΗƮ/JC��:���k���ڭX���ڃӗ�6�9��&:��پ
�e�C�b�^_=��\Ϲ��>)�z�{�>) zx�u�����lRVYc�v;ȡ�~��Ka�b3xxT�r� �F���7߼����Ba����,�}�����p}�@I�#غ��frۭ��x�A#��5��pCm���[���r�MI�ں��w�䧟��/�+�{$�&��ټ@�>!�8p ���]���}�^>|:��,���%�i��=���C{7���l��-�g06`��ϦmfdZ����X�ر>�r1�����U01]m���DA��yrz*�}��<h��Y1���b~��ݱ$KMOgY5x[1������1Kn(�b�����P���|�F�,Wg/����OIf�H��ƺ8a�r,�*|���b�����9h�Pd0A�ł�c�T�j&� �`,=�t,F�uy&��q���+c�����*��7J�&1Q�!+xx|$/_��cج\_��[ǁ��c0���^���3y�浂�c�ꚸS<��k��|��=�E���6�=��ٞ>�{�o�>�KF�j��=���~9�Q�d'K��H��\���1��?���%K�t�I��������}�z���A�{�}�4����:����|��	��xZmɩic|^���ַc̀��;o��}��w��v?�C���k��O�Gݰ��d��&�7`̍B�ež�8I�;{{s2�?���Ĥ =�����h����{X�xN�Nr:�Y���^�D����O��`�M6��{�7#�޺�[��#J����zl77�,�_��խ=�ٯ9�HU��Qdl�!���X1�������<��T�!���O�g�%$Q�2�}�7g򧟿�����p���~�or{�!	�����V��Dǚٲ�yc���{�~ǭ�\�5��#�4���A��,A�`R�SPT�ZY- �x����'W�Q\S�κbT������G��p�M�JFqjh�h�M111j�i�J3��]e�U��"(�j���a��?fA�J8ţ������2�� ]dIQ�K�P�ciRvк�1�cƿ�YI
����-X%�=��P�R�GбM J�v,��C�E �����������?CoZ���E�f��6�������ت,,��v��Yq\�l�#��\q��|�Wݖ��{m�o+�u>7M�nr��RC�dz��ةÌ~�P��@��*�K˝�݈0r%�����ݝ��;���Qn./4�SP1�G�FO4��ꃉ+~�����7dd�d:�;���a���b��s��e�.��}"p���y�V�2$��p�p��o���~%�ִi�FS�gg��Ἷv�ol�a�9�} ��fPfv�X�58��r8b�koal͋�/�� ��������z;J=����]�`�1^	�����}9��;{vf������=Jw;y��˞}��SY��X����/������ȱ\nȮ���hƭA*��-�m�1�@� ~� �M������#?���u��0^(�G�!���5:���C�iH��Scc]wC��:������C�rPf��Q+ۀ3HF��4�g��L޼{�NAݬ����3�`mK��}t�hBº��'Lex�� ��pOs�AvJf���/���͝�hįj�����t-/������d��!3 ����=��X�3}{���!���lވg;I��͟k�b`�i��/�"�6A��8 C��=�'
q����em{���s��k�w�c}��П.�&S'�=!����Ru�V�4e�8��l+��A�<u�̛Cҗ ̌����5����G�U�֪_Dqe�aLj�ر�{����=^�3�+������ T`���u���N�I��d �Y��A+^���#�[Zx�d>A�f�{sG)R�S��`���\⾽]�s�d�i��������!�Y��Ef�+y�_�f��[��aMl"��4L���s[Q�>�:9>����}]?{d��qw���������єB;��G���_��o��i�#d4������X��	�ѓRfF���	\�ÛCMkͨ�> �u�.ڤ�}�&6v�hl���ҹ�$�^V��n,}��܉G�9�IU�������nY�TKX]YP�O���[~J�؍Ðg|��FU��gq���EX�/��Nçmٜ�j�Ggݨ��Q�{�d�}ڰS���k���3��Aw�y8��2�r���y�1^�h����Y��!l�� �^����S�CW���ϸ���k��:��[��_�� 2ԽT�Q:ﱕ����`дq��6����g�U��Aq�(7�=�5|�6~0�څ�(�L l_�I�p{%��7�˯����� ���̝~��� a���	s�5��2Aϲ�`��i��xF��aԡY�6q�P��:x�e,��6oa���ty�@b��y��b+�/ �$�_��s���|bz�<�skJ>�ج;j�,"�L�=D7 ����ə�Wo���9 �k cs�_{���"�� ��TP.���5��*�9�~�S��͛7�׿�M��������[R�G��p'7�hn��=2i {�3+f���ѕ|�t�uR<V\M��Z4�A�P
C� �������7�0fw����澧 ���'G�\��:�y��ugz>}���G�@�1��d9���(��� ��ΎY��/�����7���������������~�����F��?}b�s�����Z~�uyys�ϒ�k+��y��J�[�~�A����N^�|�@p�ǵ����6���Of�r�@��gq�o��޴С��!7�r���fT˦ ئh21��,�兦�2|���G��uGc��	��r=P�9j�S?&�5��Z@űA'�{^sڅYB�wl��� Dw�$�>���S�����O���~Rn0ͮr�qqCG�����Ne�C&�q���NDh�֜[;�MP��9��`v*�moE�����X�!.hŕ�ɳ��*�/�H��5��Z���c�#��ފ}�ݜ�g������������`�	��f��3��2��l1i� ����(�g2���)��d���H���l?�!�O0� �
�D�E�uQ+�҈�τϬߓ�b��>��4 �Z[�"fIU%�z����bJ���"{�46G҅��.��ߟ��TU�������4�M;����'�={�M�m�#���<�U,c�:�Y aev�]�܃.���ȩƒ�w��fKva�Pz_0�?�l>
���6��z��IE�W	���n "y���b
��[a� �e0E�5L��nlXkb9
Ae�������X���s�0q�#K�5G�<��M�aBi�e��� ���6��b�b�2-3i\x�m�ٱDp9(��<D��B#gdGԯX���:.gˠ��͒%��X'���ez˃������O+�A�d�qV4�?TTLs�Z����[�#fZ˼����d6[ ��OĢ��E�6(�zK�N��%?�L��"���Q�كM�����D�A����4^J� �tK�)��� �@<�]2� `�2e�>������tq��)2�9��K�`���F�۴�[2Zߞs�G� D�OhXo9�Y�U$�%�L� ��zb�I`V�N���{��o�a܉w%-t5�
6�qc�n���C=�c>W���Y7��v7�is�X�{�
��\��@0H�eƞ�M�'�ON�ڿw���Ɔ��Tc ���G�qN4@H����Ãz��2+4J�8_<G����o��N��L��\K�����i�!}IQ��=P��?�g�>�+��>��z�[d蝕��AK��k���[��1��9���/_�" �z]�K���x�� ��q���m��Y���ǖ�-X>4,� ��x,9�a+hhy;��\�'t&c��vC�����������5�����?���5A�;�(����?��~���O��/	�&�j�z���p���^�����r F�#��'z�%��ڝ�%�������%:�����ݓLl�}6�(�;���K�-��0|����eȻY�l�#�K�H�6������bp[��6H^s�0���c��ޅ�%��dܭ����@���
{��2����P$�}71F
@�I0��0�Y�/�����.�%��;_+k�X"I�_����|8�fcT?X��boT�%Sr��# O��� ��Y��e����䊀��t�Ը=mt�BG��T�kRt��ɄR��)��|R˻7/��n��x�n�Tgj�Ѐ��ώ�4��(4I�3�q�7 �N/f=�n#`c��m�2�d���f��$��ny]P�t>%6�t��,��>Q��I�E&�{&��b��c����L׀(AD�rp��sT�KK��-�dUV���
��6.A�� nRvz8�rdCKrL�YG{˴D�M&{'�S�~x|��oМ�s8�M����?�O?|��`���d0��[^�������r6����dKgݓ��m�[k�X�_�y*ZL�!Ji�f.J���j)���
����]^�S���f�Mj�#W��j���&\�|��;1��l��Y��t{��M&v28�Pۆ���l�\7�)�WېJ�w��9�}A��Bd�4S��@�BX����*���bk�������O�xKi�� ����y��>7w���sK��#I-D�(M�uc���h��jDR��XW��n�43=���=��}fa�r7=���MC���|��I�����k�.�Q�6Y��U��� ](�`���(�������v��������C����ke�T��,hD �����M�k���	�щ7��_خ'����1Q��{���3�������o���H��ٶ���=#���_%3�����d�v(�-;�cDR�P�eD�.@Z7,�lغ���3u��1upl6� k�ݷ�ʥ�t��c�,J��'��3�1����}���o�6���IL;W�1A� ������M0��S}��f��L0-�6�O��������P�M&�d�G!~��H^&�g:�Ƌ�$����[�ȅa�20��W��÷,�n���^M   f���{M�ݝ��".�>�� ��
W�x)����� ���"����Ç��?���,1	m'��m��SwH�����Ʊ���i}�.< 0���o�5A���g���_�Ң+�C��%����U|�>~�(�>~"p[� ��Vڢ,�C����)��monx=fO�9�s�6��a9��R�r�y}���I%(Xш'�Y��V��R���=R�/ ��L� �4�|M4V���D�p_^�>�5�|��zGaX��uE�����߳������ P� k���b�9�4�uqo[7:7���mx��Q�}�[�YI1�79Pcldk��v<x���ִ߸��98���1��:)����S�x��9�o ̶�Q�C��
��G�Ƃ�&,��AF�kȮ_��pK
���S�����	��e�{�t&�e��<5��\kP�g쮨�X� ��1ddAj+_�p�1"�P,0�oأ޴���cc!���K �tq|����f���C���2b�at��9ű��nK0�׋o�@���|���Ŵa�y[m�:,��'z.�@���}&M�*w�6W��&���8�wX��Vv-6�k6l0DS2n
�^Ǻ�g�ـ��x����l�dD݌���4����k�d?�ǢધC�����A�U�>D6��E�2lZH��k�+��Y<v0V�C\����lI���6)�<k-�كf��w�uy�����+��-��dڒP���m{��]\^˧�+�ίu�\o�Zrʮ����6��"��_$d|�n��|A�j"�ΌI�� �Y���؄���7�i����a�9 [�'n|���65�ay\.e>o=Ӵ�n�'��gc�Ul����t��ap���5r�1ѵ{qa�� ,3ˉ[��@�l�o�ȥ��j6�/��5�Nٔ*!=�R�0X��y��'s�fY�)@�b�7Şg�a9c���x�m��\?.um�sO- ?F�5S~V�i|�f྅�⇏��Cp�<���d��,E�1�2_�5��9l��ܚ&
�v�4� 6���}�?`�%�NH�z���-l"�P4Z"e�0ضI_{?h�Z����^˕X&�=��������d[���H�Ͳ���1|E@�1@W���{����*���~d��A���2x7�=�t���U����o?~( ��*�z��bq=#�~���� �Ei赆� �x��r����6W�+���������	�{ހ���.魒 
����z_������ޘ�����!��ǹ�m�=�Y �Ã���<d���&`W�|���d�?���o0K����R���O�Y;�Z��X%t�w��$$]�)��+M|Z9ܟʑ��ӣcyvr&�_�$��u��T�}�����F4� A���OL�)Ǘ�l�涔$�M&n`풝(5�%��^�2���S /4\���4���Ʋ��v�����އ�.PKǃ��[�2�ޔA�O��p��?����3�uZ)WU4I�y�`AE�3ѬO0��鶪ʂƆ�l�cz�6̜�L���<h�C@�W�dOq��}���9` b`�rmT;�RK�8�q���L�z�T���<ɫg��w����3Z!��z�˛;��_���!>XJi���� �#��rؤ�=���7���+9�l�16WflU\�A3���w͊�AƵ��D����A��7�f;X���1l^��g�],tWrx|*'�^��W�ҫ�o��W�m!�F�`�Y�����`<2��;�j�F�I�u�a�n������v�V�&���@r���qO��Yn��`�ez�����3vB6����+46���C�`Q�D��s����ܻn�[Փ�!���i�\S`E��y���)hs���~#���|b2p����{�T�r?�b����'K������&98M�ڌk����A��,��_]2#�2�к�7�̨s���2j&��	s5����R��nT�;��\�5^����Q���oN�gN�9�ݢ?��]���ʃ7������_+г�>��x/��w�_�5ŬOf�ؓ*c���J��Kf��
Z-�5wy$��D��ۯ�sO�u ����]hΰwX��ේ4�hp����>r.h�2��H�Z�k�#�|?}��g� �6��+ �}v>��`	��� ��y�i�<A�6c
�	��=N|�#���K�Ϛ�a�ahsk�ɞ.HD��c�0�gi#��q��{r�qgrr�����9�Q�T,M"�c��t���DR� �e(n�BkvòC�����G�s������0����Wv)��&��a���,%<�ue��HV�p�k�q���qW!��ѣ* �:�k<+ �̙%P ��n���������1�����<y3���=�t�R؉0�ŷ������i0y��O�"��r׽  �����ޯ6�K��X�����TILN����%��?c�.i{]G� �6��2Y`�*�5x�jot�H�l ���{� ���� )�a��j���\޽y.�^�h<=���#�t0}��b}��r]���7���)�r��
��qn��q�XStsd\�+_��(�Y���w�Xk�Y�}�M�щ��-:e���|���6�����Fhz��k]rFg���3�k� �MP�,�c;����4��\�ML�.;���|Yj?��������Jc7F�y�	���v�B ���:���=<�����𑵁	�~C��43τ�Z��a��n����2��� �.�E��z.�z�_��ɟ�%߿{!����Z�u����gE��_���Kf ���Q�@���{A-5pl5�A�7.֓��Svʠ���w(�fSJ�ذo������~'�O�ʍ?�^���ۭ��e#�5\�M�:���P�dj��#�?|&��P��z��^iS�������e3&h���)(�(���1���nZ�@���tRi@��!86���5Z�ϵ���ɡ3E��.�Z�����;S�%��Щ�e�ǩ�c�u�z�X��y0]�,�����1'�ˈ(�l�!��~^�s��Cc��~��}��f���`�1�ޓ�@~� �\�΂k��̒��Z��p����?a���+zO+s��5���«��CS��<,��b|����S�"ig�be :��F_�V�����`��,���趃�������?��q~	`a�|����*��d�v=Jp �XI��<���|�ߛ�*e�.�TU[�i4�P� gu�L��$��fzwc������ꆆ�(���YC&/b�Ko�1���I
�!_C��g_Wr	�[i�{��G$��e�g��k&+
¡�B�`{#t^���M�U��K���Eo�0<�P),9�6�1���Fw`��vUv F��D���O 0��� ����_�J�3��އsk�<c�o�7�A���rQ������WIe.o%�H>�6����,{�H��\$$�`�`p�wޫ�c�=�0}�3M�j�	�<�-������1�(���$ 0;�q�ha!�p�Wt�#T�a1�ٚ����c���d�un�Owh���u}U�M�̑$S�\�㉏��٧U�� �~m�u�g� Zl�g1"M�C���Q���`���Lל������W�rzz �{d� �7_@��m}�G����;&�M��q��X.�^�W�#���, [�Ȓ�O�;K3��=̂!-�-��T��<��un�t�OC�� �Zk���b�A���������֨����fe����DM5F��� 욳�������n��Q�ci�;��Eq�uepdDg�w�,ۃ�����A��(���X��'dbpiW�z(xby�G�jJ�)�������ټ��G�d���Y����.�g�?}'o_�`�6͕ߧ���_������7�1��E&�' ���B0k�">AJ���f%+P�+o[M�yߒ�Hl9_��6�	�,��/�ȿ���~�?���T�.�D��@�7Q����a�����ō��p����Sщ�<� Cn���o5���S��O=����� �j��F)	l��|����J�YP���"�'2ۃ�\�NΤ���ׯ�r3C�wxĲԚN��Y@p��Lo��s	�vhw��3�<=��ܾ$ 8��Cb��vk�y��� `53>�
�Rt&�G�$#ꁃmѵ��B��"=>\ɱfn�{�9�<Z���k��KE3 ���@�N�����G�8cq��Dդ�`qtL?.�kh���[]w�O̚��>㷼<VkO�Wh6y����{f�6O����G�',_�>�D����+]ם�{K�{�?��=\���h� ��u�l�C>��Z�k-4&��i%��Z 8�[󖃠����ָ�n{��$�[ݚ����y 8�����IX�9����4eKڨMd[��W�dP繖�w�˯��Ȁ��T d.�$"�ƬP�����n�8�{=O�O�M>���2�H��c�✪	� ���\V*(eU[�V��܇���Sh�����.�{��7�LfEϛM��pnf�G=��.y}���XV����s���,W¬��{�O��! ��?��=�	�)1}���ˢiu4md*���N�����]�cq-����q*\�#�Ua�ăͯ��k�b�\U�z��ټ�8;9�:�AExm�>GT*g(c���K��Ur_�8�Hp����y��݉Უ���R�"��v9ώi ���V����a�]�3����'߼{!/^�*�Ys|u�Y�Xg�%�W��q �/m4�u��M~`���o���Ƶ8&e=��}�j�y�Q�GPV;.A�M��jEb��o�e|��Zx��@2�A���n��e�-����>�G�ƣ��x��EVu�(���ux�I��/�n�d������^yf�<���C�[���jdE ��X;C�l�^��푼�9�g�������%�ӻG������m�0ޤ�.�.ҭ�M���dF�.Ǵ~sG=����N�`N�Ȁl�\�������n�}o��tf�x��ڻ�4=��d�K3+�(��6���00(+U&�y��Y�P����AjO�N�Q�`�&&]B���ypl?�T��g'�,͐�N؋[8���� ��vqn� �BU`Ֆd�k!E����������Z {sUM��
� b�+�^�s��a�y"iqdS���e%����;��������`�Z�g_���tOB�Z�X���ډ��B�@&�z2L�G�k�}g%����f���n���_(X���.̿*��. \0����|y� �,͂9�Ȝ�[j:�7���H��m����c�0� ����s}痢ٍ ��yO�o�>([����={��6x�+/�����|����@��(�� ���b�>�Xj[|uu�5��	�=��M�~��9$��)�&Zu,��ق�˟�,-��c8��l�f�i��ʑht�|~���Q�Ꭰ��	�����u�1Q��hΙ(`���:�O�7zNk/���b-�n�3���cؚ2���SG&zM���M��b��Y�A�� ���$�[-Ct�Õ��j	�)JE^��`d�̒	���ɦ�M>�2�OA��ߍ�ܒcꂮ9��se350m ��
��S�/�L�~{�r�G�� ��.�ą�w�gn4��^JN;o,I2�W0ާ�e^<�;�Ϲ�Y#��/�!#�2�^��m��Z%�J㈜��w&����šAz��-3H�M���@R��=/>]&�&JG{򷫼4]Jś��z�uk~BX{c�H&�Z���������߾��4	=��-G^Sβ��1	���g��z��ޓfs�?;[m`9f�V����r�e��h*1ۉX{1S9tz�l��l1�T`���	"�jV�?Vk��zv��Xn�G�����2�fx^�]�k�� w�x��%GUC���p�;���h\vv�1'�/<��QP��"7]'1{�X���o���:d����M}��T���-5-�)�>��>ȍn������h(߮�;����6L�ǂ���N���c�Q�P�B͸�O�eӘ�m����t~r$������q��t�Uc�� tO�Ol��!w��:�Z<��;�ezv�`l��1L�ݑ�Q���QJ���;x� �w�u��Y��'S���^6��4f�10�bf�[S_�6p���6�m��oب�n�	 n�7������Ť��kf����]]ޑ8��;����15^��|��\t����Z�J}�^��Q�\�yWҖ]C�� �C�vgJ�8?[�Q<U�YL�P���N�)��ٶ�oϓ�<yp{<#5K��޾���'����F:��� <]Ȟ�翰�����B|�6�t'�w ׃�-U��mp������B������~e���c�ݫ�S�< K��k`6ݓ��S9}�R^k֊�f:��M�F0��f	6�9��X/�h�Ƶ��׿���
�k+��а�s&��o��]���@p����l\�]b�j���X�QY�j3���by�����\t��Kj�(�g�o�Mz�9�)�+m=�W'b]��7r�n���l*By�7��2Cܚ�K0ԛމ���g����cVsʾƐ#ـ]���I���Mo���w��ˮ�������M��J�;��5=�lH6��:��d%*�2���;^��4�x�kb�-�(3j\�t��Hv�pb�rAN#KQ�O��� '�.9 �. K��?v~>7�|Ubu�n��¬TR� ��d����JQ	�+x-.$�5_/������j��^oܽ_|\]軂��������!����j���>���������n��.�{սݯ���IG�I%��N��������o޼b�-�:X�-�h��g�>�Q~нq�Qw�'h`��N���5c�� ��W��i�86�8������ݫ��'�g#�����k�waj������,[M&���5��Ï?Qz ���n�N�[�d�3ĳ�W
j�������`pxg�/�Fb�*���3 �et�u2�Ψ�O�L��VQ��A��q�Rdǎ"���RS7J�����D�aVZ	�0������=�0�����O�r�����ʴo�Cc��`���J�:L4�b�,�Dc�������̽��p9��	zZ����)�]�%�����	-�0�ԗ���՟���l,6?X���v��W�?o�8�<*+� �|��������]u>������{���e#q��V�\���g�p�6W��O��^�I��H,�[6(����}�����n��9����nŒ�����] _t/�;����A�NÆ�Jaa�rvޞ�/4�`��#����g���l��/'$��$�Զن[ŶdM���um�QވR��;�t~���h�L�g��lژ2������ �N�|�p�!%X� B���RO���@���Z��6~���_cW���EO�g���t�A���s�0#s� ��a%׏�X�ty/��O
dz27(������P�q��n��y�� n>�r�۴V�٘b:�1�6�Cj/o4��o��h<@i�qi����:ms65�EAxc0�|� ���ȣ�%H$"�#�)���8��
g�-�����rlp��e�q���� �ҡ$��)]�^�׿�S�Dbv@�?�ևl(�O�\�w�z��3ۅ�w�94���ڪ%�e���5ۛ��S��ȸcc��M�}�l�)��;�^�If���Z�	.)>"Е�`�-_D���|�s��<��/^���'����U�R�l�����@�O�}O��`���B��QJY���u�_ǈ���T� {��v��O�야T�Ǘ s)�a���d����?	FTX�b3@��� �����u�� ��w���������/�1N�����ƈq(�i!{g�L$o��Vɨ	95ac�� 7��7���߬lҌ�����Sk�Hо0~�$�g�Y7[딄��Y���8�Ǫm*������28ӂ2���17��{+�Yi���F���(y/��t����K.�U,��t�}����X�f�F�vȪ����{����W���h�q�C��~� H���o޾�oD�����_���es~�+���̻���|1�$!+�G�/<x�6Gcҽ$��9J��b�Ǻ/kׇi�u� |}��������3Y�������=���A������ѕ�m]����+?����Sf ���D��J�
x��>r��cW�sl�)�	ݗQ��E�&b�]��?�ަ��o�7����5�`��40���z��j�V�`&��d��^��IC�W'}���o0;&��uFC�"�`�0���\V��CIMY�g�a��g_��L�|��Y���[�ToH��1����l輱�5c�ll��	���]͹�b�U�jQv���qi#��{i�a���tJ{��\9�%� �]_������"�Yr�ύP�Z2�/5I�E9m�	&I�뚄/�o�������� -J�`{��<-����ߡ��Cl��]��ڞ��o8��J�02lɎp*Bc�1Cd���9(^����k?�I(���@�/�\<Р|�����!��H��v����&�p�E�h[姥� �3ާ��nod�t�ʃP�e5X�$�v��Y���	'�dz����h"耭�I���!1AXo}&�wC��_�����>O�+:�}h��w�k� 	@���yg��!*ށxT���2-�ao�ц;;0(�-K���2BY
!���1��(�~p3��~� ������tu��/*��w�a;�*�y�F�����μ�YʿG�R����]#W�a۷�9j��{Ɛ��U哮 M�m���ِkq@}�X���WG��H���#���Y#o_=������� l:�e�`+;����,�t6�%���	�&a�Y�`��I�ĉ�p��ʁ0X2��L\�+��%��\�ܻ�w�mQ,��W��]�{Z����=�4T��w�MUcFꍁi����Ɛ|yp���vM���H!�%������₞CT���]�T,6ۃI���OnuѳL�c��d�k^(��.��m&�����b����LA��p���43x=d��	��R�P���ӵ����=6Y=9+n:j�|��^�����9V,��c��� 3�泆Ǘ�3�Q`6h&��mz3���UWc6B_& R��u�,��fr||�)o^��xo��ל�1.���k�R�R��pF�41C˴R���=�Tl�_�M���M���(
<�s�/�IIv*�� %�=�~��X{v;���&���xllǔe>����G�+f�g�����Eև�M*��Y�3�k��^P�9�A-xq�V A4ĮM4�x@���"���y�5zXҞp��z!k��+����=^o:���}�Ҕ'JS��k�p�M��o��~��f�r���> ���ߦ'x2_6�9J�{5<��2�H{��n���nQvnh�`W�ٞ�W8���G�]��17([�(�2�$��'MdjطaL!6��3ǈ�3�5ơ���ƃH��h©���Ѷ��5?�`�m7����:�a0{�G�m{x��f'EI��}v_E�9wd�	���e�F��RlX�G9Ն�oM/���A� .��D�����9z����>f.�n�bJ����G&v�wQy���Aی��<f���対ƭ�yϴ��]f)IyF�1�$d\�Ï«�W�?�G<~�{IaPv��˟ߢ܊<��a�	�� j;{Q�3)��g���P�+/{R�c|A�<i�r���߉;���D/��ǆc�$;헍�Zk���7o_��?��o�+�T��I	$�3���ԂN��F�U6�9� F�+����(Y�M�1�Í�B�zpZ�
�j������n/�z��MI���xa��Ԍ�gL�MgL��,���g�4 �R�tfVC�Νqi����0H�`�fYc#�X�ݖR��#i����ƙ��N�t�M���[?n��<-�����8Ql2���C?�0�n�޼i6�{�j�c괱?Ɛ�e�С����4�=Y��R�z����M��-����-���̑-i�\Ă,]�������K�m)��SX,�� ��Cy�옝���*?����9�IE�߼{KT~wy-O���<4�i!&�ʁ�Gǜ��N2\���ֳ�S9;=V�����\^^����+�,ph�a�.���b̂��:t_N�M=p���������?�ih�jo�P��س�ڻiń�^m���Z0ΪÈ"h�H����6z�lh�6�����D]���G#��AE�X�X�N(5a�*��4"W��s�vK�T٦��eݑ��x���.̺��̭��I���q�Jʭ~�]���|���@�c�lYjB��l�=]e&�5�ۘT�6��Z��Rk����5`��JA�F�e���o�SS&),��0�ƳV�`oyD��2��'z�mh���!F՜�������t���md`�9��C�g��On0�2��0���>�+�5��|�ǐ�l>E[�^tZ�Ϡi �!sXK7i=�&��agh}�L�ibj�B�C���s}7�y,s��??6	��ǲ%�%�mM2І�Jf��q� &�G[��]�h�wo�O����^����䕉�%��s�f��f#�,\�H��[�m��{�d��l�d�=� "��#�K�V���JR ���  �`�|�ټ{��v@f�^�.�s�E�c�4�l��<��v�$|Gfn�gP���6� ����;Eb����������J|�ݧ��-�.K�<2��`S�yc�������0^�ף&����#� % �Q3����w�������O���o'W�-%h�it�~���rpt�j�h�{�ͭ�C]ݗt�L��� l���jI�H���Qߗ,P��5�%�^,�0��9���Up@a��KѴZ�6�xU�%��7��W�ݽ�#��Df�)��4"�3�f���\3P�����l�r��l�I�vR�e@"spQd���{��6bPv�+����f[:/W03C���7�;u�fq�И�	 h�7����!���+�	)6@0Om��� [�+Ya{�x��|��]x������i4�s�r��a�yb�����$���?�7k&���=<���o��˗
���>Cٰ^<̐�z7[vЁ״�^�;0�=��P�8<n.�����p{�!,��J�Ŝ�YϡJ>���2���g��a�^w����;�l7ۧ�MX�?O[3�.%�)
��W��x�*˺�8�Jfb@ݗ;�,ջ��i��Gf[�	̅��:mn�-XG�i˒fJ� �����~�g8�v��t��.!;6	�J,x�$���I�k|�Aز�$�[���?�-%�30D��`gD�mK_��|��Im��֍�c3 8�n�J8�L���k�W'����μ� �9r�~��Kg��r�����/�K��vs�lQ�����%��5	:��',0V�źq �Y�<rg�0��֝��YT1��	l�q�<�_ƲQd�*g�i��B�3���D;����~H�j��O8C�>=�,�Y��׌���$SY�k�ց`�@��ń�����ٔ��8���ز�e�(�����@૤���K���b(W-���L#0����PD��`��v( wȯt`;�y&�e�9��c����_��>�?�v?� a;`��K���f"1�k>B��X���_}_�Z(�Y��Q�:
��W�wC�:�����&������@Zr E����&_��3��f@�&��zf�j��>?;��}-o_?��ә`�8
�m`���̼x�N�#����rs\3�.�X�+}O0¾6D]jc^�O��ިfl�ÖS�S���<j�\�M����oدf���ܙ���M�a�VG�i[,Jnz� ��pZ��$F+3O�Rlٱ�j�$�^krN��m�����ab�QKAO����f����`{��� S��5�Wgd��xp|jo�G��;ol��6Ks^~��� C�@�11G��fɮ��6D�@��7����M��������;z��u@���{���ჷ�oҁB�[������� ߲�|���-�}�����������o���?�����#���cS�|�3�ܙ�y��� 䃞A��cp�XM��׿����/!�E���E= �f�����rj�����g�7�}E�w+&ێ�����%�)tY��W�� @���ak#ZX~���Gc@Kl���+�N��ф��Y��6��B�����t݀kk�;���X�EYa��vB�Y+�͜�����-A�ϲ��sGI��кL���m�*l8�I�W�E؞,�<'�Vs��l�O>?e�l ����`
�&�a��-(`�ƌN*��K�(;e�Q:�P��M"&�6p������ ("�묜�u���7=,A��B��\+p�5GR�-B�~D���MĿ�Q���w-1�H�R��{F�`�h�s�}��
l��0i!�U�����6ޖf�����
�|�!B
QKLA��C>o���6N�;�$;;�B�9����=�"��|=�q=���؞�یF�Y��K��$��d̼�Lb��Ԇ�7�	�q.�л���]��z�d!�f�)��^��)p ��������-��㕝��Z����o�[��hO�r � �Hz��u�8C��Ư>�3f��cd�F6�Aÿ}����l}U�d��w�S���6�Kv���_���0�R�۽�9���:�G�aJE�T�#�h����F#Ƥ���<g���K�!���s��N�X��/�#b�,vb������MaGr|4�������}�悂M�{���k9>=��ޜIG*�n�B�R+�s���Bݢ�6,�v��,d��˚�&{�n
1�Han��#�,�l[�Wx'B3?_t�Zi25W�䈯Hг��`��k�Ǜx������l�"fv���[c�R�Zj.�Q����*9��0fL����&����LV�^�M���ɱ�grx�� `"Cq����g���`�/��$�@�lgmkǜ�BoA�)�o��]	{����\��r�m��6|��g:�@`+n��Ƒ.�8�i�.Nf�h�E��X��nl� �G���$U=ˣ @��׃?\�-9�C�G���?�`�,���cv�<����Ņ�ܸ�ۻ[+\��b5���B<X�eXk�3H`����V��X��M-��gh=�\{��Xn�uA�6��g_6�lڰ���|�C�Q��yʆ1�����G9�c�՞U3*�¬��LX����F�A�X��e���p>QЅNA#`��ph�ߓ���Rt�z�_��>�>n���^�	ڪ5�Rw'�1���ZկWw���Vno�,}B�S5�>TyTO|ll&-L�ϱ>}*o����;6+)�kH�a3&q.]66nR��_�l?l �:�)�&�Ed��g��ϻ�'\t{�T	Z	�O�3�*���_��|������B�4n�C��1o��R�qx�l�M�1�6�5�P`�M�,pdE�̓3��`�3pݎ�O+���I�,\0��EI3�77y�&J���W�[,q�\MhI0��Wm,x�qN]a�(w���R�%�����H��N�,�J9�y�=k�w�,���R�<ޯ<��ʟ�*���;�<6V��q��#��6��_vB��$S�X����w__�������R ��# ���#�e�x�ੂ��7��ીT��<��T;�5�C�D��D�7���t�~��3�b"��'����2���0�?�E������8�`�{o-o߾�wo��^ܲ��a����N_����s98>����{a�Y�f�kU�x
� 73`r���=@��uc"zȟP��a�9�XVޅ�q��7�	������H�P�}(E�v����m�Ӥ�-�=���7v�BS0�6�P��`�)(5Q ��'�`���������왗����z 1_Ϟ��;�B%�-�!��k�ԑu��"�osndN��9�f������<�nK�U�Ik��,&�LA߻�/�W��p�٣	i�iזE �,(���g��2�d٨Tv����3�MSfс� ā?}��>���''g<$���=��ї	����^`�`��ga|� � �АP����i|oj��3*5{�X����{SJ����'e�.��L�1V�5����Ѥ�5]�+����]���l�9Ӳ!�4U������(`�=���8��Mk�%�2+,=��Da���h���YG�qjJ��U�L:�)�Ëk!{�/�U<>�ȇ?�����d��@���;y�Y���3ٟa\�J׍>��*�{�[)�F̒\[RٳB�+|��>;v��?��ǇK�Ory1��é��3i�� x/16���1|����C���^�e�P`8?b�l� 9�%q�����#23��p�o6<�hxQW�9�3�U6����v�i5a������=��|��H_��3Ƃ4l%��6Nr��w�Y���aO�2�4��D����zH�AMe̒8HB#�yg���"�X��n�f ���cfli�󋯓��L�)ƍ1�2a�l\Q�;�,:�I$«��\H�e���)��A��)!�0?'��sc�0e�[o<�X�h��a�b�A��1(z�ѥn�U3��NlZ����5`_��s��ZR�3dB��t<��2*���a�� ���4���~��%�o�K���hX=�����h|���,�4yd��v��"v ����;Iė��%�+eޔ}-��X�� 7#�I�)޶!J�_]�<�H�Ʋ���� �L�5�1� #B��N�֞���Z���?������7����v�R�5���lc�8rM���pdV�il+�D$��J�G�����1�Щ²��B��(�/�uـ�W�4ٽQ��4�ޗ��	1�xB�FӨ�:�3ЮE��� �(�Z��;�,#F��7 �]	���ٌl����}�S��#Š���6f��A������d&E��g��P�J-F�G��wa|����s�j�)8cq<hM�0����K����I�5����Q��50�0Ǫ����cR��:�[��:�S�?-�@��tГ����Uc���sn�4��+>����!��e�5��9�j�RdGقo׻_�u<ڬ�8#�B���6Q����g"�b��7v%���������@�7o8p�c�t+��@}��������lA'
�QF%{����k�r�c^����Α��� ��m��h��f`���f*s��Vp�^+й�(��3yX>��C����s��JA)5� ��G��v�6�d[���X�u�^v��]Row{[ɡ^�ýVf �>?���N�����
���<��K���3Ŏt3:�FO���Z�uI1�:�z�!�	;H�m	��%ܘx9k��C����uL����fOr6`�z���!X��e�S��p#�4�Id�c�H���)�+I��H�����Z��b�S�����&�zi�K��U�m;��l�9�Z��3`L�+兖���d�Ò�}�,��=�rjfƲ�1�2l�A��|���8xّ��`�M�p]���P����$e��KG��q�� �wk�ސc�T���Y wR*"��'w9�����"����-�7R��.��߀A���j�}��;��)�����,����H!���K;��{�dؿ}�4�u-Ǔ,�*}um�ُE��+XR}q�񜙾.ʾ��S�c��Ȁ�����8ě2�{�AM������y���K��Yr_� q1YD�Hf2��`WDN�e�]�s�nX�^)m)�Gy=����/ �����`���(��,�(3^��{#glo�rM�j��6��i�@g&f� 	'x�S�M\����]���=Ql�wu�TF�</ZK���t���:�����h��|���/�����|Bz,S�ҡS�7t����i���̄�3�}�V���_�˛{z}x%+����1�r�pb���pk����@�
��[vu5�&�֛�=��]���+�E	��F�����PW�)��ˊn��%�()�u��z����{R��D��7��~S�fP��s4�
vfm��,S7��7>L�=[`0�� ���Z>�]��?�V��^<{%�^��Wo��}�ם4kͪA9�>���BSh��$@�y��[kǟͧcF�4�R-�Ӄ}�q��cls)���ۓ��5շ���)�zd�o�A��{��ۗ�˕�]�98F�8����q y��7o���T�l*A"����k����+�"��5���J �@���nl�������4�}����N��eSә+t�R ���w���%�k����7Y�1����aYp>��YF�L�6v�]Oz��`�X<s���eX!I����	c�!�wY�2i�&��{����c��!��}�g�<��y�q���W���>�L�iͺR���.��8$ݜ�*%<�'a�Zwl*aI�5mR[�k�zg���u4�5�ɮ��֞GN��y�z�;�V�w �eMg6����=�5}נ�D6��ĵ@ l+s�g�s��]��X��ܞD���5��p�7�AB��fk��R��|?z��P�cg�Jt����8 _�]�����?VׂMډ�e��RM�ٮ@��_,�"��Ұ�)�y$ʇǕ)D��6L_0[~�ž#l�wU��]���R��b��jU��+�G�����_�u,Ar�(1�G� ai|��������4p�]32�f�C�"l��%)�I=�WHqP�8>:b������ř�m�<ْ��b.��y�"�:����jw]|�$�L�������7a��#l[S��K��3}i�2�BT����;��9q���@��V�p��ݡ��>�����,���Je�|�.�6W��H�KB��ƚ�ҽ�c9:}���X�Ɍ,�5�k��&���8�'Pv�X��M��ņ�N�_?����m���#y��DNO���Սl&9�{���U"��#�x�bI���hd@gf�:7�L1^��x�;1(�(���iMe��p�Mb���R �OX\�!��9�n9�-��F�_��[2�X��D,#��-rxxȇeL8�cS^�MS2�S%ޜ�\=�l�!�@9_L��1����~(�0[ˣ�>:`0�{��h9���\�l���&�)�x<du�d�ʛ@���e�άi#�&�5�뮉�t�p�a�^ق\OpΡ�����ꁁ���m�ق�6�KF��AL�P�]G<b�������7Q���X�Y�3�rh��Ҧdk����}��BO���k�/o�< _(ABK�[0�����86a!;�]�X����k�6Ɗ٠�g�zOPZ�D�	�=�Ъ���X�6������l�Ɩy7q��Q�rf�zC�`��A�� #�~f(]�m����� ���])�ÃH�e2�(-�t!��H$mv��gӇ��(v����1@��a{������۲?���'Qhv�q����OB@� ��Zs�1�H��zAb�o:�� ��nJMvZ���|9k�R�P98����5��4��5;+7ވ����1y=}�L��2�m� �b�_j���� �Ї�ź���$LI,Z��W�q�P�����c��y��j��b�`���롪�8����x�t�����Og���BcC�.l��Pg��`���'P�C��$G�
�#��<"ڍ����ʭ,� >����<#{;>#��s���1��6@(�c^�'F�KLnԐ�i�-+2V-�ȼ�^���uq���='�Ę �Q�$x[�G��_��>�b�#�B�1�$�������X��������R���G��z����`��P��m��ղ�NJD���I,w��wp�OxՓ��/�0Cd_ى��Tb3�B��q�Id���)0zsQ��z��n�3�F���_�8���;�t�(��J&s�G����ĺ)iL	q�-5��1r��뜐h ��+>����/00�ñ,fa�[�{g�@����r�_�-YΣ��9w�Ն��W�y���'�R�_:A��ռ�~3��B&cW�y[�%��Cb7?���ZZ��s�_�	�����H��YF\3xn�2F7�M3��!���M��H��_lݭc�C���x���6�s<E�Ɍr%[v��� ��?����5�y�S���n�1��FA��Y�M3Г�����#��L�j� 3�(��@�A�7�Z� =wh���A�4����|�ؗF�	�W�kj� �K��k�e ��P��i���Q=��J	�=���ޟOy|�sc^i+wNd�8���s\�V)�;��E�����b��R�3V�����&J�cI��= ~{����u�1ݽ͞%)��/X�,��9z�]UY�W�~;�GS5{ ��3�v���q�q�CMMM������N
I��B�$��L���(��4i�Sg{>ƢۺR�s�M{UGۄ�/����]َ�ܩX.�W��K��z�Ӎ3q�h٦_�Y��D��k6���[��,ͤ�����'����dJ?! 0��j�3�˪�� ��`�k2���,�R�x���	l{�g�,un��=j�`mRF+�A��i�`�4lx�F΅�~U�W�Ǵ�@�r��$��BI��;ۗ$��� ;C^��ao�vLf����̌��$wJ��gO�e�b�Ơ�l���u X�I��6�.�aB��T��u6��Z����Ek啹!wc6���Q���|����ձ�)�/^�$�w���[&D�6�R*1s/M��X7G7җҟ�y��A�:��4}�>À�2ى�zz�=��\O;,yV����������W�@���������۴x0p���03zu+"��D������Q�����+v��?E�(�A��n��i  K����}�2J�=�Ill�9l�v�`&�c�>g��;W�랜�����`��m�f�g&��ӏ#Fi�rm�GC�_�=~&����a!��F�]�Sd����.DZ���#E����z��|Ŧ�f�f,���BZ*#��dD7_�w�fk�ܐ_� ��8����<<=��.j��y�c�^�.pوZm�����M�[�m_�U�S8�����k,�������k9�I7cr��py��������p7�P�b06����'���� .ߤg��w�����KwD��u�=[0�hF{��d�NL���}B� �Ck����S��GR�����6�����;6�yr���!x��Lkm!�)ۏZdvj?K����z.܅i����69@q���� SS�A/X;�j�Qh��R�9�"Z~_��1�?,�r�x��e�1b|-��#����c��ؿd�pO����L?�6^�ɐ�?�V�x����a��Qy�?��2�j���Q�ƺ	���c�8�ʙ��'m��umDl�M���@/��U�6v�"�ƙ#[<[o[q�>uх��L�8�ckA�BȖ>��e!Ho4еьiF�i\Ph��]/Y���2o�=P�$�`�W^��P?7F�EFIM,+Ƣ�N���������=7֚�>h���� �X�����g�� >�;����j*��sk؊�����y��;ۯU�Z���a���]Ve'z���^b�BKk�qۀ(�W�{�4ה5���{5�vi����s4�,�iY?��ΡBg,���̊�l�'����[o��v��� /�iL��I
p�g$�oYAJm���c���~P��A�;��d�/�i��
B�I袬4Z,J��?�9��l�l�qh)6�x�knMm��ҍ��t�i��UMa-�r�mm�P��U�� b!��
����dNhBv�l��z�e=ma�{�7��K��:���L������[�K�ď��o����s�؋P79]�l�N�4���)�_�t%O˵JT/�VU��&r/��IAZ�����yu�Ȇ�p����)�,�(�.��.�`-�d� ʐ�*�N����|d�˛�&�pJ�1��qE����A~��=O�!�J��z�k����xb�Y� �/�p4!(A
~l�Tg���~�V�ᄎ����ۇ'� Jȭ�
��Q����+����o�F>C�cYr=�������"u��l-�M2ٍ�u����T���_CV���!~L�&�B`LvMǇ��Pi{,��L���ć�jzr�v?�T��c�����]�Ѳa��N|�`�r�;Y�>7C�,�"H�M�A#��~��yG���f���ڴ�[}� `��d&h�Im�֭�<E�nH�x>�:�	n��R_��{*�A����ǁgb�h��a^���wj7��f�	��X+��-F0;�@f�ש�[G7 $g��h6�zH��(H,(d�T<�ʻ?��S�pPK�3�V��\Y�n)��m���V��\%
eh�Qi}D{�6u������|�� l�g��b�2��Ѯ%i�*th}��e�����g��A:�`O`٣fr� ��1�1u�4�d��5ܣͺ� o.���c7����Gz�k�2��-�ʍ����4��v��,նAv�R��k� Ҙ�\�u�o��Wb��c�#�\�Զ�M�m�%4�/�fݴa$v�W҃�^J��������a�`�Ր
���R��,K�OҜ�)g`�]0�61�\?���L�{v\c�i䐠[ݼo��Y��<���5��db�K遐�w+����h)xv����ͺ��1�<S���x�-h�d7���^h�<g�R�[{���J����g}���W��w�@���ϧ8��w/�3�����=ڀ8MO.��Z�^)R����>�j<��X�#�=�ؾ30���{y���G��y�c[�Iu�՟�h�\(��R~vO�d�Z\[(J
��L�z�����7�»���E��A>�y#oޢ�qKğ�whK�GS��`��GVMϵ5D���fK��5B_��������.��.��6�n��Oo��aFk����{�?����c��1o�����ܳ���{�6z��9����� �d���Q�&��ehVQ�3� ������G�����5RN�,�M�*	�Wl���*M�(-��v���1�q�N����q~`�R�5R���TN�}��������=��y)e�)�iƺaK)a��d��s�С�-2w��S���[+A UX���i+�Lư�[��W���X�2��?M�Tn6	�ZY���c��[���>��t0�T��1F�� �Z�a*Ԇ�&�+���Ӕ��EF�WW%����74\oi}7��j��e�қҩ�ĺlǄoҡ�`�@L�FW|��0݋������)�͞�iI�\���[��!ȼ�Y�`�k�,`������}5��:LoyD@�(�C� ة�@�������&k����^�7Ԋ6��v�d*87���O� �� �.���{���-{�M�4(�VF���k�u	��s3��Hc�" ��w��*���G�l�;������Wˈ5��R� ;�@ZR�r�tٯTA���}��߷L�>�J 0}�љ��|v�W+��m�޷���E�?S�14��`$-Z�PL��Yi0H���R�c���3R�A<@�y�N�U�1��/������\b�*cqF�l+���xe�l�����.c��'���r&���+�X��~�2�ۃ4Dϧ4������ud�P0�Ki��=���p�����p�_�+j���\6�0cՓF{\ 0�~�2����{-�m�6et;������ˁ|�ث�=��k.�h�|v� ���l��uj)��?-M��O���7��4��7o~�>�ĺ4C��p/��Y.�����AN�����%݀aL�%u%�ī)��D�oS��=��9�Xuus�(�������_Pp5�ă��r���l��(PY��h���K��?�N��To=K2���t�dzʮ��
�V�t+Xe��ݍ�����͙�W�:�b��>C4I�}�L`��B���/[�<qok[S��sf��=Zk��/t�9�-�;��d��hT���<��-�����9�b����AN/_�f�$ヶ��T�����w��؇�XZ3��%DڨJ��t޵%�o �^ e�1=O�q\�ؙ;=ꠠ�@K�ʹVf�QW��z�(CA:=���ef@�Y3�d� s�*U�Uh�����:�wi��P��{��]D�`7Y���:�����Ʀ2!p�Z�8�/��3]X���,23d4M��!�0�;���Ɣ�B��S���!��b� �<'X ��lrA@�3a��n��-yo�U2��U���їܤ�^��i������qCFUؐ���%g?Z��sv� Sa�r����y�8ޟ�^{�� �q @�3L�扽Vw_\��1���Gs��z�����=}ɎON4H{!�|������a��w��X�
��L���Z����6 �"���@��!+��MN�0w ���á���$6��]�-�0R<�v��|>���Iy�0�_��ƽ�����s �	`�e�>	�>>��W��g٧-H� !cfs��4�13PηL-E��q��``��>ˤ�\Ki�-3[@�}+��"�m�P�j9���yd��FGS��$k���0���-L���+|��I?t���A�J�5V�n}���LY�L����O<�_ɀ}|J�W��:��V�`ѿ��@�]@��o��`=��%A�@��&��B��Wm�ԭH�s�l[:�seiٛ���f�M�g�1R;hB;,��qO#�)X�U=-�c�m
��e �8[l�&��f��Z#̭n��(�u��ܛ�-i�����@wI�[z�EӢ�t�6�$�]C%�V�=�:%{X�
�Y����O��Ne<�|yo����B��lT��BA߂�R�WA�#Q��M0��n0�|��8�����Q��[��HFG[nz�� 5�$]##���EMv��R[�Oa(��g���w���f��-h�1�9fY L�&���a3�љ�#�m�<$�e8�ϖ5�#�+���2����o��&���GZl�b�D:-�6��ߣ���܍��S����ހ��^�PP�Q�f���V��W�x�q_�!Zph-A����rv��c@8^9H��f�����V��[	iNI{�>��3��Nx��`�s�fV���.[�FE�zyF�6�^��`� %;�X�Tb������5<Ps���  ce���f�[T�ff5��u$��Z����q�,�XM�H���g�	!��g�Yn@c<m	��&��c����}�����bE/L��lѢ���pk�����JYV����R� Q�Q����k��Y	��<@�t��N�x���rA6���^	��1X�����@k�����L���C-�YE���}MkywK透�7�i��M
���yJ7氡m3����Ͻ�ԡ�b�����9�v��{��Y�z�uQIi�2&>��L���%Ϳ�:n��_���>펃@cIq��G�d�sg��6��*5�Hw��ka��sdf�=g�����Ҭ�����J��w@��ߐ�(#��U�8;�\��y6��­z����E�A���C�_Ѐ}j@�"ȐnV�<4�J�G��f�+��@А57Y|Ѭ;b������zi6��矛7 �ѯE���ѳ�ښ���ȼ:nH fq����vH)�,g�����i��$6�U�J�~0K	h�6���^p� �����wt�͝Fd�u~����~NM���*���k|@�*�#����I��j�
�ۻy�E�b���#4w��_hD|����)x���
�z j�T˭3�g�@A�T�
�n�P�'���)��`:����}sh�63Y)�\nL���2�v�H��ȷ�{�/��K��ߍL��|�����$�J���D�)��V[
�k�_�Uy�B�c�~�4���/�[��C��Ƙ/+FȘr���W4A'TPW�cM��-��v4���X4CE�zm �,��Z��U� �xG��{�ч�0�&��UP��vL����q�b-�(z��/͒�O:_��K�,x��
��@��W�%��4ZUiZ0���e�V�͟�������Ҁ��ʨg��J3!��vdD/���Vݕ��NƐb��,XJ��lM0����X�&����)`%�님��H�8zpe\#*����n��Ƅ6χinBy�tA�)l]zOx�5J^Pm^�d;�e1_�z��Q0��i����v
>aR��Ohܺ���-��ﯸ���B6�G)���69�:�xz2�  �H�\GЌQw���X��7_����W/���^ʿ�}~G��'�Ә4K)Nf�����X�͗_y�>�I��I�H�&�v-Xb�~��������7\�@־>�׀@?�o�I�ٮ����Ǧ�ڨ|~y!��_t>����L~��g[���u�g�z�N+�gd�E��=��3`��>��������f�W���,m�幤^�LE���.�Ǘ�Y�k����S�j�@��b��)o�m�!t�(?�Ap�~�~��4x9�t���0�F$��-MSu��Aʷ|k<R�M6�ʎ�wh��ةx�W����	�6BH���,2������b� ҹy�Q@l�] '�Y;]j���O�*���kj��jP�{R0v��G��{aɡ�Y�ϑ��#ʭ+���<�l�Z��ƈ�6 f�`[}���+��r����� ����x�de���Zf�%�yA��m��/h)��M2���y�Ыh6�f�Q�>]�YX�� \����~��4�?��r	f���l���1؂���Dc,}lԉ�&����1�m�Ho�L�g���R�)���dj���nJ��*���!(��g`:���f�>\9�����;,5@�҆Q�5	X58�SSV���s�����P���f&
�c��>_QE�x�,Ɏ�D��tU�ِ�*S��E���  @߿�-��%4Za����:T��A��U2����~����\d�ڡ�� =d:���l�QX��}S�^�f��]���W,x�F�[�3;%e����;�E�&�&�ͳ�Y�ۘ[��
��|� x�e�=Gd�d3V{� X/d�b��b�Q�W'  �{,`ꓥO�Z������b���ɬ�Ї�z2ς�iz�f ���d��4��o	�j��� ��,e���@����}���Y% 0~�M�ŌKMߖVZt��|v&߼zI6�=ʇ7?��u!l<�6�cg֊K�u}wjAPô~b���.�9Ă탞���1[��.���>�w��ݯ�4����R���5����φ�p�\�O����l�w�0�����bU��Or�T{�+�A�sJ�I��J'dC�?���N��3�<�`�r2N�%=��_�����lG'D��k�	����;��Ӫ	�8�k�*w�G�����<��'��&^!�ߏ�� %����R�o��-���#v�G��m�?��8-�ޏ��E��y�4��g�GO�E�6�-*��=x�Ul`�<X���E�7Z���m�@nܬa�j閞LGG���Ԉ,�[
�VL��h��*�D��i�\=+\��8��ݝ�~�w���Z�'VS,��k$�Ejs�)��- _����͠Eʐ΅�Bۀ�6D3��)��9bʢ�;q5��<�Jc무���I�O��<t �3\���&·���DkE���¨�`}k"]�cyc����v�uI`j�v����ځM��J��v��ZC�֔��G�
(��}�>�0��e�9-'j�����稜��� 4R�"ͦ���B7p�_9��H�JB�h���	�UJ9�_&f��]���T�C덂-���FL}a��At����?��l��=�//��#M
a.�E�F�t8�~�QƏ#2uS��1L���F&����q�6�-�I\O�|��^c|��GQ 3����ѿ4�Ɔ1���R{_��+Ǣ�u4ۓ�޿��+=w���F�ޒ��o%�*�����	u_�Uzt<R ����h@4{��2�{�+L\b�d#^F�<�Y�U��P|�n � y�}XT�ď VM�O�9Z:ƖY?=�&7�ҏp)�Y"�:��Z���|�~_0瀏��ɑO5�����/�Wbg�-�2����vV���.�lUW_���l+�9p�9���}��9Fm�������HZZ��dlki��Z2��TX�<���d����dN�'r���x2�1�c5>S�$Jh�ofh$-���[eWR�Gl�S��~�q�dд]�t� iI�`�96Ū[C��������]ab�v����[�y~�l�֭� 0>ҴmH��H:�,$��ћ��/�P|�w���Q��k)��V7�N5�tu��d�`l����w^�Z$�������#�a ���Ǳ�Aɇ'v��dq���3/	Q�&����+!r' q�<�� �
��Wy��XU�WNډ���C3�ޥ����H�Q/[��������9B΢�`���)ɭ���ۧ�t�A0}�f���Y�ZV��:�+d�hVYe�y;y�I�,(�$��F:�Ϫ��c��8K�Օ��˘�4�b��"ƤUb��Y���oBWscV�x�}`x�=�$(�#�"�Ե	�!^�)*��Rv��)��*Ѻ	b��S��nS$�]��S��}��."5�y,%�2B���D��B��#�1�0�������g����
z�� TF S���f`ӣ���l\�=<7g,h�%s��X����1�5{24�)�&������OG]$�-l,�����J��������]wR{�Σ6z���.��nB=��V\�����У��q��%��(pLj�lL�9y�i��6��5�u)5��A_���Y��@4g�9O�rr4��v�t�.�d~ˎ2��x<�}SF����	E<��`��כ�Wj��|��Gz�g��V�K�a���E�{�Nߓ�Յ��YS5��?��M��l{2��dH����ǴW�<���U�f�G�>�f'u �I`�1��a]�f�՞��,(���׾��k��sK����бbZ������r'0��a�X����
0| U�L�(Wp?` 0f���f����^fQz"ƭ�H7��)v�*�1W[t$�7ik�S!xĸ�nG��`�J���g4hI�x�|�}��O�ĂI�i,M�܋��>���������s���:��1R;tI�~e!}��h�j�XY�f;u�B���ug�b8|#�յ���/t~����j���\�\�P�Lɡ�}L+�eV����\��P�5d���%biL�WUza�	�|[Z	;��>\���V'�ç�3��"�}� #���C��&���F9;;�>�&�r�3fF�:8���U�繂?�(���,#������G�4a�Ĵ��"lT������3wƶ{hN�A������ )Z��Tr�r	�Hc�� ��h>�I}V�؂Ք�2f=A,;�>L��V�ڧI h�݈Uf�q��Ap�^[k��龰qYAE ��W�=����i��k�v�S�n���}��{�<Ӓ�7�����@�t��uY*t�3cQ��Ӎ�G�S�(��i8���	To�
՚��������Vt�Ƿ��$҆�Zi�7�f0�3���Hm��O5��f�e�HA�T�K]�6A� �������6q �7����U�q��L���B�O�<����䄽���VQV`�0]1ֽ@��E<4����6�7Y��Y{ ���2�a��d�'q��r~<f �m�`o���+������F����|���r|rf@7X:,��q��heU�����b���c&#��ޫѠ'/.��9^xK˛�H�S����vG˵,�s��_�c���[�e��yf���ѰO�sdۣ�,��f܇��f�Y�"��vi�n�VI�۪�鵺�(�������~���+��pۯ�<��� l��R*�[)�sW܃J*o��B(_�l�7Ǧ/]a��1fL�0b����آAD���!vw쁼��+�%�Q�˵e�P��ϵ�3�Ǥ��[�gO�Y��e�b^��+��lS��dG���'�����؎����+bi|����3�J����C��3�/_�>	�^��Ӹ�n0ؚԵ��Z�J�!��}�%���mwҗ����{e�K��f����h��߼������Qe#�4J�j�Ķ|�U9�8+E[_@[��גqcD:0y���F�\,*?��6�[?lryb/9�G�����eHo@��~��\����I�7��d�G&�2m��Hoi�4p'm����i��W���Fl�~`�G�&���ҹ�����Sٴ=�n�ugl���"=��#����M/�&Lܼ3�����=���ڻ4��ր�� �װ���V#�j�"c��ZT�f���:`ȁG���=��& ܌��p@> u�4W��.��m���8�|M�vL��Ls{�!K[{W�hc0UV��5bH�A[���K�Y���B�5��Cu�V���
4�d�X�� Csh���|6��ٓ�`륒�<�=g��t?���V�k���z1�uJf���h��H����}�#�*#5��:DW�Rz�5�[UR�>��W.�GC� �|���+���"X[��j �R�aG���zX� N� �0�yi�э���D�Ǥ't�pva��g�3�OU��O'�����f�%��d� c�'��6K���9G ��m)0BЇ>����<,3��i�u���27\.ٶh&�n��@{�/^<�����tH�v2>�g����W�N���[s���= ��u��ߺ�.�fV�y
24�{4|-�ۆ5f6߰f5Nf��|��+�@�M�}j��]�}�w�������d;���.��b����X�O�������������gub
l-�ڛ:���t�Y���$�F*z#�WL�!��pDI���L�&:6��_��FP �XU�D
�6�>�;�ٜ��l�۞�����Iؽ���3ưW��E��"4$Xn�����vǱwIF�F�8	P��X�x ��l:L�-�w���^���i����P!�@+INMO6���L���7�[b��u�q쀯��U����W�ܝ~�����)�9�I#�T�ic[%ѣ���N�TP���C�nU?0J+wb��~ѳ��#��U�X��CW�QHl�ޚz����'���V�H$X�Z���Փ1�ɞp�hD����=K���ژ��F�j�u�C�Ǽ��uh���2q�;Ӌ���Q%����d��|m�Y�LZ�������yg��P���V��D��?O�w�.05MC��\��
��f�n*��43n�l`T^��E�zh"����)ڛ�]�L'}�4��.�ct{GiE�	�e��`:sc������16n|�-2��+XqG#�X�Yb�*�:�!Ŵz���,G+��kY���z>�Q`�6����|4��O���TN��u��ʡ��-K��������߿_;Z�[ �bLaC�Xِ��W`t-�7LiLzd��Fp2�Y9����!+r�ۨ a+��>>�����k�#ax�L4���+[<m��?���M�߿'�;;=�R7��鑜g�e���<�ײD��7d�+ث
dDNO����L^<����4�l��X�i���le�)�r��N?n�������[ts��k�[���;��z�t�?`A@�Lotl�=/s�7�.m�V��'�)pM�������R׫���4� k�cu�5�Z�Y TzTR���ɻ�W���7���d�Z�ʠ�<�z�`��jg��3�I�'�.)�KD�$��f�v@L���/�X�f�? �DZ���R��{��C���@X���G�����K��Qj4�����$@g�3��Nxdޙմ0ߝ�tN�tL�iS��]^t�Z/�,@�}|4����F���Ky��RǺ�����ǰBT����t��fk�p}#?��������6�:LtWy`˼��`��L~�n1��o%���}(��b>7{���l�֧��k�I�Z�y`�C[T�3�Cv+�w7��WH)���+mv�B$�L��4�v9��i=�Ԥ��~'|�L-Wսi��{�r�e�|�RʸEg��L&�3᱕��8u�� ��Uԏ�����M��=Em)6�����J�j�)��a{sT�3��u"n"��vej������S_3|�h�Ɨ>����k��	(�j#�1�K  
��AkY�Bv��5�b�o��U ���{���mũ� :O��3`i�'�����!6��X�&]�IՒ�NS��}l�������7��<�y���˼�����'�l�b��M�w�)X�]���V!��,c��\���褎O=Ҫ������ؘ�~�ژй2pK��:<0_���`feE�V�[��h�����fi+9:���]VmF�z?�:��Grr4�W�.�˗�
��ɳ�3`'��݀�f.�)Ѕ�݇��r�v�=ث��TY�¯��AT��( ���b��ê)/���7_����/��G�D�`S	�SI05�<�=����@AX_��pt:���cn*݌���潬g�,(���yR�5W��2�1�[+gL�H�t:��}y�\�P�uy~��t�����L�@v3�)at�_�����=���kG��`�̞@y��7�K��1S��>����@���=͘~�-�c��'��S����r4�P�@ �����:�g��g��ܗ�#nH��YA������#�=��^�k��Ҵ��X�!	i����g����o0��@T]��;�i�}�סWb���}�o?���?�C��4�h��{�7#6�r����.h+k���ox� I`n��F�}�X_Ο=����z�J.u���CG0������=j����J�~�b6�`m��Z��g�����AEq�"1H1�vmPGg�:w��7��w�ϼ>��]z&1�|a����iQ���iqE��=�KK�J�O�
i��X����8�9B�j�8vx+�6}���?[y�{��N����-���.t�O���^�ȭ�� ���Y�'F3.tp�������t��D}�͉���|4��N7��=#Q����&؅U��s���aa��a鯥d��!X�DY"���?4-KN����'Y΍"g�@�{�-uC��zt�G�i����Z&�w�� ��ـ�"5Z0C���z��0���b�|H�:ah��GN:�W��.,�n�M�S�N�T�g �[hd֤�:�&1|�Z�?����3��>7`����MHR0��)'�L�	k|��6�� Hz��+������z��4�RF%#�hE�t�SLz7�wp��]���~>rx�"�VE�=sc��a7�+J� S�nK�F��b�ۀQ�ecHI�����D�Aϳ���J�	øF�"�g���ͫ/����|�*!�o�7Ҧr ��b)�c�/���c����
�9� ��K��,�w� Ṿ׷_>�9"����K���I��w�`hov|T���X�_�*;W��^Aߜ׊E��@b3�������V˛�p9{�9�(����W�����Fr�Ꙟ߹|��rv|,�ހ�x���֌��.�1���p�G���u+(�gzw�tkW�u"ۍ�):i ���Y�k R����;�1��w��4�u,����ϋ9�{z~z�Jţ1�׀��UNڽ4�cI�5˭"U�Ѐ�ȓ��>\Ƀ>C�Q��Ctς�Hٷr��<K?2��LZ��H����
�1XJ��׈�������k������k_/�9��^- ����eɧ0x{3��ܧ/��0����Bpn��J.t,��N�>�I<��s�LF$8>K�3�b�`�v1gE�T�E3���ul<>>*�[p���MVg������܊����~��;b��I�(v���_G��`?�j��T�f�J��\Ϡ A`��P���J����]�h�H*v}�I:��;�N�#U]�ͤ�q�f�e��"z����>nVp�F��)m¡}{'1�S�Rk��B���5u"*��U�U��X�E����K?���r���z��ئ�4���=p��G}TV��
�����㓂�9�-�����Z�A;t�@�U�0��*-u�A(t E,�G���LF�)-#08�������@m��}�ⷦ~H��r"�}��w}l�}=R �H��ƣ�\�&{������)��(WW3yZx��uTI�����{&k�����^�1�(%���B� �����.:�$��ڕ4�BѦ1u����i�	�鰐c��!D�����U��r��f���8���sM���m$���Va����s�Uĭ��6ǆ�.J��Z��r?���:(�?*X�[����`��CD�$[O��>�R��
vX�d%�>l�f.O_S�K"�"��!�`,�Ntv,_<?W �B~��Wr~vҸ��1-�����
^R���7����	�
y|x��"����L��/.N	�c̿�(��hBAp���Y:�a��`=�(����h��cfL����-����ʌb3k�jVΒ��%AE����!�?��٩\^����1�-�]�U�2� 4���!]���7.��t�������!�ϗt͹l��-Xw�R�Ŷ�3�x+K�pm4����:;9#}��B��t,G�~���L�}����R�f�c^�	�.w`�Pxas/�=��2����S>c�:��"X�u|`��p{�qw~�c�P%⾏��D�����&��;���S�OUR�4W����ixuӕ�R�	�8\m$簤��3S���H#U����{���ӽ���U��;��;/2<y�����(E��$R��3�-�μ�7�Z��:v���j��4�tM�8NvV�wta������=�հ�	��|)��$�������f3�&ޘ� �X,���t��t>i�u�`�j�0�!����C�8v!���h�C�R�GQ{'�oN%�x�=�6�   �����P�y��ڹ��}<�S� ����q�(�}����#ոZ>�G�Mds��u}{#7�wL!�!�^�@@x�4�	��fzv6����as:�Ǜ�������������FK0 �W�c���iD�����,3?�hb��d��������'���?�"jztL���ޚq�ۿ���B��[Rt��&�.����5��tzL p��!�ԍ��t*���?ɷ��FNt�O���Fz_������ӛ;yXV�!�c~���ݘ}̤4X������� "ֱ��C�8g�ٳt<���B(>a ���^Ǐ�XT��( ������/hL��+�Uñ!J�|b�����LƯ�f�J=0�d=\�g"Nی�ъ��2>'�����������e=�*�r�A�
���Ӈ��+��� �m�\x+�|&P�F�B��5@s�-��F
B������x&���|���d�g����i�خ<\�D��(���B��BA�D�諗�)��=B�����"@99=��^Bsrj�~L�QP���!]R�R_j��`� 4gR�O�<�"��x��StW��4v�y��0?1�
(��G2�~�
�� �(=/���5��YD�|V����	{�*���*�E�F��������暕a[�4hr൤�]?��y&ձ+cLQ�FMXn���3=������|�J�]q�aׅ�Ll9vJ�J��eF&��x�M�f)*�?��>k��wb�J9�Ֆ���C���CH_��X�6}(;M���{��Zp���?k߾��7]Ʃ�':�f_���R�KuH,����n4i��L��4�X�W�u��-���� �QYyZ6��P��H�,�A�Hb�R�\���+ ��1F�|*g�4B�r\n����{-��3y�i �2Õ,r?'� l�{Ƈ�{9;{�a�heE3tO5�$<8�c��]p��i�X��<t~��t)X�qF+�zK[ �r�"S���($�yKf��wz�|��7~�wى:�U���e�>A�}Ą9��=����ى�kE��J)v107Ԩ.c���r�`a��5)�4Ԥàu� :Xl�X��}��!=111uL
T�W��}�ԍ���psê'c�z�֣����X�f_�g�e,_������nZgt�~����Tl��|-�EdE"y�%�N�gC���clW}>\�i�驥�Py�}ۧ`�D7��y%�������8q��(~z��<�Y�βx���nHF����2=W6��m-��@+r������* ;;?��F�h�:�ʛ�Pg2_W���u��FN�ҙ�����}�H���6 ؍xv�[���mO:��ck'�"���樖�e�~�(�h �|q��|Nݵ5@�r���W���ƞD�~���ml���Ѹ�/��u�1z;+S�!������Ɉ����w�qʬ�L�q�	��Ę����Su� ^Tѹ~#=
L�4���ՀX�P��F�O��\�M��߾Ԡ�9uW�b�l�WhH�!���x~}�7��p��>��U�g}
gOs2ZO���NNLO� �UʬN���\.V�<1���F���lvV���^1�3@Zt����sj\ ��x����1�[ ��cT��\s.a+�h� �'7��xnM����o۫y�A�x�.��#�����!��Z/d�s�A���[�3?� U��h
�1���h���8�w*�y�=� �w�}-����7_}��@Z��5K3v^��d�uBꪑ`؉c�`cn�3 D\Ҽ$��Y�ZO� ����e�&{l��v)(�����h���&������*�}J�u���2i�&�xu��Ӎ����K_w�n�|���㧶H���L��4����7TS�ؽ�H�/w�뇌�h����@ώ(��l-�8��f��+<��@�Kh��#�:Z��\��Zq]CZۖ���t�x��Z��T.u����i��Y!�
����Zvv����?���x�>��Ke���W6+c�K�'c�-IZ���]��8=~��7EϠWa�,�Df;�6�؜����k��iF�4Mue��~�ZZy�@EK?�U[�BlҀt�3��[Cc��h�Qaf	���|��:�և�h�B�.�i��� ��[Υ^���$��� f~~�V�_]�9I> ���˚w�����~L�`�E�H볣���ǅ٢��h?��, z�J����م\>;՟��-��.	d �&
��n�I3�[s8}����
)'����t�����_`��$�X���y��%���>,����EO��<>=0���}��BZN��Y��YY��jRi��7�L0�Q1�,�v:���R���v*b}S��,� ����5U�h ��[A�2��.k��!`��#�^� ���8���!�V�Ɩ���͹��<u��Y��liSu]-CJ��Vg:��Mx)?�pδ�r�쐞��{��}'���fɉ��5���P�+1wU<;q��j�Q�=��_<���������t�_ɻ��:nf�0�C����5�5�C{���)���hO�qsvzB!��-����s�S����ͧ�i6c	���j��Ȓ��q�L�)�� &�`����s�����3}���Ĝ�|��9��?��OG���#��p�Ṯ�l=�GG�O����M�������fs2h˥KԼ�d���@����5r�0�Ϧ�1��zy)��_���~{/^<�[�F��R5=����~���lA;����?͘Q0)DN�����G��ﾕώ�e��������>)h�[꽜C�����n��UZs{��΀�����	CX�
Ú@?g-ثd�h@u�vu����&��6�*{j�}��@�/�}F�{��C ���]�.�I�U�H�p�bɺ��7�! iǶ .m�dcj���g�i�2߼m�k�3v4�v|k��3c0�����V^��I�,@�QbO!��[$�^����d���_�,u~Fy|�Ql�ke��]&
�(����]g���߱*��7�5�c���ڊ��d��%>�������O[d 
)�?P�Vz�ш#�6�8)ݳ4"�r߼<W��r-�{7�I���x�i:���ޚ;#�������{������-�/�l>��"��B6I:��SJ�q1U)f�Fs�"�����*"�f1H���f#o"�=����KKQW�`�� ��jZ	���Q����Jnu -�%j�>��sȦ�R�Z;�ښ��C#8t�� Zo9�ۍ`���!=����grk���UJF˭g��/^,x�"�)7���g�c2����@� �ՠo�n�P�?q�L�X8g�"��b�����H�������mC��̪�Ě��o���"$O�֛L h��yR]`d/��U���8�W�)5_
�9y|���Ĩ��$��8��P�z����}2gt�sٵ$�&���=$f��aO��M�WJr�A�"���c����`0�ˋ#y��L7��\��ٴ��3ołEZ�ab�;Z`��dƦ��NR� �d:Q�����l*������/�����G���Ç����Q=E��&h�þ^l0P�ޥ�Y!�'�o9��:_(��n��@L�p���t�+�OOsZW�?<�+�������J3ť�����c��r4�	�?;�����<�hͬ� A��/_Q�R�C"z�Gc��-E����{ �<�~��g����rusG� su����ghR+恆ֶn�������5p�V0�sn�%c�{���V�̠ˁxY�(�洳@E% )M/ �H�����J���%��Y���`���|����鉞^+�����Bp����Z�7p�è��Tף�d"�g�D>��/	���:����87 �?|5J�z�V��3�;����%�^�Ғb������>M����K����?�|a~�B�u�O�é�1=��0g"�����P�66o�5�����5I�%�M.LJ�	{)���؆U�S�`T��>��P̗�ց��I�9Z_i�Ö�)Q�.�E�s�:�+���+�SA���v���9�w�W8��Re�ִ�h�dm��==K�R�v�3�?XG7��@"�u��L�u�"I�R��܏ DX��2`��v�؆b��F��?r����[:�A�	|�r�upQ�'Pl*�xV�YZڂ�j�r�Y�0Y'�_�%������y��D�\l�#�C�ܰ�v.�z+?��N֨������y� �t�x��7i��	ݵ\ad�(�*i���p���U"���ۨ �fۥ��HX��lױ����H����>�[�%L����:"�0�i���Q~�y�BX�zgO��Փ�UY�e@2���pvrB�1��;Ȇ� �dܗ��Zzے:&��FB���]X[�_��t�������}��N�:���Eń������%_+J}b�M�_./N���X�m�-U��d�����g���:ٮ$���Ú�)#;��_ؠ9E�-�niNۗ��9�'��/�n�s��D�9�x޳άR�Ңn���&兓���Ab�*��Hm�ܴ\��_����D������_�_��|��9]���%5%�œ|���!_3%
�rtr��X�L��Ρ����شX��C��׍�CVT����(��IǴW��庺���z-��?���v���Bd�����a�5:�� Z��O�~��F�2H������8P01R�3�.d�>�z3Y�f�����OT/��<ȿ��������<�"u��% �5�W����`����o�&l-O��cZPo����-"�M��6(}���m��T(`�e�@HyӛP	����U�ޫ��� �ǇG=�����^(�7W{0���]l����jS�ʸ��3(K��?��~��9+2�\ceX��1IS۵9$#��>��������!�j��W����b+��{큯�k�������`��1������a������6��"������בޑ�c�7h��,��3����A��¼F_a:���C�r�ә�C�[c�o#��ګ�Y�A���'���ދ�Ã�߽�%9S��-��FZF�(����h(�T_��Z�@R+��%�jb�:o�� t�2�K��z���qS���{�����޾�Y?�Rۮ��E��|Q��TJ�����(�x����ש�M;S٦�F���U�|QSU�ߩP���\^�t-�s��^���w{z���@v{�7�4��Yg�ҵ���Q��]��e�#�>J��lZ����B^�y'?��ш����%,ָ�#��"i^a�N�⚹�N�4u�;��4����uk�1V˭o�K�.�"
��8qc�\��ŉ�4Fb�*� �^5�yk��L.]��Br���&��Y(�����۠���~�,�e��,����ȼL"�#{>��9�z0�G������m!8Y�t
3��ʴ��P���4W����8�����'*;$Ƭ��<s~O�L��M�-،��e��櫵���4Ax���l$� �1�Q1�{ t�F�`\NN�>�H��f?/���g�@�(�{��)�/MT�X��]���͵�~�����i��9W;(���%�_2ewz4e�B�[��6[�����3�ф��`�a��b�`��/�� ���(tE;��F7 �o�gSn �bV��ooi��Ï?3=}��+ÀǶ�nXI�J��Y�3�[�o�k�Tp@��!{G-Gf��`�1�3�4-������\Y�bq�ޯ���+��}���'�!D�=�{:�M[����)7�������H��=S��GC� DHq�ok�m�
��(������������C���x�3s�޾�ׯ��N�$���A�U�om�&�n�c8gg���^}iZXGN�b�S4��Rt��t��;��^ӂ��Hf�@i����R��:t����~����/�_�~?�1p������c�3M��z*J)B#éiԺV��d��1� ����|(@�y��%����,T��۵��Kc���tЂ�z�歎�\�q*S�IԜ�+�^��UٓDO���w�2%�^�c����"р.%(� �5ւ����I����aQ�1���ּhZ�'�����{�s��ƈI�Z�"� ��xVM%�?��S0Rw�#�p[�H�\��R�h��+K�ʻ�m���Gb嚶x�xR֬�:�o&rtvN#K8 7�4����Ԟ"�>�D�g�v|��'��
BV�ׁ� �q��7����7��A7�2(h)��\��lt����[�XCmR���yy�%�����ȸ���܄�p�*᯴���W~Y�PW|�5�5��6�5����zRш�f�\<
����P�Q�����~|r��&̼�֮a�SkG���6I[�(��)b�}���[�c,%� �]e�(7����W�^��퀯�W���T�kȬz�g�pU҂ӯF�Ubj�Adz�#�x5�����߿��׷a��\=׌͵�� �K��(f@��̘�m����i������~���$;�nzu~`.�ӡ���1��K�߁ئ���j�G<��D�0x-=�0��X�AfՂ `�+��Cm�M �����]p,e��e�Jl�S?Y��=]gi�ϚUۈ�i���rg)]`�a��ݽ~<Ăy.��o(������9.��zyZ�� ����gK���+^���!�E�i8�T��(��O�.�뜩P�`��Vv_���8�K#z�zՔ��2v�Ґ��-�%�	��x��y v��>�1k����t����@�a�����p_�*�bE����_T�bl.W�[2�- 4���4�I�&�g�]�X���7O�������?O�>���&�c��z�뾃YJ#�4FP�.�XѺj���L�!`�>�a�����!����:�>�>WAy���h�j{ٞ�:�$0�ڸIp�}�JIL�J�QֱyN�	��=���-F&���{�c�\ż�t��l���sNm�J�4�t�Ρ����O��_����<�����2[�X�v%�-H�`����f$MO�<z"���Z�mh\� �֘�V�SFf��J[ն�+�k�C���c��H쒊Umbt�L�m֭o#��g�tMÛ/�>�ѣVW9�H6Qt�l^"�^2�uMQ�_����A�M�E�lQ�Y?E�$�\Ϣ7�QLED�B���T�;�ǫ���B>�����7˄�4�E~�1\��~��凟���|'�w����b` :����}�Z�5+M�N�.ܟ%�MpQ�>�4P���h�$�k�*7y�nft4<��q�kk]��}���i(l � �`��	гH�.�D;�0L8V����燴%&��.X
m�����ca�Aϲ�X��TWG�G0�[��"������C������Z;���m#a~��u��mt����vG��\���Pb��LA՜��`G� l��T��
�N\'�
o޼��zG��D�.w�����3�h��R7u�Q܁1K�Tx̡U���A?�1(Z|@�]tdN�r�M�_��q�%ǝE]����Iw�xx�(z�9�E�)4d�*�i0M�tX�*�\�������5��8b�2��3R0yҳ
��4C*#7�:��d���"�d�R���Y3x�M���s��7V�G}_f�D�i<T~rt߳-��Z�?���9�:���m�1eX���`)�mI����?6�a���ζ6�
L;8ܡ?C�'��+���%���]�@p��d�Ц�p���EE�2�|��@Զ��\v`��u�Mu�����~�ػ�p7��R���Kl�2u�[L�^�l��	q�{\s�M/Y�-sW��4#�Xv�CM����I`���I��>���,�!�j��^�q�~�װ\���_�7��s@`�N:)i��t7���I���Ys\<w����9n1VйbM-p�ӳS9ӏ�x��}0`�g��L�®*�n������N�:���c����x2��c���x�Eo+���!�sc��_\H@��x*�ф�Q	��Eb{n�j�A����~d�@@P_ν6z�kщ8�4�sb��~J�w���V��7g�@"�j�1p�� ad�K΋^��[���/ "���&�yE椶���`lʍ)b�3�pn=�(�A�Ҧ}2� *K��h`%�0�2�n��$�RhM�cm�X���>q�B`S����@C�=�X��f�$e|SNa���G���7�ۏo�i�ש�I(�z�c���:�ɄA����Z�9o�.p��\��y�� #@ܿ� ��A�ɪQnZݾ͸��W�(I��upG�K�^7h������|T[ �)K�BY�1�BщR?�l��f���H^�s�0y�l~[��``"�T�c<7wY�&�\3c4(�������h-8���#�j�]N��Zg�k�k�(Pw�:�h6(˚h��HyFv/�pN�়�-��B?*�߱) /���c����|U���S�PF?��M&=173����ez� ��Q����\3B���+4�E��,!�k�Hܲ�3Z��X�%�GO���6���U^��	���"Xf�1��2����:��|�W��5��zc������?n��������|��o��Oɮ���3Ʋrs}%�٭�g�0n X�Ig�N�+��6��cu`ύ�7kL�xFkT^��"_ަsi`1��)+\n#]�����8�k�5��И|b���h8�4�3���+������~���5v)E�y�Vw��*�u��h̛sh6
�rn��h��F�	�c�2��`���:P�_�p��=D� +4@�l��5��kR�W׷rssOF�X��:e@�*IL�J����}n�Q�/��T��
�+m*�=�5o1�S��7l��*F_��ZR�^zG����^<Ѭ1�Ҳ_{|}N������|�X�b��A�!�׏��æ}JWv���55�YZ���z�/���D{%=ؗ�f�O�밂�ڏ������o��ﾑ)�O��$z�n�i��>�1\�Z��4�G?��ݭl�%] `��?���H?��7y��'ZUP������;m�ȸ}�5�����!�źEY����eű��!�l����/H��c���k2K#�j��6 X$x�@l���\vC�Q�/^��T9��0� ^�Z*�(�n1��6#U�`6�\��eyCf��U�7f�|�9XT��X���Kc2������f�'�3m���j4v%�*���>bV!�^-��]<͑�1��47f�����.�ְб
�"����i%?�������凟o�Z��z�* �@sNi�&
VAqn�&�Bo�'�4��K��n��ײXΉ�=6��P�>��ܫ�)ٌ�bVq��&e��J�n���B2|�D�ٷ�8�"Pl�,�o����7}g���C�f��L�3F��K��a`\��0�q�u�hag�>�MHo^^v찷�4C��|u�6]W^c3��2��+w�&l���N_:V(Fg�<�q�`I1�mfV	miW�{�TT���T�>�L�����m�h[ɓn��͖�
����l�x��W�ZM3�6+���g�L���gHKCl�h�M}����>Z_h����ġ#����Uy�Z�ta�q�湾(a��9����s�櫗r|tn�?^��Xe�W�s{,�ŝ<T���;#mJ%�EN���y8@aBV;(6q��G��(g�D6)@0�^�6' "�U�7 ����##`CvK�V�㡋̓�*ۺ-7d�r��ܫذ�(X��hЧ�F�ͥLȚ'F��8����딦�ڞ������ߓ���x� $�Իm�gV�A  �v�6�\w�LZ�۬L#T0�ȼX�ұ� ��0&f���N��z�����#���Z��ǐ��,->�C���H80��LM���@��W����?��R���Jk�G_�f����Yf~��+��l��ƚ�l�䕹:�����(Zp%������]�^Z�*�'G4�'�V[V�4h��[�Y��䛯_�r?�Z�򌙮�+�M�|й�=h4��~	5�}�8NBY�6+��T3��
Y�Mk2$e��Bd���1k�>�$p�f�e�[��w����!d�[ڱ��)3��?�J�W�q�^ڱ�:=:���b�*��K(К#�@���A�g m��Mq�F����$$���m;�2�ظ���33V�D$h�|�t��t=.��3E�6�up�-�\���i�,n2{8�Ji��������?���W0&�Dr\`��lH 6��=�� _XLR�n�ۈ�F�`���eT�*�;[5�Yy��42]s�!��$ӣz�<�ߙ�73�8� �E���� ��h�R��aԠE�n{`}5-*�U֕/�� <q��՚)~@�1/hgD�Eɨ�@�9@�ɍ-3�5�(8-%Gt�����òQ��a1z4���)*�<���/W_��oS	�9�D�}�ʁ�V����8�9��pO�W'>ؠm@)}n��93��+��X���n�9��#��V���c���]�N��9�|0nouCDsw릷3�AI#�-L�v �m6�׺�Uݹ9E��fɈ�PP�j�zk˩�<6��d@�	��N�z �.��pn�>颊��2u���ݧ����mN`�0�����2��= <���^���uNnhb:� ��m��[�cHi ����e0��,�؟��`��0%�Up�1�A�x�1U�n�`}5ǰy��Cի�W>dLu�n..��K�(RU�~)��ާk
��XM�6?��<.t����(XeE�z�X�]]���������8a���! -�=�c!�ϑ̭Mp�=8��2S��k'�SD�`�,��k�X6�Px�M8VGk�4Esn8���>���<��}`pFmKH ��U�K������}/�7�ƚ8��1���;lN
 $��n4��eƮ��Sb�C�O�ާ�\��������)�j���g����c;3XG�mf��E]���~9�?9>�:O?0}!����� b�޽�8c���-�z��d
u�x?T�[�-	dz���L������{Tp�^b�"�����oo����򕮥z g�k<2���,���)��0��`�}����ڎ6��w���e�Rp�T�6vX]+�(��X��7�6m�J�Xద�
�yaB�%��Р ��Ԡ	��#k�6��}��Z�^�FG������$�n~O�R��`�����LT��֏j�R ���g�l�>�
�Q�&ɹ�63�p0�R��֊��^i ��{�՛w��׿�(�፼�~�:I�GzL ��G�`��L7�MU�[�Q��HSY
o8a��:��Hs����x�s�����6���s2���͗���i,�)~��+9^���w�X������|��'g�6[~��.02�8҉F@�5�>Q�Pyj�}�E��VӰ�~��q�Jl��<cXbAgO'6?I`�YN[z&��5Գ�1H#o�^�o�Ф��:N�4�����c��h����j] 董�>��h�go2`L��ٚ6����x�,��Eʀ����2]�H��!L;9��c$S��#�I�LU}�'6P�CWs.���4�*�=�.vև������SЫ��|=?o|_�=n5�/�QL����y�� l(�⽶,�ؖH�>��݈��K��c���L;�y�������;�WR�QG2G�7�L��{�}c�Q_e��+��I�x��`�,=W��&�G>�X�K}f���y*>R���u	�a��k�\�)�0�&�]��G�T�����tv�m�o�,��
��@@hcNώ^�͇���O�{��|�v&�'�d�!�/k(Q��e�Ҏ���+�w���\82k��[���� �<�#��EFݫ�T<�V=K�, ��z�B�SL������} ��u�����fh�Mߝ��|�MZ/�������J7�cӟz�e�Z� ��v�[���� ��{�_��b���J?~��)�ءs邸�hţe	d�kn�3`�����[���w��B�=q��'W��t��{ ®���^\n��>��б^��bVV�c��`�������=#��B���>�|����u�����6�-�n��h08֯�\(h;B��^�L"*�+(X�6k��:Y|7�jĭ�-�3]ݴ�ݼ�b��:/�g*�w�MK�`Ȯ�ʊt�
�@t��ߌ:̻�G�K��gR���d���V����g�$��.�Ck��d����	i 4��p�����ˢ�/D�3���""��W�V_�F�b��I��l7����6k�́:UG�2�Vo?������*��\��|ôc��K��F����|��`�#g�;�K�{l�vb��)�>�`P( 8:;���F��mz`d��13ɑ��j'�_���iʯ�>������.�+�o����7�h/i�&۬0�h�)G0��%�
vp�ɋg���7��~������������00 �B�R��b�M
3�����ф��֙��,�F�!؆dƣF�g�
ΫS[��6�X���΢��؄���)H�rK���M,�
��E#y�����?Q�W� �w�����N�*Y�+S�h����u)��A���C�|%�
���� ϟ�^#�s9��F�����1޷8aԇVz�����j�������1ǰ��#�P��$���lsݬ�����GY�8�|���(�#0R�DFc��\M'hw�gza]<�Pn�8�^�2���H�?�޴9�$����߼g�ut��֊�~؝���?`E�{����ʬ�8��M:��f��� �#�{d7JXI:���T�����]�	����ޡ�|��C����%�Qv�t���Vz�%�]���Vϣ>��{v [V]����eA�H9�н�8�'�������Ȫo��M�իSfhVI��4���'���B~~�A~ֳ�y踾 ������4��9[���_�)X��؏)Y�"�3h���V�ľ@'$-Nt����a�(�/2cw7���[�9pZ*t��>k�=����C��x~9v�&>G�m�AHP���&�E��
�V����ֈ)�<N}�9'����$��`�L;��9������S�Sk5X���\�5M������7��� ��ݖV66ӓ�b�{4�ܾ\��C}�@f���������w&��;�1�iu��);�ɀ�{�/�)�R��������;#k�F��Ȝ���(������B\�k�m-ߓ�S��c�'�[�#�./.�??�ȳ����p|�|q,{�����a�Y�=;��F�)*�1��37ﯺ����������t�R��v���I����ʻw���������ՑTG+&g�:�n���tnmZF�M{�Ԝ�'�D׾ӓj�}�{���%�e�,@�&�l�N{�]<��[kBR,�&����KJ�<�3�(ͭ	�Qץ��6BQ�>�u>�Դ-�4UtM�:v�R�VJ!N���H.����%��n-�Xb��H�J�L��*"B�օ�Ǒ�xk]����խ|8�����A~��\ܪ���+Wt;'�'�\q�4~L+�c��e��x_�v-�o��M�lsp0�p�H�r6 u�Z�s@Riv�K̼@��C{�>��:�Z����H��߳�18����3[�dXIrG�i�+:
S'��FЄM,��iY�a�N�"��k��
�6.��(٬�s�J˵wC�Ͳ1�]��o�1tRZ�#�(��q2٦�eO%S��"���M�O������Y�:���L4��n=���2&��.��IE`ղ��R��S��b�2(�m��z�>����9��~w����0nB���?p/.�B~Po�$�X6N�çKV1��a}��.m���^�����lcz��Z�0xD��E�ٗ(�^�\��85]��y��P8q��ް������������͍�ݎ���OS0��P��a�ǵd�k�P�~
 ��aD��AY��0�k�BTy�����=aOràh����z���j%�z��ܤH����f3m8s�s�Q�"Y H`O�F�2��"�ɑ�b�,��Sc_�������'�wǬ�5(�l]��Y">�F: �R#0�3ܢ�X5gW6���E�9�Q&୳mğ!���]0�m/���&��@8]6`�&��J�v%P򾺑����B	���s0;#���(���4�������+d��@�x�R����`����dүd��<�b��C~^���b|y�����[�ɡ`�Kl|���x�b��r��7v��I�=9a���Kt�Oc��	{`�w[��hA�B���&,^[����\r���l>����ѭ�tOA�7�?h@����#��5�2�{�������)���[�=�WYm�)Zs���t�\KI�*���E��4ϺACL���w.�q��|�T�:d����g�r�|�t���L�,��_k���D��ř�h�󴾧�*EU�*��u@Q3�0B�+'���������7WG����?��,�_)�p�І����6tjgTU�{&E��U���md�Mk�ǃw�ǉ��g�/姿���ߟ��Ory��!Ҝ�6�%#�x\�t�Oͯz���f>�5�yd �/2h��!�%AHmZ9 4���L-�2`��h_o,�mF�r�א��\�x?��^�|E����)���$������c�.x#��2W��..|���g�_\���\������@f7�ө��b3Z��'�b�RB	ød;�C��A�bb~��ljc ��/��w�v�k!����iREY:2��׍�Gz�p�_�'�$��y����Vv�]����nV�*І���W�����]��Ɯ\��G��EWQ]��.T׽\]|��͖�>t�^]^Pc���L�U��ҳ���o\� ����]��lfA�r�Pۦ��&�ֽ颋C���%�h���*�CZ:�c�����QV��(�a����Z�x/7Z�kZ͠�RNO_���-��0��C����H��
_Wj8��A��AY6�o����C(Vruu�n�f=�b'�7Jp�\�����%SĿȴ�=��(_����dCAϴ��}��������?78F��C���Z4��{�M-�;�n�2�}^��3�l٭Ͼ�1a� �www\��]O������%�C�?�}��z{�0����ۗJ��SW˶��|��W{��0��̎4���l|�W��m'���Q�b�&@*��T�n�����!�����?��7ݯ�smѥ��g{���A�+ų�\�* ̾��á�?���yy� l���\�ɗ&�� [��9\ϊ�~��Q����-��}�s�7���_�$�D�����tsM�1c��o�|u�l� Ӵ�~�3���y����	����})�^�b@��#��-�c2�4�Ԝ��� I��>J���N���@�^�#SX���@�_3��Q>~�$G{39=��������B�z>w<a���芮��l6��$��P2�/ɢ�_�{	1�_��"E�J�dW2��g�X?QBg�ϛ/[�HIA�_t6��6h�ި�z��1�2���m�tf�� Ktʦ�G�I��D�r�`�r�îT���K�C#�ñ��p�+X�U��݀ړG��R{����lG�h2<������ry� �
�r��Ԅ ����Ժ��B�s��]�{V.��AC|��!��1!�n%����� #q�!��p8�>�� �Ĵ%�\�	�tv��|���6"����V$u����"���yD8NjF���?��=<2k��z2�1Q⼼����k�-�����:�=c9덵�G��5� 3�ED:�s�";p(��*Xw֦�!�)uaTܐ:�p �]#WȄ|a�3n>�X�E�[��5K>���	KK���h�{};`��lQ��Ǐ,��8� �5A�I��ނj��_�b�IF��jҎ�hz7�8B���є��*O!�f�������L������<m�FV�'3�����y%���Ɓ�$&*Xc�F��2=�hM��3L��~8��e�+����hc�;J�W7��pwK�|�0 J���}��~�x�i/3�C����O����8��YZ�>���v��.n�:��O�5fJ6~.��W3�?�`����l�刮Y�`�Z9 0i�ֳ�/f]d��E�0��vq����;��c�-��ڶ4����#�V{4�ؿ�5�x�=�pKE�FR��!�fe��ݕ8PE�bR>��C��mdC���u;����*2��+��u�|ڞ�8	��Ec��
{'2�8��$�|P����$;��<:Ҽ.��?���g"�jLa��pK1I#��5N� ���u�q?ջ�,���"R���b��JL�z�y8��N㦁�o9˨e�_�gU��d3mj��*�Ũ�������4��b�F4P��@or�(X	�1_6�4�P�e��|8����#�GlHe���O��w��޸8�u����y��6Q[�|�����G�Yo��nRO��5g%S�N�r�-HJϞ�=��t��Z���^>�3~Z�Ӓ0��QZ��'�Gm����h���	(��A����p^���<���Н�"��=���4%)�ƽ��Ew���&��,��,(��^�❛�Z�rR{�1JB}6�}�EU{���Z}�����Y�T�����;}pP�V��[�g�\9M��bJeG �����h���~x(i0���>m{?�3@��Yh蔚( ���Y0T���/Z}���S:��|1�w��Ã�i���V�Ł0�ŧK�ޟ����]4�a����׷alj�g��<(en7&��_��b�:�5f��.��Iؐ����K���b��D����ϱ ��JN���	��ۼa�3�H
��P������Gg(�.L7%����1C�j�
�jyITf�����w�r;�E��S�A�M�f�n�*�7�B%�;��Z.���7o�p���į�_s_�Hf�i��r�{��R���=�'4�P`X������6I�F�bڸc�Yj���I�쐋�G	/���C�Jw���u� WA2��g�5t��+�V}�X#tv�Ė|O�ؽ�0��=n�����iK�(���?P�F�d����u��6H����0��(л��3����U�;+���(����|Hc�,����I�͆ F�W��r�ױ"�2���-m+���g��;�	�g�IX�O�Yk~��y|lY�@V�/p4Ƞ�*|+���X���+��K!���A���e�x�v����H\�W�:P��d�~6]�s�P��u"����Q}c����]�,Ye�m)3[|j�q�Y`���z_�z-Vs�7�.>��۰s����|\
ff{Od\`$����O*c����2�[`�f������_�0��Up�$[uC7VN-�U	��J�@�3��Adg5�sY�~ �����V�9�O6�9��n5�@*�0*�u2�9�J'v<�Γ�d�Zf��r���q�M�Ѿ"�Ğ0`+3G�A�Mi��+�	��빂�1��D����P7 �>��Y�bT�6�sE�}F���?�4'*cW��}�E�{�j�){b���\4z �"΁-�b�2�l�<���Lc��Wb��6=�D�=mF-����,â�'ц�d
{�m�`���Р\�`T���o�4����L/�5z|�L&�,��h�K��7md�:�،��G��h]nK����4r'�ۈ'zf+�< �;6	P22@7�䮮��^���u�/a0r�<DU1K��k��Y% S�U)0A��ZY}DƋꍃ��䀚�eJ彾{P�z$��ו�X�j�����c�zqʲ"���Xk�>Q��LW�;.�6 7�/���9&#%�qww�����:��sQx�՝�=>���[[;�L�<Q�cv|�'�S�t@�����t��&9<>b֠ser�y��3/u}��R�%-5� Ѓ�J _���+<��C9R�2o��`�?!0�b����l.[z�y��\�5���|*�DU^Idks������ze���D1._]R�ɻ^b_'
�z��)
���L����[p-�5J%����B���K� E�]�i�,���2~��yS+q^�D,�gnXRd�9��?���(��\UR$�¹�r���}L{����rA�`<��B�� ��SE�8$.�0@�	�����Xd����:�Ѵ��`���l�u�t s��R���{J��y���g��n�O3) d��]�V�1�@V�-����~�⡭�r�z���6.���ͦm]��
�����}]���SCN&��ѐ�ܵE��ߟ���Z�#�)(�QS	��ʉj,�Wb9���W������B	c�z_[�!\ݘ���9�<GPtI�=&�ףy����*~�X&� ˷Y3��`�4W�dUS��t~_سp�U�g ?�����.�M;6[�w|�2@eȓ$o�3�e�2�X�ShN9:�B����o���w��|�g�����8��h=
�J��?y �_ˮ23%��+��u/��>�a�sSY%g�<O�?����u�!���L<@ܜY/K�`o�:�um;ʦ�� 4�h-h� � �-Xg>��{d缿����֒6ȞB�)�xi��q�j��	J%�a�q��_�U�͚���ΐ�5 V�<y�3��K�g)#p�Pρ;�LYIȅ;l���	&�ؘ�X�C@���.����O�uo��X�Z�u����=�
�v�����Z���L��?7`mj��(�`���=�ͅ;�Q����+���պnXdK�5kF�v�o(�RcU��E�k�o��+֚����5�3�U��@����7u���8ܨ�1ː������|:���o^�����Vx�;�����~�h��Z�g�7�����/�<�C�1���gF��~t�_ɇ��3�R�>���; ��Ս�z�F^�yKeuf����iG�_U�JG����͑	`vYs����/XJ@v��~-���䧏r���ig]�(��	����������?���s��S�̿��{9z�V�å<��|b�n&����(o�!��W&�/�%y9��CY9����ZD׺֐Z��@{�d�\��S��x4�[lk�O�N?��� s=���ތ�;�.F,6�7#��}.�j����xf>��s¦sFy��d�-Q��zsK��_dW�X�R���ceoe�ˤ`J�ƿ���\\�%tt���͖���V޼xA��������'�q8v0h;'4e�܊���Ą�6�g����棕��At~8� �[�6�
R����{u6ۓ��Cyyz��`���V0�a!�ۆkC����3�����x���о�5������{^ʚ���*Ŏٞ^\i���{�W+y�V�ro^��o�{-G�{��*��t��ٶ��Y>|:���I>�_0�j  	�S�mR�Ӧ#ײw���نi�b�x�Y��^o��h��]��Vm��͝:Í�ksn̾ѹ&��昤	�zs�B�HA�����{�5T��gtu}-�
�+ځ"K����h ��k�7۸,�}O63˹�E�vw��z��3���>X7r�"��M�%�����;aF��`ƙ�Di�?4_�,;d(C�6%*�]���P�V#��R�gR��"��/�}�"�1D�E� .>�@�:d����XXM��f��A��U�>��YIE�;�6#��ȴ�Y|H���֟��joDr��T\ s���^����-9��*Ҏ-�F���� >%��Y06�d�@-�/��� ��L�S:�Zڪ�����a� ��������B�wv{��gU�l��b�p����]�7�ȷ��+�+V�T4���P�VQ�a��+�0�h�����B�����l���v��lQ��;�}^��� �Gڟ�7���"6 f$��y��:pKe������1�l�YYl��#���У��&s��:6?�4Z�|��n�+��c�0�����n-���T	��7�R�e��}�w �}�[Y,��޲� ����C��@�䣂HfoL�c�$��\�����T3���:ɯ��%;���{y��a�U�{f�v �u*�7S��l�#�Х�X�1k��ù�]\��̓|��'�܀A�D [����\(����^�u���g�O_����R�{-SdU�bώ[+�0Q��gcH!�&����	���)�
CZ��o�$B&�>x�[/���wQ¶��FQ3��[��[,OoFF�N�O��1�i�Hh�X���b��ui+4����������	e�4�A���G�(��yA�}h|�q�7�A�E|ٗ��-d����y��F��p�����y����߄��Y��P�3UM ��pK
W�m��8��1mA�)��s1��2a�=�cF��+�mY2dM�Y��+nW�:�~�tآλl�	��Vi>�9y�{�"#v�����h%ݛ�J��UV����!�A��A���}s���[�7ֻ�G����X^�<a�wp��g8<\f�]�~��;rZP���R�į�|�$"��g���~��<) i��%�N��Y+0ZSF��s�g��8L�'g@$��e/��8ՠ!�r�@k����{���?R��t����х��Ρ�\@QGv~A�F�>��pceD�h`S�M��$�e;C�e���|�3�4���I���#%�i�������u��Pmp�DLw׍��ʥ��4㛺:�Ձbi8��%G���GCYL�L���3_�{����w�'�~Qc~��Z%)�-9I�}̚?Zt������hPCW�N}ޥ�ip��+��ۣ��Wo^�k��U\{�A�uV$X��rd��8c�Vf~���o���̖\x�? �?�~�rJELy��.9��H�����##�3�u��/�Cqr�X��1�J� �O H��Yֵ�,��̽�鶀�\�4��	���M���Wj�k��ᐞԐQ3���m��OO�F�B��r�@=�l��L��k�i��[Ě��i�J��΢7�uh��n{��䒪��_f�d��#���֜s�N?d��=����ˑ��B'7s�T��1��� �z"�p�48�>����|>{���W�3W�~מ���;9}��Y��w-��x,�zK0�bCM3;t6*Fj)�J?�!\��l��^��D;����rr|hF4[DVG�tL6�Cھ46����N���O�_�ۿ�GtR�[�` 5�|
@�bT��Q�:X��k��hO��R��ե�N�e����L�	6 ���,&G2uǓ�"�O�E-�	�Ȣ1 ׃�	�ˋ�Cy�շ��?Pg�熦���#=Sr��4e�Jπ�#~�CĞ�<m-��ܫ�����&�P�	/�Yp/�@10HL�[%+�"K�I�����͐4,Uܯ7>:9�m�@�}��w�\��ߨ�bc�_z�w3�0Ϻ�R~7��u��-�����V
��ܰF��LXzĿ�5�轁��z@\1yWKd^ʾ>g�eف�X��cKy�F�������#Jh-�0��Z��/�,��Z+%Z��x���gyr|�_{�ʅOʖ��߱~�����sN⻈B�t�/�3���N�z���g�tq�{�徲��ׂg���Y���C��o�>�3;' G��]_�u�A�)t�1+����6����V�!a�����M|:���qN$���Q��m~mN��]�=KM[}w�����W�{�|�tE���#m<�J�U����7j/~���rzth</�c��B��?�$�����{���󕕳����̠Q��qM^0�A/�"�� �xC�ǭ��2��I�t���SG��Zj�j{p���\P�WdPЭُ�|�geY	i���c��?�Ӗ	���!���l��:@�]v�z�.;�k��^%�`�@�2=�`�O��EA��(���t�ӷ\��D�<8�����e�����rd�Ý��K �vͬ#�#8��Y�޸�'i�i���Zm��<��	o����$�뺽~�J���?�����k����܅�D�I�E��Q؈�5h*��U`}���/�I�[o���//�l]ܐ�&2e�)�CP���2���~=$�f�o�1:!^.�?�� g��&K��Vm��70?��=��+f�A3�&�H�E�e��t�XMb�kH�2�VP��{Bv���e�4��(]��:JAPr��d�4)%=�uéA���� L�[�oP. �r�p �s�(�M�ly�Xՠ��9t���"�)	����b%���罗%j	�����SΟ�]8s50�w�\���XVP�� ��9�Bgr��&ƌXs.��{����j����������3	��k�m�d�%�s���&�a�n�q�w+����Vrtn!3s����j-?����?�(�w2Y��Z*;=pB���m�lz*�rȸ<�Y�CIL��w��h�l6`��- o�%�����g ﲗO�2!��^�N��i��ғ��8�5ӿ/n��\�`�)�vO�/�o���K5*;w򦟶se�����-�a>����@!���'>0��N'�N�l%:��
 �i��. ������꺟�qB&�8���,|׍��[�X�0Iɻ�|$F��?x9Y�/���qc�C9�i�Y�X7H8WdJQ��@���4�]�� ���D^���M�1
���*g�a�����)�0"=:�&
�~ 'j�4\|����-'C��I��wC��v}���w�<��][�$:=Sr���m���\��O��3�tqɬ�g�4��
�v>~$��\�f������٧sF� �W�r���_h�9���}>n��s� �أu��ڐpd����YS(��2����G�I���[��<�
qNz��*�(+b$x����f��T�.d0_�3�����Cva��q��S
p����?�E��mE�����fZ���1���c>7� :�l��.��l8�J�_}�V�����&���F����{ v�D��Z��N���.��iڴ�̄A�)P���G�ܬ�3�k�<��m�UE.��}�Kܟ1�r,2����qѷ�yŦf��������?��#�`l�e�z'Ʒ>��:�����=G�
�!��{ c����X���7P�E<Qi�P���g�&u [�I{��|��W��w���K��;�z��v��,J�,�dZ������߫O��r��ʒ��w�1�,�!���]9]P�A��	���`��.�(`j��DF �Y��Y�2|���H)C'�MO	9 zը�%�)�^&�B���ՐW�F�KzP��7h��ŀ��"��/6!��Q��@�F^_�w��
��Ƚ+boR"t)7$��%H���c?c%MO�z
и=N���1��d�Y,|?���N�̈́������=y)���]�(�J|
��@�c'��I��C��������ӿ
{�E����W��?��wj�N��!E;��.�ͺ�;S�ǵ�v����_�;��!��I#���7H��b k='�q���e23��贫��>�zb��\�����՝|�t!?��3�3��?kds~q�r���E���Ȭ��?f<�aУ �v���Q�:P����D���T�e�9C6������c��̮H�=�eI��f����
r6�<덥�1g�%�����|ˬ֭Fk+L^�qE��kk�HV��~Z.��͛��������ZJؼ�����8:y%��!`�A��gѶ���Ϻ�Oz��M�cN��S+
R�Q�왡��
��*ٯ����y�^�e���y[�RȖO��㹮����	2�N�kP.�jo6Orsw-��\Q
���F4��fWfN��tu�#��LC�V�-g�]h����j��/o�L��#���(K��_�C��/./�`_l��s�Ё�o���,��gj�z����끙G<��cȹ��'f5@8�� ����r�������y� �hz���6�q߱��ӧ�ޯ_q�e�l<d�\`72��sTAw8���Y���325�3`j7𽋛{څ�A0J���1���;�[��l��Qk?�� gh E��_��]k�W��:����-aC�1GY٥�vE3 zO�f'4F����}��C���I�ɻ>���xl9��!�I#n��H�|��������q  �G���1�4�[��"� $]G~߻w�������U��U��؇��{�$���ފt���C�<�mu�7�@��U)��-����b��ْ�0{�DJ.��Y06{T������۷o�����Y���Y+�G�A*���>��>����z��}��A��L{r�@�FW�cs� 	��k\�V;S�4  ��IDAT��H.�čS�l8�W�7���rS�c�����|L�g��i�� .8���6�_��r(+ڴ��ĚYhr�s�F��%q�k^|����ʑ>qh����Z����I���,~ϙ��.s��$�B�lk`!�&�I�o�N@~u���Ԁ�pɬ����JWq��4�e0���1��������e�����R @���yf&R����2�/�˒"{-��ߧ��6ݚH4�lElv��j\�U���������� %�e�l6R�(�6���g�U��ԸA�q���`5��I3]����2�*����Hj]"�%��g�h1��F��V�u�̑���L(�-X/�^Ûs�v��a�sC�s�~�)�>[O+8;�<>|���~>ӈ���m(��9TP��� �����-2S���P�����������98>!�F$�Bs��Xl/+Ӿ �\�o��h �(�!���T󇰫��=�m��e1@�_�(�Z�С����Y�Ƹ�]K#��!����08ƉD�1��U�t�,�d�2-ϑ5S+)� ˵��¡�-t� �x֐ݺ���.C��ь���Ip<N�����[c��ҮΒ7�Ig�g\z�o��&o�^��A���Xt�!v��� R �K�O{���<cY؝�j>+s.p��W�)�@��{��ʕ~�v�T��:g�g!��e- �������@����o`(5��hԭ�ussM"?���X�C��A
�������Z�+&�,� PRY�H��
20��"�c�D�.1K���s#w�Y�˚��5A���?2�&O����XU{��Y����ݝe��Qk�*��Tq-%�>^���@�+[f�w4�u�2��tО�i�q+w346혭Y��Q́D��i����II �E�J�<b�rU5�V��
�H��bE�'gn��&����F���� o�z��A�
wl�  ���xd���g�Q^_
���!� ��1��xF�kǆ����z���~J�q��X'p V�����Y�Dd�h���F&�Q3�9�
r�gAѯ�����=�Q�)�\p�2�](���L��W�?_�&�U�b�o��1!F`�����@���ҽQiA�jkõ�!�ӵ�������@6i�H;�c����,���
"?gL�G��A^���Y��b ���T|/����l�s��e����LA�Ϟ#2 _y#S 0V�j��Z�ҡB̲B3v���������!m���eu-ڸ3U�{v-$AD8�K�u˿#��+6���_���!cZ&K�e�|P���Q�eI��G,@�0Ĉh�&H���K��л8\��z�4�9G��E
\,{D���2Ї�޲���ͺ��v-�|ƈ��F��_���{�5�%�Q��(./���3��B�'�ә��ʞ�����`)a�zg�zt~������b5�5�����4��<���/�������Y>k��2�#��ɞ�0��\��ɣB�|�Wi'���5M�Ȏ�^�.p�`D��}���rt��D�v{�&k��$)���Ue����7�%�^I�|ʵ���d�#d"rg<a�;i�HZ�C#���D�C��D~d�66?jJ]V'@�8�|`\�:�������9 |�� ��|���� U�UG�Ӄ.,���}�W6gg�~�'�{T��L��2�'� ��%X�4��d���������.b� �xV F{�)�_K��9~�k������"8fh�-4p��5��/����|��^_�(�LDʽ�Ri����|x��c�z��{�H���C%l�2��ˠ ���,��\�W�6�~�g��\r)R�Y��.����.�u(~�8�`ɃY��]�o���PDӁ�����a�	�(@�K׋��lXr�`��_�I����ąg�jӌj< D��	D���	�6��[� �V���8!s��BZ�ٵK��+��ؙ�<��.ȌAE	����o���>��^�(��a� NЅ�F����33g��������g`�?BCQcY&ȧmY��	�VH�k1o�X���W�����r�⥂�f�p�S�5�R��+�5�����O�>��oR3 �wPj�xÌ�x���ٳ��������½�՛x����d��g��Q���]�;���S=h�Q�޺�w��(@
2J��C5�RL��F<Ѧ��b��5�����k1�d�jo��t>~��c'6?�ְb��b�\��b3�?3���o�i:Pb�ag�$�[AU�g�VG�G�䇿�U>|� ��(�p`|]�UN���$��"�Se����;����y���O�8|��^�\��$���V)��qp�R�|�,���Ff�5F\5dqM���"�n ��2�6vVf=�v�{Km#����<uO����`iP�V���"X�W|��L#�5a!�j�2��s�<��� 0��_%e�u�([�!���v����3�q�Kc��B�I���L���R��R�[���:�-9G'G���2 ָ ���[��{�e[9�-H}�� j��Ŗ<
�*�R+$� ί��M�{vR.�S�Wjt�Ր�h�L 0tI�%����B`� Bh;f�fE�U��YbP�e�H�/�W0.f�<P�����,�~�?~A�p��v�8"pw�ZD��\@y�(�㱪���#��[�G�}�%��ŁM�xY"1�, �32�q.�iA� ��lٞ�� �J=Mgّw�ޫ�������G�BϘ)Bfm�P vt�3s��Q<�;(���6�
f�n�B��1U�)����ڳ��хE�QɃ@ �#1���0����M�ٳ��]��ߣ<�k��S�Ĳ�ô�<�[2pB�@�Mh����;F������`�sc#�_\\�1��j4똤��οF6T�GL>G�����b]Q��1���kkX�X)�fd�BH��E���.�V�r�����hH�^�v���4�zv��CF.##j)$N��0b,3 "�2Y��A�${�Jܸwɍ��������]Mo���1��eV�-�}�O)�j)�Tbc�Lg� ��V%�w�S:�Ghw7Y�/?K���(�{;!� \�$1 vL�ު	t��� 3�g�C�瓣m"���G�aN.�	:��#��������%)���@�zK		�F�~r����L�7.8�ם��a�U����� r��f�{��*G
2N�SPv\ɝ﫟��RFB�� C��^����(��&{��pϳ�q?��BpD��}L�����󿼼� 2�*�v`S�,�V�Ha�~@�����҂8�ـ��T6� ��f.���)����Q�L�0���5�pWlZӞЎȚO�&�x�A^�#��\W~n�|0� �4a�+G� )�<p�y/��s@6�3g^��i���vh��m��&2;%�M@1����<��'*�7S���Z��	�[���v��Y[����HF��;���TY+t*�V6�e���n/WVΝ�J%S&nȫ�-Æ��GR��9�<,X
�W�Lʵ�i�ѿ��^�fg�GKVΥq�f��'	K���N�ν�J�X�:E�pk���i�>�A�6�ۋ!����q6��bT��3�9�Cd�(�f��&����uZp�0�hK&(�SΩ���L�6PO��ъ9h���r_�Y��b_�s] �Rʃ�#��9t�����TlĈm���6��:`��jt��#�\\��Y��gewt��` ��Q�Ӭ1���8ܼe�:��M�<7ſ����#��[+�nצ��Q55� H��k�Z�t��Z���#i�b	�l��:���/�R9�=���)�]�xWT��Yv2{��ДG28Dv�S�%��� �uZ���N��K9�_��F�b�2�dwX��y~�*�"�pO��!f�:�n :e�����(�>lk����EVn���;�Z�f�z�)[�];��D��\����Oȁz��qJK�6���k��ml����vq�Q�+U�i���s���~�&����9�EF'{@�K|�nY�����`���Δ�:�I��XU�泪�-h��$���]|B1�G��gg���t�P2��]%Hv�o׼^�i8��2�QO%#d�� ;A�ω���q^ٚ��71n�up�,]]^]�[���"���n�La�)q}��4 »������0����g^RzH<V٨�zb�+9�3 t.�K��8���<��N��83yk��_3��ӵBG5��a]|������&g�~��G�C�������ÿ��AD���|�Ohk23�����7��8ss0]mu�'�[�M�*������L�n��NX�`����H��=���Y6���ؔ�m)Y��͝�{R��Ͽ��o��w��ٖ2亢X-^�(����QC��w�W��#C1���G��$��O�{fy�+�9	I��04�D�E���Jzl��Er!�c�p�H��`XI�͍G�>�A%���M�B�傖 Sg_82��U�e�Ȱ���La�d�b�	s���|Qh�k��H>�9�2�� ��3��6�"��w��G@��p��^s�`X�$�uL�?�z�H*�D����h{��ȡ8 ,�@[gN�6
s��6>��|�6\�Sk���$ȂmzN/�m���*���0��Q��'�6�?��`�]���E����2,��ڝ{����� p*��L�b����.y�q�����es��L�x����+A��?�f�m�G������M���UMG�x~M�^�F��\hiz4G�И�Vc�����=v���z_߃�#�`�M�dB	��l�u��dC:�^f��C��$%*".?�_��������V�[f9JG^����}bG#���*�kV>7�����h��=ۆYD+��e͋z4�*vo	{�GO5�Z�+Oˇċ�Z�1�� �Y&�M�k��-�ܔJT�����`���>P� 1p��\j@0#�g��0��i��ng��pPu1佟�΄"�I�y�xhޔĉ�i���i��M��Ujs���2���x|�c��y�!�ë��-��Q;4��)������5+��Z����v̦�T\������'Q���LX�Χ�\1G�Xf � ����u��`��g���u V��v}yC�d�����qY�� ��d:`�s�$6��N��=`3ǖ����`�dj@f��Y0�s�P�E�w�D�l��/�����r����cc��i<k�{SJ�؏���e+�Ṡ��؏�dÇ1 �rt�S>�S0����'%��Ӡ=�R�ֺ�	�=pI4�����N�习+�|>/����f�1=�l�lg_2��.��b�<�Q����=��ٰ��G�;�������4%�mvG� ��e���;����@·d� ��g�8p_ˤb�+�}���6�	��%��S;�C�ㆇ�g��2�Sok�$q|�b[�D�ɋw$�w��#����q�d��<���/P.1�M������,@��(%黺�.�� �����I͋�3"s8zC����wE�@���S$�erZ��?�Q�=c(���i�,�[�(0�,6��siP��V�٢�?�0��7q�\B��S� h����T�\�:��j�nl-����G��1��{sF��%�ɉD�Wg�r�8���n�`P��e��F�⨳�� ؖ�lD׏��w�z=g�ݦ n,/v6��.`��X��|aDb��;[Rߕ�Q^W�3�~2��T�Q:�2�,"LJ,`�Cf>�zQ ��0&�(��mIp#��
�I?Cܙ}h%/�ۯR��'>�g�ؘ�� YN���<M\he�?p-�Qc��y6�x7�>���=11`ξ5s�� >���<����Im{��iphV�g�����_R�b�()��C�x���R�v�X������{{r|x ��G�laZ�m���=pВ���9;�	l��0qQ��X<��sg{�3�֟��'?'_���C橞z0N�WB2� �a͑��⾯}ZDo�*-��
*'�F���c3� ��X:��MGG��2���#��#{�6a"����Z�!�AS<��x<�ΞT��4X���b9�ݻ�2C�l-p6�j��g������	�=[U{g!�ݧV����5g��L29�٪��W�W��&�'/���u{�� 5��Z�<1�^��+h
[4T$�v֡K��@0d0;�p�lA9��I� ����¡�.f<w����0%�`����%_��_M�7k�����L�H_f�Z��s�l�H8�'��7ad�Ud&�����s�A�w>U�3>8�L�TU9��%��ٴ��Xj�=	#v�	���;�dd��C�@Rz�S��p�`E%mdJ��`/;E�G�w�J�$a3��yI�g_�*�tڤd�00`�4����:���k?Ս���:!#�)��`��d�ߒ��\��3`�7;���R�n2�á��ID��C�7�E�X�"G�2_�ʃ�71�׶B��Y����#o<��ۃ0ğ
�G�K��^�e̉���� �#HW�^owS�2�R�q1+@�7XKP\%3������l�*2U��M 3�C� �W첏m�r��dZ�l-��l��}X�M2F���M+q*��g�q������L8�p4��h���@TbLV��؛.*s,���w6�/��Uٟ�"s�|&<�i�q.Nv�H��_���Q�/Y�a��P�Q�6�� fv/��"�T�ll��r���?���}����ذb�J6��5�4R����|��������%<������ƳQ����~�C�z��V���g�}�z��`T&c�������e��d}w�λ��[���ܞ`�%�4j*��̵�O-�<ʶ�����G��H�g�m��ǜ*�a��FZ%\%��S
�>���!��_�o�I|	s�Ƞ�@7�Ss�%E�n���c㨩�
X���v6�R~g7��M�d�n_�\� ��a�Y�R@�
x�\����k+�c�w�Z��p�F��ʫ1�gyךt�y̦f_)�\�s7�7�+h@V��%u��z�Ɯ�FI�Z~
�Wu^p/��
��E >�i�d�o�.���d���%>�VLS�t2SЇ�oK	���b���ne��h���T)�u��#����@0M�M�,ڶaC���*��t�9A�6��O�Dy���e5?f�0�]x[�}�HK�2��8�6�Pd���8�~Y(2�Wkd������#I]"`��.I�g�c�'��y�����'r*n�r�V�����MA"I(5��d��N:t�kz^]����*�-�B�.5�d���������S�(5����Pj���b_��ߨF�>vX2l���9�w͌���e(�c`�P����̂xg�`ݑ̊���/4�W�J�JW�v�*_�E�8j�:R�I���S_�rt��*M���~h���,R�������ޭ�)ILr�n&�QG�q��k+G�T��!�>3��Ǣ'Z���t�@���D�ë��W28��I����ڜ��G/����,���1�37�A��h��w�:S�a)Yr��vݰ�9i��3p~�z����N6���q@h��������(ˌ�~0�s��Ǆ'��4�IJ>��]l��l���dRu^z�s̀�.�:g�4Tޒ]��]�6�	!��2m�e��f�t
�,��3�����
�4���fQ��k��ܖ�4	ұz)8���:=х'Mݒӈ�c��I�������H��N|���ͬ�lG6 �b����2��2,UgːZֵ�(ctM�)��YD 0�BH��� �q}2u㥴̛�,��|���+sz�a�ʈ,%c��^��e���=1Bl�@�Y��@���f�wVѰ̝xi�;�[�]p"�h��?d��rE��7d�&�cĹG5��c��f����;���t5�N8Ѹ��� Z���T)�N ��L'��%�W�ސ-�&^u�ω��r�7^�hAf\�c1_��ފ2+(�Vl:�P��&y��9�����
2���{;��ǭ��r�<�	��ߍ����0qھ�P�g����b�ٹcٵ�`w�h���W�C������,�iy�~'9���5�̏� u�O)�a�����\�|�mT�*���>����ss���_�O�K����?c��r������í/^���<�6���R^�ܞ9�ʆv'�m��\
ʲyM�B�#߸�T�u�HA|}����(~�Nԝj!�X�����[��D7�xd?��zrqA��` �X�T��?/w8�<<��f��cN�����帄�a)KX1��\�d�O_�sjW����J~�F�d���� ����%�����8'Q����w��g "f�<Nʱƣ�� 5"��%J�d�0�{
�<�m��Rc�Os�#��ϱ�����V�T~<�BB� h��A�+ױ������^��X&,!�#?��܊���F��A�B�&�;Nl0�$~m�K0Hݷ��(�Ȼ�B8��f�X��*��3X9���+����PN��+�$�3g�y8.�2h�����x���`0���_�_Bj2*	�w�ƞ7טΔ9X��6�ns('�3֑%M�#HC�9��2m��8hvϽ�ރ�d��qs�f�� N�3���:�9�O���
�v�����<��Ֆ 
c���}�[�%#[�Q'��y%<4V���)<=0���8��/�jˉ�ӆg�`β	������V#;�C�ڹsłxc��<�P��{WF�^�|���lw<��w�3�B�jM?tK�ɂ�%���$�������,�d��<��jA�$h��M�Cd<H_�r�Π%)W�Ĳ���ۚd�����m�uò��c|Al@�`�dX8&�1>�%�5�[��6 V���g����ga\���8���YY���l*�� '��  xr� ^�hxt�zuæ��ً�w�d��� �Qq[�8�3+}�H�I��6�A����++�]�G3HΧJ�- ��h]�	��RY����-׭b��]�~C��X
�#+�(����.��o��b�wb��R/e�/��<�FyQr�-��_����Y�LMp(*��\��[�g��=�Py5�ї6!>'Dv\�B��0�o���m�M����8����O����;E�"� H���F�F�CEr y��U���;�tehH���峪Q���0�m5z�9�%^�.88}
6�Pj�̑C@3Fbh�2I�>ϑS�ka�e�y�}� C��fo�?��A��$J�n� "�~�*^F! 
r}��0�Fq��R��|�_`�@#s�H+�;�WQ' ��IwԹ ��ΙC��3N���VP�T�7�Ü|�v'��K� '��M��	������ls9е2�WG�w�mEi�^%:�H�B��Rf�+�EA��%Y`��D����#$���DQ{$W�=��{��S�h@�rk.h�D�P���{@恃��4��r
�x�A�<I>�T|g��k�A�h>�	�L��Vt��V�[� :FH�A��-	��em��VP�v�����^R#�p{��i�h�>�DW ��Ȍ�#��I��ހj����A��Ӄ����*h�͛�|��TO�e۵A޶���HH9F&w�b��vS�[������W�}X3�&ئlPU�����ס�<�ꔐ�ϝ�1�sr����n��Oe��//߼��b�"�mv7�5*�=�T�Z��Z��)�,ֵG���Pů�̬J�<���/J��28����g���e�}�/A��f��D���N�����2���X�@Dm:7>>���-��o��>4� �i`���_�?va��5E��A�D����ԵiT�g J���r_)��x�	�Iݐ���Te�ʦ���uU&�����Y�.���R�,��<B�r�t�N6z��jK&DG��n�y8y�'6[���З�s�u�JF�t㎯�Q���6�$kseCbU�b���e��(q�8��D��Y�,��8ѕ�Q�J�%�r�0�����Iy�w�&�y�O4;|@���(cRF
u�������_�΀jSd5|�㿣u-π���4^�A��<U_�q��Վ�|�'�
���,�,\���M��]�� u]ߗ���g/�u�w�âtp�a3��J������3q,8�ρh��S�LE��ؘ����sόi4�$�!I���yː��{��A���-�YlV��/r,���y�u�����^���F�2~EGPǕcΡ��m�ԡ�9ޫ5���ֲz���d RY�H���V�]��8�W���E�/q {���5��oX������k��Xc�K2aJ�X��4-F��QPcY����n\fD�y�5m:�b��jo)���rt|��e&{Os:��!�7���;I��~��Ā���*�Y(���j��{wv~E1ш�Ax�����������(�7֤��:�)0F)�mV����ٛ7v|�'+�kh#������Bp�_j��"Ƈz��Ǉ̂��`~�u��%HQC�A��?X���uLk/�d��M&[�e@�`%J�,i�-KS����>9��~-��^ʓ^�+��5_4��*��V�#��)���k�py��p��
�UJ^+�Ff�O�	�f(hG�q��n����������y��a�!�!����RnÕ�n-1x�	 �r.���N�L=߷���.�L��y��;s��.y&	�D�Y�bc�\K�E1�1QTf$Q�G��v���5�&�h��T��2�LNf�\��J!>��}p� \3��.����j<��ڬ^0�
V��ғx�3�R���Π?�C"���w���Y)4IQ�������8�aTA�|讀��1�eo9�H7��7�� N�d/�9�y�PfL癨4t���:`��!;8X���S����5G&�?<r�E���/��J�U�����YhE#�:����k8f�+?�g�z҂��3<�x:K$u������Xg��Y���~�喔�J�w�Ɓ3��(;e'�҆_���.*l�4n�7�</Ydgdq�JyX�!�7vX��/ �sx�G?��5y��������\�ڗ��^-�SVA
x�n�|S��#_|b�Ty�;@Ud��C��־0<��ڔ��K�Z�4@��f�/k���e;�~����~ b����� 0�|>[��:]K'�5���Jju2�x3���Y����;����If�X�P�"x��0V;��ސ�"��c�ym����'vC�V��4�C�n˒�{������F�m�R d��u�Ա==��J��ˣy��H���(��Z\^]�_~|'?��蘹����t��F~���	f����g�[̓TC������t��)�\b6�[�_��Gy��K?w�u���L���Y.>_|ͼ�ut|��>��S82Q0w�.aӓ���Vίn�͂(+F�@��͛S�曷��W���u�Q�>��O���a�_��D���뾑��߼~��oA@��^�,����bO��ɉ�|�J��ʄ-�z
�pnS͌DxO��?}<���+�����[�����~�е/n�Zʧ�K��?VNȶ���޲�tx��˿8ޗ?����.�o�����?�u�w6B�6�:A���7����#�>�N�ۋ�ͻ�����[�o�}�Z���7����5�W��ܣ���EFS�)96��]�ݨ�V���9 /7����K�-K��W^ZO ��N_7�ͼ��-�k���2@�T�H�;VҬ@����sV��[rÚ�`�� �V�� Y������>A׮����@<d�TYC�	w�	�ad1��Y1}�)tzrD�u��Y7�4E����LX�(��22�f�mN/�'P��iD��y���D�z�J^�:����_�E.�%�<��@��	v=zV��H:���Ԅ3g:�i2�L�a_�<����
�O	���o�_����I..oe�h2l���q�A�Ro�Q�aӞۯ�W����e��D�#�=�����ǀl��ê�\��{K ��I �~�)i5D
}U�X�>dy(�!􈺜���<��%����4 3��9�-��(�ϭ����<hI��j>���l�<��h�_���r��
�~<~������4���W��8@�(�9�T�����3��; ���eq����Ҟo���<@�_���g�Ϣt� ��gk��E��ˡ�.�+@X�_�Q�3f��������@3%o�C�|b��B�)���S0�/AF����ۛ�b���;`�:Q�0±��&h��a\�2i�;��`�������m��F`Ӱ�y���n(_?{���I�%�f�����������}#G��Og�j$�4~#��jJ��r||�n����f$��͗
�.�w����ĚS��h_~�o�o�2��[w)��?�$w��F�����ߓ#{ `��mi�Y��8�X꥞[�y�Y�.�y_��M0�@�W
n�����~q�r�D����R������
�~�Z���kuR����	�1E��zA���J��pO�2�b4����V�.(�� ���+h=��YP9�{_�����^�z������w8�]�a�[{J�s^"�+�~��'O���߽���)�1kz�˿��s���#�V 9s�ߥ*�=}���
캬,DG�O� z��cI~Ҏ��G��_ɫW/)��A��ٝ:�')e�8��� �&	e���B����������ưFcĭ<ޯe�l����,?����9A�=n�g�l�I�l��K��ȁ����&�)��(���T�������AWMy�;IM���ӄ@b���?3����Z��(�P�!���H��,�V��}0��5�o��>�������R�����l�.�+K���V�"��{�gᛯ߲���O�K���@u:����?T�~l]�]O]a��h8u�H�˕>�k���2֧'��ׯd��l�r�?��uc�'4�P�V�N�Ԛ�Axx�0��Yp���?|�k�C��b�]��`��gE�@����Gc.�nU�lɗ��ڌ�����8bE�\S��3��kS���c�}q�2B��V��eF9�e����-�Nq��h����x��â?� �����/����\r��p��{�57����.|�覞�-m�����>E������|�Q�6��\�W ��\�˭���k�d�r!� ĩ�r1B�(d'�\�w�e��8#l|�~]�2��e�\	s�D��� )���?3�]�� �z�x��W�2��	�
�6���Ջ'ꀎ�cR;��7���L�>�� ��?���+��;}?5��NY�������3�������,Eh����,n��(M?ګeM��!-)1�5�sA��[5�_+�88P�4�(g�R��с�#���f�C�?NX��H��8����̸�sp��}�\0C��[����L�`�y��P��EB��;�s�v�� ք��Zj]s�>��b���ƌCt��}� �(ϵ����7/_*x�q] LN_�ț�/�	;8X�Ȥ���x-��FZQ�|A���"�ں���Z�}2�2�w�:& �!���ބa�=����:7%[���FƤ�hK�4�f(��r�����\^�\��^�d�?�T&-�(H[.y_�Ԣ��N���NF<sU�Xv��	�u�g�g��3��Yة�>(���{S���b��K�ԇM����'DN_����G��>g� ������LnP?(C�:H^`�*���A@��)i� ��T �Op* Jd�9���;�q]@��9���=C�e���B�1� N�%��	VSw�';����}��6:��b|�{5�[�6����}p ���~��J(����+0��{dh�olmTZ�����KygQ_�착�W�f@�[6�p�V0@b�@����%�b�lc� @9�J��j����������˰\�,q�@�25�������{�>^�3���Y�h��"�X�E�c��0���j��c�����KC�I���=�s �����Si���~>pp�\l�)���Q�Bݱs$63��y�̒�8 �fF ��X�&S���X��g������%��Z���E�����Mҳ7~����3#/S>;2�A]�ׄ�R�/)}�Ld�]C9,�/Tv���K �<��R~L彞i����<�_�Ry_�İNc�]�k�;��Y��g�EĐ~��)����������ت>~)}�y��˗�Q��G�5���Gy0_2\�u9�ua} �"0�f�����g�ՉY���l��ŕ���(t�����7b훯�w��ZN���a`Lʚ��Ƥ�( X���Z~����7��l�\��/�������=�rs���͚�c���h�b�f��̌�׳9Z� a���_��`O�VB��d�  �������tY���Z~zgC�'N2���٘��)B���H�{ )��Q
F�L� �ι��B.3��B�� 1�&����m��eR����2TȢA�	��C�z�@����9F�4�Ig�G�O��l����5O�~?���P7����󥗖L=����M�\(������D��t�)�@R���UڿKV������&Kް�}3(���[N�'��3c���@�><���X��į�+ 
�thM5�!gâ���x #|Z��@�N�H�� ���i�LZ�M��,�S��{m�e���{��|�ݷ��j�̲^=�Y)X]p�(�YG̚]��}�,?��R���� *�=t;0ˆUE4��x�6���s'K�:�A�u�phb����N�f�E�l�-�oTQc0y2
�Œ���
�O_���|�J��5�2D3�U��~�8��xm��X��E��-6�:�3U�y���QFE��"��1�o�<��� �P������fm*����!&J4<��[rB�t_�.o����%X���	/��r8�7.����F���Y����P�z�C6�x_����%ϬߐHz��#O���ͧD /�,���U$r�ۮu�.M�ᚓ��^flS�r�t6���
c�F@e�)>!�C%K�?c��ؙ��E{2M�*�������q\�M�s�ן�僌��Z�������~����A* ��O*��H-A�'�!p�c�g�h��_���X��fF69�	ْ*6� ����7����"��4�k��]�Y>1�@��R��̉�!?A�O5�K����|�ա�o�J^��c�ѽ���[����<(�x��a����j8���������?����wZǤ�a�Sqw,�k�����UЅN�Wo_����7�������#*�#}��b���R�_հ��8G��*ࣛ	��� =��|�쏷��f����d�)�#��	�@\+$@@~X+��k���A>���+ �O*�i�=���P��F�4�y�L�Qp�αL�o �/
F6�� <!���X�O5Ҟ�S�hZF�v�':tN�L�X?=2�S�cO�\��%4���T��Ӆ� &�
Jp�
Pz��T�{ �O��G'���賽yA�V�~^��������֦�,
"| �w?���:,-�9vSf�l� ��8���6�؉p7V
jY��By�|/����W���GHSy�����3������T`m*��qF��4��
'���޾���I�Ċ�	�z���P�'��mFnc�Ls���p�<`�%=\W�
�s�-6+�_|J��a����)�(P@�(@�BAE�g֚��%Hf��uJe�@����7m�$ˑ��̏���<*����Wd��"��_wegg/�KNWwUe��q~���*�g�Y�FOLdE��]�
@���h�e�y$s�7!��⪸���}����!S�Ɓ{o]���(5�s|,�>f��M+9;ڕ�ߡ����|�I؟�M(�ֆ��D�)�{�'A��p}�?�^,Yzd0��<�/�2�@p2���0����H'�ߏ��n�ʏ���Vά<���M9�N[v볜:�'�m|��⧍5Ĺ��ml��Y5��ɹo-�+�~d��2Q��@X;���eŲϘ�g���JA�?��6�ǻ�S���h�w�R�s�ҽ��H^�|J��Ƌx�LJ���+d�.�!^J[��e�9 R�pY�I��p��\90����(m�ַm���Q�W3���lX����k.G�?f��	���������1#�+�9��U��v%C��6 �C(g�Ӹ/RR�E�X�a.#�_d����x���3��{���7yw[_��|p!v�yإ*�oͶ	
�^�1T������P�{{����OKٛ�ʓ(��(O�3�c9j�ɏ8�ٍ|�#�����g�1�ӣ=��\^�:�x���F�ޒ���~�y\���ry&�v���JR�jJJ6�S,�b5�V��3¶�� @�Z�zm�	�"�1����>�h׫��k�F5Ʉwq�T�{C�a䧧g<o4B�"�N�;�4�*�*E�\F��R	W7��;����≃�m�J;�D�I\�\����gY*p@�M��:(}�G�	�:��1�kB�0�u���8gf��D-	2����r-w�6=��b!3t�Q���V�7J� a�R��6Ҫ�e\�u�鹶�~��4>~�sp�> <�D
���Q�2��U8֡������V��A���#A��d�2S��ˠ�gd�Й7a&e� NzԶ<'$�

g׋�Vf��MS����I'�Y�	��D�5x�)3q )̖j�%�0[���]2�Q6)�x2�V*�V�U#]%e�Pt���ftrt����,�u[W�<�U�L�x52��h0������zpr��5\�k�Y��/v���=<<⚼���ۻ[���3A�%K:��\!�#(��[���L(2��]ԖmG������m��.���R���$�=<Pj�����M�n�R���Ŵ����=��['���9o��N�)�+v1o�H���S�9a%�I�7J: �뉐��f�*������Ov[�MK`���
h����I9�2�n�{�x�!�˳�p�F8Jm��I|}�Rne �^/+�u���u�������rX����������%J9� �G&�*\�\^����x7�s�R�J� ʙ������<��J^�y	��r��5����O\�0���;5x&C@=|l2 �e��-�5���\�H��C:<�r����;�A@<	�k�Yf07FyCYm�sp ��p���u�lV����x�D�X���!4��||���.I:Ei�X����+��v�qM)I�����m4�ì-e_'�WYq\�]_�D���J(4W�f�*$"CqCCW�������5�g�t�(T��n�����]���4��,f3\m�����5:=9��o��n|����]t��qଘɪ,�����7������R�!�.���?�*0��hdߦ`����G7���h@��l��!���:N̯o�LA�zK����v%E�B�@j�2_vB`c�Z s��1]%:!d����d� �55 ��4�窈Ӻ������Y30�<���ѵ1
*�º5��d�����k����<;���.[)�JTp��İí��Ad�(�{����0�
L�G]l��.aN%@@P�|:���lײ���%�ZFg�Rin�ϯ���K0fG6	3Q�N����ԛ���]vE[��\����0m��h.��Er3�;��D����[�J�5;7+ޯ�^��T�S4�O�y)k
���cf�j�X�F!�&_ǮDj�A�C�ӌ�c�h̬�6�7���_\^K���7ک���C�W�Z���Ϲ�V�G�����k�^��;�ځx�,h���J�V��g��4��N3�|�*4!�y�����;&���#r�:���x���R��X�d)�Ҫ���$U9�~K�Z��;���|��)��y�Q�H�r��@�7��lÃEw��b��WɼXh-1�:�t�=�S�0�G�o��{��ð-���WOڎ��ϲ�@��_��o�	�|����� @�^���
��:\�ɧ���T���+G���]���/�|~~v�=�+�2���6�:��7���I�q�������XE��o��U��!�̚��5�2��LB̜ð�rkQF�
p4�e�p�a-��/����:���B���" �kC��{�����fE������쀿2�|:@�]:@8�CϮ��,2����e�>گ<KY3{�6Pܮ�pЮ��*F��D\ J��j��+ƈ8���	>���Ȥm|�@�rqf)f�URhч�k%rg9���yR��\,��&#u<�h�#���4^�T�% i���p�ᘜ�N1گ� .��)��Ƈ�Gk�f��Z�qX]­� ������)S ���D1��<�p��W6�ѡ�(�ݙ����]u.^�U4o���Bp]h)�HnSK6�h}dRr`�YRE��p��}�c���18����dB %f�,�k��c35�T�2QJ��c�8-!�\���S��yW�A+��3F(��n֞%������~����TD��D��(��z��ސ&����H!��qq�i�6�#9��D8]lS?N�K��g�������.8ϳ9��h�����6!��m<�F����ݵ>Fx�>�;��
��h\��9B�:f�Ak �;������K=>:V�'���A��7�<��k�7
���g��7va����3Y3j�`n��D���OB"�lBw���t�x���]��m�Aؚ�/45�>��i.e9�
a���^r�-�� S�ppF�O|�����\��R�H9� �$)������zY�PXJd+|E�As�Lc�١*.%@����}ֳ�2��noʸ�m`�n��-c_Z�*xJp
�Ɔ��)�j�pg�(<�aơ~�ֲيĆWj��xD	�h)����M ��u�����T�/R*k�W��|j���m�i�1�x�������B�8�5����F�{
(S�o��Of�WbU Z`ٜ2��x��O]P���·K�.Lw9O���od��c�@>���lMC!�]�+�!ȫżA�~sU���_������ޯ����Q0W�e�|U��!���A�ef
��l����Nh���0�؇���L�2{x��8/ϡ���/�Ut^�x����pu�E���{�N�rm��f�R&�R���&�s��L�)�:oM�	`6��-8�|���`�������d%�)	�8O8v��k� )���9q�*T��T^�
� �� C9���a�C�g���%�I�����L��?����_�?�����X�_j�9�k���.������< ͸���*��>�A�Պ|������$%��Z�!i`Y��tӎ��fd�v�ۖw�����g|L�ㄚ��=N��i�Y�������u�c�0�>{pD�Pjt5v�����9-yjk~sP�;NV�$��4�(슌�O�e"[5������%u�R��=f�{�L���X#(j��LT5�\EL=�/�1μ2��G4\^Z`��c�>�ߩ�yfv�����
�K���Ý���_�ݻ���*�H�ZVm�uN�^�9<�9r�������]2����.�]��_7��{Y���AI�� KL� �R��3� FU��Gy���׈�5f��z\�@��`�g.�s'݅�3�Ҡ��������_� _T
=��?�~�~�%�a��\B�ʲ�A�W����!(dh6+� 6�r� 3ep�M�Ȁv՚cA�G��n����������@\�]]�!�.�@ϴ�*j�Qj�6c�%=�������=BݯrY����^�U;k�Q17~��_!�<�u�B����f�؃�_��/�A��R��w$���סo���`��r.�����<21yޯ�;��-�WN��I��_���"�㟂p��΁G���;<��I#�\�\� @<�e�l�H��{��F#whT��g7*��H�	��2�=�[��&�7��{@���c���99Hp4ˡ>�' "G�D�K#Ao""˙������Ĭ f���t��c��q��Oz@�e&|é�u���ŋs��1�����'�4�F�ޥL��
���=yz��r�0��0c�'�1)�(M$Tԧ��$��':�j�L���$��+B	e���9u��ps{K�<�V&zۘ~O�16�%+��(������2�lFϝ8� ?����5���}�`�[���)��2��> ��Q{~VЯ�c[bp4�b�8�򿪒���$1w4t��i"+���5b����P�dA�.�5shl�9���;!��d�\R&�,���`(%0��_�l'ݙ�.A��\^) �A�� o2��`��Y��l��qͱO8���.���^���5+�i���U�lB��mv���6s`�D�����0��Z2��:3��zm�Y��8H�X%��T.R+�zr�W������+�ٰ�>���3��� ����{�����A./.��,���I��g�Rr���(&R��~o��8 \��
�P���®��Rj��������|�+�x�]�ވbM?���8���L�R�ހ�U�)A�H20�h�^Խ T��2( ���w�f����#�2R�����ﲿٴ�	�&�(o݊�"�e�������i�e��E�����@�;fƔ����ߋ��a�O|�He�&��\�.��3�D�ӒX5�S�R9�/�uC�`i�y寁V`�4�)�,8\������������	�o�<Hso�� �����PP)��`� � �d���'�����M�!)>aH��wr���ZN"���U������5=x��i�,�J%�V�W�2�(�`3X$��m�A�Ue��BV#E�� �Ú�D��pZ߼���xf�_��b�K��pri]�n���Ӄ\_]�|�익b��k{�XU<~�.��!�2��?M*��"}��`_����M����Q�?���a㜤T�1��	PF`FN�9OH|��[y}�BV�؇���ӧO�L.�Y�lgwB���~�,����gG֢r�������	��3�ob�;��3���ug;,)B#l��O��!��G;{SfW����� &U�Y�ʩ����n�g��cd�r#���8~�	ch��	t��e�FuD�
�V�8��9�s�]}�p��7�
��1X�%.*Z�||�d�3
}�U�1�4��$Z�g����G�L��e$Xn[��?�=I����.��f
�?}��;�B�?�E�>�t���y�f�- Y1d�B�|-v��6�z}�z�e�9�t$s�����|����;e�ޮ��}�燓}��u]�~!���w�rqq�`� <�A���!�su�Sf�����.s�Go[�Y�af�Y�؏�'�s����K�H������r����#�����<��P�����g���A�����ã\]_���>����m&��^�f+�#�[y&���G��� a��i uzu#?~6/�j�+��-:a��S�D���}A1����Mz��a�[����`i~eYN*y0b��d`�*�ݧm�̓���G�gQ�X�r3�������@��2�"|�;=��-}�r���:ګd�[�F��!�$P��*&���T�ecB�^�C��#��!F	e�: �x�.�ކ�9�m�뀨�].�t����<-�����~q��.��+@"p��D�>V�uRs�*9Y�R%����Ή�玠*6MyYO�+��3y�Y��T!���e�`&>k������!���_��4̹���}��0ǝ���qɩw����x��1��S�������|��������FX}���P�N��D��;��Ucf�M�����gĽ�qGɵo4rX�x��T����T@�~x�SW����Kh��`o����a-^��a���\��(�sڎ��5]`����j�����.�]���������:���х>�7�����v�P[v���Ƥ! ����r$ �
9��Ȍ֏��5�Z���сYս�v��QF ��$@�����J�3����+M� [h��>{� }(9@g�"�����zf@%�X�=�L��������1SR�:0�q?����"@4s�-m7;�6�m�~?-Q[\=�K�,�Eݳ�8aMmrs�� �Ѓ���x�d����}#���S7ƣC6@s�ex:��4�:���i��q���C��G� �5�F܏ �ϛ���s�>���F��s���f��a_6����Ȱ��2y�0�[����lS�|�����8�m&�<�d�QD��M���.a�&n p[/���JO��6���wЂ��r�Ә  M���a�!��R�uU�\�)+���sF�~n��ɉ��p�a���X�Ϝ���ɦ+�֐u�|xg�;um��>}Ӻ�l��Ÿ����Iml�v��(D|�e){�)�qG5~���ip�� �<�pοp	;i5��1�@;mhg��@��a�0������Yܚ��d��-�r'F� ����6�Nښ�V�"5 �@}PȀQ��uP�$�a�(ҶE�[��Э��{ �e0�
������N�x��|֗}���Щy#2�\��}��x�òc���H	����x%
�_�2�m~!BA]�ז�T�Z�s�t�0N2܀G�=���X�q]#���Wϰ7�[%����@s�v��iD܊m�� L+8��[�b�3���W+�X~�� �����a'�W��a���rN�
k?�  �ɮ �?c#P�P��j,0
�	-	ľΒ���i�z��g�Z螚�À�`�,7j/mx�Ʌ�6]��[[G,#媌����=0Nu��y�n��k���T���yy%'{�LΥ�1� dA�Y��p� ·-�#�ch]����}y��l�cy9b(%2���!�$����>prSJ�M���n2! S��s��߾U�wn���tU>?�볽3nSem��\˟/�>9��`Ӽ���3�&��0Je�ܯ1\w�QaV.�ۍ��u�7�����l���%�9d�3���}wO��N1K҆y�y�+ �� �]lLv���VL8<�D˒����|�`WvN��s�(:/p��=ܙ�������ͭ�Y�k>ߣ�	�!2���_r�%�����\�˺�r��͚%+�g��Ig%mQ�Q��{�i����#]7�@����
�٭�n��'�� ܫ��7�9������l�! ����y�ѕfb�бZgd�9s�$Ƈ-������[n�n���6���Fd/���=�W�m�K�gL^5&�|Xd�0��Q''��n���;�#{�\�8���������m�����w?˳�i �5+J�=KM%�=X��T,�Է;��l��BU �*���*�N沝	�4�*�d��7��h/:ʣld}� �G���ll:�qIPS�Bڂn��K>ŚaZ��(�,��&��Y&���,��$<r��ZL2��l��s@�A�M��� �(�'�HrUV̒b��I/�vX~GatL�Wu,����A>+ {֍���X���f⋶�������7d�)و�&��Gj��a�fQd�W��8 c��RNm���ξ�o:��ߜ�ZC�]{dz��Z�����o�aB!�C+�"�ђ,�V	�'՗6�����)������/�\�9��|R��#~)��:<�RQv��gT��%6lo�y8��W� ����Ӹw���9Q@�;��ת}�0!��
���V�{��~��p�W圙�a4g�8��ՐղWc�)�r�0dJ��;�.׌�`|8�v���N�稱�;˒g���beI� L��wa���C����F)�3��^Yd����H+s]t��l��k��q&�/ײQÌ� �]��r�E[�5��!n����+Q�xtdb�(�҉9��F�
D&� J����G� ��Qm�e+HC@m���I�Ō�yxpDb|�<�f����RY����&.=�6���f���m� ����r ��=N h!rQX���D��JHl�z>�@�gI�R�`�G*�K�M�mY+�Ô��:��E��ASr�äu�����Q�˒2)�.�u=k ��xef�����ށ�J�ox�,���X�,��$dY�SR��*��q�����h�`���r-`���W�嵂xL#��~|���G������N�3=�1��v�7�˹^?	���ă�`U��\/�qE��v�\,���I��:%���°��}d��c��2�w��p�� ��x�/_����ڱ^Q�BL���>	"[	_��O_0�|yqI����K��+)�F�>L�5�𪞚����#��3p��wٙr}IL�6�Pg�X��� $�`U6��u��2��$�<K�3]{3�C�@W
^0@%����;�k��5F?[�J��U�C���&�{��e�DQ��$),�y;{c��t׭��7v���*W5���1`�נ((.i'��vK�Q�Q��hk���A՟�P7K��+��Xf��"+��iy6����ʌ���5Gꛁ����L�V�h�=�*�%*��p�b�&���AK�U��	:4����X8�����`�Y,�H���Z~d�JP�J��ϫ��Z$���9a�w�[��\_Q�/�u���C,_�O�eڂ�l��SYH= ��;\^7Xlzk��T�:+#�ft�G��LI�L6p��n(�f1���[Y8ǆ��:ȶE��$T��o�C�vk~
3��Q��t���8WL�8�-�	����6�k'a'��I�n��#����y��J
�nn����L7��B��*��G ���{� d�*k�K�]�Fⱓ=v�MF�n<��I�)r�[[��Á���av�EB�=�@bɮ�c����aӄ���_oU�D�q3�����ZF�P���B�.���˕�{����|�Ϟ�8?��cd;f�.>�ںe_F$�RA�
k��]�k�p�!{|j哾�����|��}}f�I8& ��J��ӽ���>��;rt`|���1[\�	J��\\���NP��0p#�Z�9@~��~C'o%�LN��1�ƞ�kY��s�������J:�.�)�0�P�i:�Ryh"�-Ud	��SX�Ԇj,#��_�w�3Xq���&,�m�s2)��|w{(�w�,?A��T�i_~��C���3�c6�;���JP�x��A� ��V��(4�A����ɕދ�&���)�?lbL��s�e�N��I�8;�W�dg_����Z�FXm̹��6�)�8bizUK]_�y�s�ޡ[I��]b�ןt[I����:�Ⱥ�^?�¬�ya�;���Zf�<�`��G�^�=ci�G�A�w�|��7���o�R����u�������G�x��X�<-W׏ry���o�`��qL}6�Ȅ��EBG3J�)�������G����=��\ ��&t��#�0�d6A\��!^���v~�ĉ͑ެ3����W�{��s=a�@JN:Tk�>xژA�aC��<t�F��j7A�ͧ��!��BD�4����X���nP��	���z`\�t?C��{ER'�·�
���D?)��f���;`#���������4�i��Z�$�q�a��1�:a3��7��&fH���}޽(I��V�X�\�uTI�&җ<	��Ȑ J�9��c�A�ip,
�ǌ-��F̈yM�D�A��r�">�(�+�{:���OC�e���_H!��E���t�o�)���2c���ץ������<.�����l��s�������/��A�cs���3�Eu.��9�54�Z#\�3��Al�Eq�3f���2�VWc�c|7(�A�aM�r�n�)b�d���ُ�u�8`�5�|s��-Y��d��Q�	�*2@��3Y7�dL��	�"g��j>��ƹ�4���qP�C���씗MKtM&q�n<o��� ��47è6� (��u@u���9�h��ӹ �$�ɮ�&yԎ�@��M@�����v�ԙCM�s#�繻�L����L�0�&�n��%9VcqT+_��f�:�H����6��02�)���'�[S3��o��L��U4��wԹ���cF��GCĎ���>2aJjj!����G�s31be�t�@�"�Ub��bI2�q�V|��e͌�IRd�=���S:����eg"���8w�ZX.�
�;[U���K�vG����{
��g'�pD��r>�X,l&l���r)�:Ws�k�����3�HНݰ�����k=�5�����[x2QP��X�QK�eC�9=�3�A
21�"�G��r�ˆb_���g�h� ���ϫ�_tm����V��g&�]�neK`� ��ƛh���L6�૪�������+$��1ު�qAf�.������3�Ӊ��>;�Y����0�� @(W�����q�M���-nW�^��z?'���߾y���^���}&�f+/#r�xJ�"ǵ����y��	z�����͜��i�xF��|ձ#�ld��&y2H̷�R"k6pTGd��̮�ٺ��YHP�Ew�u���5�Fߔ��=��y����S��0*�WF�j*�e2����H�m@�y��� ��3|�eU�� YXS-�D�y�rzԨ���ǔ)b8���TcN־s灴�.��	�FJ��,"qu���S|�$O���x�,�i��Ԑ�3[��̌\ň�]7mE&he��R��&����wdXP+��ŝ3SM/6�)�>u��%�[�g�5�m.��f1d��F
�pQd����� ���W '�����(��8-����vf�t.���):�j�@ �C-�6�p�3=8pr�m�i	�+�l[\Bd~r�ڷ�N^�k��s����7��7Ku�/�,�b��H�{��b���i!�i��ʥ L�	r�Y���c2���:����l�O�e�!�uSڿ33�R2���D�2�����8PԺ�i�V׭�@�S��H�k�{G�(�`sC,�a��R�!q;�\ �Dv^�Z��EJ�q7*\ˮ�,��Tq��*������F�տ�gsf�+�v3��%��Ũ�=Ź�X�_���8e6���Οsk�d�0+��'���>���l`��1{6b�|&� �}��Mh�j� �O�XR�-m� л�7������N�MwLc�u�,8]�S98�Sg�d�k�`Im$8(��.��Y����,	F�żÓ�#��w��7߼aC�+u�B��P� ��:��a�q?	�6��*���^�ŀ���F�:������3f-��|!�Y0t=������ �p�6�� qy�L��ၼ<;�?��w��7��f�c/��K~�}x�7Օ<��s ko2��^�����v�����&ϑ�l���^M�;*����}F������\�>��Ò{3���8ԕ7_t��8lm��Vr�0ˉ�wf�ہ���t�Ob��ܙ?�9���ӈ��\�R���.!�@��@<N�)ɺh����}��q{�Y�etp�u 2Y��v�3�f�j�r-�)3ۉl�Ja=r,�ݵ�?���	U����������������E�Ѧp_ò�q���0��<H��
���&݂�.h�%�0�c�k�c2{�.�k{&|������\��7Z���*�;��i+�����Sc�e)1 ����gQ&�t�5�Z1�1V�1C&L�M�A���+uR�Z愭��&�&�F6^�/�G�`צ�d�l9c���{����|�/xq���n�񷈄�|�	[PL�2��Vͨ��覮Xs�h��bL�/A�{ʬ�}j�K�P��1�6�s=�ͯ>�#}w`�����3Sl�Aؖ��6��[����R�����v�W�.�0�"�E�H 0�}�\� %��5�Y�;��h�ĺB
lM�#��Ze%*�N���\S��|��C�u��[����<��0�g�����v�`O���7H�u��ֈb�Tk4a򿳍�;��A�PR*��1g�%��#��,/QAݯFY�s����11=)�yy�kӚ dd]���r�u��ՆeO4�3Ƴ�h��y�h�P�"H ������|"��"G��ʞ�AZ�0��F�pg/^ȣQ�SM��"C7�aW���Ax�4�P�D���Cf�H����7���f�#7fڲ|; K�)���y��u88, �I��@��xo_�y%'gg���G��%���zT �1Qأ���l�u�<<?���95��΅�@?���Ń��%� ���l���w���݉�M'�gz޾�FN�'�8�1�'s���H����5 �&�����P��X k��$�4��ٞ:u�;=��q�nFP�3S{�׸3n�p�+�w��9�8=�s~#o4�е ��r�Z���ý����3�޿)��>u�RS�e	|�͵�� �C��ɼ T��H3l��ݩuâ�bkw�b�=�����MOv�l~��ɀ��<{Mh��ĭ_���䛈OB��h�Iò�����,y�"�'奶��Q.Ld=6�E:���g�q���(�!��08��j_K)�f)I���]��'��hm�;��N�W�_�]���'
�rݍw8�����Q/N� T���͋��x��D��w��dr sqq->\���̤.:K4�#�Y-p��ײ�`v�L���34�j�&Њ�8>)]��b"+H[T*t^���y�Df�^b�a欂���R߈:��䠷�h0�W�A�ڈ�����,PZ��ms��3q�V���w��"�n� Fc���h�<�(8��@
J���r�A�5i���ʹp�
8+�w�X�m<�~��4H+��˞U�E)�!��]Y��lQ�ST��d׍����ʺ�89���;�aSc�2 3��E� FK(��R"�����f@��2 _�����;�7^��s�+��,Zp����q�� l~�V9�����\2gP�J�j�({L\a3�P�~�ɽn.<���9:>V�y �C��̖�AKN�����+���|=��s7Cb"��;v!����ӆ��V7��\�H��4`����v$C�R7����5�N�����̀�u+�i�w�,eO/�x_���f��Fq�������񣔟IGP2�wM���F)��|%8D�n��0 �JW8F�e(W'u&v�%�Ί�}���ZP&f�`�h�7���*tD-�*�b �����N����X���=�g�o�
�N�����{px$��?���r}+�n��LdUF`6e"�ȒR�kg��>9F9���	+ ���
t���	`0����P;M�����.�/�^�#�Dǝ\�J�2�
�N�NN�i�����ܓ���Օ~�����׀�}N�
����>W������w�}Kǆ���V h��ԍs[��q_�j���9p#��S�v�%�R�gb�˭��ܰl;r_��ޔ��?=?=0c��N�����hp��_��(��\H�k  �������><ڽ./�4�\��O�,8�ѝ@͔�� P�>8���,�r{s-�Y>��Q.�ܰ1������Hﻮqr-�^�y�2L���H@�vJf�����^�h.�ƹx�^��l�%�򊍢�=��Fu銌K���1{���>c�.Ǔ��eM�{���S��U(E ��m|rL�{���wݹJ~�J&,�ȴU��qRXGXOt觰�j*���A��<sfD�8d��)�l|��z�&�5x�fkQ>Q�-���C����<��|����'|�v���L�O�t͌���!�$�<�;^�����^m���8�1[ؑX��_ˎK�G�
�:�`l�{�!�2�9���fƥ��\_�.�y֕K[ٳ�]҃�6��1z��XC��X,��Y���8�hF������)$cTӞ��/�L0������a�!S+k� �0���%���hC<��G��^�&��n_��󽺞�˿�p���G��*���M[��l8i\z��#qU?e�Aߚ{��4l��a���ףa4�v�(K���D����#2����y }z���(@X�>�W���5_}	Ϙ���SI��a�	��Hn������_`��&�B�h������Db;2A�7���A�oo�I��8��N����F5��~R��6k���np
4��y�HYGZ��jT� <&0l���vG� �0�`7��"[�a;|��p!��lMGg.V��aԗ(���a�Թ��������\���y�b�	_����yy�BNO�l�Om��ΐ?+�9��3��;���B-w���pC���+;� �A��ϼCg�:D����B*{�~�F���V�&r~�ϒ2"cw� 4�^��h���ip6�ޮ�������QD C\7
lP^�� s2�H`�R�|#�Ŋ�Rȸ�8�gG""|p�w"b�5Z�a#�.mXt��#`D��؁(��'H��|���ÅF�7r��h�9����>+�����謗3���#���7�oy�ߛ��7�	��'��y8��� ����/s=��k5�چ�`(�p{/����_�s�q��eFPj'�]<���� T�����$��â0�c��Z�u�t����H��q�.`|7��;�=��#�0��-�@W>��Zf>|�g����N������^�>�����=�3'23wJ�P2����{� 1�p�����!@\4��@��-�}�f�����@�d�D��4���<$Vs�)��b�ȵ��.�ċop���
���)�� �(v�� �������b�cd��А!�a762Z�`�JG�W9Ήb����S>e�������t�X��	���D��k�/.6k+�Y��(
٥}Lw�S2�NV�µ�g�Ɖ�&?_��}'?��^.��)ݒx���wb�1+�_2�\�Yk���krx���ɾ�lX�k(�p���l�۔,O��<_˜�M��x�k[�x0�^; ��D�	�CX���=�^���Q����>�g�A�$U��X�~��r���M��m>��V�w/ҘL8�7�*�-�r�����E�d�R���*�ǌ��cǘU�{Ԍ�o�����at�1.M�rph��I��'B'�5��OO�n��s�8��^{��@���G��k�xm��05��=퀇1��r���Uq�N����ȀJ?`�_}�_|��5Pg�4��:�l�)/?J䌆�dx�j����H�ٛ��G%���1��깕/�7r���k>�g���1�+���]5���.A5 �Ƴ:A^���y\s�Ԟ<�<�t�7��qbl�+�{�^���:S�k��Θ�C ��)��Cpl�S2�}�$�^�r+��/_�H?��70�����u�,mm��<W���:�Pd�ȩ���1{��{N��H��;��;ӆ��� �~�^.>}�\ ��Ý|����o~���?/V�FoU���y+��� F}ݭF�/�������g>�(q�<Uc�*��{�w�]�lMӏk��f��/��'u�P�������������#}N�������O�0�=���gdT����Ay�Zb
��uB�Ɛ����3�����a(ǈ���NtD�?kp������<���;!
0������Kg����0��;��</�ά'���	��O_���w�?���⑆Y�)2�(U����m���8�O�Y�Ae HlF$�	"�:L3�=�0�`��Zţ٭\��J���,��~d�L��L��������?/�߿�B;x�;�XN_�r���
l�m������\e<�~@�ji®�:�X�OS�0��45��؈��!R'�-��kL��f-��&wd+mw+Gy�$���G@L���~Z�� �N]o�<��K��l.x��M���X�����ݽ�{�;cVq���ऑqǑ,����R_>k0�I�������_��*�`3Y��\�=˿���>�N����:��Fm��u/�����2߱ZQ��)�%[� ���r\��<?.���[_?ˏ
�n�\/�2�ɛnZ\ `c��Vz�A4�!&L@$���y�ꕜ����������~��L���ܶ�%_���b.g�Ih����:rXS'���֩��M6�\���dc�[u�Z��8����LzNИD#K����ีR���ku��Ռ��f���kΉ"B�w�	�j�pd�U�*^U���T���� 6���L��2$8 J�bC_-�0�{5�� �A�Ǆ6
�.f+�U��p<���6�7�p�G76�)C��tY|�8v���į��ڗ[K�{|�Gi;���xc$�r�8u�ڭ�ۿ���8��g���\��ȌY�����#y�2��Һ�,��w��s�ΆDE�Y�̖+�ц˞@���Ov;SX@��%�U��Z3e{+˥�Of٢�Ȥ��7:UеKn���,�����y�R���FR�7�۱�-�	�<Z����2���
 ���7pe��uc�5yZf�Ѳ��A3L�&X�3*������A"��V�����Ϻ��Qͧ	������ޝ��IQ�N*��s�/�v����9� @�W�q��˛G����h�rv�/�)���(����H,�`Md]f|ɹ31+#����������~/?~���&��!F9R 0o  J> �Zf�&���s�$�V�a���֚�-�vu��ԁ|Ҩ��.���	��2b� ��6�$f�Zf# ��u=�M  ���%��'r��ʱ�	 \~�r�����9߰4���X2%������g�tu��jE��l-��q� %�тEu��u� �3;��m���@	����{����{�3��O����#�bF�E�l�7t��g1�0Yv��W ��l��$76�5a�1�#˨����+V�� g�TVg˽e�b�d!I�ɬ���M�3{�3����|ɺ�< ȹ�a�GٲJ�g��8֕=�SG,*c�Bf)�����2"eswfu)�`/����F5~�/���@B�`~v� >�/��+��IH���~{���������e�R� $l*�2N&���8Gd����I'�|�Ҿ!;,{;$��YM��4C1����u����-gKf�0��y�n��/��.�ٝ�ה��Y�6�c�&��;�Ĺ���S� \�'g�����>3�lʭہ����n���+���턯%���Q	�R�0\f(#W�5��]B������)����3ٸ*}��h <9:�໻G��{.r����}�c"u|�./^|Gm�5����j�e����X�i�s+�ӓ��i)R{q�N�_�F�0�8�Ì�I;��I����B��N!v��E���W\ _��5��1͛1�d&5p5*�F!T��]##�ؖ��a�2�o�kEĿ���o��?�A���Wb~܋����� ,��kʩHDw�o�'����ʜ\�Jڐ{@�#�����[��%q!"K0i��ѨI�F�f���m�&��R������]���Z�A!��������8{R�v/�r� ���I���L�I�H�<4,����©��bM�-o�t�H|����u�̊��U[ Z+�V��g�:�H�����r�MG9�ϟ�P�	�#��@��w�t/��7�.f`aydԙ^���-�(��_t�,;4~�tl��A�Ɠ�P�V�v���d��D���Gyyz�6��Q'��{�܏F<^�gĮ�Y��]H�>��<�	��Ņ��/��~��]�0�;N����3�� ���U)��ٜT2N��NF��F��F�W
*o����I>|R���fY�2�@r���� ��w�g�dάq��a�w��z�AVz�s=h��N�t�6H�d��wy}�@�	�s�b�r�ҟ�}F5�G����SmPK1W�8��e�q���s��f��B�[��z���zv�(?�S�ɱ�Z8�s��/ձ�V�� leJ���vc��>/�@/>_��왷�zu��)Q��(h����C�ާpk=1��]�T=u���=�<[sz�	�&��h h�qp��E�Jw�\����W��� r�Р��Zs]ד�5�/4&��t�(�&G��?�����Z���m�Ql���)6+3&�o/Zxw�e������F��������^�no�ͫs9���������;�\� �أ_n	����м1ed�k�Dmg��6o���lvy#�/�HzG���3��/_����w�o��]+����`M����0�q����@�w�?ȟ���dN�E�Y�)�#-Mnj�l�0`o�3��3��������w�w߽�W�^(9T�3epQ�&M-���	"����jV�f_�AZ��[B����x�aʲ�o�zԺ=�y#ۍ�Ѹ�D�xFէ I4�@�?�`�8$�`#��^tv���ܢJ��P���=�{.�l5^�B阎6�_�=���w`����s��u��R2��Fhڮ��aT��=���|�1�#s�lO�,x�/����P�|R�����~�j4�ԛ��6�<�f���B6Utb�}��kx�_�geJ�k ������W�/o/��~������*��J�}�ᨆ�8�m��g��(��m%$�L���N�8�QC�qR옂8^
�H5��K����r]1F8rr��m ~u[�g�$$&)1d6D5!{�M���c��e�[}J�wJ��,�D��k�CL\�~G�^��έ�B,�5~�	��F��u�œ�޳�X���i���ˍ|Ԡ��枿�]��586�IZ5�¦2!WD���2(���e_�����8@���G�d����J�����O�ۻ��?��۳��o�Dw���j�̆u����qt4` �??=TA���N��GF��� �	���7f���@_9y;Coso9;�Қ����U`���5y._�������Όj����Ҍ��_�k��3E��)����˵~�LF����{RPy 1W7���vl��R�D{�}�Pv� lE�4� �JvR��� ,PF٤{����-���.�s�;]c��+��j��V���o��~��<i`:[��ᐥSӿc7Ym�0��7�L��
`pu��+y��3��X�O�XaV���$a% Z|&J�^>�<��a��F k���?�c��Ջc�c>����n��h�O؜��4��������'�ޙ�<S��@���ءb���C���ܾ��s*P��&-�6���dbб��+���e�G��h�B <���9��B��䐶����Q��4 c��&0��z��0�祄r}v#N��(�C
(瀇>
pCJ�r�HJ�X��L��u���H�9t�Ƶ���B�|�b�z��_?~����,���^���Ȏ����̖��z	�]<�C��o��?����o���R-_Pn]�I�ܞ8�+R�����*)��6��3���1B8�����h��z$�*�*��%�ؙM��!&�*�;�j#�����ѡ>���u�T6��W>vh�D>2�rt������[�P�l��_d�b��_��4 `��r2��'�aQ� �`d/E[(�����`q:ͦ��h��h�;�_��8���^i�t���Z��|)���g��'�.i4��ф�M�'6��g��i� ��/_�`��h��/��F3��'�����Rs�y� �}%r���+Y�˰ ��!$=HrC$U���đ=]p5�^��\���������7���њhorP*�>��[��h�������چ�C �?;����U����J9�����}��A�G�:����U��>��yDT��r4F��ٍ,X`��7{`l���,{�<�����aNE��34�,8{�!`�� �;5b����� � $L��.H$=_p4���aIx_;�V����H����)�6�uQ�g$��1K�(��|F���#�Av�ț�'}�%������ڿ�b�M&&�a��HY�s^ƚz`Oj��ľX̸�K�1���P��;��^������N����8M�{��-A���.[+;^|��?��Nؽ<*"�/���1��2�CB�A�IEq^��l���K?@���AԌ�2W��?;��6���;D��_�8c�`�Q0�j��Cg+����>��(=�ZTX7+ʎ �5�&�R�l����$8���&Xy���K��;=�eO��Qet��Qr+P�t��{T�5��kyF�罼�t)gǇ��8��3^V�x� Q~�M�^d쾨�G�N�foJm�%)�����G��+~��G����2/�Q�O+��CU�Pa\_?�����+E}��?����۷
�����������(�%��>�?����g���p�AZb��SP�y3t�.�1�X�ֺ���Қ�#�#;���)����F�Ys�Ҵ��tʔ��k�R��%�e�Ά�S��l�s� ht�r�A�\���k������M�a��)(9>i0��\v�r���[�'r�X��RbL�������fEP4_'���K��iG�w����g��1;f9�V} ��Ϻ�Dcl2p��Vؐ����Z���,�c:�u��L�I��������?�᭮�C=�OLm#�6��5P�o�1��ƻE�! [ s
v6�>�T�%:e�Yq�L3-�s�����z�\���E4ǔsT0�Z-)Ȟ��=�¤��\��7oޒ6��G������"^������+�@ǂhc�l	�H0�W�<g�
1�J�8M��7��f�z��n(װ�Z����N��F&�F�7 hv[4�:;�.:�
�>]<j���@�O���L���Kݴ�tF��t	�����١���:�l��rG��r� A�K���}�� �5��PY9������B�U������������f��M���¥�,�^�H�#��c]c�w#]�^�l<�����,o&S�(�4pYDo����a����kg���[��4��ݷ6ct��P�f��g��0 =�����=�_=��F�Xw{u&����8�a��a8S�9,h�!�F�g�(|_T�Ś���I�s�L���yޒ���Z��<�9��U=!X X[��@� �
ggz=�q�q�Q��'��TN�O�=��1��R镝GG�(a��2�38��3x�:�s��3���?�Ӛ {4DI���I�ٳ~?j���l'ʭ�F�{
Zv�a��nh�@����L5pzR �Q+�5�x��ۙ�og���p��%KzYn���;����^�"�U[�u��3�
�*�w3�U1��NTܟ���t
�8(fun+4��M ^f:y���}� CI%Wpg��R��AAؽ>�5���"����17��nUp�`�[���o���H�c�Z#��ﱌ�'��s�u�ks�kgU�qsaOfZ���r��R�#S�;4�e����|N�@�φf�y@F�e����M�]mv�o.��1� V��5QXv�Ö�;��]~�7��/�X��;b�⠰^67�D�.$�x��}T0�Y>^^�-��.�r�	,Y���M7"�����a7Ep�Dl*S\G�!�H\w6�2[&����x�6G�f8{�}Hp�G�C��GY=/Y�=�^�h�6��������c��u�TR?����aFE���[ &��e��a��z�wO+�
�B�k:�<B��]@�~����nlx���g��Ǎ���kd���bM�������?~�߿�o߾���Z���K�+b��|Y��I]�l����9�;�,�'K��4�Zڤ��Qgc�LK��; ��fo,4@^;�J�ح+<��i���b�9�0!yH^`ܙ���<���s���a�3��c�= c�G���G�����H��d+% �ۙw��b\Kg>�B-Qf(�Ed���ʋ��\�k�iU���'�F�2b& ۙ��19�8;�hT�G vz�^����ߤ�|%��9-������v� �O���L �y'S�O��~�+���%�����!s)�4x�'��v��;9�rl{_~���1\��V�1���j��쥝��(� �PFa�5�{¡�
~�i�P�g������d�s��<�Y>є��E�)�Vq��xU� �č�qP�XRF�O5�d����yZ�������y�K�\O��^7П�{�'�5i:��6�cd:2j��� ȼ H��$HàkiŬOK�Dg��d���C�e��Gy�9��k�ɨ�-���s�|ը��r��|��?��ى>�%U�_�|%��$���X�C\M��A������@sd��c�{�cM��3�p-y-7���_��_�`c��.�AE���ق�Rfr�!�X�"=���
"�������o~#��^�����ם+�;wHo:fr�ѱ����yF�"}�لU� ��E�Y=�wJ6M)���)�x��gz?�m����h}�,2�m3�YkY��*�^�)���y����[1�hc�> �c�Ք���2c�ܫ��� ,�Y+�@vi�1kȖXpq��[=�3v�"��l����>3:��/-��@M� �b�0�\���Q�Gv7��q �R
���(�ISL9�Q�*�: a(�K����3d0-B����_J����@b�	M{�7Վ����!!	��>�����������ol�_Zѱ��Iㇰ�e6�.��d��n�Ȟ_��i�L"F|���aJ:���7b��"���(m$`��/OLϐ�	r��sM�V30K��W��:˒1p�왐5ƒט��!��ڵ��������?�L=�
S]��9��KXp ��ʏ܍��<vV2��缴&���t4���Klz����79?P4/�\��-�
Y)������k�ir5bB���j��zޯΏ���'��[�"��Z���Y����輣-����[H�� ̲Y��	Y�`�R�U�`�\ٜ\N����)(h5�33�Xu��`6 &�p �� �A�##Ф�������/{���$��)�Wtg7{�'�t��@}���;kU�,f��j�Vn	Q3s���iU��g������H���%��O"]k�#27k��Y��:�:ב����u���ݨ 
یB+�qS��br}Q�� w����5����;ո|�7��N�a>&x�V��_ �A�2 Ud���5x�XGj���c`�B�S���d#��1�9�{�Yޗ������A?`�Ʉ��;{��s��!^ýIy�5xR�y�32�e� A��}��,(Ӏ�uV�ЍS3ZŦ2��ڸ=��ʎY	@�^���&Q�lE\��g���ǗXC<�����&4�Ⱥ�涑B٢l1{�q�&��Ǆ�)�q(���(����gř�yM��T�t1��6R�r��72=���2g�q�p�7� Ci�������w	��N>/�3ʲ}������=�H�<��B�B�/{�:{��-H�7Ԙ�FJ�m�y���M��o�t�Ź�u�j����4#	�:׊�!d+�nP����b���F����^�k2�m뙲&"+!؊�8� FUKPg+���DQ�m�@�Q@�X�Z�(�-0�
Ĺ��p��,�f�B�@pչ� 2ɞ=�:�E�`��ƌ}>�������^#�2�2S	'����6��xͬ�b����#{Z �<ZɃ�r��Ӷ��5Ŵ��c�`O�N�C�@��e�^��'?LwD08Ym�T~&�M�H���ک����W
�>_~V'��c�*�=�/jM2�Շ��껑×|&h�.6�*ٶ�V����F�!���2 I�c��U��R�Ӝ��� �a��)�}6�Y� �4
M
�C��z�{� ���Z@�Ղ�r;x��gk��td�ɝ��W����iGnt]yyޅӳ�� ���2g,��?FK��q�Dl�cm��oc;)[��}��6��0� -�� ;[� A �wGI^���~����w���7g�!� J9���3��$2�~�����ɉ��������$�w.3$x|�ӓ����l��q9%�|�4��ݒ¨l�.3�Uv�`ϡ�!���D�סi��c<8������ڰ7 n��y��j3��XKK-bRsh����;�= W��W�姄Aw>#X�.�4� �HQ35��Qe��((���iƪ�J4`�#�����wv�$�B�׃#���o2�η�^�k���L���������I�®R �s�Q�kբ5r��E�;ytî�H� '��zD�)3�ȿxU����_W��-�Vr�	۵�@�=o���g�H	�2�]Q1�2�	PRs�dB�x;��6�YEr|ܰ ��\]!��G%��a)����w�p�u)�.� �~�Q"�g0Zfy꒽E�{�?��g`�����Jd���ĬQԪ&� �}�
P����wz��<dK����5�j��?e����o qZ��� K��2�o����d ���f4�%�i�������Z�k/;��R��l���ԯX��M�>"�`�Uc��umݳ�Ek���R*�����u+�xx�J�Ը��@��ӧUK������~�eN���5 `)ėS��s�*/Y�� �5�S���uɲ���b>.f�b /�L=ή�Df������i�^3F��uT!S��yW���V~�؍��� �C��kݵE"�Q���%�ߑ��y�Iy\q�"���4���qM^>�YmL����$��;�mP���TB]q/�Df�r��ʜ�!(ɢ�t�kogwl���L��2���R @֬y�Q6�0vm�p��}C�#S��٣�s9D�E�����%��oi�3&�_s�S�ٚ�d��O��V>EŪ]�h��=���k��v[�<ĉ-��Xw��YCUܧ�]O����u}�Q.?~"�	2)g�/巿�3���dMsd��Enl2F�P1��ϴ�l���<�yn��_��pj����%�d��F�-��& ��f="(��]=2^���A�b�nt��B�z�_O>���Z�I��@g�f�K���b,�a#pg�?��Zׂ�r�Or�ֿ�������o���md���(���;ѽw|��8Bx26
�� ~��o]�(s�>�{p$�g6� ,�h��m�	�\)���%�k��5��bh�+�4h��#�
e/C7ӝ}Ya�1d_l�2f��M�������U��K���h�%#D�8f��E��@nW�ǥ��	]�c���;ty���6���]����1��c�����ma�Әu񎃑�t�:�hu�}>�������7�_�q9S�C��a�M��z��es��C���L��uEr)K�)��������3}��Q�;�����@��� ����ʢo,������}���mH�W~(��nWx��i�lps�FΩ�� �tn>�Ò�)���w�э<���2��Q���B��"v6h$+�IW�x{�	&�V���.��Zk������2.���Ά�W�#�D���!_�Ot�V��U��ԑ�Nܲ1�n�X���#ć�;�Rgb��#�,m��>����5�*��4���lD�yk��N��P�0t���$1[���t���r��c ����5�U�^�2rg³e���!�|�x�O��h�d����0Ǟm��lAD�(w��H�A��r��)����#YYD".
y��פ��o�� J���]�,��8 궉55d�蔤)c��c��ʜf�R�)&��Od��Fd��c	3Y�E59bf��)�MP*�ߋ�3���M�4�2����(������I%��%a�vD{�iM��몵��7�	f�,K���e���� !�\?ȊN�����c��V��k̻�4��)K�]� hz�e<�!@
�V�6p��>I �;��2e�����=5[�q?Yg��Z�}	�:@3㏷r���]}f�	�P�������jǙુr�#,��8N:y����!?g�C,5�~�AaV�:��y�~�-$�_���(*��7R�-���4��b�z/H�E� ���`���ώS:�Ŝ������x�Lk�x�X`m�n�������|��+ٝ�ZCиZ0sE%.�(Ggr���I�.j|�z������+"ή�����[���.l���4��ג�4�N�f�+Ol�΃'̠4����ή��Wz�G���
���J"��OG%c�`�3� B�f)~SR,#Eb�H�7+���2t������X���vU����Mv9� ۓOd$m\8ҍ�C	��E��/_r�:y\lm6Ҡ��$뱊BWðb'���z1���h΄�*m��(=������S���E�ot�<�Ti�Z��
R�j���r6}�*;Ȉ&��+,����Z��8O@�!2�q���^1@X�Er�o�<(��Ԕ�w��9]��2n���<�d@��x�ɴ��T[~j�+��A�l�!y��џ3郜_��ˎ/K�t}�0�<6�`5ժ3R�K^��P����ы]4B&2&]�un5Z������ڌQ�s���C;"a�"���xI�K\�ԍ�I�|��O]�j�W�e%t-Q�,��6�RQ�M���ߕϖ۽�}'N���I� ��k2��3�K��Qzή4ιu��d{��g粸���Ǿ;�j���8���[絑�m"�G��4k���!�j�8���\����=�ו�c{�=��g�K�w^�������2E"�G$מqȱʣ�d l�|���!���~���V��T$W�ў�O�ʞ����n���:��0�FF�Ul��O���
��J= �|��rq�b@��H-�k'�@ �BIG3�^�egY�pu_  ���r�G�w��F�;̂^�<�5�CtƁ�ӚD��������ͳ}�s�V]�]��<�eB*f��3���i���Y��}�<���;�sy����F}�,e�|����<�05:W�晠�� )�M�,:�/�W��	�	*�	x;��|���[d|"X�k��5f�&���q�j�T�m��T\�(�{��'��\������M�$7�41s "�:y5��3;O;O������vW��b7��UWf��`�gf�@dUQ� �"2���>���2����O�C�x6۶��-�丳/��B��#d �y{i���������ً't|x� �w"�b���6lK�����J�Y�K��.f��]�_sȤ$߲�)�/�3 �,��|�����rZ�.fY���Xc"���PG��兯�ޚ:������c�k�&?%�3NZ;N�Q뵊጑{pשj4bV�7���Ԡ�,W�</��.*;m��j'=	"hs�r/+�8J2سؚ��۱|ΑoD�Ѡ|�i�`�فU��N�N���v���8����%��r�.�b��9Ib�y�<W�_����@��/t�,�7�gz8�i ��ZD�0���4��<ؔ~�Sw����;�zH$&ZT��� �	Ƥ!8�+H�l���`)���k�����V��x'��sM_E��N�	w�LQ!��8w�����V*��-Jh.V᜕�7¼�6?��TǀA��E�����6�%E2W#r5��' � �<��ժ0_g_���a˼j�jo�Dj`pU�;Ir��#����dD�-���R�C�l�~�~�Aت��4X�����/{qA.��I�e���P��$WS��<��S` ̏TB[��l&0
^��[&e�l���7&	�%m�*(~��؄L
TF�!doӑ���!j�F��>���B]�s1�3���i�Q���%G&���x^�5K2vU��8��v�g:�
��M�N��q@� �ť��x�o��T;,�z�0�{����M�:���w���]<�v��R�t��!(� ud�젪�FC� "��ts����3�� ;V��	���UA�Dg7�o5i���8P�|��ӓ&�aՁX�8}��}6Z����9��@{9��)��QФZ I����T��M��Hh�����p����b�k�=�9p��|����4���j��Lr'��Bx�LK��+G��yL��k�=Ēqn;�ע��zD2e�7�W�5r����g�9�T�Gr$��R}_�槺���nuUPެ�Q��)���x6�i�������/��sN)T鎥P�e"���b8�g�}� �f�7��#6��N{9k�O��J�:�K�������㸢�E�5���ؠW�N��� B��b�ti��ӧ�����:�XZk_|��n�׃-Q؈̶���od�2�O5����ꎓ[�Ya '�|��J
�԰�O�)��N���^r�=����Ex/�ų����0�].
�6�(���;9i])������$9
y�����N��M:Αp��s{=��_�������$�ۿ��޿�_�F@��/'�/�!��� �w{�F�N(���E�R��64# v�-�E�ջFc��'�-�ㄭ�X`;is�v&� $�(%��e�g��uè�i' ��`¨ތH;�Ht� (�'��ɩ�Rt$�Ks)f͠�ZL$m�C`�k���cj�&"�� ��P�I��v�����?<4|h4ox�U�x����%H��A&E}@b@s0b���pj���zT)��H�M��M��La0P8��vG����s5��K��e@&�^�'[WHTaO(��\�1�H���LY@�$�|6��,�kfQ�2� خP!N՘�Jy�3�);[�� ��C���(����tGd%��-D�HNg�j����a�#��¤!E��g3y{�F57(�LX��ǉ/;����`"�e��RǕ|�Ϧ��y�T
�c2���*�O�� sksiL=�"��ޯ9�9;���}r-���&R�^sv�Ö�#KA���&���,U�&U�UQ��`3��&f;ܥ��8m�-m�,��RfIBݏ�1 �/�j`=�����a v�G%@@��<f��i��p_��
�WΦ���A�j�0�(a!��砗̩@۬i�kP�v�Y��	���8&;	��Һ�%9Aw�ɞ�ۆ��Jtd��� �m���`u.�t��	���L���i+��Yx�t��맷�O���G�{窽�8?.�N�<}.�[l�.I�+ҙ����+= ޾{��^5[ۇ	��Jg5����6v��`�#�^������v>�A|J ���]��T���5蟌jG��7�D���^���I>r��E͡�*Ƀ�MJe��D��q3�ȎAYV9���_}-��YD9Z~:���!� �ӿf��0s�ҍ��^щ�s8�q^��,'V.�mx8Z�����"�A���+I]��g9EHZHa+as�߇{��xU#�U"�krW����@������k&���qD�Sռo��9��I%TJ�T5���80+�Ӆ4CMD8��T� ���0 )�`rʭ����7Tz��Q��AH����
"#��`Z��Ò�%\+Z����} #����h��f1���0�xv"�Th�S�����
�XRၘQ��f*Щ�d8&
�<g|~��;x-2��H�̘ʕؠ l��l�Q��k6�Y�^P�Ëہ5�7��,�cY�xg��څ�D��٠ ��@qM�^��C:g����Q���� ����E7t��{�wxC"��:�$e�������ܣ����jfZ&e(�������d�7��!lke̊0��28�)�l����S���ͻ�n��/�)��mV�K�I���x{e��7�B V�iH�����mv��'<�	�eMp��N�ά�&˔�<�#Et��(K{�!/�Рj��Fh���j�B��4���$i^ޟ=J/?{A��� xF˪'C�R�j��#xf�C�]�}8�c�ȼ2��!��X��6�~��[�0����5�����w�O������38�}�B��������:.��(���_�o!����gH�m�g
�,��u�W�����_�W_}&�����NG�C���o�=���N��r�~&2��p�����@��w��[}����8��e�6�l�$w$GQ`;y�`��u�(���&�QW�y�.����,��UL�jn�����R$7��ŧ����B|/�u���&�;s�(ݬ�d��/���^~��}1�d�x�����-t��ۧ�\FE4�(u/�������bc���3���O.3{O��_��\����Ы_�	�a9�����R[`����	n�C��M>ھ�8xBH'Qs0�zv]ģ�76����8K�y�`�����{P�|��[�%���,4W%9�A`�
+�A�Ĩ���$�/�N����Ww�E��w U��+�7.?Tjo,-Sh���@3@�0�Qaj��&����V��h+R�O��S��* �y���S0#ڞYɲ�IR���6G �����bm�󫁇���A���L��0��!��Az����H!��"��j���c -PeR���IR�^�s�В>��"�1 �}��j6��C�d@ Fi�d�3����4�A�!N��L �4������Z��#w C �q*�԰c�=\��V3��f:����}6�ǚ�r�2�NY& Lج���3�b�R?���Hm!g�ET��~_���<���s����Lk�];��&�E�u2k[��nfb&Ru1��J����`����m�x]j�ۑ�ΎS`��Ӊ����o�����߿���^�2?���<������5����Mp�N!�>�t��|��0�T���G]Cc���,��;ݽ�_��~��;z���8N���c~��9=�~j�k2�G� �4� #��Ӊ�I�uد%�DH���.b��Z���~��z��ZV���9iXM`-���kKQHjs���%}��`װ*Pl���s2�5Y|�Q�K9wn�C�p��A���Lߜa�^q���f��M�����V`1}rT�ͤi�xIl���(@Ɇ���H�� ���?y�B�^~��&p�h�.�#�e���a��.[-�YD"��ϖǏc���#�D5%��0>�Q��D�~��}�͗����(����$N�d��;2_�-�	����i�t�]*�fi���#��I=��ݝ�SY���c�p�@��#�Mc�1���f1�(RTET ��ǴI��an�Ül�j��f��3J&��b�su����I�B|�@_�D�7`��������+j�.�`m���x�9!�Um����|j��H`�!��8Ѻ
���g�@Z�Ӝ�B��{[ǉ9F� 3��a�kL�l.kAX8)X�[f�
&?;�`��xY_@	���l^V ���Щ`��;�tq��.����3���k���3)���4������X�yl�3(�I���!�ٳ])�}�գ�	f-�r�z�uhL�T�����ݥd	
R��BZaԩ�r=��B�u)f�)��M�P�p�)kC�aɾ�6(8D{mV��66ּ����Ԡ�c \E'�B�T�[,�
섧j}�)v���G� j�'v��$����?�\m���6	��|A��;2�;Lg���}10<�	N���1V�Rq{h:��1�t>��� )����N4/UVO��8�8�T�A�Ҧ��p.	�%���)�����:M4�5���̦�h�Mf�z�f����K�pX�E��Z@�&��tV�~}/�\�Zb�GC;	�`�[3��jj��o�f6�n��$��adP�·Q�Y�.V�<�ƥ��Ѳ\iX,���k�8p�Z������7�#��wَF�ؕV�h/ ��+օ
��E������^�����>)/6��E�g�_;3��aw{��sd��Aw��b����B΃�r>+���O�ѓgO������/wt���%��zVW9-Id�A�(T:y���W��D����$6/��J�sb�˯��w߉��]��������_�v=�7��E<�X��l N�2��O��W�պ���p�B����kg�.!�/{@Ip?��ɍ�����P�&�$�R�eϰ ��0�/�8��ٿ5Q}�$�c��ɃpB*��UPP$,r ���ߚSʙ�]�#}���S���l��kΧZ#�p��������8�J�jd�0p3�ݓ{-�C����L��䓶�3�5�͓S�<�XT:^� H�t���[�-��g,�<�?Q��0Y*�U#Z`!b5 &�qS��3����l�wPIo���l` Jq�o8i{�� �8�U�*�cS+R��eeY��$>�t���!Q������u�\5W髄%(�c�-�AB7j�A���p�!���}Qu8�4�j5�$�R;���l]������ B�ͬ�T���H�u<�1��*=��3�8%��fhR�B�w_"�bi���Ym��,q,y8J�Q�B�8%,�[�����ś���0��Er��f�[��򮠝A��4H���������3�_�&�,��ܪ�}�RC�p�G6D�3M?�6t_��U(h�����R��d�f��1��@�W~,ɣ8<����e|��VT����r%0�Dex�DT{�p'���b�����
m_�._EU������&IqV>x�ΰŅ6H�WkJ!M�;�4�����C�-�рK���ى��>J^�3'Hf4x��)����-X؞���O���/���K�� 
R.'@�:�DV�ж�\���q����,����eI{yrHNQ��?��~����?Q}��`CQ���T������T�S$ȲhF�Xaq츜�^���~}�=���?���70��.m���h�q��� @��s���we6q;$QkT	�W�#rp�2�� �$DG�[#4S�P���@^.�Т,��ܕ��)p�j�ae�U�S�@UU2��$.F���K���Ōc�h6^�.͹f�H���R�h�91F�p `?aCT	����Ų�X��nAmu 㐯�>&S�2��t�T2�4r@X�����|���I� ��.�`B��f�=��8sG;���,B�4q4I���G�*�XN�� &;	t������5 g£�B͘�!������%J���b�VL:�\���-~�c�`�*�ϖX����zFj0W�)�9�M[W��<���D:9Od9P�>��1�w���l�D�Z��F�1��a3!��<7Cݨ���,H�g+��Y�f�e{�uhL�c����i�W����ܲ�~"9e�i2a;'�(��3�6���0>!�w
����b�c���Sp�T`�AmުB �e��j{NQ�"��28M�'�3(�)Ƌ ��y��y[�Ci4���08�"p4L�0Z��+	�zus%���ő�9{��Xi�t��>x�fRt�Jw�e��R0k^p���t#�E� ������K���[fC2�m��d��2=,[��8��Y���l�d=����� f�9OK���n/�k5nN�Xn���Չ|�Cj��4`�=S��_��
��x�g�̼�g�J��׿���fY��7q<�W�� l���P��q��ޒ�KjUdQ�SN>���������ǿ��^��J)��������������}�=[��cWt��:{'�����?�[%�@�0��4K�Kw��:�D��E��-F��ⴰ+�Q�r)��
U-�[]R��7���-o=�ʬEb0*�����h3�� "�Qԭ�/]� ���l/��,���{})��d�1ԃ�� � �ah�̈}�I�ιF�|L���ݺ�viH��Q0�����ּ�2] k:%���N�����5����>�ִB2.t��K�[Q�( eE/(� ��Q��9j��(}g#�KT��&ݢ��k�9�vem���h�i7�6���n��z[�vWf'�`[��$U�7�8=�I���h9�,��](,�` [,B�+���A�d1�f���m���F ��P��\�� �,h) � Fq�$��BC�<��=g͊A��$��������$t��mia:�Ty¼�����ھҔ9y�8�ä��l�̃�_֎����C�Nt���o�ӻ��$��:3�x�>��H�Y�i�J)k-��i!o��פ����'��M���b�b�1foYp;�%��0�B�+��{1=@c��)GK:�L �ʅ��&�?,	�Z������`�/����Z���T�b/6��aG���;&\5'����+�$�*�h� ����|�bLۤC���hi�$Id��نb-��y,"��!5H0T4����n9��v������U��ò�^>F��|��H��^9 �JÔ�1B�F(G:���$2�h�{��MwD�����[	�!����ǻ;z��O�l/�q�,���^x����D���D�Y��͸�	Z�k�HH�ىr��
��Nqf�Ӽ��M��ߧ����D b�[)�Q���?w'�� ���1#%Hi�(U��i�T"��� �`+V���]$"P1���!��i3�^C�����������[�@r+�[�]�-����5Х���w:��O�b��]��W��� ƙ�u� �2$#�4�c�u�N,���P�����<W���Z��џW�����nM�Z����_�Av�Fos{��Js�?��S�͋�� �rAɉܡ¾�`�Z�p�gU��;�H��Q��=P����I�����t�fsV!;�L��3"��at[�՜^�}qO��(N�����Ьq�$������ǉ�8q�QK�Ց� ]�K�s����{��	������!%`|0O���0(1�T�ű�q�X^'�3)@`U��(Y7���TICs��������F�}�^�)�B�it:D ��l�YU����9Bd0!�+b�m$�xm�ø'n?Ri��ݛ�r���W����S]�����Q�`*G�։�k�Pt�s+������|�t.�q"�=�MՃnW3��-���c ����@�>���7�nr� ���%4~MC#Jߵ�:ٜZI�+��q��v��*���$��#^�$�q�MR�_rgu�H��ԫ�Z�dX����j�Xi�'�,D��ӧTP&�K�޽��גjp}4<�$�j��n��`@�vt��
5%IgA�C�P��b٤����b�'/��_�x�h��@6�	�WBUmI���TsP)%�au�(�]ƺ�)P�!?Ic��%�xs��_ �*j�Y�!�x�S�3^���:H��(�4�M��s�3�P"���qA��B帢
0�5���.�C�郍B��\g�4~���@%�Ayip�X�!�P\͈��X��F��y@�2�1�Mƽ�����5�8A�*��k��W����њ����,a�d;̙��[���j�"� h�C��������W��1)�4��n��'��~��H�Or�v#(���h�l�}�4*����)�sx�`�z��Mb�iKɼ6ٓ�J�xq�:���@�o8�ba�ɣ��Ѥ~�ꖜ�UspJ��A��q�qM%�*���X�@q�����CO���u���o��q,��w߈��~_�[�m��r@���xr�v�z�p�&0]w�r���(;X�:�����r2}¡bo	|�g8H��߂�m���d}����	��)^,U�Iʨ8� ��*}�3�W+++�WWv���f���&��ATz��a��q�Ȣ֏ �z���t����&�����#���Wm�!�pJI�2B̰��^W��0H �YO7��W�Z) Q�E�� ���O�|��@,rm��bjR��̖KSſ���������aI�jAS6dwWV���+N&1���z�(luHI�A�($iu�g 	�#��lQ5� ��"����i{B-�
�`�u�$�7|�� *K4���8��8���X[5��j)|4,t��6 @_�` �5�7֪���R ��d����5��������>b��{	������-∕�e�יp�h�l�IE���7��.���)?G~ Ҿ�1Nx��N3=�+���`/��L��%Hm��o����f�:�(�ҹ��^��|0�kC����R�'�j�������X3z!��o���'��*����rЛ�m�M��eiX�ٌ��+�OS4�c)�=�`r���JǬ�]Hasċ�ЩYS�-%���t�lTϥqf
���I\"�XO�UU�ɪ�!��R�am���l�7�����j7�X( <kb����>����H��Ir ��J�V��C����ǘ�H��x신��/� �+��^ʂ�VK9=; @0 *=ɉ��������䇀v�ǾXm��*���Ԍ��!Q��#�U�XBZq����F%oM5/�G�W��o�cE4K��φ��a�;�O�$01��2���?����$�[n�]�z�(_�4T���؞�Õmd5�(��YS,���x@�A�ެ�����']�TP�
�+�ޕ7�{�I�,��_~Eww���;��u��}F_���B���?Ѽ�-{e+������B��9y�����!���_�[�*t֐�׌�ť�^|j �H,"�{�d2�������.�,���}Yj��AU8���ݗ�F	pU��
c��4�M ���&�%d:㖊� !��k7�P�[**_j�*�ь�\�qPG����A���5�Oû�B-�c	��=��z:$�ddE�5xwj@�bF�8@D˵U����b� ��>e�d���ȁLb2��P�{���,�{$י�j�].��qg�P��U<;]���\[����SnJ��0|L	l�)>h[^[���,,�GJ7g%�n�M5U���<��(�� �������l�T���M��L�*�����D��ż�!�����a�-����i�Y�LT^�8Nq d�-3� 'r%!�X��괁|�mSZ�~"ܘ�Zr�η���Sq|� i,�;���H���'��R7v\Xx�ì1Ύb�V-o)Y:.%_������צ�-k&̄�5IWB�<���\��F����v�+����c�:������U�+ ��k�w\u�[dU9�{F��iɚ)�v�q�T*�Z��[�r4��u�{����1�-�9��+�����6Z@c'�%��8S�܀_;KD���@~2��wa8��KV�lF��dga�u���>�8i�[��'[�I��E�͛�~��������W�{O���D9~���W_���s�s�Bۺ����.�)6��Z��P�h�f�Z��b�!+�yH�Ę,��fBj��Z)q�v��}nN�i�0�\pri�Z{�|�c�,R7���j�R-��%�굚'��7��=r��s:;���+��T���&�a>ze�%${ K
<j�U�!f��x[5~w1�
�Vb<��CE��I$��Ġ˪�\/)�����Zh`~�!���#�6K텽�N(�((!���� ��C�L	;����c����m��Qc��r�;ԍ�KSS� �q���ۧX�e��P��`\�lT[^%�q�2���;;��l�CA�����`�Z�V	 �k&� '[d�[:l�������+H�f��0�`�l��*M+d�ɵ:*�l.���&Ci�����Gt  X+��	lV$���ǉ�9H7��T�4\�ʬ�F�jV��H�T]))�P���$���0P55��&���8�B@7�9j
>V�H���QI�z Xl�g�������+;��U��9�&�B��+�r��PO����]���
j�M���,ɭ��*��a@i���)�
��]O��r�m�8�a!Jմ��{�U� Vܙ7�y`w���N���NiY���ㄉl�3~bL�@��@���]��Y���Z ��3���?�Kn]ƈ��>yrK�����+f5��d.F�&y� �hQ�2�4���`��1�0~��q,�~1��0�"z~�U������R��%=\��*hB��<�FE�1���;���*���eR/W�b����� �f��6#}JX�	IuU�m}Asj�38 �^��-�"�q�!pAF���c;Y\6��AB���o���5T�Z�\���܎���@d4�um�C#� �-�H76��z����jk� �]L�kc������Ђ�-�V#7ه6ѿb���~��f&F�lD�~{����4�����B=L6VM��ZJ��@kX5�JK�~���]�9�$6v��`6����<�tCZQ-�X���<$�j�h�S R�������Ɉ=��*mz�쉔����������5*\��h&$C�� ���)�&Y[���Y:�U$���%�	b�/>��'�����i�[.b�#�xn��~5�U�>�QiQ���]��Җ9��O_� G����u���;��9�"��#W�@��5����(9Ϧ�܄E�����YT�2w���6�XGT�>d궋/ۛ�(����êS h@�D3c����{��AoM-@@q%�˃�$*�ܢ8i���I��+���;yi�+��v<r�բ����k�*1��!WX1��@i�Q��k�\>E��;N����In�Y"���8��RS|8ء��00R��>3�Fy�z�R�/6r�'`�7BC�нRl����T��|��Ԏ�.�i�c�:��`�%�i;�^~�6�tGbr%����}v���`�9��U�U0����8a��t-�R�܋�����ĥظ� �Ьnj7]���/�-��D�MO�(���B����BƷ�Pd╥J-���YZs����SH[J���������`H��W�WVs���ǩ}>�MtTK�L�-�Ǵ�]�eC]�v���Ad�\�4��_���a�?š$3��ޝK7O�I�/�[�Nhk1'#~�Φ6�`8���1kңx���}��6V�`� �.����>CG@�p�Җ�}Ȋ��%d?[�3��ȻY�1Gsc�$�@���I����P��؞j0�~�0/��7�E��� ��;Iْ`{Nա����A�j�WF��ԭ��@D������GI8��_��ŝ���k죿6i��p�=��I�L2)k���6f6� LL<O���L�ֹM��p�.�,Ӿ�d�?�=����%['�����{�h��)���1�D�.�%���L��e��$:Y��Be����H'n������*q�]N9��r/��r���$�f D'm��ռ��p�"t�t���y��l�U�rJdC��tbS�"8ME��l��F1��i�9�4�� �Iަ>� ##�U�&�����ˌ��䀅ܳ/��[�96����$a!��4HUz����z�WfH��!�iYN�k�V��nT�XQ�%'�2�0\nB���ڣ�4��n�1F۝@<$DR����3s~��C����G1�P3&�D�U�Ge	���`�-��7>��$龻Gc�6k5��s�ܼ��5�)C��m��0����~b����c�5@�ǯYuA��Zپ֚�%:)��֕޶qH���7:ť�Ŭ�ǽ�+�Kg�� T����C[|0F��V�G�ZMb����,����9%��>�$�%�sw�q��?pT37�|�	���7�3c��[$�ϕ��%҂�ٲH��l�V5��N�JVp�:MCQ)��x�����ȹ���C�m0�����W��E�V���l����I�Q��s���B���J���ү�����I�s~N$��fN���(�ռ���lbl\i�m���W�0�:I@s�b�	� ���t�u��X�v(m�سk��Zo��4�lß�O=�A��y��s)��ײ���t5���2�,�=���'�/��x*�EQ��o	1x��¬Ķr:��S���Q�!0T��橷���D챚��� ����Ϊ9)��)c�� ��Ĉr� ������D�HSC�1mܒ�u�ާ�4���՗*��a�2Pt"�1�7�X��J�œ�!�B���5�������o�(OE�)����u��!bPQ6%h��QM��~�̍4���7/"C����Z5r�P3u3����K�x�0�PR�n�����[�R����&���Ur/|9� v�J8��N��J��t{���4��1��l�$b~������~��Eo[��*��6fz^�kK@��
�n��cI�zz����ƥ�֭$��pFA��+��XםZ��3�J��ď�����NM��uM�TO�F!X@q
:-`3�F�K��W# �vK�&>�\w0� ������1s�~7qE~�l+	Id!�}��X���Y�K9�/|�p8, �^�ϧ��?O4_E(S�{ʼ"͛����
���^��@S��5K��I
 l2	��N�"�}�@;&���~�7d!�5q���*���ݚט�^�x�L�pĮ���1����V�����G1+��v]�Ӭ��8!(�͒07$ �+���n�i�,��;L��{�I�Ԉ��j�M�����E:t'����7�8i�c ����'�8%ЯJD8�v�����������$	�v0�$;^J�����VqohG�5H0����6d5��U�؆�`/u�I)�u�ޯ�ۃDfh���������'ԣ`�.i,1nD�܂)\`��>Gi|c�F��Ѝ�PK�����4Ot_���m�np���E絕\D�3���1W����+Y�������&A�1��G��~ �|�>��l�|�`�_ZI��Tj�E�c0cL�$u�C�
�ll�Y1�}��恬��������'�C�US;W�jřo���b��K��@����m��aZ�]�e���+J�k��Jy�Y�.]#,���k�?�{C�����j���s����,�a��N�0KO���@��?����Q�tZ>�h��Y8��y��!F��~������4��I�<[=���e�6z�+�jj�I��gIWx�~��l�]M�88y`$�8rG����\���p�ԧ�d�~��/�I��1� ��E�x6���x*r��r�[v琞�mW�Dg��?�����PIԙ�O�J�l�P<�3$�tKb !'� ��|�~*�w��G��cg�a# 5�-�4S�4Ƣ0�o���'�]1Z�����Q֔�mУf��q:���W���\�6���GR/���r�.�	�_;����n�tk�&�b�ۈHl���U�*䌧Z�;�M~2Ds�i#�"�ab싗�*us@ry9T��M�#��ǆ��%>_ ��W��KZ�X7�Sk�\����Gݨ�`��9��K�Y�[�l�C+Mt)Zޓ`����=<�^�\�%�l@_c���e�´�a-e�ݾ_������uss��%ݓ�C�\I�!��3�	_4��sM���%٣{m��l}�w�^?X�6 �Ľ: k���*�.����^c<3 ��NM��o��".1���J$&<*�{8�����'*�D�Áv�{���,p�*���7���bf�$�պ�ڠg#����-���P\� �1�E�N	 L�%�����&ֆ��Ƽe5A�6�v_ԝ�_;�J�˨#�I�W��j�IQP#��M�=��bQH�������2w_JL~�h�6�����O��!�x�ӄD�E��|/���D��I�j�4�ސR���,�Y=z0���s��`��~F"�,G��u��S2&%�L����A��j��٬޸�c>���ڿ}�e�	"ނ����_���~�k��R)�u��������{�H�D�_�5��8��ewCZJ{z��,�^�O�M.����n�a6�/1%�Y]+iD���@ێ���dn�Ӛ%|�����o9�G^;������]hlil	\�1��X�k����@���k��l�/ss��+��h����5��.�1�����,��t��[!i��7ZH�S����bo����&������.Ӹ�g�:��.�=X7ZY8�� �N�3�[% �<��@�Q���4n�ṇ��8gzww���1��L�zb�2�"8����ٺ�K�8�.�������<{��p|�Uǹ��z`��Ý�d�%�B�ɀ���:�%ߦd���$�j�mڈj��(�=�(�U>���պ�D��q�d��Mtig�Y@J���L4��I���E�������1�O餳67E�¨՗��t��F�s�L������vb���Q"����f��X+���-�_+a[~Q�"��9�3^[ꮯ��2�"�����	�:#�	�6�
�Gm26����ݪ��V�6�,��ރ�����`i5���^�\�D	'` �T��U���"%�Y��j���-��<]K�������-�����,�ؾ�����<���\l��I�ق�5�د��j|7�x��k�`۫�mĻqT�t�JS����� kkޢ���]/��~pnе�z�k}��:��/�o����[j��@Ÿ��:�E� 3��L�|y
��.s�Q:�B����=���(���㱲������\���w�뎞ގ���̀������^�I9�����	��#�i'٘��	H����5��  �~� '�W:ivg����	��Q���ql�v�:��;L��f�g������%�+����:[��=�ik(϶!s���'��fh�)�¬~#�&h@h���n�瓢\����8ב~��}�������UR��<�ڠ��#)�^uX�EA8�&��XͷH��p�&HI��G���}����{�QZ��w�����Jo�>(��T�DnHI����������_jC���	�1Q��� Q���y���(�RnG��8�͗��$:��j�-���4�ɍ���;���xf��}��B��������|�-���nշu�����H��l���XJIsp�=[�ؾ�՟���],�z4׻�!��Km�-�_?�F���`��1�k ��s���Z݀�|0O�A�K�Ǭ�[1Ν��{�q�7�Z�o���۲4L�fZ4�ь�Lb���Xe0���ݵx����[������L�zX��R���o�1���Sb�q,_)����Ѹ�hO��K�9��� �{{h>H\0J���Jr7�pv8
O�]�/��PR���9*�e�^��ϟS7k��[b9�4:�$Hr��
�d�!��iW��$�n��Yc����aز��%�y��na�9���-f�A�N�\H�ʶ_�����|G���{QCC$�%E�ΑH�ě�Y#zw����X�TKx<���ڂhª��h�Z�z��H���������0�0�߷ʱG.�ն�]��/�b���G���KlC�۷�$Y�q�x�{Z�2������.����V\�$F�*,QC� լ�m�Y�7�?�u���b8�k����`>x&����2~��F*+���?���)�ڞ~wr��v �X�����)�M��*y�����!�HX���ԅ[�n6�o��#��^�-�[���oT�����үv/��*<k�wSVh�Z�Sw���W�F�wrO�1p�T�|g�s����C�-�)���P�zV���6�%�q
'F:�_�k	���O��������l��'R��;���^�t<Kڧa���u�:s�B���o�j�9+��Tcǒ��%Z�r�O�O
���pb5� ˓�i5[��/}���TKտ"Cڎ�v�J�w1Sf��
J�V�d$��Y: �0@���f�>�be�xZP&�+GNG� ]F�Ot���"��BB�bnZ�Qnl'��f�7��L��ƪY�c�ׯ�����������#�v����r-��&����	,�v󋵗$���w]��#�&r�(����A�3q�m冡���y/�v��=T��Fm�e�e���Z: Ѓ��&0����][R�ͭ��"�4��7W7�7.���O4�]��T�V�K7���ފ�Pk?�f������0�h�����)��&��w}:�!��Xv̱_ݶ��i��W㗹C�ܶ7�
������S�ȏ:lPbJ	����#{�(�^�w��k�,[�æ��x=�ծB�x��|��*º"�i'@��v�Ź�$��8���_�E��JMy�^pد��SJ#r�=��� ��T�	��c]`�]R5�H�HBM�2���7g~>sb���;v����q8�x�3�ގ�/��{��>��O��v\x�J������ۅ����5K�n��g�=�f͂��<&K�L�5�N"���R�k�8C�e���ի�,̅����>.�[��x!��\��- ��i�xGT�~\w���o��+��f�N��I8 C�S�����h<(�s|����OJ���ҁ�p�&�v�6y^5e��1����u��x�8O�~��|>�۷����H��������_,�]P핼�ݵ �3{tL����r�
�P� $�Y�0n�=���"��V�#F��1��P���26	`b6 C	��V`�"I]��6���^�d��n��- {þ/ ��;49�#�� ,�z��R�Z�!�\����Ȓ�f>�d)��f�޷�z�RiΥ��l�lz�������-	�����۰�,��I巒V����L�!�G�έi����Ee��K}Z�!><V���>J2�sMb��v���Jsܽ��ܨ�?|n�tcoo�Mu"։�O��5(%����-����!�/J���'��%��m�2����y�:�������Z�&"A! �4?4�!�N8�~G�~��_��gODj�_^�N��9Yx�����̙�ʋw�{H��4��ܶ�<���j�D 4�d�09�L�E�T�9l�rjb;!2�:�l7c}��Xh�<��-��?��Nq���8�*[�ݼ8_�<���Qn��'��`L���, f�i�j�~v���\K�J�]a|� ���ۣ��fz��qV�9�ԇ���������O�_^����׷�]&�x�4�����:��R@���kA�����~IDޛ��V���=w���1.���w��OMؤ��M�@P�e�M�:����B�llp��i�[��7��w]�;BDv5�I[CU�V��ޘ��?��4�nKS��khNZ|>�a	�0�����͏��%]�ZK{��~3�jϥ�ׯ�~�|z{�ϯ����>T���y<�ZR��V�2j��Զ|��[�I�t�S�h�Wi�[Izi=�J���ƣ�۾���f���O4ચ,��dd�E�w~��M�G�/n��_��pc}�')�0�����NCQL�N��|�ѫ�_Ӌ�����d�93C5��A2����P��|/Ұ��^���'4\])�3�5[�5�b�N\Ɓf�űHc�b[����N���JU{' yS���H��$$�[�ubA�Rް`�q�
W���{$x�hqN�G�2�Y����d�TʼI�^lT����%IC�=��l���IU30�4k�Ӣq��8��R�$��I�k�j 'M����PD�Y�2+@d��ĢF�tx�vVm�=��_�ҟ�������|9���,x�f���8z� ��N'�.Ϲ�$Ő4t �Q�c̒�=K�j>Ɂ���!o+�SAT������pP�|��%qa��t�Ѡ���A�[�{��b]����3�D�;&����~�:�I���i�pBC�oz�R��=�✆�E�I7śP���j��\�	\��h�m�.��~-���Aci��d�es']馡Q��{Zf�q���4������ъ��X��V̓��y�� 9KV+Nk��KG���W_XoJ��0v��;�cj��v�v��{Z�� �܎����n��D'�f�4��>��)
m�}]/��%�{хԀ����6 y�ά�`G2q
�jܓ:g4��]��q�o��#]s(��r`7�[�q.�I!�iq�>5�9��pϠfl��PJ�ޔ9���~<���A�B;�-8<{=J��n�a�}ȱLծ��m���	\`�1&*�シ�q܋�$K�D"��;�FlG>1NN��E0?��AB�%n��҃zZ�w�n��J$i��IP5��R���;�us� ǥ���%�`�Ӭ�g���;U�&1����F��9��r����Y����w���|O?��f�+�y�v�O�A��"��륝���n*�	��|�(��pb��
�R���*�h�D�@{~�j!T\�]16#�)�M3��oh%��	�0T/�ZIfJq�LM��0��{ܟW�fd��rj�H�MuKi,���T{8\X���{�V��)eu�,��z�s����P�X�?�-`Դ��h	��0ޒ \:�g�n��B[�?*[�o����@�{4���j�[3��)�?��K������d�`��m0��?�6����+�vv�H��ȴ�vb��4�r��7W�UQ��ߙ�~D;u��&o&��AUCՐ��x�K�蠛�߽6�P��175��j�o2�ڇ���a��锊��y�yR_H.; 30��Z ɓ�/{Z����t|O7�#]￤'��8* c@�%6I�-���~������L�k���h�8��n\*6[&� {Z9�~��
`R ���j�̚��b ���p[]l�6!.���b-k��}�ܾ,���^p����u+6b����9u�#�w��UU�+
��t1��zz	�/;� Tד�2:�#��qgO�'�~A���W״���t��e�e]���5!��Ig��&������]����{a,��>Uz�����������w���o���D�5��gʾ�YNA��C�s���f�`a���Lg��p�������)_Ӗ���KK��$�1ݤ_�C"�ا�
tS�	X��K��s��'�QG�0�>���`��&��8.|�W;U��$Q�J����'l�ڦ��k ���PxX�?Vc�C[g��=�N�ü�`.3�v���������j�|�3ͽ=�ٺ'U����iu]Ry?<��J�����47�KJ����K��b�a������۞�R�4ёP�S7� ����|h!�;^��i?�:=�Ôl�(��Uћ�=7�	�ã��Ć@������2�\��ѵl�!�����ɢh��:K��q��:��:�{�@���*K�~~�+��ԗ_���D����غQ)#)0�0L�
Z��{'����ow��~������٪{�g��0P���9ڀ��Y#�[���~HNx-1�>\���f����7ؤ�Z�v,�a�� �Qg_/��"d�
7��<{���qA�Z�ҙ�{�n����׸Z�$���,��3{�}�0����b������{������z��=y�tA����4=�fF��L؍�(w[ߒ~s���A����x:ʊd��^�����3��O�.�kA�{�A�v_�k� 6 �K`V�S�f�\
f�<�'�,���F��iS`#Ue�A?dIh�N ��I��+����\����@f�+�
z��Ji�J/m����$��`�,���L�9p�����h|�j��a��@��$ �TDN-���}�87|Hv_�t�&(�j��M���	ںo�h>��g��צt+����_*�`^��?vm٩�g�E�ڼ��~ͷ�4e�� R?�ף��h�Ǐ�>_����U
��W��s����qzb�䛛v:��4%Փn�\�j��ﭔ*�j�JIU���^����~x���̋��HH��Q�81�&����/|��q�|��+zw�������zwE7�O�;h�t�`�$��*�q[{�z1 ��k�;0��$����3>5{��{]@<f�\�|�+�ب�d��������W�lߦ�Y�{�~��w��T���]�$��#��V@��Ie0#Fg���5��c� L��O��l���OL9��3BF�I���$�^ �Y�I\E�����lx�^���EO	�,�.x����j Rr9Mҷw����O�П��w�뷯��/�� �|Ց_�Z>{6����V��g�[�|7�k���y�m�t���@ _��)�}R�. ��ۊN�؆�Fu��+Z��!~��<�@$U��)lpb��R�v�������^��?

Z0��h�H8��~�g���3�4��H ɹ����������1^�wL��=�����{6���֏����i�M��,a��A�m�)�gJ�C�oK��u��ɪ��f�����v8S	뵽�XZ�}�DKw��%x^�jkax��mH-���~G��z��G�*
������F}?�3�
����ѫk�!��68wh�f��uW�N�2T4W��x�k�-=����r���JԜS���@_2�Cx�ςd��1>�u��n��(ۈ��3�@?�rG��gz������>{~KOn���$I�r�Y����av�Q�i�+(��Z%�|����R)�F�Ici
���x����o��lV0�Μ��rNc��'	-T�� ̥���Q�a�Ș���o�ю���L����N��P̳������؈�r9
2=- L��ޛ��K:(�`���֖� L���Uƀ��:@������=�{�Z�	X�	��:���e���]/���%邖	���ǃ�ivc��G���/������������^b���d��z��v7Oi\yv�~��l^R��E�O��ͫm[c��>��g�w�!�g�@���:#�a;I>OJ"�K��j�n\��F_4B�����`?'ZM��d)bH��k�jH� ��&�d�g�<�j�F�ӷ� X*-S�?[h�bB�;�����KgCR���_��C:G	�)��Мv�"�q�a=��	��ħ{�s̹hP��  ��IDATU���N����4�;=Y��n�}�-�����	ܶ#ҏ���Gm[|�8�m$L�v���TEa��U��F��6J�=�%u�%YF�����=\�1��Ʃ����k���Yn#�W�w=l�����i/��(��66�=��>*�,N����Ǒp`��������7+�BH�j���gSeFaNu�^F[��T_cR�8���k�a&�e5��M�ʗ���� j�Rg��`kl�b����J�aV�=Kî8��Y�V @��.@�\�������������k���_�W�����y���������$�8(P�����,Z�Z��)���tP�1���#�n�{�,c���U�uM��i�}�,9��ٜ�Tpu��xhw��DW`@���[ د�,,���@�߽ ���K�(�U<X��{r+�U*���y>��%4V9:I���v�;'�i 2����lQ��s�(�OUb�@�:Px!��j�Z�]��h�!-��� �eԝx+@���{�����O��?�����:������'�X=��F�_=oH��Xz֝:b��-�xY���VD��e��
�\��G�����(�	Y�K�T�|�(ͷ  `�^�P�4�O�q��?o�nA4����9E?�+wrI�ߟ����,�i#9�+w���Uk�km�B���\�^i{���Q�Z#�m�Z����g����1�U�}&z	,�4��3����p��Sӛ���+��/����u���姿{�F���5^�Oe$H�׌�l�~5L-�����Z�2څ���vk���l�R�[�,�_-�����QDܦ�@�jH���Ȏ`6;����5���zi��� =��z.!b4�1�p�Z� ��־ݹԞٗ
ފ���$߮B�D3�b��:_	H�`��R[��?���W����H��D�����gz��v���,�Z��(�y*��̆K�IY���f��\�b��6�ɀ�i���U}i��<���i�d�O��������fs$�i�^V��}wG�^�  l�����_�zǱ�Nt~xO��z�K��ݠg��|���0�=I���T�pm6�/H�b��Dg� `� �9yTdY�#��/�s���a� fA�����k����`��tX+��i'��r���o������ͻ:�;$��SQ?��Փ�_^������ª@DیC�-��o����
`�g��!tk��m6�
۠`�Dȼ^u`kG��@��O���Ww���
AjC�>�㒍�%;��Zn&�k���d�	Q2Y�V�W_4�<�62$e�,�k(A?ʆ�y��g�]���cݾO����g/�iϠV�L�n�V^��c�ٲ5���ԯ鏵�rF��}��hϑӁ���%3�K�o����T>z�}��~��ZiƱV_{�k|�_M���ގr�Z�c�����Yn��� �$Q~���ѝ�rT�>j4���o	����+��������� _��,)����v`)��i���QŨ~�l���$�F��>������_�Ͽ��?|�9����{JO�\��El��DJ�]�˜���|T�B�5ި��"5�'5R`�C�	x����,fC�gB���0fN1Na���'��t�� �������oN�����g�0=�q:�-��;��������y/h��p4=,?��&ޫ�j�r\sή�䂐������@T��d�@*�?@A1�
q+D�dbV�x=,�8r�w��y`ߊ䋍�i�U/���l- ld ���k5�� r'��z^�p�`��|�
���c�:��o�vxZ[=Aĉ,K�J�ɦ���+D�8=ĵ��W۴u�	 ��|���ڃ�\T���G�������+�3� ���SZM][���ݴ��o?��+��s�J����8A�Xm���z���^F���W��_��h]��y�a��������^��u	T�Ǡ���v�J�UQ�1�O-��lZ�}�C�ό:��<6�^�(�N����A�/���o��&(�=2[�FE]�hs����`̻�������	Z�� �|d{}�Syϕ���:���50R����R=rPUӴ�����+���`�1�}*i#�*�da�Ŧ�C5\�DI�8l7%pm�8al�t��@�wr����~��������[�� |������qTA΋��l#>0�9CP��^�6YR�N�,q����0��YABm2�^͹@� ;�U�����������YVV��?���Á�߳-;���p�����޿}-��l8π�ɓ�쳗���Kz���R�2X�ú�VC����aQZ�
ƕ!���DN!X.E��Jl���Ε�=��6N#'�`i�n9��ai�O��a]?��3}�����������G��[S7��=/�q؉+}�V����kR���F{X�� �f�K�3���T#m_�㚑l�ql�d��Ȅ=����M2!{�?6�-�II��1��4r5,�)���w���!���r+��x�yKD��������4�s�e�sm?h=�vC^���D�ɴ-�hS%�7"�6Y�][R.g	e���ؼ����X��)���%C�-��/򞬫G�s6�->�.�H�$l���d�C$C[�<�$e�@�G�x�x���81�(���@�6���je���!5m��Զ9����o҈�"��sz�$0���ڶ)Qƃ��&�V��BP�š����ߥ4�ذ��ec�|9&	|AL��)�<4Y2��W�P�϶t�A�������x������r�_�������=����/�, �9�|������^<#wtu���UW�QCR�ڡ	q��ҿ�r��͵���N��� �?�c&�&A���HܱݨX@$_��u��Z���P>Ntf�PR���|�_��z��W:��5�0N�7�r�Y���b'v0�A@V�lq��>|c��k�Y#��;K��TA�9^	uuhE�1��=[&��X��q�sM��{�����w��?���Ͽ���_��{�%��]��`���������� ��4�������7_c��i+>$6�.>��&}�ݑwj���E�`�P" ��m1Z�{:i������yϠ}���t݉z7:�&��_�������o��X7"��d�U���ZI�|��<��7+��~��`�6n���@�&2c_��/�����E���3���RQ~�������� OƝ��P�Ps?��e��?ƶ$_[�o][�����&H��,����o��,l��m���oH?*rY��<Εߧi�m�?��J�0� )��O*x5��ڋ�~�1�af���l�̖ɞ�CZ�Dzq�X`���Uh�k���`|B�3Xw����3���$���Vvƛ�D�糄�8��-`k�7��ӳ_����wt{}C��������%v�NT���Հ�g�PA����Z�l�ZT���>��3&�s�W��-���q2��K�8L�ҏ�w�O�f�.�r�\�v�@�1���$,?gg�*���/@�<�!<s��T�`0�G"��ڬ+`� ��^�1��g2�fൠ��2�zB�;��p��EG�%S�N*Ve�����駟�������?�Z��� F��aAͷW�CN�u'�k�b��F�_ 8�Otu֠�n/ ��;vj`���=e��S:�a���Apv92�l[^�kʱs����M�(����ʛK�#���@꒤�g% i~�a�u��G!>�_����^�:�:Q/&��t]+'�[�7w���y�1��o��u�[���+�aK�1�fu٧\��K�L������z��Z��H�n[��X����l��I�.}�۱��>^z���m�W?�c�f���[��P BP$�O�7����T>�U��N�I�0��'$�
�$�"��q~,@Y-���Q7ny�|�$���Uۥ|�B;T�N}��.��Y��[x*㉙��Y^�x'���]��:$i�NtX�=�=�O?�I
�B�w�����$�vI��b�j_�~,�BU04����t�^h�xp\?�cyƝJ�v;M�-Y{��FE��c0*���`���*����i��y�޾{;���r2Kv&'�r�(R6	���0_����-C��R�p��FX�W{	������$�f0���#�x�b��� �z��_�ի���J��~-��v��Dr</��8*�b�F�IU$��"5��Ćs,���Ic�ل(�	�՟pUJ֮U_إ�W��.���qM�e F�^H㪿�����ZՒ�|����#ĺ]�`4��\E���oO豙�>��1�t�?��#utEx�o�Ӻ+���'[�]ۿ:c����|����&_������{�c\+��J��9��G��\Z�G�����܅�G����WjM���x�����*�}�ېl87���aZeՃ����Ǯ�P���Qi|�;���h��7`m�^	�d^��s��6�/D-$���]�>��R'���o-�f��*���"��V�{JV��W�X�_����A��~paB�l��!�Vn˜ؒ�c������-@l���:.���8�8i<�򽄴�VUN���~Z@�$`N5jGr�������%�R���/}i,�Ɏ\�:�ܮq�Y��:M�� &��4�	����2�m�r� 66����]=o�
�y8}��[���A��p���S�L3���f�wK<,���Kҗ��׍��p8Ed'�=�)a�[R�z�����p'�p\ $�ǋ�m�n�_�N$l{Z����k�<����'"�b/HN5�t[l���B���o��b)M,��ۄ�T1���!5�9��G5�V�Ƒ��U� Mt:[����ʰj�y���ɲH>d�0��=3��{�Pb*'�M�ա�K'�K�Grp�h}�B1݃���yj��@Al.�ej�u�uu�Wc.��C��Pɖ�D�Q���o>Gv��^�ѳ�{0�ͯ�J'�8O��O�4�z��̀{v�tq�|����0�}�a��BJ�gۥ�% l����n��t]RC��/�-���j渧����=Ϋ�s9�Fy9��mЏ�X��1�VS��Ki��COJ�XS���dhփQ�m��̀��1�!�i uS'_x�Z+�<�hl��BԖ�
P̵x���zۃ�����DNV��\ ������,���N�?t:����$��c�J4��Z��% ���hʕ�G�N)}TmX�8g� ��<����K�Mɚa�]m�J��-8c%V�
ɣʞ�l�v}#x�����)AF�%t����kɵt�K�t�ދX�x���;+ �&��`c��+��XY����1���Xd��p�,:���H�P� SP" �j�2����]��ͭ�.�ܿq�Aa���}Wn� �z&�_�f�%_��Ug)%}�6 ?I��,|���I#6UKEp�j�U�h�za���g	!bPH� �*�
y��w� ��>�2�V�b���N�=�ߢ����X��Ɔټ��%�	[`��u��L��1�<�^�3���-�ߺ����1���g�/k����Z6����X㝤�n�[�����cQt���t?�%P�r��<���HXa��YǚA�̜:��岚{k�[0B��!�.?���c�[�q[�^{�4�µ�����L���{�5��Z� ����H��B-~ݢ�m���+�X=�MbD0(Q���فm`5��'5I�d�?G�j�حJ���d�.��6_8엒vv"o��h�$5g�v�j�����&�9:6a��*L~J>K��A "׆�\bl_f�W��8 ��g�9��$�3bF�H��,��*��$o5�*��˵d������`3�~.γ�ǳ����x":�!:G�-t<�4���M8k� xF
���X�d��4�=߰�t���2�bϵ �QC`hN���ª#�K�fú�Ǳ���9bٸ�c��|�D;�+gf��yNW����P�%��H��ɞQZFC�&kǀ�#؈�-�낔S�ƒ�հp �JI�@Wɘ�b�/�:���c@�vT؋߶N�����;$t�������@�${��7�S/�#����:c����T��h�t�A�~�銂�Q�|�#�A���I�?�"�7]�8,WR�������X��YW���R{7������^W�ѽ��8~�S�ǀ��>������z?���.����v��~<��@�%)�O��
>i}�j��� ��d�TK$�"�,����2�:�5�CNk¹���yD��a�88-�'p��؉U�-�f��1/[������p��N�{1��2��A!�spZ奅4(���[s؝ϖH[%q���Oe�ɓl=� `�� ���PGkI4>�s�$���qZ��FL�*ۯ/�" �4�8sŕ���u8-`ly�`��$~����"h~aQQi�`Xl�Η��םE�����{:V���Su ��$p̂��PN�"[��"够������#�i����?�d�i�EN�\;�զ���s�`��ƅ�\��fg(H��I���+:g>��D�E*�<`\l$JH\��6�5���5a+�s��D�K����v�� �+�Bj͟� �ю�)��D5?bG��ت�����m���=�s˪k�W��a0��	��Ճ��.(�ڊ�h�WP����}����h�V���B믞!nH6늯��\}j�O�|߷��)o�<Z��m�TG��&�j���dN���t�����^x��hP���Ȑ)���\n����d��n������ǬC�Ľ͠�C�]�5��T�uj�#;7ey�'�FZ��}Î�d��Nm�b�z?�[�����G�7�"{4��Z6q�����L S��ʠ�1��ZL=*�fq&�����(F���aO�7X���SBhp
ĥia�0{~�ޞl�u������ۛ59�$ibj� �<��ꮞ����>P��������B�{�gz��23" �����T��<�g�*dD ��v��~zھ�Iϔf<��f�å��zb�b��V��M�T�)�:�9~b@Ï�&A�|�7W��8���:�a!X�����Z<]�
�� �I�n�Ez��#i2P����$�������果d��W����x�&zOS�>t�H.q;(�C�`�jA�[�.R��j'����ʂ8/P���:2S0�q � UK6�X���|sx�U�{�����c�j��5�Z��-���{%�(���9��3+A�����-,�.9�n�p�2���>>������%k�gH�޵�-��r�e" b!�� �����D�|Q��i��O��/yѿϡ���[�ˠ��럿p�v�/{�)+���k֯�ܽW�UF~]|��A{�U�y�H��:T�{?Nw�/����q���%���B�_��-�]��G��`#������\�1Q/��Y���UL(`Q�;�Dn�ue���j`��i��brێd�~���bg��[�ɔ~��m��d�K�����iY��^��p#p̳D=&����t����g�EOO��Do�+5b���f�8P��jy��(�'d�N6�E�%��Uc����� �N�i��;���ր=l���>X�0ə���&G-�A��vǍ5��@X��i%.�S��'&\>�ݔ�c��%-`X����l�5�>�bU��~^>%}1,��L����e�VvYj���ݔ�"��A�m)`?��m�1�h���$�Y����X���9Ĳj����7�ex|�ՉuK@���ͧ�cd� L�b��2V䣶^��A���
.�P+�{�E�#�\b�
q��/xe���C�
��?��Z��in/xd?�xu��B�w�!�U6�Ww�"�92�;m�w<�R�m���,��5+��[ǎ9&g,�ח�8|�5
͘����$E���u��Q Vi3�X�����t�v��kn���m_��t]s��k�	��\����ק�,1��^A+���^ џ<7����,n���|7���u�v{�n(y3~�u��c_��^1��w/?7g<
`$l� ����U>r�[� �����j��Y�l@���p*޺�=Y �^ ʒֆ��)�JtN�'Sc���
�&���nd��qs�r�,���jȀ�*�;x�Vޔ-�ҟa��N���O�)�pU��Pl��5L��O�����
��q�5�u� l�@m�ȭIp�t���V��d�21�tF\u�z���:}xz��g*,d	�p�՚M��a��Q�4�4M��\bB��H�D�,�AI�f�G2�T�����7���L��o�� �RRbu�!A���p	*�b|� �sOg��E�#9�b�)�Z�5���b����H�Qj�-f4�Ez���_%0���y"���w�M������kA���Sh��k�/�Ύ�~�ұ�$8 ��}���ψi�����Fc ���Q7���'��g�v�%ּ$��*�4V�Qv$3}o1-Ƌ/26������{Y@�/\���2/b쉒���%)�� �gY���]���.�/Ǔ�)���u�y�x��U{m>.Z� ��	��Y?v�K�]�l�������l���͒�as;�E����ة8P؎� UbW�����K� ��>����[<L:�����{�;UH�x%�k����щ�>p��P����#�=ZX����u�]���H��Y���La���+x��Ÿء����Z�D�����e��u��p�Q��B`(��>W�~�*0,� ������߃}f�d�3��3����̱�����bPĠ���jth�S
�eA���B�������m��L��7C��`��}`"���Ǫ�Ue����(P6� ��f�@���Y��*m����}ǍȦ6x[r��(�R���� P�A����X'&P�+b��kY`O���u�z�������W�Zp�Œ��FjD�����[�w�}is��ɶ��:ZM��>u���e��E`�پڀ4 ��2W����^2�kZ.�����5%\j1�RI�|مB9!�/��̅��5-�饨����Z҄���,h/�SBt���
�ϋe���q9�-ۏL;�j,5ߛ��Zt���m�\�B?��R_.�/��&�-'����}��˼KA�s���\CIm@}�������N!ppsA8������l~���>�793;�s؄|Y��/9t��`������|<Ϡ�����vJw~��-_��e�Å���V��yi �z ��9+��q��"W�#�N':����s������۷o��A,0#[{gv-��he���֑�$W���#6�+�n���& �����RR�G�T�Ca�!�j� �|O��0��|E*(p��Q�'gT�FjZ)�y��z��^�D���j9�j�W�g��ϵLw��R{"�21�����>K�ԅ�63> s8W1�=<<4�pCǧY\��Y�3rv��ܰ��)�?*�!Z�f@6W��U_��+ˎ�8�ُV��>+83R&I�&5;h6�R}�L���2C�U#+ eb.fU��8b���^X��8w����r"��������ny�o����B4���YD%׳��J�n�x,��4t�l�S�2������k��}=�{����o�!K�We�YS�zA�0�7�Z�mv��b�['qē��V%0�%BX!�kS!> _$�!�f��=��a!�z�$k5�SͥLv�eo�)h-I"$0T�j��M b���s� Bl	�6�&�31g��B���g��~]�K�G���8��S��Z<2�%đ�|}?_�	�x����k{"w���������zj��޿}�9hc�e�)d����	�6���w�ݘ�O��M����jMjM�_`a=�+bY�v%u5��<w
��Z �4�p�f��7y���M�ۧ���UV���2n�Y��ea\�qܱ���2���>����_�����1L���k����~E#��������/{�h���cНy>�/ª��z�_�l�4W�>��)����}R��C� z��j��R�B,' F�V����V�+�D���Ha��W+ؒ�N����y�K[�Q�f�W��qAR;��q̤p6B{s�R	`�)��g+I4�&	^
;��d�Y`��.e���o�$(��ip&���^ؘ�%j�%�(zL�6+f*�p�`�pӭ��u��G]�"UІ��+�5���( 1��Y�&x�����>�h�����{z~�'z��F�|���@��n�nnha;�,��z�G��q�Lk�_������/L��G�	�W0$C�%/�;	�K�����A���/���MC5}��A���,aQ5F���3L�8%�����~��l����&ᇱ{��&��Q�#�OIV]�2�����"v�b*iZ+伏���2�|*��ZT?m��k����jgI��c���>N�s_�|���\Wl*k�]�'
��p�f����]�y��t`(��9�ղo�"����t�9J���%�bQ�s!�.o�h+X��c/W�Ӧ����j�Mǭ`UM�&�;ZN����M�_�޵�*˞֧���iX���Yy�z���f�GPq���_�xrB�2�wn7ym��n>�=T�(z�f�Vw�ظRӲ(�S�����6�����y�X��b[A~^U�\Wu��h��E��ġ�E�d�� K�֗�k����$U�W�[���`�|�\�P"�be����}�q)-U�%�0PA���1���J���)�L�c�˖�EWL�5xd�x v-& M�����J�؄j�H����<���}O?���K`l	{ܵN�����gd�d�gvs�X0�^�rt�;�^��b�H�]��_���赍�pf���w�8 ���W�~�ml�L�v���F�8,���AFZ7޽�QK|�8�w̾8�P9��P|�lǱ����E���a���!��v�^[9R���5�X�.=���6�!�?�U�rx��<�^��KϽo$J�N�z��Z�/k�ℾ�\�L;hzBm���{	<ޓ�^�/��(�?���=@o��3��Jn����k��ח(n�s_�\���s�0��{�Y�$����V�~%9_���@s��禼�Lo_����>Ot{w�3S�O��=	�x��\�X��7K�X�5��=!5�-��S ��nM�'��*%T{1M��=��o;��V7�"z�(�����qJQ��+�)��^)K�W�-����i(u���8w�P#�׆`�z�rF"�s`� �����'W-� F�T����W
��-��l�_����v~����C�|U+W��=�K�Hkkоy�vG!�%a�n\�-ڮ���Rn�.��1/-�7�)�wlݒ��F�v<����ؗ5>g��*?W��TJ@o_��~����.Aז_}��%���%��~!���	� �[-�)�@�Z������y����@�j�u3=}]��%��K��W0��[	�u]�������ߏ��~N��GY��L�DM��W����������7�h�wmʺ�p�.���_S}���d��ǵ��K&}�7�"h��6�bM?)	��p�� �r���ʌ�
�.��ݡi��t+A��|��3��u��AAs��������}�ru�����'����O��K����Q��-���U��`P��Fe�����}{sh��8h����F�@���,:����֫[~���{I�����y��^��CH�q��������?���.��c5�\m�8;c���aO#�[�&Ƙ���?1��e�Ŀ�U����"�0~�C�9�ʪ���g�J���`�J@��X,� �T|n6KD�`jjw�p��b��� O�#A_�3����Bp{��Ԯ�66�Ĭ��Q�SN��p��[��K�-2��]�X^���{�mü}�������v�-q��}�g���CC}�יP���-�J��OS��n���>ŷ^z},���+34h�ؿ:�`0,;��C�����#.�����g�.i#���QO�#���y�1� �����N�����@"��Z2�ݮbP�I��傍R��ڽ�ϫ�s[�ܤk�8�՘h�et��%�_�'C�w�?�(,϶z��R�f�k�o��\����-��Ƹ.�/��V�m?�?sk��\���f�?K����4�l�����\��˧�un��~��#���_������{ė�3�ŏNG�Vܷ��v  n�6Q|��"�4�ohjreyb�}#]gۼ(Q�%����ާ1%OԖǢ���/�b�o;�C)��y��H� ��Οeܬ�:��vY|WS3xxG�˳�����eY�mz^�X���3���]S:�d��C�އMI�N#��Q��1���!��,�OW��UQ͞�j�ԊQ��JF?A�=�����S�%�i�p%)`%0נ�|p(
]�|͐%�uz|ʟ�$P��atDD*�`�����Qݽ�N��|t� o�q�̡�[�L�OX���;�f�\�%~�ӯ
��
��Lk������_C�j�	<��ԇ��Â91ꞿ��^��yu�7�]t>�d}�x�X��t��:�� �Wh u��hwF^��x������_��9X6���1ve�Jj�� ��VHܛ��,� �(�=��%���J(�Cv�\s�m�o3��f��^&��K����` ��,��F�8�"�p_���,���F��C�\nram?�� �/y}��l㓽5�M~��*yz�w���E���~���]B�8-K,?C_���yY���<�K)�4J�|�ܠm;Q�*�q�Һ.�:%�����NJ�En���R��&W�R����|կ��-f�{>���^���� ��r�>k6eCIu�8��-�Vg�����A��Tkf�5�S(��N���ĢF�r"�x/��9��Pm�� �*�W�n ��k��I�a�pWh5>����y�#��^��KQ�VA�u#V\�\��č�.8��
����|��8��͵�w����#=��m��'��q_�TR�0f	��*1�,buV_�^З��3�j -o��OzeM�X�Y���b�h��{��t�zIU����Lـ��`���[;�����7�s����<̒6��)����U제)L�9�}g�[!Jճ�J\ܱ)wW^J+kB����2�kb��֢uq�ƺ�r��gp���c"����tm\�����������KJM�k=-���j
ە�?��&�b�\��r�Q�M��S���;��l��Bc/z>?�r�oJ��Kb/�]�����zl��V�D�s �s�!���������?=��d6�ǵ��9�{9�y�'?9�2+�������
�D�֞N��
��Z��Sw�;o�	�Y�}'��`����v�/����������K�w�R�F;�o��5(S��D�"b�:��k��9��{R?�k
�`ŁJ,��p�sU����+R�s�ʥҵe7��iC�B��m}�_QH.�U[����oy�8|z�S.������[:��p��k��tj��A?�x^�N�0/�z!Ⳓ����/DM.x](�s�ߟ����L0#�y�<����ʓ����/õ��kq��Zj�� �Xॎ�t��a0Ь�+xo*v��Z�����X�l���'�L�uT���� �>�5��k.�ܿ�o>�J�}�����&��<�����?%k\<t	�n��o����l�k�q_�#��u2������ �4��z��]��-_�-^
rj]�������X���N�
 �O�����E	����X8�X>��$�i�[�X���癤�@Z����h_��U����R��)�絽�N$Ao�Q�S��EY�y���K��U=�[�Kfp�� ����JO
�[���d�J���{zMC{�	6�
�N��nU�5�>xx%(��0Ĥm�Z%��[��Ֆ�;"�����q����~[���bȥx_��be+�3�J�]����^e�}����X͂g�2�����؊�z�����%�p3�M��x��ؿ����
(n]��l����$��ݫ7z$��y>��a���;)����,���Y3�]��\���e>�\�6�[�v������_W�?n	�eJ���e�e�]�e����6��<X8�ī|��=k�T���c��H�G��sR��$2�#��?����Fз����B	@��ك��w��4��9̅�#%����4���{^"^�-�e:���+��e\׶�3N��E�o=9A���X��-z�?�|O��dLE�U�펮z�T�wsu�6
��$�(������v)A�5���V�����+yI|_���?^_d��u�����0D�S��ĥjZ5��p�{	�g>�Y����9�����hh����0 cY"�|fY�J����D�ޑx���^k��,z����~*%�i����i �� p���,�."�5�J��Wο�*{�a���a�#���e����l+��EӔ�f�bz��yւ�l&6�>s���I��:!��씙d�2�;6E��X<�e�!��Lx����N��;���f�"ȏ-�w*8d���q�� ���^ }�ۙ�z:I�>p��gv�����vp���x&�[)>����)���ܣ�I��6g��LN��k���르��@X�C��Ŵ$�S��!5j��r�*�Gzs�������#2⼲��4�mDed�O�){Qo�~��hX����Y�E�������?��/���<�4�<��Y�g�o+��W��~�8��-:g� !��1�'�U#����"(<�r�7��y�?*_���;�iXJ����=-޲��Ε1w�e��NdI\�V�/�'�x�Tp;Rz�:��tr�'����w��Tzr�w%]GPH;�J�H4d�X\6��X� ׈���ZEb���nv`Rl}h�dU%�,���.�*os�æu}u�D�<�^�đf���0!�D�\�9��"�5�c�w���a��"�-_�R�-l@�ԿJ�\�$�e>����#�g��j�r��>�@)C�\]h���8/g�b������Y�h�K)����tHV�.�P� !C�_���u�W�� ���Q���H<��eweٹ���ל������5>3�zl�vW�ewc�8�q�.ғ�k[��7��Ͷ`��&)�iI�u��&�Ų���ne =$��K��P�K`����������^ʊ��NoM��n�gF��%�7�#J�d�d-qhe>��Y��432��j�B��6N�%�*ИE�w-u4�3��|�gf[%!^��l~�LE�
���6{Y�Q��[P6Df�mt�6]��߽.L3��W^�n�������u�0W���vS�g�^r`�6��rxi]*zq#v�nί�Ӽk|��e��%@�7(�CY@���W�b?̫���=N�h����	@x��<���������P�rt�L�*�a��O�)O��u�k�U���ԛe�������]ނ�ݬ��`Fݜ�L��]p�w�˼9�b�f�+�ST7���x�\\�]vt,1u���K�w�2�XqU���J���`Rb�<�A5
�dU9�f�긫��u�bV2��O)����uE�V�����xL�`^%_TS�W1��� ��&�aU6X\D��.rd��eB"���7����|[���K5��0.�Vɋ�qAY�ś�z�c_3�ħ���VMw^�	��7���}Rا�r�%h�5}�����ʵ�>��d�{;������������	f�꺢\���4���h�E�
ȃlj �uE�J�Ӑ����N�Yd�<o�,�|.G���$0OĚwn�����λ�ֽv�+�7����_�P�^��ڗ�(�>��S� 5�X	�R�~���� �-i,X}L��b�V�S�g�c�{)Ծ_��Ӫ���azP���>����-¿z����n� ���g��3��;�����MG>�~�u���b<۵�x��W�����#78����ҷ�'X�٪�`l�rG.+��/v�5�}1PS���k��
�8z�J%���Il����9ї��nǋ���g�85 2����C޾yC��߇��T�?x+��z�q�'P*�U0�������+�� ]���1�H�"�J��>�z��>a#W�>�;Ɂܒf�A�k���c�����u����&�I���[
�J��,�l�b�H�'�� =�� ��ی�V���n�9�Mn��K��C���E%�Ǡ�v�8��Śg=����*����ȱ6૕�W���� ,-.����6>�l���� �(�4�
����3����`}���;�`����вE�}�d,�@_c|},RH쳠�h�M(7�ͼ��C�k���V���3�aI�5���b�9�N�	�N�&`�� �x�>|�����|��8����=��#�P��4(4��"h�\�;M�F����q���u�ᘅ�� @�{�ߑ�l)���V�&�u#/�%����3�2�`[�$�'	@��O=jq�����G���Z1�����K��-����W��&E���ī\#0��k�o+<+��5VaݪJ�~�c%�����%B ���*��s0,Ʋ�$Q!'����n�>���M��X��m&E�((��?����jW7���e�Z�����>�D���j�5��ě��F�Ƞ�$S�9��]��y���e4O�wc~:as8Z�������U]'���!�l��'�k�A�q���`%��-jzXeGØ�(����I�E �1	��(�k=��>�[1��y�7#|Ϭ�+��(��J�L ���c+$�Ky1ԯ%.��ME^�db>/bp2�L�<�hdX���u��ܷ�I�e[f\��?�>��Z$ N�����Q�d��׬� W1;!{@(��B�L�]՘&�a���4yXp������z���L1���N�������Y�&��Gנ
վ	��[}��W�ml�c7k�׵��y9b�����d=u�	��!m_Iqu�ȯ��=t.Ú���ދ��q�o��V{v�;��>���n�&�őٌ��i��^w7'%wUwW�[CjZ[�7`�8��XX���?�u�>�������c�  }��n~�ԒF\�ꎃ���խ�zòVs�r?��M	��c
�L���8��}i�/?.�w�|}{�c����
g�(4H��]2Z2F~㊰���G�������]O�\`-�ZCue�0����e�\�p�]��� �sH܊Tv_h�P����ǜ�I��eWu�J	�2�Q,f��u���	���a�b=î`��uY)V���	��̭. ����X�oٽȉ�\��4��k�}<�ih��s����5l,&���$*	0��x��h�둡{WI)�~�JQ��aL�`yL��nۘ�+���ϊ��=o�����j�:0�vu�MX��_h�iޮ��c~Ք�zbJ�O��0D�jw��ށ�&�$ϧg��J�����S4����gi
�@���`�l����Gaq�
=��v��F�7�+���,�/�L�O�U$@��	��7�U�y�5ڌ�v� �!��4���t1�-��*�'��G�q�JV=���[��(�6�lۏj�Q�(�S���B��R���5��5�wK�����.�u����»Q6��RR�3Qn�^/y��m�L��8�Hy����u����K<*[���e�#�vp$."-��_��	@&�)���Ҷ���q�S����l�BI�zd�,�*��^ě�g�5h��?:��3Zc��Dx{��t�w�>�e�lc�z�d�k�`L�@L��"3��LV��J�c ��)�bd�h���;�Y{v�ǭ0Q�D��S��YN��o ,�ŰHd��]�:w-=/��~�� �D�[k4%�@�jqq�E�"�C�d�q�5\q�F�����>�ARX*��F\ӿ��m�����X�˗�`B�C�G�Q' ���h�׮�kӤo`Gj%]����R�$�OF�+�A(�1ڥq����p�Q},�_��np�j�CC���g�\��(Z[����Z�p�&�n]�e�����y��	0��wF_/��B@��py<y��)t��ޭ�m]��p���f!@2���,����o�ߩC���[%ָS�j�߃B���P���l����sn�߅@��r �ǳ�ǚ�_�̒�ݟ'"�k�
�us�VY�2�Z����{��^����]�<)�c�����&��;܍"'W5ZH��<tJP]C �Q��`��/�]���W��l����=X�V�qf��j�C
xv�f�D�\}9�$��m��/cx1��ӱv��B��#x��O��H^�b	�)���y��4�Y���ž`f�|��m�]/3��+^	P��q�������@�$s�|����g������|�$�]@�	�T�����+����BHD���!����D���&�$kT�(]L�@Z����8k�ۯ�� �?�j�k5K%�� b>Q�-Y��Z�� �`��XQ)�����0bZ|�:f^�q\�B��U�.����Ԧ|d�p}fJ6w �y=�� h/� �*�ݳA���3�(e�g��6��I����Z������B�gf�s#H�l��%�Ṳ��MtkOz8�~��胝JQ�X��	̱-l��㲸9=�du4��s3���X�w���:w�؅n�&� =P��*P��*+@ŭ�h�$��t_��dG�l��ْ�y4��2Y0Fs� A"��/[�zp��3X�������L�q�J��FQ�#�WL]Jj̉�B	���Sk�@��+i/�V�i~��������N��b֜�w�û�����c��Xn-��������|��@���Km�^kt�V_������bVS��$^$V�mDF��Ru���w {��n��ށ�vLn��>���L��������6�F���2kF��������A��k>��Ƙbv���"���D!S�M�h8�w=�Ed��d'
���rRZ7u,�Ү�QD@t�N�B2	,Pfc��8*���ta�����)�Y�AJ�K���[�A��y�18 ��05�lS�`���`��f�X�X:�#�ُ������+g��(�Q�E"|۰�
|1J�x��;����3Z|��g�t2�CXEjz�K��h��O�������(a:�R��V���W��Ҩ���d�ڶ�}m�xx���3�g��(P��c���kW.Yz���i�E�}�e�&���v8,{���5�V;Ķ&��C:���C�7��q7+>����T��x�n���2+K+�T6�;��Y���o ��ұ'c��z��{�bD��L��m��n��kjp�yͭe�����&�Q�������R'UJ�h{H*��{�C<k��x1�E�����d�����6�eqb|i禱�X������vɨ� ���/��ͫ�%��M=o!�#u<p�+�Dj��=x�O��L2ӕ�AE���{���|��$Ƞ��)u*��S��TC�S��;=)�� U�V�.�
bj��e�63ˢ�O/"�t�x҉���*�Ɨ�����<�c'1�8;[y��sd�G�z.M�d�~��:=�܎��ō�x�LM��&^��S���
�N�c;�z>�cw����q�G����B�S�	��58?�-��*�L�e���!����RO�7�h-c5H��U�5tmH�FYB�V6x���S^kȀ��x��w���sV2�ʦ�����eT�fb���b�?J�NI@0@��M!.�5��o�YW���`8�Y�:��_�2�w��2$�Y�\�:N������A�,dَ���L���hf��|>7z<�;@6�Ӌ��@�BJ�rk5�Z�,-su0�����y&�![��gh��/:+S�f��h<+gCb��E�b�IAo��O���kg��Z]<v�@��e����Z�����F�~���<ǭ�6aJ���V��H���t�'�/Z�ZBY�?X��؂0_�T��=�E2�PԔKi�%�=,0��+<�Ԣ���f��
�9;�oc�.�	�u�&�i�d4�L�f( nP)���݅���<L�����r5��	?^`�����������1�
�������6�uV�(�)�
�bj�0p!�(,]$y�J�h�����ȁ��^�n��ۢ\<1P�&�Jj�.&�d�p1^V�ż��*��(���Bg�
4�2��E�d?�F.�UӨ����:�f�V���W�=>ԜيY��i�ݸȳK�4���8�a7��ni��@��F�1`�� Evܬ���5��g:>��/���܄���2��ʚ�
�}�-/k�l]�R��q02��bi����3 �C&u�'�k���d&�D�
��,E|�j�3�nu�^�ˁ�DY��+�PK~w�d��(Ő�*�I��h^�f[RVs�ԏ���D��F�~�LB�^|}�Im� ��^.����6�İ��F��aR�k-���'��oP�T���ʾa� V���h�jNpqa��.8,��7�ҫ`bM�N��>fH.�q]b�|�Жm�����nȞ�J�Pk��R��d��P� dZ��j�,��Z�9)�B�Y�_�sE�N1��fuhA��@1�w�W<#ȴ �u2��ݚ6Ok�GV���6�{.�RX��Ǭ�Z�W��,JO��+���
�u�~|\��z�D�H1���9�C�5���˚_�t��}n�b}��A�2}��_J`�_
������߿���������Ӝ�k�X��䕃��g�O�l�x��dIJ�#�fc�pm	�i�J�d�����x~�H��?��a<� ����p� 	5�1��U�f��`����ĸ�,���MV�u���:l/3fY�:^g�����XC�9�.8Y�ײQ�iה6`�L�p��@��H��������\'F�& cD�Y��G)��)Z�ϊz���EP�r:��N�gl7��P9~qQ���dζa%�UƤ F|Ң���t>/z� N�_�9�V L�ډFŋ�O��a�*�,�X������q��w��д�����3i�\�������N�1f�%�h�k���n��[��`�/W������q���b��+���o���z��e���I.��a�2t;6�;6h��'@- `$9��o�g��n7>�����*1�kU�)���Y�lY0����s-�����a���|�qo"�j��Nw��R@���{��o}�=��ab�*�#y,؂�r:�箦��\O�2��*ծ�����b	�=�%�_�aѠ�=b�Ђ5���R3�v��
���N(�G�5�)Sk�4�Z,���T-� 5�\��K dV � �Pw]"=���0�N�y��[�_'�eA��Ќ��vQ@�kWeʇ`e�5qB�K��r���(��"!�l���d	J���-9�W��ߗ�.���_q�6�ت��� ��������d��~�P�� ��a%���K2~I��g8���~F���s)����5 <�x����@�vU.N�@JO埅�n!c����7:�kxB�N��d��}�F[�"�	� �5��+�ȭ�.����֊[��i���,^�j<��0�_�y\�<��v���-20~��.~ֲֳh��|Z���L�����fj� ���vl�6��ޜ
�������Q�[3��Ufޓ��.VPP��j�J��@�f���M W�g��H��n�,�(O1��-a�>Swb6������տw��_#���UɃ�M����d�eM�BP �1!az6�@���Wv��~��+����X��Wo�ɿD���QHz<Q���+�R�٬r��C�L2��ÛyYg������R+��_����
���i=�i
G���ѧQ��� ��4��'�(�E|+D^�V\o=��k9��;T;���
��~��%=A��f`�P�?H�r�B>��ј��{� ���I��5t�Y���N6���&m��VC�/|� /f�����N��W���2_'�;ңА����`:���b�)O\ރ����cw�0��B���@2 �A�̿�G�.���6v�y*b����_�"��A����A�3(]�H���!R����q���^�%�=��P<_�E[m6n�������w��x��p������u��ɜB~�\2tPRVK�0p��?c����5��-f\�� 3עd��zR�B�{�f��������H�U�X�Ϣp�\0-U�AC���=��V����Jq�cj l�_E9�2b����+�yh8j��~��];�0�Y��eVS���#-����Lg��.��r;44��21��b�s�x�y��f9Sj՟��eE�=�agC����b ��KE5�M"�a\G�P`���`�	�A$�bRH֬o" KT�G*����]A�-W[������4��J!B�����v�[ms��l�F�Qkn��^�L�@?����T6֤�x�d���}��� 9bՋ��f2��F	����3���ڦZN�&B�B����sc�*,��!�GZO���f�R�d|���(q�s�ѐ����Η�V��j�ܔ1(V�R; ��23W̖<�}M`�9����Z@vֲPq���s�(�ر�M�,s��
V��YM0���ek���b��	�O�'��e�A(�T1#���b�H��&��E3�xT�Ӿ̬���wE�ƠA�`N��`��l�D����e�d�oq�+H0��L�ٺi�	W*uQ�_&��LaQ-ju�z(�Y�G{_�(��-���Es$����{��01R�&13Y�d����Y^&���Jo\r���)���RE����×/X�q���K��'o�^�u���S;p-�8� �6o����������
�����*\%�`|@�Ivf�*﬋z$�B��uyVwb%ZZt�����a=�&C%C\��j{�<�[F� f��(@fy�ڦ�R���A**h}5�Г�^3M�����1al=��߱|=��uyl�x������Ӹ�n:�=����qb��Z�7S���޴FM����6A'E�ӡ��� �<+�۵gcz~!�ÌP��V��b۹����_��X��w�C��C%.����u'�(ﺓ�P�{��t��u�l�����es��l� @��� Vk��Ʊ��"�K�nDg��`�d-�ڭ������Ϲ~�����-��Đ6����@�\K�l��s<@���0��A���$.򁵮y"P�X\��Fbn�����6��j}i�K��~��n��坌��E�� Dn��)��]WX�֎���A�
�0n�:src�(aj'd��[c%�s�=b����1��2C_mq4�l!�\r��,�Gd��UV-�A��'j|��BB�cY���`��1�����X�-VKI-`�Nv �g8�� ��NQ���Ͻ;ʁ�F :��'��JU0�"�6�w�Ϛ�W �S����ɺZɳf%^�  �Z��H�p�r ˥(�p�˼/Җ��II����9��v~�t�?��8��/���,4э�ȹͥp�h6���#k�x�H�����60D�^��3S�=���)�Z7cٽ�#�[Lq[5�\�8�=�j�����`|�����"n�"a�x��Xę���!�Ԛ�dp��yb�5����=�� �0��ˠ+�"��a�����2���>�9�ȋEp�rj;��p�|�1csCg��K`��#ڻN��T�ٷ}qKbN���Z����O��$�.����K�NTgƖ�3�0yWRO�ƪX����ZR����%��J���`F<ie߳%T�g!����ҀX�:f��QTs峚�� abc
V#'���@�6��f���	�(��c_%}�N�|�F|!M&a�`��-�ZM�� ���z
�]���	��Vo���T�otK0�����`�LP�������)Pt,��%�X�Ǚ��Q3Y���e��'�L�l�il��P�*��eG7�M�9�q_#�:5Z?��Ƣ1��
��}kH���-���F3TQy�hy4�6��{��D��aR��e�b2G�)�TW�;S �EB/�c�D��A2�Tj�� ���%�5zQ�l���<�� ��E��&[�,�c���Z����*8Pqac�^lYs�cd���� U�UkK�]�  �#��v�	�����
/�X=�,�q�y^�p�b��h�RF�Fͫ3��5���x��p��%��ǳi�������-צd�VŤ�[]�խ쨽����^_`���|u|�%����Bj��d�Ö�J���$�8%{��X���,Q�_����S�(2ps&n�&E�_��q�ת�}�Z�r\���1u?���I�Y�O��G���]ex}xu*�N�|g�qT,<�7�����3&%p��y����d�S��$�ݎ�Bj�Ж��q�nV	ݚ(�Ir@�X�
�3��a��L1@�(�Pxn���<��b��1zB�
��b,%�X)�Z%t g��KhODZ��)���C�=#FD�093�p��D�P[��k�̉��0�����R������8(_�$$	��V�u��<#��Y�iC��%��p	�Ee!�ˎ����&�pپ�qa�F�/���}�}��/v�*C����3_1��oh;�, �
��e�@K�D�����167��#A�L�m�Q�V�QP/�V�ǌE��9
r`�ea�{ך�7��g+3�v�^2�s���6�ݎ���^��x�[躎[���wK�8�f���A��(���)�_R��e�m��g:>���{ZOg:���	4[���,�[f��F�� ��4gAX�$�繘�/�
�ցyW�j����%؛�%Y�(H����;�©f˼�4/jA����W���g�1����W1���D��n_XgY7��(����t�c�M�(zB��/�u��i�c�����l�j��!%(�W���U�-�<�P�X��&>I��	��Pj!V`� ;ًMiQK�3�ͯ�+9a��^�;2 U����I`�c�hhH��������AW��h<�I.;��RӮ"���;�L_%��g�e�>tPS�x؀#A���F����sSvN�Tq9�&�z\h���Mc·��)���K�>܍8$/�� �����(��ZLQ�͗��*o0���"�s�I���-bԒ |���Z|�3{>��vl�k0@%�W}]*=3]��-�'ط�����1e��j!H�X8>e.Z����l�ҭS��0�D��[�XPp �2��Z��y�&�q^&	�[�s���f�1���
�R�]�|�#!P?��[K�.i���5,�->FB*��������� ���-2��A��
H��T�k��:�Y/.���f���pm�����{���� ���V;`��
����d�P5 ���jZ��@��rr�hU\��0Ыۻ��� �g ��*�7'������(��h�Z��[������
��5z����o�Л￣�~���z�ȵ]��4јXA��4W��s�\�)yV� �b1;����<O�x�������9=���Dm���2d��3��*K���4i��p��>���_J� T�UM��KPL���%�!W��w��Դ���@77���������g�=�;V��莁�����Lϣ����y@�X_���;icr�]�o�O��'��5�ƨȑ��]��- wfY#�j�/>�geM�qG]SEa]S|͒�r�/�&K��p���ᆦ�^�.{><>j��tc��Pnod~��,����"�Oa�8aV�Kً�\���,��e�q�Vx�ܥuL���~�V�%��g��#`��J���j����+�s�e�,LrʿQ,�F[J���1a���>�b�a"�q{W˾���W���H��d�?K�,q�����LU2�-�>[N���v��CSJ_?ܴ�-�j���W������E[��<X��d�1�^'�iM�R�#���ʘ*S�*�;}&��ga���v=c��>лw藦��B{�j\]��$�25M� ���Β�x��ݹ�衟+\�n(B��}�x���^�B�p5�c���8���������'a�$U�d�3�uVM�4s)�c��$.S]e:�ݷvۻ�.��,�]
�U0׌"�*�uٌ}D�%r�-���z�'��gx�{���#���E�кn�٠���dE� �˯,���K_�5��	Kbu��G�$�L��(lG�Z�H|�?�1�(Q�n�6�~W���Fz}7�ׯ�0?���P]}b�M8�Ͷ��"p�Q}n��iw����W:~x��A��6�������;�Տ�ҏ��+z���4m��Ƃ�+�v����+u�45]���n,�����U���������ۣ�����L�ѫ6?��*���Z	n��i��؟���}1K�
�A�KYvAP]�X��3d��_TC6� ��}����w��1 ����΄�e��3�����i0����\ +')�(�c�o#GE���&�26[	��39ii��?C����H�ײ�Ei��$��kS��(��o0���I�����J.ӴĢpӡ���X�ZߧQ�6��M�z#�X�*B綁ֱH��c����0�X4)Q����Y�q�E�ZsKtV�%���G��=L�Nj����US�IkK
H�9 gZe��G��}P����S�(�
&w��zqC|�D�>$#������?�M�&�<@��]��]v7���]tÁ����eB:�&q�-R/Qd2[89�I�@�Fs��X&�����fl|w/����������^�~�7�_��+`\$X��E�"UE�E��23)�k �[Xm#�i׸8���10xc����x^�Gn��.Qq<���_~���?�"�.0<!cet���EL��Ot��Դ�3kN��Cƕ1Ю��h������ L�"�����`�^�Z�RI<�rY�sx�O����9���MK��tlL�6Fyl��H�ޑϱ\���M�56�@le�n�6�����*��$x�]�R��dA�����t���V ��U�t��]�<��pM?���!\c����Vl��@��;�ՙ�.�m����U��c���.Aݵ��b�>qg R�0�v ��ń ��R��0��U��[b�V
K�?�rFѾ�}� ��7���X�D;��7�f��xCmS���3PM��i<2 k��Lݝl4\���#:4����[�����o��wo�� ���H���)wg�5ˌ3���<kVu .�gҼ��cc.�hw:ҟ���h��Л��L;�BX�L	 0�h'Z�5[��{A�+�:�^�bѸ�aAe�hW���{����#��w�{�+>sl^�Wd<n����C[��j�I������2��d�9ù}N���75� ��`Y�!]�Z��ĳ�-ɮ���KB<�yM�L7�FOlAۻ4fK*0��+�8�V�I-� a<~�~1�yz~�?��L���?��۳��jJ�������I���U?���U�*�D%���â��y���N�*Xb5,Q�;-^��1�
\�ŧ��K�DE0l�xh�����U��쫃trX��l]L��2Q�,���-_�1�}kih��t�Ś�hQ��4 ω|�q��6���h��V�]���nO����������@�|��nnv�f���Ų�qW�-�8�˦X�8�K�|��φRC6�P������,��IE|�}�+��L��O�����'��z��̧��e7O�"�R�P��ό�Xü�߶A۴�������h��E˷v��RB =i�0���y_ܨZ� � ,�h���>3rm`Rd��������L��}{3{n����~��=����}~j@�Y��ź�ֽt� ��b�&�����oFS�H}W��u�@뽭�v?�U��sz|�C����c���O��7�YPP�T�w�	�ǹ�iW��zqm�1���>W뼸����/�&G f ���4�$�ْ�����^ҡ�ZvM�rL�|�(Ǯh�^���	���@��^�t�/th�(;��%1����%��XY�
��ܾ�y��	���X�x�Ӡbln�Yз~߷}ߞu߄����B���Z��<l&����ne^p̗1]XI��?�&���l�os�^����ٞc;kЧ�o����v*�$)Pd�g5�.��2�,QL��k]��60%��"��m�i�䳝)xQH4	l#8�g�'�����&��l�,.0m�V�
��a@��<<X����V���1i�����)"V.ag�L��ed���mt߄��-�7��r�k�
�f�=:�Q���k?p�[m�WM�}�ھ!��͢`#�+YT��ճ��j#����<�ob�;�<�� �&z>�}q6k\U7��k*P�f��V�HI5h�׳d�Js}X����;vJ�*K�O��Jr̀e�R/y���U����{�>�̀"�5��|.r����s0Zk7��i^6-����n�bk2��W��pnXcl<�-^��W�~��w���~���@��$Z%��,v1�[��_�8s��T|Js��2kQ�Z5֝��l�ƵR^�)[rۛ����^��ׯ������t`����'���g/�u���y�5��G����i�~�jY��kZd�̒,a1�i�����H'_<&i��G�)��������� ���F�_�6�y�w������7���W������D�O��p���Y�v� ���G�j2��mT�����*?,F�{�,���!��B�(�E`&I؆��C\����@q!\��,=� mĢm��mR�3�
]�����AX�??�P(��L83�cZ4����t��$�Ί���6c�6u{�Iƍ0�ev+/�^M�|ߨ ld���hLcW�R�X ��ݿ�k��(q8��`�Uvfay`��8���N�{:�~i�=� �S{��vj{�>�hy~ߔ��x4�8��iE}1��0h���	�� �{���ǬU~V�����W�΀CbOt��i{���mB1PX~)�a��4���6%/����������HM�$�����暄+!��j� �e5��[訆E��F�Ob� `��9*�Ws�yȀ	�2�Y���ǂ�"���m�^o�&��*b}�b�G�6p}ǹҮ��}6|z�����T�B1��}`d�����T[�ʊ�L��?6�}���o߾j��״�yh��u��Ю1��\=�����R:`��Ȱ����C�{��_}-.Χ�I��˸���=�����h��]b J+6m��{�sA}b660���s�[l^�gyo��F�>�5��
�q��b�u��>��-�On�R�w(�4#��{-w>ër�i%S����c͟Z����
����$`�-\�V}j����#������������o������>�]�Un�|>6�9[��fi�V,C�������������H����L��������Hi��\c���c^^�gQj����o鷿}�p�.SN�e��|V��� ���nOw��y��~�ޯ��<q1��
'jdM��"B�Z��ꓑ�)�ֲB+ң�f	�Sa�2��c m�M�15��j�N�{�k���^:L�|��5}���^���?70�����~nL��4K�ؙ����a���šb��=�5�Pi��h5pt��66J�^@ܝ���|�[V��]Qv�l �C�_f�*�q��� �5��z1p��vF\�������
�?b�ε�߉�TԞD�����{������o��o~����������u=�}�h�ih�noؼ�k{��f��yg�� ����JZ����}3����a!a��ց=�N�>6�[��?��	0��˶%;V|�d��K�E��^������u��ˈ�����9�)�b|撯Y�2�^P	)Z%�$����9!Hǀ��Ԡ�����X �P��p��Mzig���r���}O��7:X+>N����X#�"欷�&��dF���Y���-݁�F~xvq3/+(���e��D�@�}Y]��	N�IٹJX𬃶�3i��\�t�>��][����4e�ݍS����Ċ���zAMV|w�R�Z#�����=}����Ʌ}`�%��f�j��88���Y�JU'�%�@�������o����M�>>=K��qwC�������O�=2ʾPa��;RױVPh��sI[Nӻ���������P���z�omI(���������܃EXS�,m�"A��g������J\���!e��� V|_��%X,ق�n�=�^�|��)�3�7���o_��������@���;���+Q�'�����J�;���݈��PxL�vwp��/�d���`�s���U
y�[,��N�p,��ϯ���5agj�����_� ����Ml���4K��I�m�ى�j���_}Oo�~'Y<s�ܟ�8X�lY�RYKS�u����Z��W�]�F���bO�%_ǶT�kRL���G���� ����m�ҧi:HL /wb��tӘ̏���ino�w�#�����4�������Ǧa�.G�;���Mf*�UT��#gA��³C���kaFO�B8ƥ80pSqN�>�j��L
~Z�Tl0/�9�F)�,D�,�t.Dy�:8N�g�=.7y_�_���3�`"[�Xu��m�����!������3n���Y�H�����w��~�W�����~��[��ى�x|z�_~�Y2�>�'���^K������� ea����������I��`�}6A�I���H����ه��,�g�"�`i�\�n%	hߙk_�
0�5 �Z�ؐmYe?ﱶ1�	0o4<����>��[|=46��bݷ�rP;�Kn�۰��8�\��gxG;#�(���4k�m�$��%�|V+ݠ�VʑH�U�f����̆�t��,VW���T`_-���,�1g��ߍV�jF��b�!������u�V��)�r_��s��%���8*ΫӍ���&�w���S)�a���9�) �v���Z����{qW�6��ʁ,(�[��{�[�X��㞚����+z��[�{x���F�����	P�uh���d���T)?��|��bsV	�o
�}�ww���+���q1yˑ3�I���le���%�#���s2����$&X����g��� =�.�s���%�7��%��_�!�oL��y<	䈻`���Y�F�'"s�jR��KZw�HS�9��-�����K@�-�؉��$��n�:?5^���@W�o�>�����o�o������h졁�A<�RF�ĚZ�}㺈��<?s����ȑQ<I���{��'9���L?�~�,蒑ɠk���W�~�b/qd��!����F!��5(鞝W��9NZ�����J�ӱ];ѫWoiw��ߧ��C�L3ݴ����5��{����]�Y)���͛uP�*�+��|H�F�<�a� hZ�� 
2�F@+�A�����-�� �'X�f�j����0�E糘�HOgv��>���-}�6�ۇ����^5-�n7�?6�����=��~���^���Y��3�	�h��+��2�QͲ0���(�T�W�����ɰ�T��$sw'j�S��UM���z ,`�a ��1!W��D	`�K���~z�u|��a��||���:ϝ'�:N�#+$������i ��1 �,�;zh 뗛�gSw�B 0.[�V0��SjK��T�Xu�k���o�Q�������|�q]���įܐ���88>1`�6>wW$���9s؁	ڴ!����~�4ga#��k_�ΥJ���2}Q슞�9[�N�a��AI��Z�#��fƯ%D�"hu��I�	G/R��-` Q8��ƿ�0�1@��^M��d�E������ΧM���1	aO�ŉ|��9vM���ؔk��?"�^VPv�gL����.a�fi��d��)m�������8���j�Y����E�~��k��Lx��p����8&X���m>h����ʵ"9 Z\���#y)RQ��c���y��ot��S!x#���џ�5�7���VXQ	J��iT�o�:�d��L���t;n�IM:.��ߋ��ݙ���S(������>(^���/�a�e�%Vhi�2-�k��G�8p�>'h��J���-�Ý���w��I�N�)���b��a�������|C����������w9f���Y܍�Z��ŭnn�#?7,�q��K���Qb't�s�VYN��Y�
b��4 ƀ��k��UA�����>x�ҘF�RX�{���)Z���2���A��I]�|͡��+�C*���������xv�L��Uv�<�݊ 8/o��l�R��	�-�ȫ#]ݑj�<H�P� \-�C�-�l�(�}�	�,G{����t��{�,$0�Q�\Z9uu0�/5C�Xp���q!������Ĵ�������������M�O�F�4�*A�T��`�i�e,�F�4X���n+���I)>����X7[�zUq���܆��Z���gl���F�e�(�����#n@�o�̤�nS�@�x�����9�s��˯�����S�=���ꀪJx��%@S�1Z8�$�kt1�~MwM0_�K7�{ј�~Y�i����?������M�:�~�V\�T+`�1�G�)��Z�U�QqMt0A,qh�w�݉p��L�kI��밝� @�� �.c-b�`j�q�tjc��u&��mѿ�x�i�9(C��dI��0P���U���J�ԝ�y�R�L��\r��Yݱ�k��&�Y˕:R��8�f�8"��&n�6�~��ed.H@(Z�gbFn��a1�=$�"�I��V塺+O8e�p�<�ܩb.pĪ)��4v���Uսw���������z$���,|���Ӯ�X5y��� u�Ɛض��	�Ya��$;���3�u؋�?I;��V�Ac��Y�A9i�$o�S�ҟ��ykS�����Td�non�Bc�sD��;Vo�!T�V`W����\�F�((��?>﵍��8�/���?���:+]�~&�?��ٞQ��B�jlp���'t�x<d�0�D~���=Ux.�	i0�~�X�j�2 9ͬ���x�����c���2��vx?�Gz����/?�����������"�x���j�Gm�ƞ:���؀���p{�7�w?�7�~#�-��3�3<>~h �$%�xW1�a���mB�z�n�Dٝl^�"6����n랺ق���G����,XCx��{�C>
8<g9~q���#�w�}�����od�0�T��z�J֎�OmϏ��ojg!I�����@~�A��G����ڱ
D^�o17&�힞O2�q8��֯�Z��2f2l�X��@��80tZť��VN��~׀�dl�����Y������G=������S��:�mbB�"q�*Z}l�l�)�R�L5qVC�Oֺ%���s�C�
�UaA�Վđ�{�_;>�:6�%A����i�����/0�k%^�.iS��K�<��t8�]���̼�"�&�W��3YI鹰ٚk��xn��{-�������͆S�+�V�Q5=��1Bkŀ����� ��P��Jh��������%x�ok��ԭ���k��ߘ5� �iU!��)��Lf�f�"5��[�ʺ�o��̩���	3G�&?�;���Aɦ㘊[-�:��gg�U8��Ĺm�a؛-�
�.JG\g�=#�X��t�ˆ��d�O2�(��	A��[{hS��$��2PC `y�|���i�Wuָ�"b'i�y��e��n�5�[Vk�� 㪧�.i/��#)��������4Fe\\��.��h'�1����Lh�HD���6Yan{�[�V;a�,��8b�B��%� �m�[�=�%����W�R��|�}���e]��o�����uKH�XE3z�Ty���	R0.X�dEW*=�/ʀ����X;{�v|�ԕlǥ��D������]_?�7_�j�^�Ā��
�g�r�a��>�9A�i�����ƫ�衽_�yM7�gJͺ6^V�?|�@��������i<b+���ѭ���@j,V۟�m��AU�OUȴt� �E�j󪧞h`5KX�h���������4޶14�����X��D�@��y��~nH�Y��̼npa��To��!�<i iD@a ��P�P�.�jq_,�v�"�5��U9f������`��Kh��ąc@��.�'�!�⁬2�e����v�:&H	�kc���o����׆�_�q�?�������r�����zR��h������VZlM*�gG��`#��]�*B��r����K�whS��5qY�[�Dl��"RƏ>o�����UlR2��2�������bp�~�R�� ��DkL�5�@/Ԍ��4|+Y�ߨ ���Z(t��Ș����^�j`����4jB�<�E� B��f���bJ�dF����Th�Z�BcMs�,bxA���~rvK������YB�ck�W-�J�������������eP��%.]2��*4k�M��4��V���[�?pR��AU���?Ю�gA����1H\i�͒�%mBX�ۗ���%�z��"�J�~�2�b�TI�0����R�
�$�:f����
�V��1��Zq����YՉe�>j��N2���}b�>/�W�Q������㌬�I��"��P�}�q�Nd��6�X`V��*�Vٹ��ay��f�ۨ%����bEy֘a�[�V~��\�\�`ވ����)��◎�y4�C����	���+~dq8����p%�Y�{��W�����i�|�E��~HXE�#�<�D��r��,��Q��,����]�&����B�:_Sbk�H���;w�B�Y�B�O�9=5���o������_����_ݰ�J�G��b�f-��I���n��|�x�k)_�r~/?o�o���I#�i6��yn�����~�s��O�����Ӈc�K'I���[�wS�\	&׭�����	�QC��p[��(����>��o82����I0��a꯴j�r�և���|ʹ;X��U7�V|�k<�&���
2tr��m-��ã@��5|.��&�Mw���	�܋9_ۖ�h�gw��X{�&I��JP�=X���d�g�8����n������t"+� ��`�TM��Ξ2S��̪ ��23������S�t%9j�\1Y��N�`�	���~'`����}=����׷�����E�+Co�s�5�+��&J k�(Ü,�8ltbq������{��ee_w�������Y+�Dy�*I^V�5pl�0u˱�ڰ��F�xDb���Y�
�|py8jJ��d�?�iCS�ύ{߆~^M%Wϕf��B潂�F� {���h��ee5k��ENasg���Cg�W8�ǜK���*s/�K��];�f!�-a�(uVJ� )����L��P9FY["��M,S��E�W��sBz攔E�(xxx�(tB�)f`G8����i9����e��F�D��z���bX%'R&l=,k�|)��	�=����*�=p<fk�j�L�P7u+�4d	rJ0^��f[�C�	'e��.�-�,�aܚw�"��I�g���<�����m';y�JgQ:
 �v�L����<����+H���NHi��_�T�	Շy +�8�y*ޯN��u�Y4�G�$�f��m�XuB�Ѷ��*ĵY-��V���8}T�d�+�/ş�|�K))��y����*��������f3f�'����O�>��1M�f��G���ɓ�G Xrz��U����檟�u��_�qd��+q��-��5����������+v�WB��$�Lv�52&L	௻�|B�_MO�>-�x�2X��iM6�N!*�g O@��0 �m�#\hU>�-�M��YǞ�N�Mn�ퟎGRmyƬJV��1�)���H�9]>yJWO����H��P��PON�Ň-���<�T� ���R�=[=;./^��n&V%�H���oLy�U�ur'%A�+�3�HA��خy�0P�ܧϟ���W�p?��$�r^L��g��{����rywG�߽�bb!�$��g�(�)�W����?��gW����oZ���"�I,yTG�v[�Шnh����g64,������<	�ZB���V:ii3��X��������d���{���N>�L��/����G"�|a�.����o9T 9UD�ߓIY���C[JTc;���y�6��ypc`FX&y_�֯E��!Kj5��1�*���0l���Ya�A6"���3&�8a��O�5z���F.R���Z�}5�ۛ�9wen�M&$��`����sJ7��0�t�Q�ǖ�e�yf��dM���ľީT3�kSI�h����q���v� 4BS��5�dX���K����w�-�ȓ���$ٜ���9�\����(S��k�c�4�	�;�;��R�V˺HIZ�-k
V*����){�&�x����-�(�,RCؖX�P��0{��'��	�l�K�N<hJ����ȧ)�@da6?e�I�p/���(ʎ���؆ù��[��6b��c�fʜ��Ok���nJ��)�5B��7!��ZW_M�}n7�������;����C�I+�)��~��Z��DA/f�kD'`?�Z��h��y��ݮ��U��T����Oٓ{��Uw�L%��ۻ�p����r@��Q֭���������/����o~��@�r{s-ՙ�x�� &���qGf^����=Ag�����em"�0�N�`�M�N����fEO�۬�i��C[�:Y��;�$��=�zGΖ��bܣ���wZpՓg����3:+�e��-�U�#��E��K#���s���%烕��e��A�~�NO�Cڳ'�˙՚3&l���n�,y�2po!��Io��F���ɳ2I����^5�.|�5�]f!-$ʱ�k[n�{&��;N�ó�&�]Jʙ�]B$gg���o��ǟ���jK�QA��f~&}��˨L"\�����\�6�%dS�j\_u�)Mp6�vnic�XC�jɛ���(�����\�/�<&`Ah�a 1���`ǃ�7����zh=��ڗ�_r�G?i�O�)7�ʗ�V+TC�9^R�p��H.���̈́��~"t'������1o�W}�"j_�˽�"	]
�������c��*��Y� ҵ�r�\�m�Ve~���)B��͂�9�����J��V�dYZҋ����9���6�K�����(A����{�N$4!6��)i�`#���2+/���*@���u;�����n��:?�>z.������4�� Ȇm/͂�U?9 *[y|����{٧�}5��R���Ӥ�U�Ҝ�7�I>��{�����ENKhP�����5�tִ89�P�T����s���Ň��k�M0�i��HSC�F�-�٫��u�PLH-�l���}���9�=�r���\�p��<�~�x1�,Wk+�u萞,O+~F��0�O)��
���o�e$�2�F0#z�_�]V ����}vy����}���?���o�z��pPh����J�����)���5s�"��т=aTH^��:��9C�7|`�M�p$��䄶�%c�5����#� �%&(��)i��P#��5g��@�@1J�..��Y_�W4]���萮 T�(��Fq�N&�+!!��d���=��W'�5��J��o���7��|�D5$�q�t-}�\rrF�|�]A��
j<�2e�I����c\�M[-zX��ޜ�_�We���1�9����L�7}�$9U:���˹_�zF��ʸ��_?ҧ�6�	CUd����۷ʯ�9%���e�|��7_Rw;O�sl��RI7(Թ5��՝j1
�9,Ƚ&ߓ�=�o/�W`��1V�h�ζ����LY�jw ������?&��C�W�x�B>Ur!&m�Z�3��g��d�W��=�W������L4�&�\5����V�jMڦ�OD��MA\��ޱ��k�\���yU��>�ï�^P7<,F���Z��&yY�RL�D�ȇ(��s`iU�d��-N�N/+�(��p���1�J��v���Ȝ���o �\s˧	i�oE��#�-K�sn1U�2��������z��v:�^*?��,���ߡ����a�����=���@6B��
�lx_rt�hm��)��u,�6���˖?����8D#�� |��Q��^.F ]'	7��b&��Jh����^"r%��gbP�8�v�mW:�����2�3�]�L�S��0z�E�A�!t.��V��C�ÍV�xږ�N��¼C3Qm ���5�7<E�o�<_�í��@���W>��{<"���O�8	�F�z�:�D����l�8W�L�X܆׊�M�s�jr��F�e�ע�;��۔{*��=�ϧ������)<�X�[^�{���B<$���X���L`g���]J�rVGC4ի����*�hUԋE5*IR���,%��ĉE�l])�m�`	���P�������|(�8����Ph���O�6��D���&s��{w;)wj�) ��P�e�D;%���u�l�,�@s��R��J���͔��N8^���W��Lk������T��*%�D^��PM���s�[���a�̖��J��NC3]������n�����o��fU.M�Eв���3sy�y�X�>��e���a:s��,��5����Vw�h��p����u���B/]�"���sm ̾g(�(@�m����Ŝ,��l�C b�.�+���D�ߤ��8��m������_���)g�}kB>U��q:7�$���-��x� �f���V
 �1d���Cσ�L:�X�i8�z���?��G��d:X�r	�IU�M����	T��x�3���Bu��t�����`N)'ܫԷЯX�-cTE�[��Qs��KR�{)2 �Z
i��Y�f$�� b�x�ޅ$�Ir�~��{��z�>���=�
�Fג�f-(* �y/t|
��01V��U�,����ɤ�j9f��m��v��s�\-�pE*�4^Z=Wyᘒ�۳5�-�+�RTX��&��Yq���x��{Z�Vj����*��e����]2'X7�ջ�;��ͷf��1�#%,��Q/�B�n�_��Α�E4 Y_��K�@�c����j�A����ES��:'���&(Q_
�N���N��Z�C�^o%t��
C=�9�-�9���X���*�r�+pNƢ�:�s%%���������)}��W��o^�,��*�ܩ������H`G� ���K�����x��r��Kr���-T3�y���0`V�#̰��c�v'�^�S{vxH
�/./�����|%5~�����Ozs�F�l�]�B�DATAGRM�ƪ��Xg�)�x�$3a�T�q"kN޶b����$������.��ۮE�rFZn���z��0 OT�Ұ0U/�VJ�f��9{�֫;X}�+{�Yq~�7_���{���B�XP��{�!�8q/��R���H"}l�"9Eu⫎WE��
�a5Ry��ꤕ�ыYb��ٴ�$�}/$o}�l�A�7u�F �!I"�XK�aTM�(R�TaH�ׅ;�G������"�0:�[��u\�ˊ����w]�Yr�(��1�2��K��	�3�z�ؓ�mH���.���h�:��ydr�(QE�'��k^�(\�x�j=�p2D��^���ɋ�R��i֝ "PRLz�r�g�=�[�˄����*��KZn���
`	���ŋ!�y*���\���Y��r6S�T'T'k�^[���`����d�����:`z,�;f�r�M���Jiǟ[���+J���q͘����:���=�r����k�L���Gs���-���&�a�͸�2xx�6�ȥ�"�W�a�l�U��z�v�]����9-��Ɖ�k��N`�Zp�����r�������W♕��-�\��®M9�z�sb�	W�M�-U]����q��Xye��e����c�� h�?��1��#�%��<�7��>�ƐiV�'�@I�p��'�/���C�J�T"�p�x4�_�h��K/Ͻ�<�Tu��U���c���y��p�1�I�q&Ӹ���(b�"t�1	��~E�	��HG HS�:����]��<�S� \�d3��Zʣ�B�:o��`o*��IA���Xk�Qrۥ��7�(K�^�E�0��M�/�����,9"���ĕ��#�ډ��ߤ���$a�6��^,v�G��;�$��T:ɂ�*X��4�I$�={���*H1���%�}۴�ƖS�+�k�0ej�����ʄu�)�c5[���V{F~Ɣ�Wg�~zyF�)����Z]����]P��b�f�UN�F���ͅ�6ѼV�=��D��xM���T��B/�mU�p��h�_�zY� ՟�`�<�D�qb����B��}���p�����W�7���������V�dyNJ̷�$씸�f�-XZቃGX=>����EB�` �\�g_S���Z+W���2����!�i$�Ǔ��$u�m�"�l��u�9��4�Hed�JZ L�. -��+�Τb�:�̬�Q�ؙ T���A���dF(���� I�P$he��K��@k_�J����};���a4k\�N����h��52�6+9I7I�^��PRbi����@�� 0X̒Կ�<0��e`��@��oH��׶ p� vd�B�J�2X0�ʚ��Jd����P�7���k�\dHـ����8(�����<Ki����H���84<�\�������Ý>�Z�'"�M[�Aź�6�@Z=l������T�c�I���|j0���S8���`>�\��Bul�O٘GS���P���e�|���6��r�u�Gv�T����׹�i堰Z���Q�zL!��i0��n��6Cg3���-�}���`i%���#x��eE�W7����k���8a����ÑHIk[���;)��bx_�"�zɵf���ܖy#Qp
��a�3sZ�%��'�6�g�$���ƴ殃��
n�+�oH�9�N��p��9ia6y0턖�v�"`v��/_��ӗ�.|�@��)I�@xc�dz�h��i "�7��������r�)��W@�m��T��y�k�e�>~ɋe����D@�֠�p/�r�Y uAۚ�S���Z)i^J�����,�O��xvR6ɴ(��=]��� e����8�z���\N[,�F��N�a�rE��&�7y�{hl���16>!Q7�	O��ɶe���&�/������tL<믃�w��f�c+�פfxV�5�c��d��w}��i����\H��u`�ή9E[�%ҋ0z��$��+S~��{x���h�Ae��MO�����4�$)m���0�/Ϯ<l��Z��Ġ��1�yi�? ���T�	����7\�}1xnmV��W�6��8����D_WSx�y�=7PGjǔY�&�@w��S�z&Qi����ϲ#	���"��4�S�'�2��cɳ�36���KU��~ٵ%�h(n��2�Ri�H&��F�!=� �S@4�9�����4�¼�L�k���a]O*��kfB�r�?}Ԛ�D�͎��t/�K��:/���H Ѧ
��6���t�[�u� `�";9=K�}u����]�~��˺�1zlo�++=Ea�F�zH���,��|�{����C��UP� _���O�n���û�k���޽}��T�����s&iErp]CY��FM�h�\/��u�Q�#�=co0��:uR(Ŵ��r��E�o�_��7\--�Z"��x������>�5���(��Va�	R��V��$���$��
�B� ���F�ͽ�hsqȄg��tr~Q��1�U�H|���//�����gL�����2��YlU&n� �m{�V�sf�Ε��8qm!1�r��O
���q���*��'�@_E��9��;�qn˰�V[��+���"�1`Ir���Ѽ��W/���G����x9��3;R2�D5�-�d?���ٯ�>�sW��b��`Q�LY�bY~zO��D{��\P~��7�����i���P�B�m�jIƶAU����VW��ٿ?���cuU��=:|�{x�F�q�w�LÉ����L�;d&s��yR|@�Ʈ~���6l.�֋'R
2�x��4�<�{�a}1��U)³���;m�ß�.9 �l��!E0�\�(���mEXN��Dj+#-��N�<��}���,��E��T��6's��-Pt���5�	˒9��@q�|y��S��b�m�o˾(2� �+O���W� x���8��uhC�`�Z��r�D*"s�C+�I=7AG���vE�j�^N����+�wX�k�2p2��J�!�d�����F�0+�5>�$�I��㼼/�G�3/  � �(�5���ҐS��c5�yM�ٽf��V�����O�� ��0>$�#g��� �u��Su�T� (e1ٛjHx�A���*)�^k��:?.�>�F�{v��>8�ٚ	���H� ��1w& �b1��r�MO��/i��eE��~}By��������iD��'�O�y��^l�U���\R �`x�={rV��s&��\qػ�5��e\ AH�@>�p^��C�Tm
�nH�6k!��ßs.*ٲA!����̅n���*�S��-
�6	ӯ)��
�r���!Z���p�q�E�h9+��0h��n����a��ٙr�$�f��|�O��1���&(Q/��(�.	7�b�qd��?�?E�T��8ˋʂ�Q�p~��/< ��;cR�-^�������~��-ݭ�[�iD�;�\�	�u`c�ޓ�D��ʅ0F��b>���i�\佾������g�y�+m����L�͇�4CI�;�����V{�)�[X��MF�p6&*g��UH�*V��?~K�m�4zm������?q���<��>l�S�A��GKcz!�E�˪��3��������Y�ɓ./����y��D��삶Wk���
_Z�fU)���Gу����<$T��s�4�[�Z���	s�I���p��m�غ��+z�?����2�j�V&$��� G�9R&`�J)Q>�\ӾX�w�ޖ��#�?"��e��Wഗ���+c��K�������g�~�	�s����H j����B�nAu��no����#}z��67���d/�U�N2I�d屲~�\��	�<*����|��4vM�؟+�0Pܩ�n�[�0�
����N���>�BL.w$�C�'�ڒ�3V�y�%�N��˺�;�[&�����|ݗ���s(���&�ų��fjXg6._AF&%���3 �T�*� &S^�7^���{L��Y>�>�[�}6���ܣz��"���E�\'���<`}��M�����?9/k�<E睝��>�~-�`��(g��y�_��j��\��5���-]ù����JMtBx���T����1��)���BZkq����vCӹ;8�[�;��Sի����G?Z��n��ёI��4Ln|�3���Y#�Qr'����|��|/�j	� ��M��S�,C�ر����!W_�z�k����SN��q�T�j��}/������.���s���c[!n�y���^��=����&<����<��-�?���V���9���Ӳ`nˢ�½c���bQ�����䂥.�J���fEO+�v*s����暮?|��]����Ǽ�t��%=)���9�+'�'cj\L-�K��#���r�֎Y�q�<���3}_ƕ�.]?�|���!�z�o���n'W��5/72�:�j�F0��9��C�y���_IhG�V�� ]	 �r#c���m^�
��& �p?��<�0�ÿ�jL��qxRЩ�z6�K$� R峓�K:��[z������ot��KJ��"����!�I�-�3��Wk�|����V	,0�V���-�LU����� �r�n^��ӧt��7�����￧��7�mR�\@Cf�Ζ-rVl���ݚN
���K�����_���{��/��4�5<I"��~Js/^/�$
L�U����>�f�Q�¨���)p�e��y�rX���Ⱦ��i{�w֎V�x-A�Q��m1R��%���T�1j|���ȥ'ҹ$)��t��m��[_��ϑ1[������ҁ1�_�VW>�9<P
����F`чn!��j���F$78�˫<|��e���v�˕HH#���O�9��4]+ m6�{���xSxY�@�cv�V� ��I��.$��q����T.<��]}U�s���߳x�ᩙN�K�<�9S8L%�*k��؃�� �l��6��~���ɆA3��Q8^M8]�d�m3e�x�v��NQq����$_v�vX�#G�A���dL`�Ys�U�G��,\$�� |M�bBob�xD폀��ރ��Y{�p�:w�a7��^����+z^@#�$C�*���W�d)�U@�蒄lH���ˢ���H7��[6��L���6O�5Zr{�����o���m�24ޗ��7�u�ˠ��h���:��Tc����qY�+?�Y���x ��s���pRv1�&f�\4#��_h���#$�+��e��zT�p_1�� `��w��٫�51I˙�HY�	���;������Z�hK&�2lR�#�t0?�L��g��6(��/��'B�9k(T*	-eDz9C��~Z�h��_}E_�������t��	5ggeĆw�H��ʔ3P�R�@����s��g�/�~,�]��%�ȓ=�$��J�AN#@���y_��?���}�=-^���|�i. �`�C	 �i���L��?��ym�|A7�h�R:TU�I�������P�y��3�[er>�i+��;ٛ�~�=!v_�@��*�@�����~�޵�r��),gګ�1�ڿ��Fp��\����>��S�(A����M���e��C�ٳ>�q�������lk��޲c^�
;�}wmߚ!׫���2}-x�P����HG�wF�;�y�I���a�u���V=�}����;|��#h"��W*k�����<�{���M��J��̕�-I��%���C�j��2F��E�GL���5�RV� wAu�lΡl6�8M��(�y�G�x�Í*���2=c�Ү�a������se"����y���I�3�� =�>�X�� �� ��7���F��&�W ��AH	��f
n4����l�9Lv5Rz6��a�Y/�ґ �"Oy�qOT�Q,n8Wl�xH01�%;/� L�S�`���x<[��ݰ!�lv���F/�Z�pE�2O�j�p^+֍�`["�U�j-�_�JF�T��}.���x/��1D�x��36��e�.��4|1��,JS&��U��!��K^�̽�ڥFoX���<�dfR�O�L���bJ��k����<G!�I���ƚ3 �/���~��N����>M������y)�'q󲫞/d��D�8T��g/_����~�]|��'B��V��[�,�.˭~.H��Ҁ-E��;Mf�I��!�����g{R��gt��7����	<_��@��\@��/=��(!���\X�0)��&o�К����NBݞ�[kK��(�M�۱��x�k�eT d79 �ڨw ���YC�9��M�������L�������>|�� �N�P���z�Ì'�t1�E������x���C���=�x\6UQ#��z޸����D���:��(&*�{xc�}�g���Q!ٽN�����lymN�I������T��H���F�7�?�[���`Ԝ�D��AU����?�h	�ER_�OI�\˘`�����7I�ud���z��{7��a|����J�d���덒�h��LJ�38V�=�2ī:�焎>�.�X�X 9�)O"��d�p�
�|�p�X;��R�&���h��O�:�^|Xb>&o�B�6��5-(^��!	au����R��M}�Y4f����l�6V)�|#B�ŕ�����E�!�+3��q\=Cc�'��{N�5όo^y
��� tS�'S�.Si��[�c��!��+xB��䍠ҭ�p�4��zh�Y�=xk��o�#tS݇���#��J�����8-d��X��m@�;&�d�YK.�T�4е{SL��^� ��:�|�5K��
?�ȇ��F�� ���.�PZnB��^,��`�>9=���==��Ot��Î�j ��^�9vHx�1׿���M1�e�D�����?������;}��e���/^��W�}��=��kZ��Y�O�T���]��ùUm�{�{(Nh�˗���~�xB?��?�����0��p2�Bd
\#�eOy�x(S�l�-*d7G�Ou�dW�D;kc����y�^��}D�'d�v�+��>}�. �C�<w(�Bg�	8���3N7�67{��MJ?�7��هB�֎�I{5$����Zȡ���c5�;Uv�{Șs8^=�o�����#��ߵݝ���~yS�,$�h�7M='��A}sC����sF=;��m'����5j��>�s�w�����&�lXOVajs������^��-J�3�����n��k���m�l`9��>8@���Co���߽]��U�9xT�`d�iQ&��Ü�jp�����q���i��`aą]?��3�4�`��9Y*�0����d8˓�9^N8���vL�;��Q����?��l� �-�b�A�w�HK�VG�P�3�J�<*��u�����q21h��|����{�oV�BS�iC�ey�f��e�t��oT�64��
F
<S�����uR�K��f��c�����_*����6��>d��D[O�/��JW:�#�R�9|6F�/wǸА�F���T��ė�W�MZI�tP*h��^��I�XFj�����L���}�#}�mq���%߱_��B]�=�m��E��ϟ3XB(27���J՟X���Hʹ�y1��r�Nhrv�mDWW�-o\��+mP�S����%���w���O/��=��s�Î�/wJ�9�i̲{\�ڄ������ؖs]4S���$����������m��� Tea�3Y�=�d�����p�`q�뫃��}K���A��X"�42%	=G#�I������5��-9��t�;E�>�����@�Yr~ւ�J��xT$�z��s���dS5`G�ap�4~%��W� _ٿ�Ǳ��U����?�pLG�v�W��{T_��8qy��,J渟����	�� :-�9�=��☢Gv�f��AV�����ܰ����fό"2�>U�[�l����ͦ �����\�a�⒃�Ǡ#r5��hjcq� x��/rOz��A�M�B+�6��M��1���$�t9C����=9�v��Юa�=�Ur�Ѥ�b�}5�Z=2K�w/�i��p�:�C�5Ɩǰ�#*`��{��q=9�dS��%��\�ך��y���+�/��$�/F�x]�;�t
�:��|��+N�Gr���Ϟ=c��$$o3m�I�~m���QP����sT���D�岍7��G����#`,V��z<�Y~_�aMrAT����I<(��S_A�5��F��+�l��je�~�eҍ��А��1l��U���׀�U�k)	��I��,���v���v�掆sg���BքSkY>���0d�
O 1���A4떑,��03{�����٫>UK����������?�-�?�^>Fg�-�OuQ�Ӛ��\�W޼z��3|b�o��<���x����+�+ �[���0��?�* �\�_U��7���7it����懙����lظ�!����n�;��ik �8�fB�m���v����`;)�	.D��#T�ז���l|��Fu��$�P�h ���0E�?��?z+n��2����K6/:�c�=8�э�����$?v���:���`(�ŦI��L�1��-��'�35Ǳ��u{��Z0�C��u�gE�����uֶ{�s��b����7s�c�<�+\Ry���&����S�p���Ct ��֜e:mK��	q��`7H{_�z�'<b�h�_����j��=�Uf�\�np�#I�����傷� �x�O��d-I.Kk�xv�	R锎�m�rR���3,҃�G���g�^�GIj��%�MA�Y7?�`1�p'"z��#�����.b�۾$
	�x�l��⦞W��j���P��dΖ˦gU�z�6!'$���3�9��P��c���/DG�c��1�U7S=��x�9�-)"ŻO�Lp�}��k:�2���H����$�vZ��6!���!�_x�9a����i�G�
�fx���艢
v�=WZ��mơ��@�%�����I���5�$��-�|�s�'����PI��C�@��D�&��~1k�Ƭ�P�3�X\IU B;��f֤�x)�땳v, r�� �8��g@V���꒮^����w�|�s0�Zo�
����+ʠ�,s��kH������@X?ny���$��ͱ ��RE����X���꞉U�۞�@���	�<}��9�?b�3_Rb:!I���f��q�{��^�>5�(NP�9~up��D��;H���c9���4��6�8�ѩGjȮ�p��?\\�t�%ȓl�	�qъ�!�U����9Mf�o� �S��\�H_@R
���C�u$�3d%��$ �	�gx�����w@ֻ��zS��9�u�0ș����t�ۗ�.�"*��z:���ȯw�R[��+���2�9��HJ�06.����b�2�Ӛ��ޡ!b���P�D�8����̀�g:�����BW=p�P�[��1o� ����{�|���/�L�xu���g!�e�I>t�X̄?-�N��	*/��C�~/ �c�c�(��
x����������0�D�lP��������7=�1��4�� ��~~9%M��\���B���y�a��t����RJ;;R1D�N�SO��Y i @�cc�,3�9Ti��[/t��<�rd����p^���&V����)����4�ܪ��<(�Al�#�'m�۳Pe�*�N�������� ���WW�q7�=_�����ʃ�_ͣŤx�1|U{��� Q��t5��y��Ȋu�	�Y繂t1g�@5%�������)ȇ��Xlz�|8��s*(���3�A@�{%��LF|ʝ&��pl�+$� ����p�_L���3�v�{�x�nOv����0 �9M�,�^�Ѵ�0��~�� S�G�F�lNG7����`��&��Q�#��G�U���h��b��|�H6�+:���ю}�[e�c���n�3��7���V�`m���'�}����Wa9lT/-M���r]��Z�^[�p�@���g=�[�,9�c�[�>\Y=�z.���(�7=)B��׈GR8o�6��<Ǯd2��������сU��<J�MO>hW�K��W��W�x6,�s=�=0E��
�������lͳ�z��^N�Va��+�L���f}�����٨�-t�L3���,��^�~e�X�u�{bҮ	BKgE�6+ƭ �44^��2���<�H�����聲��[��1�I�dEB,��F��Y�~̐k����N�+W��`'�[��~dx�{IUM�5��A�)W\݌�rXl��RUɹ��,s��'���s�'�
�=�B`vpl�>ol'm��(�BS{���i$��|P�銲���CQCc���zU��\��~z��f&}�z����I3�cqy"_v}nU��gί-�D��"Bo�/Ķ�x�2ȓ� |L�����=h� �ݚ�Θ�Vdx��K��������=������K�<$/NO8���H;)��r`GL'�m��9���/x-�:h�k���~E��;/��_���F�!C'����}Mm�V�d�g�?Ǐ7���I]�C�ڗ ��?�Ƣ��say�l�!�Bt���-�)k��Z ��F���1��}b�&܂�x����z���Y�;�خL��\T�`�w�j��݊A>{�Q���yǍ�Ԟ�ŘR���	zΥR�e�`5{D͓����v�}�ƹ<�qL�/��3u�^D�;��йJ�K�C�O~��WE!ˀ�d���pI��4��R�^s8$����>>qǆ�����+׀Ye'E��E�rw�� ��E)���-6SNL���i���r��K6i,Y��>W5[=�ٓ�@�%Mkn=���}��{y�{et�m� �
��Z�Gv�a�ͮ7������̫M���/�_c��G�SC��+mSx[�����cc3쀓�|��ܕ�?#kS���c�Aɠ8�n�Vr�-�m����jY��KF%`�7Ϗ?���A�� �o���z�ڰ�}r��������].����g�P:Ṃ���p��۲ozmĞ"n31὇�_���T�������������q tΞ=����N�ʫ����G �<o�Sa&y5hl�8g'�Hx�xN����~����@Nӓ'W����tV@�Oq�4���ڍ�&�V��lU�4�H:y�n�c�;��R�붣��h'U@�_��
��y%* �j�<YRk;8�N/T���\
:m���vԖ����l�����;a!��ޏ��a�V�p���]mMP�+6e(��$)[����#��uޏʨ
�l~	:�|��4ܗ��~0������Ǫ���OL�S)�E�*�'h�Rd�vW+�yV8PhC���uOV*�?U���Їb�[饒�'P�N��q��( 

Ǯo ����'�SZu�lўyC�'+����ό
T���G����|��$L�DM�0������^���,�z>�Zx�7�3�U� ��嫅�n`_�����d���:r�v�07�uCj>���q�䉆�wC��m-�9���R?w/,'��W�=��A��j���T1��4jo������Qk�́�s(D]f��c��Ѫ���!��*����DK��D'�d�槙e7��l�������V籙�w!X�������2:j���GM�߱0�ퟁ��T�?*Mͳ��`2�K����|_<Q��~&�m��gL�S���<HWի6U�ǽRSU�Ҧ
&j�����U��[��/��_?̥S�8���i7¬�tv�4�:���l���(bX�D~��~�������AsQ��/_j��� mn��/-��M8QI֠�W�.�cJWk�)�x��Wz��Ol\��:����0���a�^�w�a�[�r�5'�aɞ�5\͹���i�&��(VN>v/��>�I�;�
HU�0f�����h���ߨ�}Z��%��=�Z!ӞL�<aH�Jq4;����6U�dq��`���-�В(�Y�,ǢŶ�{�(�9�^��]����ƙG�ynܟ�=��G��#	6��&���S#�^�5ﴓ{�L�9�k�w��Y
���$"��6 ���E�:k�V�%+D��2w�-�/���%������ ��b���nKF�, ����\{�a�N�ѥ7���|G���u�N�1��@

4�e�cOݾ<Լ/� ��nNP�t�L&�uxÏ_�)n�(�4���ԅ7�ƪ�Un�	&k�z^��Q��/kmϏY	�<�MB��zC��y�������=��޲�B�ާ�sK�f�P�(0�j��,�X��2��%���-խ�iI'x�I6����ٞ�ݫ�ܛu���(a���'4�hQp�9�4�q�~'��� m�Gv�����#r(�p����)Yqf��$�:����h����i?#k�A)(m<���zR�^x��dk?%��f�m�I�*�Bd�3�Ĺ���妚O��I/�p|�;&�d����7R
{��J��" ˪t�Ė���(��I�dVqǡƮ�� ��"wD������Fg������?�����{��dFl�1.��R�����-s���	r����}Jk�gBh��
V����"q�ڞV77��_�Bo޼�;��kCk̀wƤ�Jk.���8w���+	-��$��fV 1��pTv+"��ws��h��0[=s��{}m�9�P�\dT�n2��|!�+�P"+H&0oh��gz�=s9IO_�n�g��^]P5ma��2`�����i=�x�k��%~T����z����I/x �������Q<d��jP�Bq𮆎�����¸��AX?����%a�Za�`QX�f��LV���a��˹���fH@@��������:�/��[��▀�U)B���������¿��<Y/��i�X� x����Z�^;\�Sτ�[ڕ�?,���53������ؘ2�оTB�/ƍZ� �
2$MR�Ϳeih�����Ix��e�c1T�h�#0��^�M���O��ni^����}��Kg�{/�HV�T%_��=��$$'��V�΁���S ً���H|��f^�����ٴ�y�s֚8����)Vi���d���`)G<|TPf^�~��-�/t��g㭩u�� 5�J�}	�=�p}���ѳ�2�?��N��;V@ f�Jҥ ��mz�a5n���հ���	~8#O�9��_sk�v� ��3����ࡹR=�
<��#�B���q6m!T5U���I�AV�C�t��||O߽����iB�V���у�# \�E0���	ʜl�+p��RO��CC��Ak���Nl�P]���~�ᦿ ֻ����y�HۉYqU�QQ�0�E�[R�4��
f��;�LN�h���)Q�����t��\)U����d�#c1^0�|�x�µ(��b�����(�����>�P݋��;D�� f���k�B_�ڳJܻ�$h�	�?�ګ���P'��˅���?~+Dk�C-(3����_s����#�G�s�*��,�L�h��h���0V�.�'�7��ݸ���D�eTe��;���8�)��D���PCjR<8�tb����~Ka�9�7�`������É�ػ�^/i�Y�'l�e�:��s�m�S��<��$%���6lҢ�:������9�U-`�Napl�kX��j�\�6E�&���)�Vs�F*4v�ב�=�)�ǒ�3�aR4 ���2^<0��޾���޳�ϝ�ӄ�u�ɜ����{�O�O�ـC/ɐ��hƋ�Sd��9Ε󄙍��T��d7�6vp+v7�q����%JQ�D��M�>8��&O�B
���Y��,�c��&L��q)��ac�=&�k�p+w�Q�"we�<E�_�����Y�Ó����A��|IK�� ���n�ۇ����S[1�"����2���N=�6�<2�m'�d��c��Gx�'yB���nuMs�N�2���]\]�l1��fҲ���&�fx�`��� �hp��r��9�A����_���k���_ʱN�8ؓ륐�"����\��ш{q��� a��} wyA����?�z%����ap� /��a�/4^�wz��z�MQ)+8{��oL��]x5x�ސ��7�R:l�����C�q�����<�$��Ȇo�!	y����ď��b�ī�*����;y�jȳ�3���:�����#E���Ұ4!d��}��/%ʴ�0�[1��#����uD�^~����b5xꇫ �%��"��� 3C��Z���e]1��z�ߙ�����w�lȲ�)U �O9��4����f~���&�w������ ]2zR�C�_?�����^>=�b���{M5@�ے��bP���v{�6f$Ge#*�6�#wOAi���Bu�v��+�����D�� T�]SS���yJ4�#KzR�H�_>JyL��5l�� ��H�j߮9�êȄ�}3K�hR��*)<S۱{t���T��C����12�x�t`�|�6�z�k�g[Y�˂������G
�dQ���Pܬ3IR�)S�6��ƽip�:(�z��q�^Z��u�fb�9�u�̞�e�Jբ#"�ٸ�E*�s�{�*>��r>��c���X���a�L��x5i�_��z��9�����\�
*B֙�W���UhZF�5�fkk�!�tO���g	���Z�iژ���x�O���ѩ���*�}9~'�C�k�h7��>;s�WK�M�t��2�K�b@Ӫ�|R�W�~d�\�%C��;���LĚ���d&nhr��Dr�	 � ����u�6\��d�W�^S�����ⱑF��H]���a��K�
��Q�ht,?K��&7i�ԯw����k��W%,��.-��xU��*o����kxJK�j�!"���y?�{�)��A=0�M���s4�p	�~���T�8%�ȁ��|l>��;� ���3 @
8�Ȫ����<�2���}��ɶ
���c2A�FQZ勖�ܛ�]={����;No�[��uB�x�M�?����H���4[1�[��z����.O�ty6�y�.9�%+�^j!`.�g�J��n� &�hףw�@�ȿ�^`��4�"ɻGĕi�������ܚ�U���$p}�{WyJ�q�v��"c���$\ ��6a���'��g�����9�ڴ3��϶�-s�$(�� l<��+r<���:�j�"�wh%�f �+�'�:���/�}�xC;:aB�"�|q��v��}mNj��>M̙�4�~�ɑZRL���+'
��H�iJ~�ny�ʜ��m��盧�@�@�g8�� kb���DC!�y�c����e�C�U=w�}��:C�P֋f��w�s��mrx�[l�%�~/����@�v�]�獊�!x+����(2��I��7����`��<	M�-�ɸ�,�勧�(� P,Y�K�;��B��o�J����K�����ܹ����feq:�*��E���D�lE�����ީVյY����i��yh�=�!�J���_
���rd�]^�W�}G�|�-W�19dC��I�ڬ�ٕp���
����\ڍpa:�-ћ�N�u.E^��=0�d�ž+��5�;�di����Bz��^x۪J�V�﹁8<��VHS7�t����<�����"'���E;T����X9�%߶��c����[�q���g�*��1�K�D�xΐ|6�Ń�t~{qꇊy���0��1��� �tC���!��N���si���c����I�))=�4��O��sg��$�FѬO��y��3c�`�&B��L&��ڄ�5��Cc_������W[���;:�5���:�Oi��=�!��ܯ"o�޺5��@X�	���q���b�26`��P���-�s���agi.(_4?ߞ���e�8敬�+��,� �� ��.h`�TEhd���hǱ�%{�p���(]@�.!���dؒ�p�¼r#��	�����밢<�����}�4���݊���2�%r&;�Ҟ������>�����(�EQe1��x������b��"Žr<����	�^�:��	�kw9��7+k#�������V�8$8$#�������������Ňr(C��?�A���(X%�^��1+O�8̍�U;�u�����*Qj"i���I|wkM�.�H��ޮ�JQ�hu���7#kH3s�$BY�����J��cn�jD����Ԏ��r��x�@r̰����:Y� ����)�WF��jE���P��t��<I�|B�Hs�*
=�jXHIM1��^��� ��Fmu���v�1̳'�sV�����|��R��䚽v���!����1rD0v~�"`�#�z=��V�2t��� ���6���Vڀ-o��!�ui���g;�k�
(E��pV�z6�q��|P�,i[���v���m��ؘ��� 7��X�K��gO[������k�<~���`X�u8|��:8����&�#� roZ��c��Ƨ��X�GF�R��l�pɖ����{����Z�%�;Z/bC��\�0Iz����q�y�&2�����E�PAE�`<��(J�]�r��S�)r��͒޽�Do�}�i���I.�@+�Ux�u_q�-dD�d��(t/.�߯�Iv��>X�;�W<̍\���� i+�}͆b�����\dn�|w�/e�_���3kG�8�Гf��)�'Q��w,3ha�7Nf_�y_.���z�N*���%��D�g� b����a�! g���+���J�<t`P�ׁr �a���a�07�WWƹ[���iʛiYn�_~�����[�]����>c���0Y]`�~l�=/�d֓�ɽ��^���QuC�w�B�Yד	Y[�4�v��DJ��(�h���;/�;�\Ày:���b:|���1[�P��w�pH~욎)դo�GJI��V�*��l&Lލx�!g8�K��Z��R�7���X�l;IR�8Q�����:I�}�l}�]���|�.�������M�n�S������_����F�G�"��W�{��	zK5@�P��nSx�gh\@��C�@�zQ�Ai���A�1������$��Y�4rcɥ�D<�b��jF����=/ ��g���/����d
L�˼�q��"�>��f�����������d@^@?5���*��c��R��9o��I�n�vJ\�����RiX萑{���P1�&��h���@4��?���ݺܟ�?��{�I��d��|U `��l���P�*{���<��/IQ�i�yL�0/_n�bë^�� �J��tc�Lͅ��s9Pp?�B�|<�Bo��1��K��t?Ô:C���@о�����NT�y�H*�=��$���qL�8�Bβ�l��&���c溞����܂1@w�� �!ST���yG�����_�_�w߾���EY;?p)3Yr����wY��OivrN��K&*7����]���w(�vg%Q��
=L�XZq�����x_�x)�!0V��pv0�?N��K\���	=*��yrv.9�(�h�5#���9���B��-B	�W���{ID�B^�ꎶ�r�~9��*��8��PA�k2W���g�0�*��?�fe��j��ɂ@CM��9<���2���X��EI��2ځ�n���ӛ��˯	9�;&]�/9e ��)/2n`�1��R�XD�{���$�g��"nPp�ľ�)�,���l�;���h���@Pb�]Y�~oU� �}��<axC���z��[K���I2�UM(u+�6��Z7Ir��%V���0�0v�Ӝ �wڕ5��*�Ze2;+L�V^�9ƾ���2fi��s��M�W�mr2��f��0}�[6��#�_�׏���a�U�� O��a��Ҥ�1c�z�=���o6�+�g)KC�L��k�_�B��JmS!�8K��Vb�6(s������6�C���<�a1zއ�{�jR3�s��D���=[CO��-�T_�[���V?<�z�lu�� �mS	�̝���1K.,�.�9�ޯM����ԜNB�s�\/�Y��Q�|D޲����r��
 �>ZE�0��a4c�sH���kǲ4>?���ݭ�NZ#�VUX���Ϩc�4��y��e�5_G��M��b��z^��?z�}�A��Z&��W�ʮC%י�^Sy+�/3E[E8P\r|s
x�2k�΋�A!�Z{�ve���o�_��W��� �ph\�{�3���sn�ZP��?3�������2�VU�,|흤<u;���h��"c�n�Cٽ��f:%� #���������QP4���*�s�h�$�ph�Е&�U�K����m���K6�;cu/�=H�3�c�(�X�2�@�6"py��.�1.�L�������k4!�]��J�$��9O���2F�I+U�Ed$�b���𱀯[�J{ϡ����ۻ�y���}���5?+�s�.�"99�0$��^{0���uAr�g×T��@�	����r!����#�A��X� �@\ �#�Ib�~���f'���zA��=�����]�>�����Y��"k�+=�Y���f-[,��+�,���ȡ?�����W�W�;2�	W:��K������+$���+�Ly6�u:�S�%��ra3P7@�#uG���Y�� (i�H�knEfTs� �7�����/���ꂦ'�iylu����Ss*٬+��2�l'�4ENt �l4فC��)*���!e�N����3�(���½���?�#���(��S0·��9��2`BdJ��A�擳SZ���,!Q���ަ��W�։!z��Z�g�L�O5I3W����*��}��=�%�u �4Y�3^������]�����~O��7B�M��6������ u�1�벡��w�z�D징��~x�������"RO�Ko�|��7xsln�j��w;Bej��'18��GsM��*�d}���r,�����M�����(;����\I�S�A-��a4���oz$�!���c#�s.`��I�U����͋��*r�O�X� L�Qڰ�|��Z�8?�%ps"'���x�f��+��{,3o!�Q��l�U����9���c����;r

�V��RY�s,i	�5���~ٮ� A�޴$#ho��D+�tٳ�LB����3� TaI)|�����Ď��n�ܲ��0��y�䦪�4UK.�E�:c�wt�<a{�`�]q���0�����őzl� C(۽�����#�/����?�޻�[#��o����ǟ?ЇO����� j=���t�nPp�Y�X6e�|��A���9�R��D��509p��ym3g��V�0=�x��T�E���0��z�*S8��q���u��Ee��~14�=��p�n�^�\���j]�n�c�W�(�X%ZH[���L��L�_�r�H�8��y���k^��ro���"y`��5����x���y��c<��ڄ�He��z��gn+3������g\���ԯ�p2���)�:�������Tw���r�FT*O��D�����f�Ţ.2�݇w4��^~��]\PS#�b|6�ԛ�z]Z�d慔+d�t�P��|hY���k�Xr v@�`��b@sN�NV�����P�ZD-2����W��g# zY���@�)�#<��ږ<��@f�wk�hp�"�LuB
,�
��R����wB l9�D���ZɁP8��ኴ��4X���W��s`�D&��):�d�+�(J��� ��-Y`��t����ne`��UNE�3��j�O��CY�JV��

Ƿi���q�g��\&��US����"�L"6<�V#f�G�������Ǜ����:_���� �&�F��C�)���I�� �0���.ˎ�4�$giԫ�mǸ�ieϦ5B�L&�M�ɖ֐kkB]+��5�L[��RDa6���p�L�݂Ӡη�s=���lU>;q~��ת�N�'3SM� �� ��RO35����d�.�G�ə�!l��.l�`��-�U�7E؝�y��O���D��Z�+����G�Vh&���-��n�!��5p�z����[����/�/���b}O��:ἯԊ��$�E�tHfE^���h����1ڻ�)(e>��3k��)�#(KI�>��ܫ�J�����K���Ł��z��)�UF��&�n
b'�ύ�7zǀ����z��]p����$]+�����<��b�j��A�J���%[_B��qG�_6M������o��kM�L�{j��DVʘ����F���v�oxD`=G�]��$�
��<'�"	B��Jf�+{nʍ���ѓ�!T��)8G�3i��%�B�e�wB+_O^����P�@��ݻw����ʹ�g�����3z��5�������>}�X�e�o�n���:=?+��T�dQ��y>i���H�Ep[0��*�!
1�t� ��ҽ틣O�&8c�15-k�¶|rv~Du�GIr0��T��:	��l��XoQ(7�-f���ۮhyw]��	�ʺ;=���ײ�G�r��t:��0s�ĳ�T	([6�'��ɚ���)&��8g���

X��g3eQ���5+���a����4>�+%8J�X�?jA��.P5�cU�lMd��Y�e�h�>#�d�Z�F�E�Wbr5���ʿ�U����>g(��D0؈q
�Cr�=�j�d�D�"��U�{�=W.������j����N���Ô�(�Ym�M�[>c�����;+0�o��$�r>+�"��,�g�ܭ^S�x�"٢�g.��,u�d��TP�.$��P)�*k�
H����	��-k�+�ـTz��v��6����ֽ]��qS$���z%���}qn��q[�~՜Q�b�w�"w��UJ���s�I�8�y"l�y�I>�#"���ji��X!Y�dԎ��;M��[�����yC�����-B�3_�V]Ll��X�R��u��Bρ9;٦�6]��L7FT�����]�����n�<�8%�j�pn�Ƿ��{H�ǫ�0���jE�J:_�<���:���J"�ü���g+����,21¡8L��1=	H������i��B����(qe��y+�pJ S$���*�<ٸ�R|�8��g����'W�W���Vx��>K|R�&_�Y�q\�Ĳ�{�4۽ʙ���/^���+�{��v�ˀ2o���) ����_��'���.��(��ϼ�/��7�VjZW/|}��7L��s��b��>|�D�����/V��D���^���_s�j䶧m�Z\@3��Y�M����/�4#UëV�b�Њp�ip#�?#����Ǧ,�^Eb 㵝&+Kx��|/��A�Z��tN������?���@�If�b薹89�>��|"m���O}�:_��\�/���j��=�0`S���Pb���r�'޿����^�v���=��(a��y̫E>5u�*�?���E8�q�h\.vFC56��Qv�"~?����sl�}�uaI��iʭ�R+-ɸ(���Fd�n[�q[��nvy~JWgtU��|֊'K���t9o�r�s�m�j�{�c X�2�;p5v��,6B�0�E潜#KT��>7�%f@9xM#)���E�>��h��{5[���*�a��o~)�mtC){=��S�K��tb.;C���]�{���I7I��ڨ�ƚs>�y#Un��3�I��gY�q�O���Z�;ˠ�
²F�3�A��a��yi\�J���p�l:z�������
 ���}�/�o����R׀nbF��ǜQ��)�������Kz�pqg�.��	��'���a���������+m���+r�R&�u�O�V�����笗p�1��r�㌿X/O�p5K�<}�^�|���A����&xZ��Ny�mA�R��f% ~:Ge�d�p�ޑ>�jӫ'Ӏ�����n4.�Jq@677��
�s�cӐ�5�.�{.?��)����0@3��q�rr�ᖥ��^ֲ�4��'�~�+�0,��+��������"��ΰ+�	!�UYח�����|��7����S쟳��WԔא�z��]>{B�O����ў�C�������R����?`�O�����H�x������=}S@޼ ��Ty�:�;W֦���lo�nk��R��m���©&�s;12Π
L�ʐ�2U��2%�wĘ0K�9{�5�*s�Oi��F�� 1��e"��J�I��W�l �x�+����j�h�,��^�7��	� ��K��z�s�<����<��!����2��`{����ums��Ϯ��`Apo{S���! {/e����^8���v����^�YA�̥��2������z�n������J:D[��y�(D :��E�佡$���F��d��2�3{�������t}sGgz��)�.}EϞ�8�p2��)<VL��붫f��+rU:�⹴,3p��#�:%ٮUǌ\s/���9nT
j��؊wQx�dR�����b�b���o��P]���`�˨���o�t1�$8X�\b�#�0!(�a'I��7��O/ya��%�*����$w�3���Me���:1I��[���阾b�!Ѽ��Û�\<$����q�n�V&�gs
I��K�t���-��Ƿ��Q�xC�<tM��m��3���0���\�(l
B�*����+G����dsd�v���,נ.�$�}cT��Ǳ�r�Ó?0Kre0��駇��9�g� 􂨍ޭ>�G2�s|���Kg��a�d$�T�a(����p� W����y3�^^$��N�KB�5�GQ�!�^U���L��@�H#{��+Ty�D�Vpn�)5�D������N=��u- �k�Ղ�g�Z�	�ҎN���fꦔT.�� ��
�C�+u�O�/s|��m�-}��?��t�s�E�)����z������O'�_���j�T7�1n1ϯ.h�t�>kr.�=����H!��-��ȇ`c���s�u���i���׈�!�#��BV�f<�ǔ���XQn��[^Ɂ� g4�ߤ�0��Ođ0	@1q/�[CNɑ�0E��6\��$T�f�I9~^s��ɉ�{��eQ�ohy����V&7@��f�GX��м<a�N8�c*y9d2�Fkl(|yڿ��O�i3�b)�x���z��:�cn�"�k�B%�&!������\�n�c����츥*�j�ر��nW������>��!'��S��:?yp��h�]Z��ME��J��+���)C��o��F�4�x��V`��E'�n��\��v��\P|v��t~vBgtq�����(Iy��E��5�CtC��̝t� e���Ȓ�\vW�ȨM���d_L�c�R]T����b���y���Ӛ�V5���@m>���Mڔ��b!m��3�uAq���j��!�Z�i�fCf�g߃�잴ԕ$����N�_3F+�@��[��7��J6x�X`�))$���,�9� )��ٛ�{&�����~��=},7aG$�Q;�}#��(�'4Y\��FBݶ�i$�/�Bj��`D��gtQ���4Z���W:�4k���TjEF���pmSFa�Iï����`���߯�=Ǐ�fb� ���K��UZ���^�����u�x��&�H��_���/\o7�%:;Eg�i�PR��Ȕc�s<<�����z;{K��&�u̗�{�[ޏ���0v=���$���!Z��h�_ �\�~Ev��Z�x΁���	Ij��\4��Y�m9�C��\X�/_>���o�����=�%9�,A�H�TI�$��9ۻ����|Yq�9� �(�z�D���kv��#��3g��x*2��kꚜ�OH@ь2�*U0u��VE+? ��ʬ�{s=�%t �4'��ם�� .��_�;�z��<y����I�|}S�����W,weI���[�!Ɍ_�3�eT�� -L�c'�:�&�X��S�z@��c/����z�)��W59�Wb�f?������.�Iv]h�{�ap!a�P��yպzΐ(����|~�F��A��}p_�o��k�ˁ�6�:����(�S�!P�^:�ժ��zò8��:�"�#YRn�H�i��6���_	϶Y׷b�����O�8]�%	�V�I��U6��AeH+�$�J ��m�� �7���)�w.:c�c
x����\��)��1�ޥ�À�h���G�`+`��'��4� </F��Q���_��7�_�������wo�Q`c���r5R��f^J��ZW��f2�Nq��B�F|��~�hkR�����C#����v������k6�G9�<�c=���'�������jѡ� �`�3+id��������g�'"vS��B���=6&k�n������+�)�\�OD[�:�V��Jݘ�|AZMyV���q�/���������׿�Z��-C�9NWU�^ɰ��z�F��UT����Iǖ�f��M��^�^|���m?�~������[��c)�Co]��ǆ��* �Z`���_K��[��޿>~-^����-�Xb}}�A��[�{	��Nt��9r�Ꜿ���I�m�oTz���
��Vޢ�95��bH�Ʉc,�J�����sa-��֊;n#&��ޢ������N���@�/č�b� 1�,�1��=�F���[ŔCX7�������ͣ�yA�6�`�g�zU����зKP��ۛ'*�a��H�n6��z[-���䤧�U[l߽xi�U��c?u���~���*�,��ҷ�W��qP ��h�o���BJ�o���b��S_^�Cű�=�3V��4�\���<0����s�FY�7c�c�	���n'�ӓ|��T�S������[�)*��p����WϛR�bo§s�z<�����=.%����$�p�������5��@<ұ�jM���>{�w�ⵖ�ί�s����K���c$��:�cG]X����ի�\���0ͧt�o��c�����iPj��-��Vci�qf�T�Ұ��s���Q[���r�ΰ��d��u;!�.�>�Y�H68�h0z�J���eh�3���
^���X�r�y6����;^ ;�e���[����N��`�F�e�.+��2�>���H{9fkIa%�:dm@Cark3Y5��]�-Y.h'�p����)F�J=�Y�A����ಝo��2O<F����2pkB�(�Ơ����w$�Լ�������0\�[)�^��V��|]:�!��T���ҙE=��c0z7v��kz�ZWl�FΞ�G�˶m[0����������兵svW�P�W�_�Oz\?O�L/��:�JD� ���XF�K��ߧ=��O1�T�@L��鐰"�����ɬ��_�����*����1�`C]%�����lI�}u�*Nq�v�y\a��0 vԾ�g��g�^���sr]�a� �q]+�n!����r�Ӹ��y�̦͐�O�|� ˛Ou�*�� hL6^^�<!<(+�E��$�p�  T9IDAT�T����&�C����(�c��ɀ���t�yc
*��E����$WŎ���򉛎�]?�dz��vyz9dB�&�D���A����[�U�>x�+4�^|�v���ʙ6���M1���2{��ө�@�,ɪ�PPb,���7F�#���Z�o��GU�|�P���~����ܨ�M��Bt�D4�
|w���! ����CM��~���k�gؒ��b@�bm��)4h���o�u.�P�BД a�x�q��/ݼ'' ��ҹө=���,��'>��OƸ>�W�I�j ��'�f-�q����G-�2��W٫ @�9!�}+��>����g�j��ҵ	����\��'��N�����Zs�^�V�|��^�&�х�9
����p�b�ս�0̻�++���m +��-(q�ʏqζg�7ƺ :^[�[Jo��<�u��hE�z�V#�p8���W�4p��(ȻH,�Լ���}�O|���q���IQ#��,�"���0��� ������n��n �R|sL�)K
���{�����\-���y������;������cUik�ޯ
���*��*�o�~�s�Z�h� &o�-l#a֢W��X}{�Il���_��f��q܌œ /6�ö^1�pp���ںR�Ŕ s����]^G��k�� ����-�������q�����-J� _kJ��iE�[�6#�{��6j�&G��v�T=?�	�k�|W¤��]�ي�`,�l�G�(K����S
m~�
�GP�/�����{3���Wj�uX��B�U#;��E��W��x�E>���W��7��[VuR\�~���DOVG���U+�7oaQA�l�(�A����Qܣ��91_��0R��?o\�G�J�Ǆ������{������-�b]i �i����nKc����0%c �P�QZ�5=�7-pa�{`�k��<YwKZ�@�u�'����Vi�(��K�8S� 2�yc�3(B�{q'�_��W�_�-(*���6��b�a��t6ހ�^�:s�ɷm�o�^�]�+Ţ]s��O�Ǯ*X�KQ��a�\F�Cr����o�v��;{����g�a�Jk>Y�IFa�/��|\܁��9�q���1��ڀxݫ��a��t��L
@��������i�,M�]�ȝ�ߗ�ׯ?m*����핼�@!I�1�B�܀��vb%�&w�%�[(r�j(����vڰ��z��ъ����ۂ�Z��2D[1�U��H�u����6#�����_�gk*�ԇ� �{I���R5dG�z4w��C&j�i.�`9-�tڻ�3Qy����7%���V�.
H�ps�<���tDm���I~{�������G���E��t���Yg� ���cW�}E����R�6W�g�M�P���*�YS
�� ��2��T]@�n�8�����-0��P�ɗ�+���\<��mְ�CY/�5&s��g��c�{��>�/�_/4W
���z���\� �����1�(�<#��q��l�X�|oS��1�w���o޼Q�~[-x(��/��Z/�j�l�TA�a�;6K�,w�jVd�y/H��v!�}A�����HMa���v1kO��g	��+�'��\+��y�y�MZ#�!��q�}�LZu������,�u��뷲{�Z�P�M 6P0���ͤ�H.T6A	L��r�� n����������I^Up���y��?ȶ�HV-v���q]:=�IV�#�����-�K L���_������G�摝z�H5pT�UAX�{�Ʉ��i�&.=�M�|}��)�8 �o˱+��a�#��k��Q�8Wa�)dHQ�Ǎ~)[�;H�M�Ca��r����Օ�F��~/���w~�js�@
SFHŢ>�������^ܶ�;)ű�NM�4{�`e�$Ā��+'�5��26��\����Ⱬ}���Rn/�K��d�{�WVp
�͏-��Qx����|��1��uV�������qT�e��:~E��8~�0J'[
�ek��G�te�W�������ko����d�����j�G�X�
|g�+[V��d���Pn�|,�No�z�Rs�$2<�����lI����;���Z��٣�%	+�� ��SV�I��%�N�*05�� �>Ȯ*)l6$`Z�S���Ŭ���Mt�c����䌚����FZ<6
��=vJ��5������h%�5��IK��b�a��Ɉ�0� �9��C`p�?Â���:��6���S�i��Ev����n��#mk��8<c1d�g�=�^�ZRx
{@.^� �=a��N�&�9���6h�)8�I��R'O����5���^�t�[�-���W���ݥ���F�[�	�Z̥�$�Ɉ�%���G&�h��υ4�s�'%���Q%���OB��ӳ��n���(�tNB�u�t阰�����{C�XAr9�T�C��KXJ���x5���}�q��|���������ɰ�=B��<!�zu-w?�U+��޾� �nŭ1��f)�5n��
��jg�JU��˽��������r������l�oS���$�M�ݣ_B�J�K�y���C���d֧����/��/��?�$O>ȵf���=	Xs�+Lܫ�O�}�o��^*LU1�P��u�6��9ϐ~x0oa�u��K��aL�"b2��Ia��&RƺR�|?�Z+�����
���u%o^�Q�0B��T��(������SC:���ϲMC(�~��k2uH���ޖ��u��Mi�_�
��6�NUQ�X�y벽��5�jk�e���u���j�>M���~4:���2dB����)�ܭ�:9�=�������_�k/z�d\�Z���C7*�=�d�d���#jN��D������ Ǩ���pд��v�A�NY��,�
�9w����vg�%��.M6�Z͚̔��HI�7%җhm�π��Lg0P(z���f3��:�݋��Өc�X�:d�kc��p���0b��w�fNG_5�M�H~� ^<��L�q�-I��5$���J�\b!J<�N/s�f�%`��@�%�V����2gn?4�(��y�0�������f]2Xv�6��r�*�3��K�Z�Gs�0�t��ʝbw�����oP�� Tf��~��[�IS�fb846D���_�� j��o�#�����6xZKAQz��?�:W5ht+�-�L�lU���q7i�\r<�ZS4d1��i�) u����?S������3Z�7'*n(��w4�c6��5&��w��*;����[Ͳ���5�&HK��L7u������|u�W��,v���;�I�P���^g
���I��?�����W��A���Wy���{�J�lU��Ƌh��9?�|if��{�oOr��A>��|��2o�E>?ʾ�T������������KE6h�e3s�����G�7r?��^�C�?��������.�~��ac�f%�ǈ�)P��bmL�nd�kZda���́��T|��
��y�[�ɑ^i  ��8�`�hϢ�0[�R���)"�HF�0�~�����O���C��O+X��Ӱ#�>)�H��������K�n��@�z��xue���J�u�k΃�b-�B�\��H+�}Y�� kU �Ĺ��߷C�k���2��8���lq`交yW�K�/J��;R�vI|5}�0�X�d�w�Wkj����\�}�5S�.��t)X�G�K�e����^g6J	P>!�~���Hd�s�1<W��l���]��;5�����B��{�:1���A�c��Ѩ�c����:�
�z�X"�WOZ�:�9>��V�LG�'�9g��g�p�$�_4��Z	�-_ wG?A��4�B��y�^o��Z	���y�"��s(�D!e����r44�U����#,J&��(eNd���ڢ ]=a3�><�:c�q�|!w��K}3�[��Ҷ��|�r_���z�����(�|O8��=���:H>]�a%��E��s������5o�������s�P���o a�ض�x|4K��o��}q�W�����S!E�ޢ��rq�$F��w���}X�rT�<1�� y�{���K6B+��+\�_$u���VE�B�W|���͇��e��G,�������_�	�eT��]�J�AgPX�&�>�I���5���z_~�j ���~'W�^T�p/���N�ϼ�򬉥7x��2���Gy|��,������sy���G�*�*X��y�ɜ�;V0��I9��s��{�����(���/���e<�d� k`O���-y����qU? 4e����̅ŝC�70t�Eu5���Z%�u&�O03\�=��T:��[��]��U!ik�ۧ��E�}k8��M��9 �0����{p/�܅�d��]n`���-刢�lW�Yj�q�O�����J�O��XZ�=���dˁ/�H�
�������C~=+�;V|fyq���B5��4ky�0*�)�����<L��.%3��Х\g��u�x/�ձ]P�"�D<��C��T�X-��k�-
wl���G��5��$��x�s���X�k��o���R��U�ŷ��q��#r���=�b��@t(��َh���}H���� ,²tT#�	n��z�"w}:Wr�H�"��i�D3U ξ�c�e51��A,��2�|�,�I�
y;(ˤt��4��''��,��_�m�������L�@��-˙ +��A�㶩�{U�F�Y�H�[.�� � �M� G�rE߃�u�FZ�_ZWt�k�e9��|�4X���\T~`��k�Ð�@H�����`c����]pǘ��_	�X�"��x���u�W���ܥ4~�4��h㩊�K�����\X����ϟ��Ub&=i�m�7:"����Z��t�y��:��ǲ%�4�� ���h�3����(}�h�@j���ٍ��~�V�|��&y���R��o^P*ؔ:������Պ�𰏵�9Q�� :N��R4�F5��y�yn4���g���ѵ��_�]~��Or�捼������_��w�3���}�,���r��[��4��||�����<�������a>+({:ȏ��k��ۗru��t�SVl�C ��K���,�4��t�C��~��������w�d~z�s3����ZF�u���V���8��
v,f�on��̠]�����*o�^�L�J|c~������:�E��;�q����V󞙇�E�Bt�"zGF��427m�FǶ��ʹU��7�7��)�Ga8Ee����*3b ��

��Dc>�߹�oK1�ӆ��������ߠh��ϏXu��N��Y�S�hKܟ�H�/�LRn���Gh��W������e����R��Q�k��[޴�Vǁժ�c�u��^��*�^r��|���m�к'd�C��ё��{�Z. ޢ����}0]��3%t1��M��X19j��C��/�W�)�G"E
<� cKޚ�'�[� ����(��I�8�X�����D=�Fӳ�>�Y��Mt��\,��|7<i�#�i����m�P]�A9�ك��X/�|� ��0d�{����=R�����ʾ�z?�+��k���w� K��p^��bB��b��U�`�J�4�����+k}N��|DðӰc�7���^D��j�r8*�jz�F��o 0B��)��x�CGf��D��Ј?�aKv}WK�\��� qN�}��r]�S�'�������1��%-auyqK�[����Z|�Yc���6��#%����nD�2�-���o4��t��#��WU����$�e�VDI�&�報k�'tS��B�׳��d �J�7�r}}���~�zv1���Z}�����_Ba�Wh����TV�V���n&c똌�z_���S���
j'y��Q�?Iyz��?���+��&���;%P9*�!�a�=<?��w�ʇ���d۶��\r��B��Ou�����"C��)h+��$�I��2B�f���Ј�<(��׿��_�!K_��Ɲ]�jN�Y:F��t9���U�%FW1U :e�V�7K��������%�� ~�C����j8e��R�b%[Y*/�1��T&c�7�=��Y����`��_s�aq��n�ߣT�}��	�Frb^�f-̍��g���hF?6%*�_��2���m �8k��Ǳ�F���P1�G���]:%dP!4Vx��z�d������� b4>	�,*1.w�3.yh1706��{V��ķ�0b�x���1/vܠn��{)�CƧY�g{���t��X9���b���c	�പ`����8o�8-P���0�F��>Yn6<�Z�ޮ� ��ϡ:��z�*���"��m_/�ɋ�����bs��"р��`�6I���:�O�p��&��	�⳽�)������+������yO)�_��8�^�p�E:kAm�~�s �E�.�ꝅ|C�8��e�-�QRY�dC�n5䈁��T�[3��K��|�����&m5~��h�}�&�O0���F�mOz�v��	VA����U{R�/��`��˽s���}��������vLZ!�&?b����>SV_��I����N�_CKmQ���|\�nc���l�%���+�Y]��*�
��Y]��n-�B5�-[6Pԫ%�r�dh���0���.U��b�7�?p�[���`����s[�5��v9I�}y���x^���)$Y����x9O�4d@��X�-�l �]#W����;Ϗ��[9x}��gٿ������Ą~��7���w����޾�q}��Y�����/�hnV:>�5<e�<��ўd��Q~�������]ƻ
bQyw+wo^��?�A�^��-�ѻ��;dnG����w�ӿ������?�M�����W���jo����#r��9"���s���p�s��B���%��D�xh��<y��B�Q̷zA����X50�4`\_�:��*�O����#`ki����L�k��f��j(�U(��x��
��o��~�P\Z�?l4�R�޶�V'��@��(?IY�V��1�&T)+q�d���:��JV�q�
�0 �+G�Vո��SM���~��.^1���]ԦL^l-��u��w��nQ���
kR�l\�Ct{���)/P�n��ظ8�I(.�"{1��{����J}18%�jܯ��8u�Q�УV$��Ҝ� ,I,ef҅`dK�7����"g�QqDꊖ3(�_S�>lx�h^C�if��<��JY�L��SM�� ��TZ/�c��@Gs�+��`�i_LM̨]���2i�SI���)/k���p�J�lMb�LD�ޮ 	�͗Tq ֬�U�?jx6���R"���eaW���A�$f��&�G}�+z1�dT��i���cr[�5�)����>��|c��
0�@X�fZZ�=��D��0�6�|�v�.D��f���Mƣ�\*�j��V����0k��{��J�8h�A��˅`iǺ��cݟ>��N�����^x����L��,	Vk�	�>�-4ہ=�<U�rY"��͟�ثc
%BK�Z
�6{��K�G�yb�&-���r<�FOFt0������~�`ts�Ǧ�g�YWb�P.@�
ޫ�!|�ܤ0�~�Xj�6 i~z�#�T����N��o( �|� ;��(��A��^(�������Q+�������!8ĳ�+P�¹����]?����J����@���)�rDh��N���D��N������ǿ���|U�'� ^�J��H9ѫP�Cr��K�x{��@�� ^�|m�|;�޳O ����U��'nܒ�΋5h *��X�Q۪����s˫J�2��z�Ƥ���z�F�Ws����#��ׯ�j��ݳ����t	@�.���4���+�����ܓ����E��W;�����"�El?�P���v�\��FjF���~��z�7�Q�G�Y��^SH��$�
�❘�O9�ݚG�x4���6��*���(;�yf�Fʡ5���*����M�rlԘ��yr6�9/\Дnn��9g�*�`�$��z8%t}[�J��
W 7��ϒc�K	�l��9^#�d�)��| 
� &fmO,�R��ybR��}ּ<)�����9`�`��+�X� $<�{�8h�֑��q{Y�	kdٱ3S@�Xq	���!{��P�� 
�r��B���WI���@��!�hAM�D;(#�y�2��'u�i/�^�\��qb��	�ú����-�f]��n�D�t�P�fk�/�@tp7���`�cX�5Z4yR�7���M*��%�����{!���.�v�36P܀N���y���ɯZ�y���@���z�t�M�4��LXCn�>�Y�dQ����҅
.s��I���Bc�+��M 8�W	a��g����ϋ�9Y����ɠ{��˃l��e������V
�����b�~"��^��L��jBM�)f���P�Ͻ	�#*��=51�z�P!}xV���G�R��tI[~l�@M"�ӗ:v_�����iT7?==��Ãz_����z/㩎�� �ӳ��A��:y:J�2��˽��>����٫������r��˫
��j���_E>?ɦ~?l2g�L6Y���z����.��6�O?Mp��7�皭���$SqSX�3v�P�̪����(V1���SW�NZ���d[��s�t�W��{z�!u��z��#���u�N�4n���yUg���8
��]�����6x�l��~��{��=SxY+�Nr��6�{vX	����*������������C$�w�e)9��E(2��2'��b:�t{[���?ޱBݜ57�x�*��d��/���@�~�*�����vWA�v����lͯ�l�P�G7�R����I�&4Ǯ�2����i-
m���H�bœ�u�-M��5O�ț�w{GHQD܃i2�X������*m7Z[��{F��m�׼�:�ͨF'�"��2 �Ȝc�e{���4iU��1��<3i�r'��{�
�}��]+���[p��@MWfH�{jj�j��U(8�o���Dف��U���Hv�cb�P"��3�����L��p�&�Ÿ�:x��W8�条`�{�#k����W0���X�����n��������B�(�k�2C;���H��1A�g�d^��7�#"߸�>y���}�7��WT���1��V
��ϗ�\��؅�X1c�l -� R���е�gy'���uR�f��y�3�_v���'�98�����-x_�dW�i0���X�\��������>�u�L��������+rkx)�o�6tBЫi�MHɢ�q<���Z�d�:�*��$4��2�
�~��˖�g�n�YT�*0�O�>)�x���M~��Y4,L  ��D�2�ڨ���G왤�>�Gq�:�(� zx|��X����uEvo�
5W�7���y1l�I�P�cD!�}���Cެ�fA���5]ω�d��O�qv���8��l�M�w&ߑ��O�v�Eb���۷��g�DNL������}ڸ�<BbU���y1\:�v4���qq��P�B�Ԥ��꾒��f��5�� '�A���w�"�-�BoX�ļ+lV߱Z��%��"^��OHh��en�"�0�LCK+|��W14C�,���<J���G�V�Ɇge&�QC>��0��峵���I���ܤ���V��Œ]����U�����UssS��	�Zуm�.[s���2|����{r��: ���m>}��d�X��bL� Qb��)����@
�a���;�a`�]n����	�y�k��`��Х����'n
6X��P��XT�hU�Nd���n�=�BxҚr��W0�v	/�LY�� �{#$����M�rx�ޟ�|�i�-�L�8���߭��O>m,�ɪ���
���y/�Qc�`���6
�F�1r7��BI��Q��Ы>:����������8�w��
��Xr�'Ǽ�H˾k�һ��W��2gj�&�ڪ~d��`�����G�F"���2ϑH���B�1�oOE�P�z�e�Q)�uǗ��{k"T��*��U�ۚ�5�3��(������B��L��|x���|x-o��{�ػ��))<j>$��0gb_q�5D�^�m�dzh���u���\�۫�u�jaՠ�S�v�'�o����,��-��6)W漨X�)%CR�N%9�����Y|���`U³U�|B^xP�
��|��E�����aT"?M�%zo�z]����ܧ�jmox����9)0� �Ie�Mȓ�8Q�=(眳=�.h��ܕ��ɝ�"%�����>�jl��V�y!�\�Ox�ul�h�U.��Q������8Չ���B#�.
� sF�����5FN��)�<��jL��G�r;�k�ϐ�)��dF�h�Hi.�4�bd��)��a�����f]�"�DM�ƗP��d��ݸH�bo��y,�9�D�A���M`����I�)_�c��v�M�h��F��&�-^�jk�����Y>|� ��{'GP�����K��w?ȋ��e������H���f�nF@�N���Hi�*��`��&�����R@/_�.��Jak4�.���{����S|*2�u�w���)�]aG��G��7���p�U�ȭ`�!�)�k!=��&�S0G㰈uV�u�gD欈�&sA3�nA!Ia[D�դ�RE7��x+�,Nht�\C)�R�.n�Kh�V��W����0z�����͓�=|��rjt��Z�m��h�/W���A�������AFAF�I�j	��
@k��m��.���tV0��vw{��v��*�mU|Պ�tp��!�D�4->u+��v;����=M�hVP̧���u+����"�v��}"�u{)%%<^�-\,>�A����|.�їF���j5���^%�"��5F��^��MuC��y���ea�z B�K:UA�(Q&}_�h����Y��ە��/"�)%�K���:R���,��_OP[�m�](u©t?3H��u�!Q�
+�|C�  �x��|���O�C��i��h~��'����*��L��xVw������=�?���=W|.�TX��r��d���NH`��,��b1����QNt�l������*����J��W�5K��T�5���ם�V-ْ�Y� V�~�>��53�e��	V<�6�I���RM�lh�â	� �x(t��͇�z}�'�y�kJ��r�y����޼�����F���t;��"/��֯�~�e&����y%��$�ɞ�����9�~X?����`Ά��vY���H��q\Mz���#����-�f=��"�WWu��d�u�����-2踫�;��5L�r<�5ROh�+xlG�,�w�>��q1���369W�ٱ�_�@�+����A�H�6�C�Z[k�M<J������:ВET���]����<=k�c�zw�:���i�/����l��Vii��'�xeO���g��X��Y��6��j��b0���'i�ſf���H�C:��Zjh8�P1��|`��B��	��5���,��0�V�W��jVR�ڭH��=)�%(��G�|�`;~~�"����<����]���k��7o�ʮZ:ǧ'yJ�<����,o��^��Ȕ����F��Q|�};��s�Y9��{w��p�����7L`�ռ����VI�7g����[4�,���C&^^ށ:��.�����W����h��ͦb�nf��p|V��r(���J���$1]F��+��4����Ȝ�5a 	�{G�d7N����+�tOv^��y��贄*�?A��qi;�%(S7�![���9Շ�����-�\����+dl��V�����2K�J�Z3�������2��H;�p�2&����U���.�X��3�x4��A4�6P����Ґě���'�L2;r��&@���\�|X��s(]2P7��x1t�Dtۨg�X�]�-x/�YS��k.YJ���-r�h����Pm}�@�( �|��
QA0�[�6�U;CF�~�R��Nn_����%�!�c�:X��`a���\�>>������p^䥹���\X��n�N7�X��|�|�0u�+�2<�Z'��l��2Yh�D��V�v���<d)E�\H��|h9�` &��H���eҺ8_V��.��*��������Q�{�����۪3��e����j��~�F%�4��7r��VT�n�*k�6� �\�s�#,:ؖ7��x��Wm�
��������zN��F�`C���&]£S�;�{ʍp��w�ȝ�m�[�l�.=��*�Ē��0M_1a�ȕ�&2�!q�9��PY���5b���r���}5`�:��o���[ 0��=�$uh C�p��Ъ��*�U�p�}�|u/�|�[�|��0s�w��"y��W�\H� �y�Qu3KS�M��<l�Vgo�� +̓3��/>�ރ�H[��|������ Wur�=�+U�﵊kF��y//��,w�r��^�4�Gl�Eߞ�emW�&�t�n:
���v�A�c��˘gj��-�R�6�/�ǧ��������ԭ��R���<�{f
���W���1�z�jJY���Kp��R��I[U�q�N `g��9�z̊5Q.�$O�t�X��C�h�9��!¤R�֪�����v�&Oݷ_:M��y
�\|�}$�9(~N�[��w����m��[:X�d��~��]6@���̱�8�9%�''�R�B�!���s��%Gbz�%.�أ~b�p��K��v�e0�<�\��C�dpooUF��mL��si�Ä�9���/W���P;�-X�|�lU��Y±��O� � P��Z`�G��q����A�I�R�<m ��*c�dT��7W�b��e��t�?~���+����´� A!xʠG2�3礷��{��$sߧ��Vba��c��� �Q�xr	}-Rh0F�E1��y�XA�i-Tp8ǐ;O�x.Y�>����_��^l�kI/ds�&*/hH���0���]��5�Iуyn�.�e`��(נ͹ZD��� ���3����B:�|0���s�0z��[-�N\�J�kG�>bJ�����i���9(͘=����r���+�A�����,n�p^RT�4L8��I[#1?6����C�;��P���7-��(|o�7o��f'/_�a��fEq���^/(�?ِ�rf��,��cSS�=�amV��,����xD���Y:�7X3�ߴ>w���'	|�Js�A�]�'Пa=�"�L�$�f�#�0�[9a���1�����s��կ��7�j�_�e���W�7.g}��k���HI=�4:2@��"`*M���n�V`T8��@����>k+��}���ʝ�g�1��&�bEQ����|�˩�X]�(67��UkՕ��!^o����^��|N���X*�MΡ8��0<g�$��I���Ir�2a��%��V1߫䎱۞'3�@s
g�vKޱ�^0 ՄU����U�J���8�Ij�H(��z5��eTp:�@���8�$>������z����R,O/BFC��9Ow�E�@��_J�f�����xwtM�T�Z��0�ba�C�}�ôL�8Mj�IV)�{i(�(*m��F���(��)���|p�gWZ�]�K.�zhJa�ڃє���;z��"�
��:/�}^�&�sc�ߍ���(J�@ד�s�nq���'y>~�����<���]�{����a��J���p�z�Xe�X����k4�I���_rbw
����?�J�	"���CUB)(�?4�}v�e�Dm�%�*A/A/�2������L��qr@�@V�sc�͕�i_=Yb�������(q����&ۋ�s�7@r��8����Q�CU��\���F��]�r��VL�N�;j���A�����5�G*��;���^�r�BF����:�N��ᢩm8V�wn��N_�*�,�=9�f�1*3S�����um���|hw� ���k�+�vh��{O�t���$�
������{y��F^�]�� ����+[Ԋ��YA��8����s�7w.��i���j���B��2�cz�o��K�y|(7�廁/�����J�C���=8ٺ�;7�4o�+v{�B`�&Q� ��nO��O���'�5�����$��Z���k��2��2I�y<J�C21@��d�A=`�������ƪp���oc��/�ս�~v��y_��k�i� Jrq6�T�����nS�J	<�aRiL$\�^5/�:�
�|҄J?�h���-u���<�z����C=���賶!����3���n�˥sЙ�| f�S��!`�Փ����g�3;�S7��X�M��'�ا���H� 	O�2�o��ň���MU������u܈N�e(��krt6���+.�(�L�E:JЩ�ޝ��U����J�X,�>���h�v��r��͗�z��ɓ�����y�	�e�)�7l�2nP!� �
�b}{��k���u���up"��zP��_Ƅ��|bn����v5c�lZ~R쩡�'��p��ǣ<>�M��j�Q���Ԁ�U�"tm�7�Jޤ�ަB�3���d������z�y@GL��� ���VOǏ��λk��
[ACn�>3ײ�ǩ<dJw�ɋ�\[�i�<q��h���g��+)j#�վ�OV�vD.$x�0k)�Z����W�}�ޤ�(�<�N��ֹ��d9 �C�9bwW0����ZB������ՠ/C�
6�c,���Ϝ���t�Kr�"����C�>#�
��m0� 0���z_걋�<d"�4��0��ͳ�Y���#�sZU��>	���o�* �!�1����~�1��oQ��w���m}����͞��?�w��M��+Yl�Ӱ�&T?H,�xt_�k�r_r�J��0/�a!����q����L0���6e�څ��p�2aD�	$8���ƽ[���BE)�:n�������t ����H�3��u��������}�C�в��Z3x�j�2v_��ѭ���u��d�c���+����B����ꖒ�XS�.<��/�M�]1�|��Ϟ��u�rhl���CP�`���"3?(���<6k��x����������{9<��cr����%ۻ1�`��-��I\o�p<�zq�ټ1��um	�c��[j�R��]�6y-�~�x�;����`*�RbP��9%��'���4T��=�E1�.ճ��u &B�@�$y7�ʬ�LZ)i
  	�<,�Jz�F�-�}�옹"d��)�*G�l��~��Fn���
�n�a!�6����h��u:zg<$�u?Z,��.�������P{�e[���P֤�a�D�����Yڲ�p$�Z�v�,��9T���$�"�����/��{><˱� $姴���Y+*����.����κI��,��B@�Vw��<��D���Q�����Օ<�����v!_3��N)7(����W6F��5g˧��^�*6��o�	��h�p)x�Xk�q��lF+(�1X��@h�F}�~̳�S�}{�va��*w�X&(�&��UZ�=[H���;��nw���sz�#4���{��~x+7w/��GP��s��x�;J��bg�OYR	�t�,���lp�İג	#M���֋NB��8����+n~Oݑ]^K �!��?Ã�T�f��Ҝ[��F�U���=�[	}��S�k-�=oq��Q��PeV� �J��`��׍\ME�v������~�y`Ӷ���ﶉy��`A�LM�˂|�IWT����-r,:���+VOҍ侒�P(�	+!���BO������V�{��9��e��tI��Bu+D{b�����*I�k`���5�J$m����@�N��:���`��!N\Θ�:HZ�¬�U@�ht��Øi�Ƣl߹
*���¦��% ;!^_��b.UZ��gX:�+���W�S㟍�&�;�<��ō���dk�/�s�M�P���o:��V[qMq�6��#u-#����þӨ.�����d�2�?��+���A���k���w���)�Ī��lڽj�Y���Q���i!��;�O��	Pg��6cX��D��H&Vˉ��E�뷴��0�����59 w�N3��mj:�S� #�T��\MօG �,�c���[|Q�f��v���5�EO�����y=�#+�RE#f�#��d��
��B�%Z<���B1�2�}B!뢳z8�\��|I �I�X��k��^-��Ҁ�Ka�Ni@�"3̖�=�mi܋PV�@@�urc8��/�8��$0΃[��A�2���Kh��WJ�͍Ddkϒ)��-���"�/���+�|dh�<�Զ���č�Q�as��%���>��� x��n�G�7Un�"$s������e���v�������R] X@��fT;�mL�{��h˧
�����A�1�~���P�L�I�%���gs ��u��f$%<��Y��kR������c����v�	��V��*ӌ��"��oX*�J_��MU�r��y����o�wP�Pu�UD*�,*'��zc��Y��ثz� ���e&���{�s������âkPk@��7����&��}� �W��j�Pr�R��� }.{T�tяq�wup��P�R�p��=3��ı70��� ��Q k���c}u�Ѽ��jH�xq'߽}%߿}#�_��\(���u�dVщ^ c�V+%���+H?9w���}q�l�<G��&;X��g?)�k����=&a8
�ߢ4���9Q�L�8ě�-pLJ!˷� m�%�F�p95pc�������PZ܅,C�%�-D���,���l�����^6˕|����
6u�]�I��C����"�:��\���mZLI�eȲ�aX�7ch�L����D��HiJ������D�GV�(��_�D��Շ��du�x���BQ)�;)��߭@a�"���Y�|Voأ��&8�ȡ����!����Q>�(?|��]_�TςzW���8�'q��!����C9b�Y�\R�7��d��g:�k>��l�1㾦��B����)
���is��ݪ&������Q&�v������e���hx	�H��٘�G���������!v�X(TGT���@C����b��ƙIϊ�
ے��A	�=<٭h�m�N�ʥ�g@�\�h������B�`�b�V�񕗖0�]
���?��P�kki�{�e��e��|���a��7�"��� �m�ՑcY��
�������Ga��R,�뵰�A�������d{�5PX�Yxq�� ���7�����\��ݰ��L.0�ٜ}~��}���'��"ǘ><�*�oQcV��\Fm��	��E/V�k^T ��
��|n��T�H�Q�+�1�'x�m6���||x�@��|<��
a%ϟÅ&Õ��1fm����U���z<+_��&9��<c��f�Z�Œ���0�G�p��g����)��8�iS�u{�k������V�k���s}��*���T����GNf���.�X_e��9�Q�⁦Q�E:��8�@�bm�ڥ��gP`m��e�h��^�A�!t���P���B�J�iHK0��,[g螿l�: @#{�b19��������!t��}�2�^��OZ
솗�O�NC�˗/�?�A��/�"o* �W=�kO���*q����ynE�' w���*Y�X���;�W+��˾/a��m�S5*�Q� ��lD"�Y�Iz�t�Ɛm���B.�'ǂ��\��̠K�c����-N����B�.s��󮺤�&�)��F�h8V�|�C~�]����q���ڠ��E��?z/G��
ΐ�^4��HZ�>�K-��7p�0�e\�:D&Z���cY߿$.����t?�5�;W�Wzyұ{8��u��ڝ����Ұ�9\�̽�4j��h�׼�a��Ѫ|��Ӄ��흜*�E���t�yA�����U?���zx�"_��z��=6���p���JS-��gc�,$5\l�:�¢p�U0�۪  ��y��
���#
�2s�ˇ��~��g�r:�ӒfKD������#���Ҡɴ��#��?1��!l"n%����X���RȀ�&Ŕ�欜Y���a��A���B���P���%'윶m����o����7��|8Z`0�1϶'S��#���C�3��@z@3���洜t�躢�����؈C�ŹކX���[Y�َ�)J4�7Y(&H�a@,�2���0�}��O���d3mT���N�j������F��:f�;�r��յx~j��>�h)'�y_�da3��>�V!z�!=(�	ʜ���.�����O��0�vV�4~x��F��P���s���JΙ�X)Q�(��0|9��J��88���{D�q�Ɋ�dt�mO7M\�q���h�lR`�P���yr�3���!HvIP>�b@^��b��Ws�7� \D�]=��N��N��l�}�jDN��/�/�!Q�u���hu�bP"��� 3��f���~�Ǭ����Pͫ�0��l&�</�	�Ix�u��]���
$�!���'�e�_�<D�_ ���K�5��.��p�P��"�Έ�@���",����|`9t)6��C�nY����rm'�o޼�?�����/�ww����?������	^��;/��|P�C&�V������VIc��|P�r���g��)}�	Ȫ�d�
 �͙Ǔ��|\à!U+|2���;���0��E]h�Y/Rޏ�n�cH���-��b�9 d$%
Q&�r�i�|�ذ~~�<�\���s��w�W�r��*t4��
�>}� �@Aca�7�"la���zL��.-���!��	���Na�,\����qHC�Qy�=_�~���4wE����,?* e�F�d�P޽zP��v(#�${⮓xn���]<�j���b4�b!_�=:�O��ۯGy����g�ҹZ�Hu���a��>��	� !�烑��;�p�Op>Т�b���/a�Ұ��v/�Z�Ǫ��A����u�<~�M���/깰�cN��cR?�O���I��9i$�gv� ��Q��������@
�|DHv�^*������3b��C���Ӏ�f1���Ɓ��*'�"(�p˶(���CH!����Vs���An�B8��dV���~>AF�>��`d}'�7�Q�t'es?��Vfް5��M�z���C0���R��>�4�U~f�% ��M��u~�֍�^�����\5�)(J ;��L[�bU6�\���*]�[HJ�Yؤ�U�|4
x��%�H�#|<?�1��Y�Bi���2�ވ���{�4 �r����9dw��il�ɲx�|ٳ���ޣɝ�.w���P��$���Gu2�Rcg=-=��	�o_݅���7x��g�����Y:y$aP&�R�Tb�q=[��s�"=�\�ZP >�@�����=uV/��$ϖ�#�<�U�����li�)�PW��h!�\�(��������9����Y��Jm�J�h�b&��3���p~%r�1���g)�N���SG=�)Ha$��9���^#A_[p�����p{s#���|����� ����ʰ�x�bOX���%r^���'�Y��p ���%����0��ݠ�V��Ydr������L�Z��,�³���
����Y�����nI��:����`�=���=��Ą���W��O$25w�fb�C��	�e�X��+� -E���YF��g-M��Z-��E��ۗ*�Χ�~��\Ee�����Zu��ol�QB@�G��L�{�Y�&hl.�<$iU=P��W.�ՆH�P(����31+�u�d
��n�Ы�B���H��f��LP+t�Jf-�7�.�i2 0���r���uO��{P�
��̐���v$KyRpͿ��C���u>�T�U�T�/�V��s	1Y�R�SI�gX��'�«������N�D^�X���Gkm֣3q�:�hɛ���K�����H����Y�WWk�=3^'�e�:(R��g�p�*� PGki��L6�s�H�e�8�w�}�o^U(Y�ܶ�xs��Cn���!����
kk_���o<� ,Cf>bN��rH�F~@�(a�Қ�ðwL�}�+(C&`72
��� qn	���y  ��6&�l��l \��$x�z�* �{,d��@�:A�����ɼZ��ʓ%8�7��袁���Y�y�� !�0����#�_Wi��t��0'(�S��֔ZT�v����y�n9%ir%�U�#��ɪV��)�����E��zU�������y�g��$��m`�}�\��2DAi1 �N
�,݄���eqV���Mj|l���=?�@�}RJޟs�
���7,��fF�q:���.��s5�ԇ�v�h��ܓ+�S<�//� ,�N1�]Vު|�\�Vp�z�]5^���G�X���s��y�
��?Ê�klU�).��B���Jk�枨N���^�.sCuC߹.\���ƿ�����;_���?{da��t[�?���&߽}#��
�`�A���g�֑���I�Kq/U��r���\[C�2Ŧ� �Q;���#̶�c0���/��z6���{�����6���%�M��m��#ݑ���fq@=�(-\���L,i^O���g9T�d���r��0����3+JK���*u��"mL)b�|T��Gs��l��K���=Q��Ą�{L�9�nqy���x�z�Ȍn��~��|�Jq���A���Vk�w�G�UX1$!a��Һ�2t-�l3�S	��ݘwO���p����6t�� yY3Co�T|�fP̳�8Z��4�&_�61�~=���Q�>� 
q}���B�W��dZ���@=(le���@���=ͭ��zGRP}[+�¶6م�	�!��q�M�(8IL;����/A�ˊ���y3pr=��DyƐ�yDA�ӡ��I��1�UY8WWB?I��C����`�!�~�t���o����&���]F�$��;x� ������÷Xc�d�,o��f�:
�O����<��ǫw6@8T�6�6ϣ��g�g�ŉ>�0��uM����Z��uٸ����0"&��37��p��l]�U7`?!���Q�ӑ�m��'.�]�7i�6�9�t	���'b �s��r,)��R�*���fF3�����5����G�I���lF+���sj�UͨL����Y���m���C�>�?�H��#�,h��X;Bf��pϭ^o�	��Ӂi�ևj�N�g�v�����.R�S7v�o�eɴo�5�N��ҟG���h���s�;t�rF�t�^4���")%�������&]Wz49�zj�޽��x.�j��l:K+X}�U�}w�Rn�y]�۪�=���d���?�đ�5p    IEND�B`�PK   (}OX�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   (}OX����;       jsons/user_defined.json�Xko�6�+�?-`j|?�m��-X�u�����D�#�z4(���]Ʊ�X~E-0�Թ�G�\^����óa[��c���p4��:/����R�.��g�|]�\����ś�����L�b��
�x�ybj_�f	���3�#�!/�E��ymR�`���dJ�Xo�p[V_ ��]�,�fx3zLv��Yf�uXG���SIu�9G>p�x�� �D�f�3�O�-DX��y��ó��p9���?� U�����a�g�ت��u's��Ფ�V��0*�1�q�h��׿��� ��Z��ܺ�Yߕi~�΅�΅@�~0�͠��<Q�J��� �E{?����~�s�jH¥� �[�ˇx�'XH��_/Uv_~�n'6\T�"TM���'��)�RZ��"����x����1��2��f����|xW����:�(�y��X�kU���UTL$;R�/�-�����B���V�M}y�b��/��VuJ��"�E�)��1a�ijCȬuOZ�苲E�aeOH��6\������p8�譿[
�Wϯ.������ﮮ���-��	�V޺Y�UX�'�h�W��\���!�V9��}�=��R��
�3{�rK�@�3���G��e�2��ά,��R1�<�3�qx�Id��PU��B ұ�z� mϪBG�"�h�K�[Gk�b˕&��S#Byb�aGJ��������T�c�[��k��v����<	~6�c/>ہ�J����l��w�Q���&��Ł��)=	����c��T·��]7o�3�2�����s��ɔ��`a��C�@F��v!uVƻ�G�[0+�1g�45�aK��rL�r�Jm��{���	(@"������5�2G0�'�mn�`-�Ns�Ds(�/7���B1J�HȄr��ao���R�"وH��ʎH��ހS �Xj����8:� ���]GKa�5#B�%�޵3�%L+nFh���\��\&мJ:��1T	�\ W�$
+՛} \�k����������������t�	oQaɁ!õ��!�u�:s)@��P���Pnp%�߯D�u���'�-�u� �4��Q��SO�:t�9�#�?����:t���t�8�Z��5�_�0m�;�6MYl��Ł=�c����F��Z�Q��1[v2g�?���� K}���`дs�ga]��{�b9ɺ���P.�޹e	Ø�/ڔ��'3"����v����ʶy���|f_��7��#a����dv�!�Wy�?J�b��}
r��O�J0��I.f#:�x;�?>��c0^u����d@q�i���g��\2$�bi�����ۿPK   (}OX����  Ӑ             ��    cirkitFile.jsonPK   (}OX��g  n  /           ���  images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.pngPK   (}OXhT���� ċ /           ���%  images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.pngPK   (}OX�Ɍ�� �� /           ��u� images/53a6c856-3ba7-48d9-b0a2-5ca2401e7b62.pngPK   (}OXإl˨6 �= /           ���� images/734bc482-36f4-48b6-9076-7f88fee16b3e.pngPK   (}OX�1.:�  )  /           ��� images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK   (}OX��n�% �, /           ���$ images/c1d4a215-2c3d-48ac-b15d-f6239b4c4b94.pngPK   (}OX5r��W
 zX
 /           ��GJ images/cccdd3b5-475e-4e4b-8694-ce23b104edc1.pngPK   (}OX�GDU7� �� /           ��*� images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK   (}OX����;               ����" jsons/user_defined.jsonPK    
 
 j  �"   