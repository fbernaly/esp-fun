PK   NM�X9g�s>
   s     cirkitFile.json�][o�:�+�W��]dv�p�(p�!J�a];P�^��_Rv�86����Ecr��83����u��[ΫU��]�خ������v���S2���_�?v��>��~��o.�V�VK��禦�˝�u.�ayY76��m��ֵl��f7���E)��M�sW�\hKsM�K�JV5�R[ͩ��&g�f^4���4'�F��H&(�UD4��D�&G�����\������k�� 8�0��M`x��F��"�N�x�H�S�q=E�^aD��L�0�~l�s�Z�:dr�~c�dBf�<��F����\�Ʌ�ua�is�&��A�Z.'���pI��$\T.E.:	sj�s[
�A/M_��4��<}��(A���1��b{�;l�Y����d��s�I��$\�).���rr��)����S��L�E%�R$ᢓp1iP��i�K�����/M`��4��k��t_��f��_�&'ٗ�s�󇅭\=�)h���/qn�����$W�Z/�Ҽ�D�[Q6�(�}p;�1�q����J��Z��Fr��YZ!L=ga �h-�I�*~��T��棈���]Vpju^�rQ�*׆U9���(.
;�1�eQ���2o�ƃ[T$7ΐ�.I�K�+�7��8�P��eI�R,�I��:�Թ���K�U�xɴ�Æ��V�&���)�]�D�r>ʢ�Qc�5��8�Y�0�)J4
eG#kKX ĉ���<"Sfte �
#:�2T�V1ѥ��J�k�ƇQ6���LJV�&�2��h@QGli��S�Em���F�bt�"!�9����l&�'nx�󱿢*��Мԅ(H)��qq���(�@�#�WB����q14V�<�D�(����?i4�E��G�M��;�R�6��(���c$�������~�����#�_ C�F�EdC��?̉B�5�9��G}5�Q�ab
t�j�=��;�i���s��m��z%��g~���t�rT���*����ґ�V�plT@{��G�P�9[o6@��x`��G5�ȁ�Q.q�W {��� {
�� {�� {&��أ	��
�؃
����p�v�:����q.p~����
.a��*u�@�Γ�B�R%��L%#.Up�Y�^-��_&��F�x��'�h���vN������n� ����Db��%U
0��$��e��z�<��H��N�v����uP���Y�be���rT��\���B�Ы(	p��8��]�Kt䕠�6���dF
`�I�����7N�%.k]�(`��L�� V�^�<E&����\L_#�lf��T�b^>u���x��*�`/W�5H�bc�W-G"��%>/�/^&P{�r���Sn�e�n�mc!���dC����w��#m`^��slx�w���� �r|�/���64������k�X`��}p4C݈���$�]��.�χm_=�Q�{jk��bd�'RŁ������:؇,�p�e�=v�1�cg�_��,�+cz���Hz��/��Io��?%�|�7�P���bJ����W�#b	C]c��${!l�W<�ǐX �1���4	օ:hx��C 0{� ���4�ȇe�pSh��CCW�U�Pv5h�a�9Ok+��F��e����E�6��x@����a�繑����z�W���O�-l�S�`�������Gvh��Ml���������i�y�9[�+_��e��/��~��x���ǿ���Ͼ��V��[�xx�v���×��2���qE�0᧘Hi���1�sn|�Kά�>�M)�J�/E�f��RjDS1J��^i����R&��-�]VkF�3�V]�ص�Y�~�����nc�-��TN���>�{��~�����7l~^Z�2!H�OLi�d�}���A����C�T���q��)�Cv�т��b�r���*�I�v��pUS^�6�����W]���*�V ?���[??=�9Yh6����&���`85Tȉ"b��7��i�:�4��o[��(�#�-���+փH�M��5#�Uh&�c)4�z�
�7�y33��hnd�S�xM��v�}*�,��ӂ?S�n�����lJ��|Á{rJ<K���Io�VC;�V������z)2�&Ll���q�6B�w�W�[�#FHϑz7)v�}gL�3����<5?B�Z=-���W��� 3����Cg��p���خ�{��ڏ�ǂ���a t,�a������ޡԱս�������o��˿��
���,�T�e7���g�d��������zh:�z��e}���Xu�ˇ��y��H��ê]��m?��>�Ͳ���lއ�}�.?>�Oon�߻3h�2}�����y����,��l{1]��k�Kԛ^�D���쇇�.���7�f&�Db��� ��u����;�Ŕ_ΘI���|`��eɎķ ��ud��8H�T:��ԱL%�I ��,���N���z�K�Bc��ah��E#)4d:h��АI�A@� �t�f��z��	L�赆F(������ۻ��_�<���q�v�d��>��ݧ���Zُ�PK   NM�Xh��3�  ��  /   images/3af811fb-ac37-4701-87db-865e720a6976.jpg��w8\m8"�A�w�G�;��(ѻy!1Z��&�w��ޣ���(3���������>s�r��)����9�_���k�k��� �W� �0Utq 45�  1���@���p�r�?W^����S��w?IL����=�ˀ� rR222Rr���m�;��w))((���PѲ2=|������X�����3�S~a�'bl\����2��b�D���oS߾M�����������&�'�$!�����{��	��������)��;���D$$ķHHIo�"P�4�-R���dtz��9��~L̻�����A�-a���#�
^>~AI)iY9�/��5^ij������;8:9������G|����5���=%5�G:$���������WMm]}CcS���޾������ٹ��ť�ͭ�ݽ��g爋˫k$�@B����[�Hn�����8�_"�-���d��z���8�~�M�<1�����>���{���[r���_H�A��Ч�_��/@���.	Aa$4 ��:X��3
��ɜ�1�ڱ|����6�<x+4�L�5|̭��x)��M��`%�������Xc�oӋ�� 6�w��%��&Ճ&����\��c����ȸ���h�t��vn:�uVf1kL{���eHQ/��WfM�s�g8��
��݂S�y<�;~(���J�d�j ��F���habՏ�t�B����H}���1�P��k�U�n���h�q�6���\�܋"z{Z(����	��cU�q�9/��_��6�0e�+��3J�(1����?x�p3�L�A���}'��-�'����}�`���w��յ�{��q�Q�Te/�溳TqH���%,0Ǎgڋ�RX>�8?e���� ����2�Y��L.I�1�Wy� ?@.�
69g`�A���/~O��/`�Vy1���T�W�Xb�8�u�е!����� N�@����*�˘s���*��������l�$��
�i��\�[�)�Q?h��#}e���Ĕ���-`;z��i����M�4�����"ɚ�m6p<֚T�.R�'��?L�L���(ŁN&�:Z�������O~w|+��T�ɴ�V��Y��(���� ]�z�!EKZ� ��֓�J�C�J<��>Ǳ�jJ襗V��!x�о�jԀ9#�>_�����F�P�'�LB�c\-�.P�:p�`3Tpw�l18�SD|��'AF�8Y�E�#Wņ3}���_��4x�hu����Y*�����A��B�p�X��|H�5�խ�!�"˧V���6I|���EQX�v�O���q��П!+�<��Qu�a�Tq�q��Ҷ`��N��a�3�3�r &�ߡ��� �d?�CJ�<e6�����4�J���cE��7�۠.#pH��7�����0 C�}��_�?�0��p"m��W�w�0ֿ�!V�i���+ΚS 	��ihQ�f�������\�T�t�0�m}������ַ�%re$^&L�//EBnᗭ�G�F7S��\�3��3��
�C�}�_��:��㲀ɡ���J]Ls�`��:��	Z#�*�D���S�$wt{�_�w�P������*c��b&c���[���#�r�'˼�����??x:0#)���4`��B�6�o��r$�`!Z	��V$p����j�����?#�n���T�)�ĥ�Qৠ���j�K��Ɔcܗ���K��Sj��3�AK�e7����<%�������A?�,xN��i��6*��u���=�<_�-�upP�-� �w���B'�M���)��5�e�.��N�{�
[���FO�z��4�9�z���Z�����>?��3f�7 �S��'�F�|�;�Lk�3�M�%{���`��7���eX�}M�2����J.��
7�������8����p�dV�m������5Vh�5��h*F�&}��yT^*�n���i��S'#�v��Bi�Y�ktx](!:��P
ɨo3�s!Σ �\��Q��$���cI� 6�뙠\H�l�N)Fe��<~Q�+��$���O-��NֳN��DD�E�<�6�#;0��r,�D�P���劭��^G�\��=ͽ|���� ӵx��S�<�2�Qj��JCf�U#��D٦.����$��q�k��.��b�$2^�d�䮿��<���8�4pwm�=C��S��<��=���R�	D*�0���W�x I��Ң��T��?h���+�Ge�-�`s���q̕r���'�~%aO1�Qg7}�$�5�3Ƨ_�J���\���f���7a�z�h�5���5��Fc��$�ZQ�\>�*]�*��օ��X;�� ��-�F"Q���}��uS���g6R�\"F���ob�n7�@�F��8d��+C�@���ҟ�rĎyY��e�h�d�Ι���}��-�^�Ͷ��	�⺠�6P�k��b��v��Iɺ�=dԐN�i��/�
�D3��T��y�n��rԲս�����CZ��q���X솅��(��c�7�&�^���ƙ���$�p���1]Qי�L}���P��㻕�إ���[�H��G�zU�~]�_�c�f�75����6��N�k4����9�����R�v�ܹҒ�}��r��^e�Y= ]~����i��y5�]�f�Jc8TVB��A����K��>ݛh�{�
9����zi��M6g��w�N�d����`*x�ˌ׷��A� ���.}��`���/S�8t�()EyY��;�-����μ�L���j�1a64U�z�@e���Ǌ%P�{��E�IQ@6�?���I�k&�j�<��Ӂn��i��=��Um��Ym���r�ޘ�۾&W��� ���Zb�)�\G�x�T�q/�FT�q�Z���fs2vp����V�u����0E��Z/��Ѐ��[�$8�N!�"����&Ė��?V�� � �����M��oJ;�
�]�S.��G��"ٛ�*������OM�JW��"��LWL5��;���c&p��¹��U�v(�kם�m�_<������>�y?�Ɋ
�X���抒��BeL_d}�p�wl��\u�ǧ�����*���[:��@��y�G��Y&.�J|F	y�R���s.�c�!�8���{�!�LyoT�����7�K�_�gR�mWKUO��L�~���W@42?��S��İS�͵���:#����򄱧?���'RÓ�S$����u8g���^V�Sۤ&D��|/�N�ΆnuU��4l��ȫ�|�AQ��ܥ��q�/�x�y�M���ng�ԨވO�//N]Gz,�0�C�"#}wB�qa�?�$�+��G�`U�����S�?{y�>A\�2l��Ghj�~==��.�I��#n��l�p����l��]i̝TJS��A<@�έ�0�ʐ{��ˠ[.O=��{rDz�M�%��$���B���Xᲆ�y�n[�K3��R�o��ԣc����w=��?���5����.���`8���M��jwT$�:(6��π!��د��x ��`���b P��o<ܷ����Q�K	#$i�N���=}�X�������[�����qӹ��D��N���X�|vn�X��6Z��1���|��-Yt�'�!Lh���%���(&�/7&�[�!�N{ |l��ơ���y!�a �օ���;R��eh\��=Љ�����=���v���X�����~t�P�Br\%b�s{J�&u���&�cH5�������K�}��Ŏ��0�
���h�}J��aL-@~.�X�b!�W�]L7��U�vX�vSk{�5�S��g:N̮�ʾٛ.��.2 ��p?V�OAܨ�s�ɤ��$^q�"t_���y�y�d����>���m#��%�!������G.C��)l�D�ќ�l�	{/M���EڤS��-5H���נ�#%�F$�c�k��U�C��Վ�Ntc���{P�%N�6�����}�ٹ�r�;�"�x�S���شoJ�4߯�a�*g�@���x��{71���C��ջ�C6c��;j>u/@Z�-F�^(h�ƴcL7�|}�p��K�,����/37:f*+�G����Y�q:�fVG
1C��g�ŌD���-l�J����*i[���E��Y2+�N�A��v�׾����zi5�κ�S���(G߅���H��k�o��I�
�Lzx�w:�@��ݸ�c���>d;k��(5h,b���ky�Mt����B򂉓Xױ���fk�l�����)�	ZcH_�K��J5�^�q�c�4�6��ot^4ף+k�<�����~�M>Q��.�5�@��w�|PN��k�"Z��G[`[6ځ���5�,z��cQ^�݂?���6A̅S�4A���Guj�4w�2RǞm���X�x;ѥe��<��=S����d��� ��+�"��v�OK�d��)����q�X݋+��}w�������[UB��U�M�9�竐*[«����h<�v�Ae�;��ǣ�?��o�<��w��)��ܥA�Op,����?:l�eᰥ�HHL_��Z�s�����z*!i�J75$��`ݣ�r�����<��w�6�2�En~Շ}�(P!m����e��ce�p����������6 L�-a�Lm9�M���O�P;,��9OS~�p_����k�u�d�kmS�~W~����wϸm��|]���4��f��%�`pV�l\<B�W�M�>tZ��K���nOM�	�*fDw<sE���m����;�c�ɺ�Td~Q���(8F��x�I��=�?���{R�ڷ��`s~�;j"������_Mߺ����]���|��Z�PM�3GJ�@�G������7&8Z�Ա�ʙ�?��B��0�ޯ������n0|�����hz�~�0����%�Z��ӱ�|辶���p<`gK0Yb@�2~����[g��z���jL?��z
|�8BM�,BsTr
��yE��g`|�}j3�pWF������F)a]��W{��C�J����~�+[�z��^hu}���n�^� "(+a�]^\��4�v_�Q"��e�U*����;Џk��A�$&ɲ!#'��J�l�:Y�.�;?M���̋l����Hoe��VDߛ�3��_n��9�A&sm�؛���ϭU��8�K*=0���71}I:��]�7a|�܍Ǣ��z��b4g��� ��dȘ)��~V���֨���U"]�c�;�n/D��n�ּ>Dƣ�=��gd~ٰ�]m����9,����fy�q�'s�s������m11o�1�ԄV"LtERF�b�R"%��G$�Z�{Jgl6U!�/��+~x�|s�Vj�/�?���R�FRU�
�j��$p �s�'��yF�׮<cǋn��h��"�����)W�$��Aǻ��8?��&�*���h
uc�1��{Bݕ�P#>L�K�P�u����&�}W�O稂:��F�3<��ؕ����>S���h��v�r]VyU����(�$���ҽF�4g�h��a���u%�ή��L���?s�լw=�k�4"W�M�ɧT���m5��e�=.-�*�]�������zVwv��|_Q�N���R���[������&w�W���8i��i�ﾱ��rĵB��a6|�fK��;��.%�Uot�T�~f�j8�����q*��H��5���\�*>%6}�j�9���1�E�J[���{a��SΦڶ�_���|*\��I!��Xrǥ�+�b4��]VO����"d/�@m�X�7��[̗0eE<�˖�S�1"t�L�\��qD�����$�8��7k5��:�uE�ˣ���� �����)$h+3la`�f6�r/�����u�:7{�]��;���6��v�r����vl$x]�<�0>.���}D�~��5Y�ޗ�[m5y�`wX�=�cY��3F9�o�+�^V�^�����ګ���b#\�{��W�^�Ht���$J�H��qH�&oTn5�ؠ��U~�7��u�t ��=V���u�Qc�����'�OA���Q�o:Pw3	�<��� � .O�.�JI��A���6��ۻ����6��AU�.,A�R�۱�V.a��p?�:�c'>E���OX��m�wh91qL�`�V�I�_]`�xQ�Y��c�^�׊F����ߵ�P`c��u4�L��"�W����ī_��q�`���H���W�׭]�������	�t�h��9���-�9>��z�W����V�U��^�������Y�Ks�g�>�	��z�)�D�6�SC��t��"�T�Բ
n2ݯ,1]6��<��������oDZx~|�N$�1̪m)���ڶ>�3[F� �D�u=qmA�9��2�8|�<i�l�k�<�K��OU}2����;&kձ�����}��(��K�WVi��H���.>�t�8�7]$^��[>�M����*���{V%�(�
R��D]��k6��m�ԫ����k��R���?k�0�}�ysۥ�B��%�����*R�@>��"B����B�^a��*OJg�|���?wK����JN�7檪VQwΏx�;������'n��OS4N	���\-�����(�'D֝Ҙ��5K�+��~E�z5��BѰ�n�^�������r3�T���XS���9|��QN��������祈���e�'7O��������L�")�?���:�F�
�Tg��z=Iwf�]��n���V���g��qt����&lu��5M���XA%��_���{4h���b�:�ồ�Y�2�a�y�Ҫ��u�t8Ϝ�f������T��2��t��Q�5
a��K�!Y�aF-mݖU�;|Jm�ъ�lL�WKWE��.�� T�I:���[!2�����l�ξ�Պ����I�vDwj<�L�>[>4�����z�e.�[쀊7r�!�����F�ڳ
<��*���T?��>�0g��*���(�Ҹ֋R}Gn;3��8,�L���O��RE��%Z�V�v�j� 9RXs��F�Oy!o�R���
�ߎ�W/���K ��'�_����"�K����u�S|3�ᵀ���ȑ��}HK�b�do� �����Tc�i��ɲn�RS;��p��̐j����*Z��)E��6��4�-V��<��3�3�P�-Tm�t�-�E�X�j��=��ӟ�D�,����p�[�=��1��c�Q鞫��r�R�"�f�>���[!�)��))j��
��{i82����5��\�<��2�^h�}�U��xH&u�U��nb���6�Ly�@cZ�WX!bb߈s�i�.�d��T���3Vp���eŰ������ec��:�(t�}A��4k�y�j�x]��nG�7ҏ�3ǸZ���ʉ��<w�]Qi>������G�/�P�S���qs�����KUW�X2_ҩS,-⵨oYbi��@��qj"�*�0�R��*p>�&�<��>-�20����3i�ז��B�>�R�����YQμ�a��w�x������l�P�,$�a9�񩾚�c�k��
'����؃��-��7������%
3�������,�?�}����z�\mB���k	EJ�F}R������3C����3K=�.\���4�`�GQ������5ya�dq�2~��Qyj���9)���d�������K:�+<���e�s��^шE����/�Ҁh�>��:�)�<?1϶�|��b�����d�Z�>������Q20�q�3KU-�BT�[�g���@�9=8������Q~�)wr�	T~��VA`�5�u����X�<���xq3s�Ԥ�;r6�g��P��+��� 2񀊳'x@��v���Y�����P��{j�bg��vq����u�3�o5�a�[��߁䗤����k}��R�CS縫5��c��a�9�[%�+ػ/�1�2�_�Yt1'�8��n~/�����׆�<��m��%��'��Q)��cq�>g���ix���+�Zr��>jk��ay��'3�#2������#ޤ� �h����#�{��#�`s�|�?V������>�TS�k���{�16_|[��o�ij�÷`�c+������d���MD;	|-�6c��}!��x���{IJx@�FI����8-����B2L�3>U.�Z8�8����8�kvE�a<SY�&�"}��i	&: ����m��U�L�D��� PEz���k�?�J.C�-�N�[�,g�'���1��M�8E� %8������+��e����tᠮ6��'�cZ~���N(�7uY�&b]#ji�!���k'�D�wӣ#ǌ�6.Z�*��;z�Y�O�:j�T��Tz��Ny(�mR�ݛ��~Q&J!a>\�L/	Yf��07�����[6P�:��.�X�yH�.`�m/�����L^�܉���=C���� n͵Kɦ�_�sc�3��j<�o�,Cx�U6�s�f �O6�+�s����N�0D?�������P���Mh������ōeM�\\Ǟ_���PXǷ���@rc=3����\�c�ݰ7��Io���F:�_Id���n�vyER�6֢K�0���w:⮢����گ�.���3�B�>�D�(�3���[�����E�*t�>��8�l�2��soQu�e�[���]�Ë@��tC�y���^���1��%��
0��n9F�B�4߮,�}-y7�7x�$q�S�h�>-eB�T!�'e�^r�L�����y~�S�iu�\�rP�������_��a9P@�ڍ7L&8p��c&T7���b��<���3$��JC�����;�Cc�u����M�.A�b�j�E~Q��V�sě_!mtƩ'�]�Q���l{�rӵ2�՚��o�ypc���3$rW2e*��w��#mk�
���yf��@�N�dì/V��0p`5)����>Dmt�޽yŹO��mq&b������V���'�{dt�Ƈ�͜aXP������Q�z8���?K��L6;���	T��`��m��e��S� ���#�ԩ)�ax��I6T���/�yӿ��ְ�"#����S��&]z�y�p�]�sj�uNΰ�+#��B�NA��W'�c �u�֣��J0?�P¯Mϊ=쒏��ۧ��ӱ�;7s5���>�L �����FBɺ��x�t~�{	zl��q�{�xm@��_�U�{v�l��֢:4�챶��٪�J[��.�|�`�}9��oR��3J-5 =˝�QRKs-��(z=-~@��+g"5]ϞĜ�~D���H�}�L��]S��j���ՌLyO�� ���6Ls���f!� 3�q��CTD�~�L`\ksP/&A,�K��0��?V��rw�qL�vxSWU�_ry����8J�]��١�]!e�$�;���r���)�7'�x�޻����SO��>��)�9o5(�u�
2��6lb����Z7�f��v�����M/��_@xU�A��*Y>Ɵ\w�Y	u������܋H�V[�Vx���E���$���k�-_�[�L��e����4��R7 *��F�x^�5z��Ř�7.���(<��� ���E�-j�a������<�������2Q�U��^�%,/�ĵ9�h�λM��x���!'�Z��H��դ�o�/�4���s��0}պ����'!N�s�}06�Z`��PK��&+ %����RV�6������}�f����mxj%�z�%�h٦���)g"���(�ڏO8>�#l[�*�� ϝ�p)�>��J�YA�n%Y�=T����R�+�%&X�oXk�w�[�ʖr.�z*
��@��?O'�bօ���UM9�W��ف����!G,N�u�7��U�ȀX]�ֵ�о���C��kP�4D�"�l�'Cw�횣����7��x�s�\���u��;R�Mw1(�A�$;"���ςɦ@ƕ��ǵ�U���r�}����S�9�H�Xd��B�B����[�}��H�D�iv��5�?�7�,V�4JA��~�X�*rץ� n/ms��'	Ff2�q�N����H�^: ܯH���$�EȩD����jJݫ�8�j-��}���s�ݑF���'�l��&Wv�h�g'?%���+��Kl	��18��0�D��=t�g�M-t��[�]��퀮-��'	/�&Sĕ����O�W�$���!��l�t���"�?#���;����ZS9b��l��R40Ջ���N���aKt0%�dF_:�'�Я�9�'�uo�R���S��siN|����h�[t.��%�@Y��L�1�a����z���f<���-�	�	[�4R2�}{ٯ�kn�ۢ YcZ�~3���(�-�Ύf�����Y���~��OS�v��]�a����̑�
U��1�\�4j˵�S�Ce�3���8����#x� �s��Ⱦ��.�D������Bb�2�*���N)Bߟ��GK˘��-�;��춁z�bo�Ņ��@��K�SM���]��Z�YO�^6:����<�R����#	����-�x��[G^B	����ִs �ћLq�R�QMQ�R=9�C"��,�~���M�4��.���Yi�����lI��6r��3j��=zg�T��Ȑ�R���Y?��<��C�a���	U״�4n2�k-hSO���49�e���?1KxA-���Q^l�̇��}�?��ؒ^I��A���{yc�*WG�)(�Q��xԧ�mw�g����u���S|k�{��D�����u��=�LR�g=#��H�aq���َ?���p�;��n%�=�����E���3sw>c��<���9�!`���9��KZ+]������W��n_(�l�2=��������;�D�r���"g1�!Y^ۋ^ѐ*C?k	+�_���!
	��9��	�cۺ�S?qJ���*�XY���1�T�$�bϹ�L����e�h i_CX��Q���S��!��,,`�q���*��|��L�?�z��W���|�q���FIO�Y,��@
,����M=������k���(I��p�݇��C��.1� c��JGQ0�_��<y`\Sh�à�`�Z�tF�z�X�w����Us�睽�::|l�����qI�S䷾ji������[�&-^/W	#Xc�>���e�b�b4F��ݶ!s�m�-p<��c�=�7c#�N����NZ@�,L�Q�����8A/�޽��FR1J��P_%�(u�P�D�"��i	� 5�8��,7�D�(�4jg�r^C� �5���༈"�ƴ��dIE�&���Z.�|�hu�����j��e�t|kDQ�c��5T��p'�q��g�Y�UҎv�ϣU��e�*}�c�-�3��6���ь(g�L���R�^Ɏ����>��#��� �ҽ��x`�D��D����jtQ��fjF��u����4]�۝B�ہ�R�*]ʬA�^����Д2+�$t:��b<K�B��2v4�$f�8��l.�2�f7���=\J	��=o��܋�%)�
*��T�Ѻ���T�/^��p���X��^�� ��4�z/�����b�G��|�,���a��r6n0�'F�_�I��t���:w4(�0�Y7H��܃PSY������P�5(�f��g���} R͏x(*���h* ��0����|��)��r��4����G�GcglA~�����m�C���l�t;���#p��9ɶ�Y����ӌ���0��W'/�x
%>��>�RK�KK��*?B��eFK�Ua/���"�X���c�Y���G�|ec4���ٲȣ %��v�h�e� �6����%�� ����A�i�]�X^��Vym��6���]�N{�X�e�h�k�
�D&�9? �\>/s-�nm�q|��r��O�TO �~7���I#�Z�|a����o.���=yF�׆i/��_��["�����߽�u���-��V���}/9�rK���<�o��(3v),�ΐP�pQq|̳mX�Tә->����%R��h�,+�Zc�"����Rel�}Ҹ�&�6
��q��L<@���O��mx�8����5��W����Yk�_&�\_�܆���}��A���6�O��792g,L���p͕Ǔ��2��R����n� ��;#+�ꘊl\P��w��p�y��^*3��4U�Y���8<�j2Tn�v��	C�T,q)�����:ؽ����8/^�>��KBa�$vJ5S+'�yU�~RƘ��VN���rj08�1��<�W��%�I���b�թ7l��k�vRQ��˷|�NpDȆ���\���LE�SLF�4>�G��zkC��Uu|�PA�8��̑C}u���@7��7d!{�'�yf}�ɐ���d7���d[�����,n���ư߁�#?n��V
a�ݜ��d7]rD��=�:灺�P�N`�<�w����p���W�q��.���>�!�pwx�=*�Agg��J^��Ŀ7Y�_�@���.p��9�ڣ��E����]}���������1��$)&�x!����:����~��{W~�~�!ۊ��N�
�.hCm4��&[G&��#�*2���P]Vd��~8X؟��0JP��\ɵ��)�?;���e����Z�[���v�ӸQcc��Jn�t�[n6����5z}<�������r�)�b�{;4��Ɠ9P����0C9�)-0giP��[d�f��h+_�&o.�=�[FKI|��+q�vO�c�]�\���L0���ǜ�pW< �dY�V�g���qV�{�
F�a���(��X@��u�����f����ˆ6ް���s7�S�T���m x��WNwèo� ��^�p>�=��g���ƠY��ÿ��O!��Ec�#��3f{�X�2�ʦد�pDX�t��?��gH0�J�Q��/`��(o�&�����?7�}BӊNg_^�~���=�$2T6��;�lo��6�D-F ��X�jVב�#�@=L�FP����F������(��&�+�^�����xwoZ�p�H�>��i��/��<D��s�B�4��^�!RZlo�j9��N��A��W��+�I�&r�/����_��,�J��T�զ�F�;� /Q����Z�@j���3K�=!�B]�>�d�GJ�/V��ۆe!ϔ�=�����P�3p����3��qO�!��;�˜m�k�2O��\g��[�L�$�v�=G�-6l�C*W:0<枋G�Ւ�u"�����UḔ;�u���-�C��P������>8]Jm*�E�_/YGU[۔�v�ъaO�k���j�,'�����s
�Y�rC:��A>���:���V����Ħܡu���^�\���Fo
Vm?�m����3���C����S�)B�O��rW=0��&b�x����Q��nj�4�9��t�N�
�Hx����:.*{��?�~�\�� c�Xbٗ�q�J���zū���l�-Җ8���Y�#=�+F�o��v�y��M�}�Z�����_�鷾�T]�r	�6�z�I~���g��^�n��nm�,zS�y�������\�M�6|�l����x+��
޻(�)&g��W���ɼ�3��\ȵ�.�����0���(�Ck�J��Ԧ2�2W�t�_��U���,3+3�f��c�h��5n��ba�w9df!C�:>�`������� ZU�_v*n�W�;�;���l`��c�!��x���Ѕp���]^�5nג��eϹX�e3���qPU27H2p;�d�]tn�G��qf��Tw������%2P80U��L85������ptm7l�����Ձ��
NP�}�($�zs!u~zƕ���.;%�re����=)9Έj)�]9%��N�X����ƾ0[q)�$W�\��j��g
&C�)�nv���>Ҏ���YOo��T;��ު���h0Ծ1��9h�)\c�I�c=Q��~���O��s#jB��0t���;;)�Cl�٫i�$Tf�w>ÿ���f�!2LQ'Oױ�|(���߮7#Zui�/v�ٺ\�P�(����	y�E:���I�����v)Ζ�c��w����T��aQ;J��{��Tݿ������D�A8p��Ƈ�>2u�q�o9����~���l�����M��'����̫Bd���r�����%�	ǔ�)���ro i���O4h�P>�����6$蹗��~Kkuuױ� ��&����>��%
��Y\~�H�G�9�Q�{�\0���,��F,�H�S2-X���,	�#����~zٺ�9�M[�sAgVZb��|�j:�p�˜�u�I�œ�q�=m�`_p~1�-��1���$���o���>��SC�l< �@�B��i�-Izz
�\aٻ3ժ�k�~/�<�SA�7s��j���<CV\z��f"^�R�i0�xYer�@U}���S�$C&��͕�c#���r<`�0Bu��۳B>���ͫK��$"��g50�F�+2(Ays-���e��
�E�1J4��T�_Ub�@�e�p�/t�� Y��{�ά�Y!�{�*-f|�A�Թ�_э�G]��4 �AiZY�:.&1FF�I ��❌|��ʝ YԆƂ��}��.�u�K~��pp�G;s[f����s��p�[��Vo-��2 ������ Wc!B�.��Ēŭ���C���R< Mt��u�VB�:�X��u@�s����N����'Z��Dm�i�Q�r��1�!�Qwh}L��&���T�]Y����ԗ_���e�g�_��l_�Ң'�̨C?�Uo9�l�s<����_(J��e�����j��t�R���gڡ�?
��5|h�轵��z����<_����uCJ���dJ���?;x���U�mE{,��><5�5��Ս��Ƣ����h8���6��!ld�M~cEb��A���E�ʳY�C�Q�x�Q1�C��GI�D� wKhb�����7u��&�\g�)�����)�O];��-؟:�*'`G�|��������lT�K����M|9]��Ef��^���Qc#�	(?ߝ�;	Kl�����Q��jr�k������bv��������$:1�[]�4=���� "h��^"6M�+d�&�j7O�u7��ݑ�g_���Z?8�fmG���&/�4	Wa�*�ƿ\Ү��2I�a��a���$�e�pQ&j��8/�̜��`8��ռ�R��M��W �(�}��Fg�U8H����j�2���>6XFF��mX�5�rI��,l<���k��V�t]r}�C�hR<��I5�g���u��Z8�9��,��j#N�q���Ua7Z���^�_L8%[�t�;��,�qRkn�?�s���ᆋ�P�բ�� �i�T��Ӟՠ�U��Dy4n�؋r������/���aY �
�J�������D��#L��$�����gsXuT>e[��*�Y�>��9�A��/֎��m���c�Bڱ�3T�q�d�����2m��|����+�ڸCۖo��`�ڃ/Wn��ju�QSlt�x@h��)?��R��pᇎ��W�������ֈp�
T�ر�Gl�Z&����%֥Ds��t���ڠ����u����LG2(������Tz�
�3��(�L�it���K��tA��Ee�JN[I˽�w�}GMD�f��僎�\(#!�r�a����v�ǁ���%i�5pL>��<5�5�o8�Μ[m�k�����t��P(j[�U]������ϒQߧ�}�4��S���nSr�|�U!�.�O<���1R-�q�U�m��kN��;���C��]cׁ[N-�C4>e��Ui������)υ��D�b��?�0�}�	R%4�"5&G�5���3����)��@6%AG�].���=�{8�d�K�B;�?�-g�s,mt*��4�oZ즌9������ipR�Rƨd�f��)��]��?��b�^��-�},O@E���{�f*'����H�U��MO��w�'G	��;6����i �����(m��6�\���e��A[3�k�Ɏ�r�R��O2Ӡ	i�����2�!�����К� �5�7�������C6Qcy���?hr�3}	3)O��!/�g�?T���߰ͫ�����)x@�cKB�&��P���$������X������R�K.���ʬ����&T].+Wt�4\��+���>�O��]gЛ��WH�H#
$��+s��Ԯ#N�;=$P�)W�k�U�EL}2u\FJ�h⼬[ [�����>2i�n�!�N�P@�佒hk��s^~��.�,���ݽɄ�]t��b	�؎���#�o�&�=�V�6h)zK(M��JT���&8�ƽW*RKM��O4g�^ꑯY����5�o�_d�Y���Y�a?"�+����b�d�� ^-�$�'���,~?��%(��G�x�p��&����U���9�Ft���K���Da�vw�����.a���4����r�8%s�Aw�@n���n��2��d��b�����Y�g#�k�r]��_��P����u��;� �����lo1��{��tJ��n�+�hE=l�U�P��}\���b���W�?�z븦���ؠ�� I�n�������!!1J�s*�2�qt�at(���) �����|��������v�8���^��u��ݚ�5��q�z�~�UW*�?k�K݄�sq�O�H�pc��{�FMda:x́�u�LF�
h/۬�5z�����\���C@�WNKϠ�*���m���bĎ���۳3���Ĝ�aU:
���ě�����|�pa��bH��3�,F�a�f���"ښ&Ψ�c�X�%a����k:Q���x�2%	�h�Y�=��,�E��zpXs[z�d1[eS�ca�F±�_�[��]5�[q�i�8�B �
��=��'�� �-�d@�����}�#����E"勈{��"[U��-W�_��	��O{$�]��Q~�l�<��J~�u3�`�����n:�B�[�����rh��&تٞx9��A����	��c�zPb�E�jο䗒�`|Tc���W=�B��D4�DK��3�1h0`�zP�?@��_%��������g\sZ.�هw��J������'��%9�T!�N�Z�Wc#j�N�c�.uO��mA��滙���-N�8M)��U�I�ng7��N�=�$:Sa�2�Š�6���iIl^l��i�>�J?�����t�~��8hW��	Nr��u�~��\GE���
]YN��f*?��������X�k^��αF�������1ȹ�Q�6���-!��Ձ��̺�o%���h[����)y��g�~@����:8���e��acٝ��ێ�LG'ߑ��B�Ǎ�B�N��Z�uy��Q�ٌL��	4���,W���y�}w˗�0��z��BQ%�I��'Eeda�1���^>�Q�+vuh	��i#�����P��X;��ɝ{ SvT
޲NG,���JTfx<l�����ҳt��9`�g0�ϛ�����?�ι��-�#�U�UsSl�f"�u��s��a��[�1�R2�^1��se*��>�����}R��~���h��lڎ=��0u���|&zLbU�sfR*�$W_�w�u�F�9�ak�4��5~{1���N&��ěg����`ؒ/��ج�������+�����'L.�1��=�d�c��u-5����x�K��8�h�9Z��O�77��K(u_�:Bس����
���5n骜�$_RN�E}Z�Z��kݪ����7r}�ќ|e�;Q4��0|#���I��ݗe��qw��<2 ���	��KR��ݭ���NT���[��!TO8z'����������N(+,]�I��-�H�����?���M�U�5��{	�4)�n��%iѲb�n��u��z����fU�������q��>P'��%5Ҭy+�s���L�y�$Ώn1�;�x����:�z�����T�
st��"VD"7U�J��kd�JJ�h�OւNK&ɀ�b�|o��uӜ��`2��鿦�Z܋ȭ���3Xw��#��w歸.Zw�4~:�l�A�A[�"���Y�lPИ&�W^�TՊ�mr��/�M����t
�ho��=����;��%{� �/ ��a�-�`3��"}Ѫe��̫�=*����>@���T�~i]f��?s�(\���@�D�_��C�􇎓��~~G�uvE��&�0��~v�V��%^ ?��M��x�5A����&�[yп��R� ,��22��0���������HOӽm��t�n/P�#� 1�6���V�9�	�:Da�aA��������$3���#��L<͏ؤU����~�>���Iٺ��F��v'�"z4�6������
|����ަ�)+���E��������?�%FK�J�a��|�y�;}�43�	��?۔D\�2�.\�o�_��?,�.�7B����	�S����	.-��dF�u�8�=	����=� W��3�M�5ul��dN@P�Z��ub�c��R��,F���!�F�*v�h=��CQ�I,�.3CSJQw���δ�8:�E,)�@�����͒��t1�����?���Z���W�uM�{��n�����"������V����6�J�Ğ���Q�>:S]�c��✎9z��ش��zH����%jd�J,�|�kW��e<o�=�ۆٕ� ����/Z��������R�d��
�r�⻡�rݪK�r��8{�j�i����X�˶y
(�>��Ζ��[��+�!�3��%2 ���)"Єi���mZ�X�(^��><H��\Rӡ�Y+w��[d��S��2�G{]гu\9�7����O�U��.�?��.�"d���~lט�4�-J��;Q�p�����w����b�)��>����j�������C��*ĝo�i�8���Pb~�����eդ�t��T�Sc�!J�!r���
�m�	C�(u��B���U���Õͦ�+�Τ&�U���"%��	]��B2�� r�_to�]j@>���\]"�We�ll�t_�?|P�K��F���	���~���܇E�"L��r����T�p*����yεx�x,���>��Ϙݯ����)ѯ|-��V.�F��`IKc�J����&h?�	��97_G��ϡ�ƭwV���B�'�~�P��D��g%�\�uMn��� �1x	�W����2)]e���*��u�M0{ݺaYkF�/���L	�neR1��`�C�ߧO�M�_�_QXMwl���F��p[cn��"����8�n2�V*%�����Qb���}铋:�<bJ�"�˨��cDl�a)5v=^�l�;��{
�c*�Z�Ȁ��dr�X9?�����-�A7�[ga���q�%C�b�$0�яr7����_
]j����6�qY�ގ"�(<�A�j�'%�8|���G���S�d�\ %-z[���#e�?(6��q��]�R�5	�|=���Q�/Ȯ
�13�0��j�U�'���/2�Gi�h�v-ں^J���r���E�F0�V���j�w��̕~���X��Ru�)��x��A�ו��p�`�xu����x9B�p#֯i�Zɣ#��n�[��Uɿ'�P��)2E�>�s�obAC�|�B9���JuO=�ɀ�6#�5���)�S�yo3>\�(�}j�1pv�*T�x:�n�K��*����{z��Խ�U����ja5ү����¹�5�y�w���Y�=	Ϧ� ?a+󀏷;`���xd�a�3w+rV�l(P��yD��SJ��7���SӒ27�����W��� �Q��� ���Z���N�j��2�� ��4� U5��8X�����W�>�? ��&���>��N�tv�J:2l�Cl������{��P���]�Õ�	D4��Eb�<jt�������1)���4|��1UA��_,�!�ԧȄ�&XL[�S�~#�n�'��{V�}��{���0\S�{� ~7�Z5`S����;"�FP��F�^�-���28m��GW玘-�XZ!˼	kj��‹aU��L{Ģ6�%E�0\�kM������_��D4�)��]����<�J�y�%�����y �R2@��Aa6�Y����޶��B5e�}gG�,A�cǶ2�f--h�WN���ig�}�7ȸ7ٯ�ᄞ�?a��X�#$�4�E�B�)��>���K"��O�)�m8¥o3֣��p�Jd=׳�DJ�X+:�{ v�ǅ�)1tT�O����.7 ��'E̷']$0zpW-X}^
�ߑ���Y
:a$���Ktsa˜i�"%��c��|�~s�v�~(y��8%L�IR�ɮ-j;g�v"�
��A�2�ɀ��"$�U0N��?vg`�*�G��CWK�<�'���&f�+���MU��A㜜�P�G-�����S}?7[�u�AJ��8�m=3�7�w����nr�%O<�+��+�뛂H9��Q�ld��PG�E��I�z��`����`�3�E��7���!��MB�σXLe�
e��*ȝw��{�w_b���7-߆/̆��C����O�a�eW�<ٻX�.�ѳ�K>�.���.��o~ �� o�d
�Z7��!�1�:h���.�N������MQ
�1~U	������>M��H�xQB�``22�ċ嘠X/%F����4"���4��x0ij�K&�q���E�J�h�C���_\O���D]0�����+�E�!U�;I�K:�C̯ƍ��^H�b�*�}�Ľ�J*͓�oꋫ��8��n�y��		.Q@X��]I�deY���ْz����b��0݆v�Q[��F���A�%*;[z ���#[�-�V�d�3_A!p�R�r~1>��ZX/)_�
��2B�w!�ߏ�Nc@ie�w�@��Oݢ�t�S��e� ��P5+�������+�K%��O���˥����4#I����p�d�/eg^��e����o� ��/�bC��Kw{A'��!&b�B�Ϯ6A�����#m��g�����W7gXR��}G6�&pt�?&��ΗM��������^E]�����(.�-�t+rl������/��݂�Į���"�c�u�H��EI$����g"�y��<�^џSW�>�/v����K������.��8��ľs�}�H����$�������TuFs�_�W�����γe�]88���/}Ϩ&�1��<6,��')Su��F_�	��\ր�׎�bg��hE���H$��h�M�J���-W��x�(�_M��\�9Uܼ�:0�Q���tc�a�C�'a����K��r�l�@��U�t����YX���P��,иV3%N����`��:��T�:}6$�����h�oJKt���s;?C	������I�-�}��l}"����9�* �+��3R�*s���\zg�#�kd@�6�Vլ"��jEj�;�
�c�Hi�!�HU
g��v�#��;�2�)vv������U�]/O���TyvZ#m��a�f�ɄA��O"|���-�uXڥ˸��C�1��zG��U�D1�WoԬM�lZ3bsc�U6���q�p�&�����z,΅���yoeu�%iqV�bz�<�\8����M�k�2�[�!��%]":�,�o�m�_H���%J辫+m*�}�-ws�.�oj,��7���ZKi5F�S%+�q�S���\�"�N�zY�#�p�s$A�ɓ��XFz+B�]]i4Ԁ�Kί���
~7�?.�}�>Q��Xn�)���+�=*�kq�K+������`AS�+F�Y�����&���,�8��������Z���]�FEZ`GD��{�`8���w���$�F4,͑v�C���E�D�7��Q�[Zl��.�e��%��ɍ,����@�mj17$���9R�5R�c��Y��ڴ$�*��.�W.�b�'֣�zg_P��2��#�A�H+�{�d�6(���nªU�'�u�����v�ի8^q ��_�U4Xǯ��0d[=U:�_b<WF:����2)�s-?�zY/�K�s$a�g+�k�o��o�{�ygH(W���Dmx��ݻ��8Y�XW��@	�C�� ?�l	h�1�t��3�"�u���=��V� ��eb�"/;�)��Q�������e��,=�'l5#b�~��6\=���ß}!�HޢK����{!�$;e(��-u�fI�DYA8��(�$�!�����G�������w\�+�	/��03�/�⊾���`��y|}���y��F��'ӯ
ެ�7��Q��ӓM�l�0�Q��U�!�����s�b�������s,�����O�'�;�	�U�Euш1�;!G�C���^JC���b%�u�ӵ�V'�(�8J��Ӻ�C�B��Z�'\�H�B�>�4�"��ȺIC{!�=���旗[T��<D��B��𐎗��5���M�2��8F�+|�Gr��B|�v�?f8QG;�}�*ѱ��b���*���X���E0o�[�ta���O�a:�c�W��B�?P���$�v�P,�c��a�T�s�t���#:ͽM�\�D2�)��Ű��w��ǲ`��k�A��ޝ�6�K<��d�+`��2�ހ�(]5�3�ɖ�������HC�9�nI'RʑC�������+�o_�'��7~�T[˲�֌�`+���槐j�`%��.Hf"6���aa]���~�Olx��5�pI�����~���-G���ӟ�!�,~��V��s����d�jv�:���R��pO�h2w#"N}�<�P�O������3����ܩ�K��O;բ���,kᦿj&vDB�H��Y�I-K�4V�P�����ܬ�n����Y���?��v��r���&!.�1[=y��v;7��d�nuKC�SwgSy"���!�, ���b��u����k�*���0ƻ���RNC(7���i'ȍCSL���g[Gzw��f΢��V�uu�G3s�/��zz��,��O_�1��E�j���
mG?��&��n�y_ �l���a����N��o[�e]��!9�_Ns�I���=��<��Hp�Ā6�I*h�N�	����6*�S�~w��b��D�q�k%��u���g`:�ys|;�����+�9���.wz�5p��|�#HRC�����}�$��,j�x������ Ջb��_�N5���[��N!;&�+� OE�f7�2DA���|#�	��� �/;��E��b��2�\ϑ{I�v-����{v@��3h�G�n��2�`]$�@������>�&}Zr�r1��O:%)����؜�[~��v�k�X�Z7ћ@Sl�z#��`����~���d(8�������LQ<��ZuUa祔��![��|Eh���l��[�9����q��(����36�v��א��$�Wp�,ۃ6^`�Pl��qG��dZg�,X��eZ����{\��;W�$��7:~d�d&�[]���Xn���xr�v�#�5}�%�m��ajE����.���"����U�m�G�S�G�c����⾘�q�z)lP�,f8�<�V풅ל�_��w�|ȗ��+��W/�r���fM+�ol��}Y�@��^X��q�\�&lZE<���\��#̶�}��e$,�׌lT:�6�Т>���r�D�C����B��2�/���+�����mL^I�+pxdq�:7HM1:���}ۡ&-z�[��z[���G׆5�p��o��QU`�Ce���D��#[o���2���#V�6"�#��v�C������jm:K�Ɠw��������i������Оf�s̱3����m;��������۞��A2�ܑ�b������X�D�ݨ�	��a�{��\������t��Z����s�������7��`�ݑ!������ߠ���6�4���fg�_�N#����ɀ3#����dy���tO�tk�*WR�"���͒V�^�ܙŌ��\�l��7��ᘰ�d��B����7��?���!�&"��p����Y�X�y'������c�������q1z�\��յ��@�3W�Z�n���-��b���(Pc�*0X.W~�vn^j:}�lV;��~�M:����i�I�]��R�S����7e��G�E�I��;�vO?������Ji�kG?v ����%�1�5`0[]���?�,�r�$\�����gkX}��s:�yl_Z-o��'�xe¨��}'��Ω��\au�d٠��[�C��ͅ�
�2���sm�1<�6�S�'����9��'�}���/b.��s�!��ȥ��ǯV��\O���a�,��h�}�E=͋�w�p���\�豥�~V��r���2�#���]{rȏ˞�VAg%m��U����B��P/m.�/;�9�h%���AG奭8gKhE��Y1�qo�Ąl�
J���L��]�S�ڋ=�����V��8:qǳynuy���?�<���-Ϊ�e1���ihЛ6��uϬ������k`�pҿ�����/ F>4(?�[���Y�)d��:.J��ZTs�Mqdm���Z�GB�8�܃�k��\���fz��?d@����@��n��=�|��P��ݑ{�7zBw���yK�vl:oÞp�2�>�9��@��?/Z��HE]�w�,���f�/�e_좼1�L����u�aY*�9c���f:�&זT��ٷ&���'Z�؁c��i%�Jn7�SN��Uܹ_����$��ɬ��XC��B�$�V[5d�m:�ɸ�h������x�H�40+}q�tR�^I˙|�R��*̪0��}�)K˹h�P�,������n����h}�qt�$�U��h�x@�>vﰢUX�p��+��g�(��Ch�s�AJri�|�\��>k��y��
��Kg���?\�����cm����!맭IC75��D��F�H+K{�W��ר��؜�,lhMg�j��Nҟ-:�G�������.-q�%�<�uH*��M5ļ8Y�u���� *ig�@�N�"8�<b�4�N?���Jոɲ�`��/��M���-�]�����XO+���*bBn g'�PY������/�o[���Kҩ�Ƥ��f�??������QU��s�R���0���<�:,��r��x����9���# xn�6�x�G���Ġ�J�:�̹����;	/�8	U��t��5ߺR��D���
��
ʸ����T����o�0]
\�,�PTww=��i�]t����n�Y��?fJ	ܜ �\h��l�qu�v����+�˯g.(�z>�:=��̙�$�i$+`�����w��i�Jtj�m:i�O��-�z#]�j�_���F�>�/#|�2]�a+Y#Y[��m����JA������Gʳ=h�X�����X�M���Yo�6�q؂W0$k�xyx;I��T�-�G?0�qֲ�׾������8�S�;`�7�_"�k1�ɥ�9�e��T�����>�Rg��j�׳V��ɰ�Z"���]��7�JG�=�O���/�!w���3������-5�U�H����z�#%Wk�~>����g}����Y*���u�I�Ec�Oc'Z�+�<����'{�*���"��F4]����:jX�p15n���k'$�:��;ϽtC��u�n {�}2 m�\m<m7�u�����C%"�Um�6����oeᯙ*�bGv����>8�,��Y�9��F����n~<s���]�VN�n��AB�'�8=��E9�x�?C��L۬\�6�xk�t*"	��V>E�6,�z�W���k�_�b��2�9%��3$�!��in�
��}�S��ɒc~}�f��R�d�UȒ���2m�5��}Ֆ*�a|9B|�4��4�:#��O�}�`9�*&��w��� ����j����h*�c���K>���@􁮛�7�Ʈ��}!J���7O�Nu����ic'%C/c�i%hh����~���U�@G��>Ed�nȃ�EIg����r����fΧ�1(a
1$.�f_8��Y�}}��YV�CYZb3>L��#��S=�~��s8~d���3�q|�H�,��EM�O���O�����#�t����[D�6�n�L�~�vꑤh�Yվ?P|��r����\cf�L��>dh�<����+��[k������x:�>�?��}��k�6��b��Ɲ�\�CG`��h�[�cn�6���G��>׫͸#}�;��U���n�7nʆ��0������ZnSI;��Ĳ��Ƅs+>qW^HL���U�N���_��]Ka�e�����r�GjSS�##	㏭W-�)VQ�W��0�|�sa7�xܷ-f�C���a��U{�}Z�w��>���(�0ݍ9|�d��Vmu�R<�R��Zb�Mx�^�n^�ԛ��wb@�]���,�9?sh��j�>'�i�nW|d�Y�I�����<�G���!2@j3G1"�!lS�ӉY�4>]űEL���&���ޙ�ft��ߦ����$���o;5<g�댽��<�3q�?��:�f�}!1�b���v�<�ۥ-Z���y�o�꼼�h��MMU���^�"§� �b?ئҺ��0�������Px��[�����~W��	�w�����~W5$z�9��[A�$��Ef�F�`��
h/��06���}���������۫��w�#��m׮+S�n�<�0e�hR�!��W�3W��/�8E=�G ��Uh��!^�{d�K��~�g�;��+m����M_YnT{���`�-�T�7�?vN~Vhꁦ����2j6+�ļ�82Љ>�$���i]�1�Ir5�ڜk�h����;��:�lI/��:�q��U�>�u�,���d%��z���j���z��߾��a�%��v����ƌ��fDS޶�]V5`��̴D}t��L)A�V+�g1��o�F�ۛ׫3�����a�-���U�%�ʌ6MbG߶�s� ~*�L��J���0���	��n�L32��L���4�u]���l����!���|>1��(5��=�kw0�dQ'���[Uԯ����M9@S��G,�Ѡav�k6X�A������Fx��n��}���b_�vI�Rd����n�7nqj3ʁCZQI?>ZNt���@7��t;\��fE�ѓm_�w���R�'.�֛�o�^!�s	h�6Y�kJ7'tY�v������,��3�\ܳ��ݛ�־�~��}��|֚���ut��@^���uP�� ��W�����U6���5�qg�#���g.d Ǻ�O ߔ]EWմ�^��HI&��I��^A�}}���,,,��|;�3���,�	��R��o��[��b��>�j����7r����!��U�òW�
�v,���#®����񅸴��+֐��i�����L�	����R?){����2�Z�ɀ6��R��I�D����i���«�Y�YA���>��3.��]�&o&J�L�m��|L18P9Qj���Gr�;~��}5u�֤:D��%>ۓ�Ow���vq(��h�����xFh�[�"l	@��@+'��&��Č����C�U=�|�WI<�*-����+�P���sw�{���?����c��K+�ОӭP���"�kL��7��@:kN��+���&�=,N����L��8u�� 0�d�o���l=U+����٤��Y�m�x�p#�ayJ6U4�j�wmdu�i������	�JG��j��c�@7@�k�3nW;F+��W|�^i§�<Ẇ}�L�����fV5C�"FcZd�,H�������wK78�m��	�$�����������bt�+�$Ъk�$��V�p��K>g�||�^$�2Az�@Ԏ����؟�� /~_,h���3� �z<��U]~2 �;r���t��8|�ߢI+5��tSH�gMf�Y�W�վ{d@�rd՜�����qԝݨ��u%��7Q������4�zl��^�Z�� z���ub.�{�5 ��z����g�T����)�B�9�J]���,��B���p�����e�ۃ�Ϊ���ƊD�`1�ր�o�+�������|���1/�����-5E���e����O7pN��G.����g� Z2�M9��Y�j��^���*]i7*ϭ�&V9��FS䉛�G����\�ܐϨ�T'��V�b�Z����7[>yZZO�"%�Nws��������A�'X�TmtdO��}��O?E~�oFo~��R�61TJlZS�l
^1�����)IjZ�5xd�9K�����w[�(��p��~9'΄i����p��"��ڛB!6�3G���o�1`p�⎶`��!��1H��8g�=�k!o�#�pl9%��_�tP3�|k��s�.-�t��Q�Y�����2c��5KU�4��tv�䀜6Zu)��030O�+�ۀJ��r��I!��s�2\�i:��3}+���<��i�(�?6�j5�#�>���2�A'��tCY�R��Ю����3S7����`��sn��'|�P̅rR�{�_	�wϔ��"�
X�$�G{KU����v�q�ʫ|���BvD�pt�T�i�+��H0�WB���{��=�5p�c�].ZK�զ�fP��Bp�J洯U+>������U���l���JF.IM����sש�^O�{��A��U�'�zZ1��ߟ�g���56���}�#�qvӂ7��=��z����� �w.A�T&4:�mR��P�1TQK���E3!_�ȳ���[���Y_����3,nI2���"9�s�r�˲i1e�ven��Zh
�eK`�+�$d��
[�/,U��oT��N[tF�����M �Q6��~��08Vf��61r0�����<�O�
�Ҏ�������cJ�ҟ��G'V��A����nF�_M��A���'J�xf�uQC�:�4d�爟]W�~��ۋ4LKy�_nqo�67b��dM�e��!I�h�.��x�CXf�H6�L�hg��?��W��MCq{z~�r���ԛ��f~�Z��FN�ɭ� �@���$׼4|���v�:^\��?Y�֣]����K����m��NG.߿����f����-���*��EK�	����N�.��|gA��v������d@��52 @v�y���֓�u������>�A���!�*�H�A+�"W��M����4�=����U�,�o��d�~j�,�{T�v����U�qy�(R��[�c��mQ����C8���_���(E5�n���h�g��+�^��}��Zfg�i��Ͷ�r�m./I�u�S&�Yc���G�q��%����h��z:��n����B���[�*�6���,�����C�C�X�*�G`"��?������D�p�+��/{�n���[�x~2�q3�3��p������>EI��)5�Y�].��͓?XZ�3�,�ɕ;{#�@Z�
�uR=ZG�G,���+7l}���q��8����Ԇ:Q�ؓ,����	Vm�5���/���B�{�a��
��'t�G�����y��v!����榍X�X�D�����ۊU�>b�O�,&�TD�\<i큝�o~���E׊%d{�7u��sp.'̴n �e�p�0?��d�X�Q����*���,�L�
��8��ë�[Z��<� �_�GY�0�h��y#�wı�xU6t_,�����JK�s�&�nI�Bλ�|K��Svw��R������mm��k)Ѝ��_�A���\M	2.�ν�ͮ1�b�/5�	7�4T�{�#]������0�ՋZi,ڟ�� ��J��p-�2L��P�5%�m���?U��e;,F�@�K�ʯf��-�;V5ج�����/�� �-��X�a�w�Ӓz ��0��h�dV�e��p���Mt=j��%Y~���u?){�ux%���Yl�����7k��nv���̀��j����ϬRߗBF7�5�+�s.K�$�r��\�? H�.У_]q,|�b]�igl��M��a�[M&_��B��_^�أ�/n�X�6�[�*I 'z3����'�-2�s���˝��XVo��_�ĉ�l�/���nf��qs%�š*K�ek��ǍQ�GUL� �T�ZY��y4�|�8��B��_j�mO�
�7���N����ェ����j��XQr����x�{QKX�M�*ts���S\�S~��W�s�
������._'��#�t|��U��������G�v����:*�F�cA��üť��3x�TK�2i��Xgگ6�	���-�9�|i���0S|
�(x������A�3%�p1��1q(Ma����A��a�s6���D	8HM��3em�y��h����N��cB����US�<i7ظ���Q�
N�_f�&�ҭ�n���V�����E��
v7$Z���k�C�Ck��?k��#$���۾݁��ok25祫��pz�xA���}|���6�*A}]�<�5w\���ـ��t�'�:C��k��Ru�5=.ڣf�`��[�u�B� �
��|�*��_�˯@�4n22`hZ6<�S���_��=�C@o�{�*uޅZ�g�a���qe��Mg1{]�owY�M(ea@7�V�����(5D�9D6�?�NӐL�́0'dF�̉�&{��SPA����q���BxBQ�8�G�D_�v����>�o���i�+��z/.�8�O"�D���4��$ԩz[��е�E��mbu�C��h|�Y����hD^	�n�9��B��XSՎ�K�#�h&��E���OCk�H}�b�z���
����R�V
3)���t��Hg����%)/[�V~õ\qk�a�I���f��b�/�?�����퟽���ʧ�(���腺���Qy�}�z㢪������+D�B��`$�Q�s�y��e_����S����
�;^A�%壂z�nY�C�$�dI�<�34 ����{xݣ���T&�������*�c����8�4jӂz��̧a�e�迓7$��H��޹�~�B�Hk�� �q���H}����E�����!.��D���S�6zc����+�R�$��ŵ��ԝ:�*�y����E��å���B��07��j�c�k=�O+���R���?J(U{7S�狠	��I���8V����=���ֽ���o��;)�����Q`�S������a{tF���s:o|Wo�Q��+?
vYNT��AI�j�ã+���E�c�f:յ�^Uo��s{���~Y�'\-�L9��j��a0�k
�{��Fd)1�g~֊���ݽ)w���\�t�,vݏ�	͑b�~�DypɌ_��4���%?��c�8n�&���q�ܟL��q�R��,Ʉ�A6�h��X^���hh�f���"��E!�Y�� fF�����B����쮯���oO,?�	�b��{\���w�jl?��"а3����=����k�o�@Y:*��R'>��ӝ�d����7l9
�~�z���uen��������\���$R�`��d��g��2���ā�B�=Ѽ	s�lu�@`�@����Hg�e��IGQ���r;��ݍ�#f�>�xm������	y�Q�l�Q�fqF)_K�P�o��l�{�]�����9� ��ґm���搢jms��w�aUy���'������B�`��/�2���+�u��o^B#ZX�=p(�}q���}\��H!=<�hc�aX|[֦��-�q� )����Y�����	���S�	�	X�"
�\Gj./���o�	�8	�IA�{6o,7k�%�40�{:���DK�9��K�8��u���%�8(��'�uwlB�����v,���3������Ì�N}�46�rx܅GkN1�ۧ,�-��Z,1\ц����Dg^��Ϊ��-���҆6�"��՟��"��
=�,�����v�ۺ��i�Z�s��gk;��MA"�*���)�<��]h� �q�O�]69����o������؅�9��Nd��tc�)��F|yk��3�Qw�G�g�,�7��L+\K��FNG���l�􅮾m�����^*-טƉب����*���}=�5j�$*j]�(�n�����s�mT���
ҋ] �Ľ躹ܐ�F=?^����~L{�ю��o�r�l�
�z+�ǹ�b�mCT1	�Vz�ZH�*moZhZ��+��d<zD.d�q���)u�dn�C_-t7�[�[�%�{�9�<b��\s�� *�r%.����U�J޴�����r�a}���؉�w�&����|Y0��V�A{�U[�Ű�����i��g6��]"o�K1���?��4�����qʜC�!�N!au�+F]J��]+�c��>+7\����X�l��]_�o��.<��iU�|�\��V���Hi(�Y�䁰�̐����h�uGf�E�M��p�6�|���E�P�����+�~>O
��s��^j��Y�����Uf�?LyvyI�x2=>:�<�˸���?hEg7�0~��e"<&8��h��x�Y�W�M!�i㽚R�7Ym�7� �k�>���֙ܵ�����c#3�pa=�O	y���]��7G'^�о�cs�9�)�r���?]�ܕ����4�Э4�>g߹Z3�]=��}|=�[�$y���K�X�4}���~��X��sQ���S�����%��7 8�c�ꋑ�`D���*�J�
�V���Y��ֲ �(>�]��ԒЁ']ă��n� �uX�Uٽ�q�G�k����ʬ�#�� P���brKH�d@�Q�]Η���|�__�*R�*�@��LOR�f���G�z\��,�.��1�D�p���yr��^f~�:�JD{��ڤ8z�Z]Ǖ��W���L��)� ������c�g)�Y���ԵV2�7��|���_kx;5�o����H���O��f��2�tc���{@�����&\��t�8d���;;/����fXH�UO�u� ��
4�4R�h��}�J�U��ݜ��^m�� �W�նg@����Cr%{�:�n�vk7�~�X�,�gPS���O*%""%�J��AA���{D�F@@$"�FZ�]:�J�5����Ӟ93g��kf��}������#����6��*�2|M�6�Ō"���= �e��\��hz+"��� ��_����lW�E�] G��f�a����kjn���m��#;���s���Z���������'��Ti\F�8��.��v�S��̙D��A��ӊ���7ws4
",�ˏV��Ǣ�Γt!�iK�7b*�f.5��,��z>NB�B��yII��OuYL��gT�I �B8�~�x󱎧�6� o��Gɗ)�t��_�퍎"mo�"t()v��J,0kC��8�E��-�F������`�v8C�;�������������ŧAK	�����j��V#�s宓^���OW�)eAM���Q�l�ןqrO|�����pmя+w�V�\8Y(���;r�u
퀠X=�6�$,���>��p��=i�r�r�䀅���i|�P���F�Yo�:�ov�#�T%��<�q�qd��v����}�)���
w�)4)\ t.�N�):4|��˩/c�R��GyH1AAmumEUv������W(���T3�g���jj�)fGV�Z������{�  ������:��Mܟ6�����Ӈ��H�^�n�3d�V>�Z���6;?�OI�	���ضd�쒳�*�����Rd�	u�����ڷ�[�+y�V���](m���6aM��߬�p���Fv�$�?Iք�{;��l���G{;`�@_����.����u2��gw����z����SBI�S⍏��=�{��T��n/��~O\���V�E쩿�T{W?���UU���T�⟸ ̣���&�@𯛓\���9~D��F����c2�Ԩ{���#���j<T���v�q�c3��<�p3�`��x�9Iˑo&j7���L�Dv��_��U��I<��ƭ�OF�TS�;��O�D�F
2,����뜙Z4 gK��Q!i��ً�O�M������񝂚fn�W��6�n�U��IH�R?�ZW0��i�qm�}���/���a��麳�A��~�|��h[d����z��t��+�����r�Z��0�ba��r|sj:�q���ثV���NC?T�j(��s�a�6�: ���M�Ǻl��|f���#�<{��ӧv���c��R3-	m�1���a%S�9�gΗ�-�������Z6(a!�Mn{X�PM��Ԥi?	d��s5��*_5k�쭊�M(�LU,�Ӽ2D3 ���;���:�NF�j,��vt��;l53�ڶK���׺�zO8�x���t`�-�/ �"��u�v��>>8��򻮚'S�[Q:KJoE`��7v8���w&��������=Du�t�EI��7��ė�=�ž%b~u#���=G@F&�Bn%\*{^��Y�:<��-N�Gr��&7�C�J�NOҸ���Z�[�OT3�.Ny$r)�R�H���Վ�O�w�0�!/$۴�ov`O���o�Rѷ\��ٗ� ������!�o�5kE��-��_D�Oj�fJM67`���D�
�.8@"Zd�����=�Y*�?O/��N���ʟ�>�Mi�z�9��詳פ�|s6���e��s������Ǜ����6�ɴ��}yV����%�S�2�h1Χf�(0)��Bh*�r̅r@SS�F�Y��`�,N�^@���6_�vh��8uF�:��3������b�2O�{�(+���i��%c�vP�@GrOc��k��B�g���e{���8m�J�ҜXEv���y��Iء�A�g@��P����h*�H8$������Z{ ��^B�AL��l����r&�	�@đo��l~�h���Ѭ��*�W������'4��X��(`��{�NN������aEۣo{���!'���3��_�Y�Ǵ u��iŁڼR/~�Z� (r+<�-����|N��q�m�O�B�sۀ�?}Uѕ0�^������������_+|�����f4��rm˥U����i�	�������aN�}A�tEǫ�՘�I�����[�*�f���(���aA�P�ǁ���%w��e�T��S?B|!!0����G�]�4j��};z{�r�-�(N��^�%�l�è1�3�]hR�ޥr��c+��ko�;A��p�����ޘw+G�"�g��9�������H�8M��F�[�u�헰���n��R�%sR�հ��~�+E�SN���%v�(�˫����Q�1��b;7��dۢ���u�[?�l��o�M[���ޞ��vXXl�'1�Z�ʓ������&���ާq,�|�U2��S>q�aQ���[HzC������H�-�&b'|�D�g��~NC�t���G��Ty�OzT64�U��>�P�<T5t���Ja�.)WH�B�kaX޹[󏐯*z�Dz�q� �g9Ln`=�;	G��`�a󽗽x1\`��t��ݱ�������.H��GY����-ؽ����O��+Ԍa|+�ѵ�N���9t�{��%����N�ڴ�|�d��O���:U������]ϡ�0 )����G�_5l���Z�E7=�v����hҮMbJ��w<6f짻R!.�A�"m�*^CD�R���^6o�᜾��i���޽{F�*������H̜��P��+��KH���:��NAm+�p�3W�s/�~����h�3�{����c����)�_L~MZ�<A^��7��eq�Z���M
$і{pΞ���M�
x��� G��i��#v�Ct�u0.���H'>�x��q�K{�jͶ�qUQ�f�c�!�Jb��6�������^�Z���_�Zx��lB�!;79���N�m������ȅ�G�v��"�����īQK�f����[�@nF��4!���)��688���B� �8B�0�@�#�`߿��N�BW/�e�V�*�|�x�m��Y�M�w��G9#~���2f���������0~V��_��kf��l�hr����)W����|sϦY�s(�J~�P��u��]Zvp�AU�&�8����%����-�K�W����o��0�Cqb[��@��d��&b+D����Z��M�凉�>r�����r�A�­ P��Q�����W<[O��B��Z�ʶ�])�A���
B�����qs�Yǎ�xU�A���.���0���V��t��I{~9	����<=z�eQ�rs�[����l�/��RI�T�&k'�Ы�ę��=-��SS����3��Tۢ�E���WX��O�^������[ƕ0�ϐ0�<rr�%��4�&�5�������X���N�@h���W�RW�mŒ2�Ui�rɆ�Z�>�<�g>^�q��b��J���gYf�>%.�NJ���ߌ�ک>�?F&����#��'�-�E֙q|�NK��ǫ��J8g"�����W�ί�|X<�f���0�ǝgV����g5?��WM�����z �xևJ���?�6>h�|��e.^���t�1f��?E?T{�C��u�P���'�'��t|<���b��r}��"��b9�+�����9���M�^�ƱRðuD�����̿��]����
�@�3�tdS�1��&.j�N�g|���?=2���58¢���I}�ە�{����K�F��2���o=I�6�}��i�4�Pj���]AD�o�[rN3d~�7�J�ߺGʊ�.���-ݎ
R�8����0L	b����}�n'�̄��mL{ZUvI�!gN�V%/�S"5OH��ّ�-H7��f�	q�쐞�.�:�l|��&�l����ό�%*�!�P�m���jE��*�  /9P��QG�?�4f�WE^���ŏ�wi�����м	�:j]ǃ�PGA�UD��}g���A[��5�c�u�0Ks��oar}��T����,e�q~�c�dTl��hy�u���ezv�NX������p��(ݐ-D�[��/{{�,r3&)]}�����u�� b���{����;��ӏ9����ԫ�(�T��_�\��V|�Ѣ�_NiV�*{�U�6��4�Qַ�Y i��I`��������;"�Ā2I�����'��H��9�ŏ�pe���k˻0�Z5ch�(�r��]���مE1{�g�ڎى���2zj�zI���i},�ח� ���[̨x�;�N��ñ������XR̪����%|��)4�n�x���?�'s��[N-�nh��<�ͼZ�л��0op���t��~�����%v����1�H)����N��߾!��\� �@�;gemXX���3��'����u���l_�����]Y�o���D��ݠС�Ѻ�i�lX�squ�Ǒ<AUmE1�߰c�3�= x���ıҮ� WB�ٕ���An��DS�䥡VO����R6�,~�m�����e�M���#to�t >ڰ�W����s�W5$[�sCC�;�Cb\�}D$�|/���8�9ڇ}0�n�.�'���
fCC�M8������
p�:����C(y��X�3A@UU��KlM�J���l��Q��K3�\��q�V��Ȧ)&��P���Z_�O�ul̘�j��PV��ù�ֱ�7:4_�jN�q��5&�4���dl"�T�"�RK����y�+�� �~�F��G>����_�e��D���byO� �#�n'Z�Z����}{Bբ�a�l7�� �І��Ij�}那6Ͽ�����9�"��_����]V��������b*N����q����7�ɀꃓѿ>q���GA8�B�<;ml%���sEw󞂾S�pĦs
>��\�Nm }C-�g�DV�*G�܍�1
�6��W;J��#=��`�}�}��qC?�:��� �]� ��{PW���
�� �*�e��gzx)*�ڡm�Z�y���|��gN�.�Ͱw*�y6�sK��2��+���{	g�j�utA��g�	�tT�?�j
����x=��t8�b2A�WoH��l�h{��3� �.#�<����,�}�d�7��qr�[�R.m|Gpv�(�+ޘ��P׎ׅ�Hn��m����Jn�}��	��*9�ݴ�:�����=[xj|��k��J�p��dO&o�iR9\_���"gL�b�H��=����W���.!9pޤ6�JyE0Hsݝ�W�l?;)�N:��l�6ô������݊��� �� Ub�^���c�7��J3���C]��0_`�\T�v��l�i�弮E����@hH��A�1����e��!���s����.���M ���7�ܵ���¸�w�p�SB,s���_����[�l�t?��-�����(�hE�j�Pt��X�|�������s5⑏�!��1��`
pe�xA�3fZ�2�EZ�����Sn�/�Nv;q����揢��R���`�f���1�p"����mt�?A`�j�w:�_�~F�ǋm�ŀ���?�o^u��;R>�5�{��qN�҃#k�+`��^���Ur���������]`�US9�3���b�Q��<��-�|�9�P9i�fx���iV� 	�R�8S#!�. ;�]�w��C��}�����s���G���5xE�k���>����v�Z�v+-ֻ8ZV|���:�$/�Y������� �Ra��k��	1LB�����ᠼ�@���'15�|bN���$�d���[��?+�	Io�B�꧐rr��=fY�� �7走"��Z����T"a�ȅ����bLV����ۑ\$��ѣ �vx�q�J`E��N���_� 썄D΍+Eӊ��U6�������K�����?'��Ż2��O��n�G��l���5�"� $�c=!2
���eoW�S�Ŗ��#"��o\9	��.�ȝ�nv�em�(Zn����1%��g�|�p!�#W��6��&�a��W� �
d����A�>�b!�rYI��IWX�/ �=�Kdw�\ 6��Ƞw�z�ur�^(Tk� �QW�1u=�P/�۾ d�P*��Sc?O�.��K�8�p�8Kv��#���y�B���.y+������
�=f�k���U\'�g��DL_za%�tS�2/��Ѩ���&ǎӭ��c��e�c���؅��8?I򚷐��~�f)���nW���|�����ep�+�XX�������B󎞩��辦��q���v V�r�B7\���x�7. Gf_��}&?_ ��<ӄ����r�Wi	ӳƆ7�˻Kʱ����S�A��"=�lϻy\������7O�&�Bz�`IC�_�=��P3�S*���Y�@�b�X�
{�z�W8�#Z�Ff��Ĺ|ү�G,߫��*�;rHv���>��&qo��x@���+��U��㘤���5EE���z�9�bֱ���wG˫��S��X��
��G�s#N�z�[|ס�nrv����~BX7��IÈ���r�^���{��҃�������Q6��y49�[+��B� �?�E4�/i�K��xQp�;Y����q`^�@��o��X������WÝ��#��y�2B;������yM�Ì�y��
�ĶO:�L��ۡ�r�n��G�u�ኤ=��O�-���h-�X��}�6f�M��{�Ϋ+��
�j���T�ݷ����N����v����/��*��\1���/��x]��Ȓ���}��~��ܷ�?���ck(��@��G���t;̝��a#�����RSv^1X;��&>M
X]����s5U����\�w��ɦ�8���+2C=�j\F�H�4<�#��3�ޞ������6`�
�>��o6]8�[�z�-:�w&���P���] `�7�q 	�����mz�q6d+@ c�����3�\��a�h�������k�ʠ0:G�X~Ly{f��<m�:�X��>Ӕi�Ӝ#�&o�w-TY�<t@��=Y���F'Y	��<E��8�&WK<�*@����s�S���E�$�Q�PD5�F�v�VfY89;rC�L"���G�`��e�Y�v흣���f����tܞ@��T^J\֮������$�R"(%��p���������޿�D��v�����)�pՂ��A�a���[�,v�z��?�歵���
0V�̣��͚��ÕF\�]�)^�|����w���z�ۼB��*����'���T��v��7�lN����/�%M���p�(���8aT��Šw��&`���m&��!����p�����"$�:��[u/��Q��Q����������w\����X�P�]퓨v�E���(��ǅZ z�$�ǥ�����W���Š�eޒj�_�ش�*�O:��@�W4��e���}�������2?�#q�a�"��T����I�n"�9yY�A�9��O6�V�-$���LQ�����E
�&�� 9�M��3ԡI��	P����8:I��s{)�C����~z�U���r���Sz��(WҘ5�7��P�@��#JB��S�t�Z����7���\�$�^q�|C��ۦ�|#�7g{q��+�y�L�:}�Qv'��o��k/�p�<��vD��Y&jaog���(�R��`������<���}TS#���OrB��q��&]Q��"�6��N�2�G�u����dl�~B�0����[ţ/��_�����Γ�sZ�Z?�3Y�����wt����a}$����}�ӊ'|:~�[���H[8��W��g���a���l3x7ƫ�2 ����d7�&�e��OB��3b���67��Q����'N�a�g�N�U:i>�gic8G��C�nXha�}�L9�J���l��c�;s�1�є�{�/��(�X�w���.@u���9&����Ƈ״|�m7D�7t�
�=2�/�_�;ܒ�/󾴪E��c�Y_�}��v��g}�r��ajfr�M����V�����g�m�� �g����}1�H+{�SZ�����Čo	��tD(K��D��,�c�UZ�� #�ZLI,��p̏�kNM�|���3�۾�:sO�����p��,��CY�#&��{��_ �t���c�B���sV_oC�?��B�2��ʩ�1	;&��RKħ���5Z_��&����͈�/uo#s�w���rp���e�I�OJ`���Qyl_�.L��?�����&. >of�*���SwT���N*���|^�ꎯz��߀��了Oɿ�Ri��`P�K/�2lY�YS:@[���Ә��V��� f攮���5����;)}+_s��d��O}|p��J����Z�@�a �){�y�ɢƺ)2h]´�|ݭqBZ�t�z������0.�y]�s*����\䛀Մ�Eհ��>���F�~�w��E�A�,|N�^��N�dy ��| �Ȗ�X�f�w�-o[y�_/!�KuUd�E7a�d����)3�� k��p��_���;"�3:�A�@M�"��e��s�>�e�:	e>�O�K��#�^���f�f��G�IC�����O��E����<����l��bg�1�vyF������Z�E�_�Ly��l$Ɨ�{ztb�S8��pw��e_V�i�؎�Y��
��1%�T�|��eM�-u0|���k;�1^	�<�ڔD�g�>t�]�.Dn�/(��EpV=jg��GȈ`X�`��er�+�54�.��:���V��o*vRac��`v�v��������w^��8iV��v�)�������c +�>}q�=�m���ό�<_��;"Z=��=ӌ/(�]�ܟ��y�����uķF�ƛ�J৵����������_g .�uko�I�0�,UYuzTg+����g�W����6���DQ��$��6�+�#���VdAp�/ٲ��5��
O7v4Ѕ�<ƔQ�V;1~�<����������*F{���1i��KV�v�>a���;�$����
�Uz�S�¹��ԉ�#�&y�=>M}T���2�,�{� �]�t-αmh�8��}������6��j��s��|����N9���9������j:���7��������m��i�|օjgv[W����;f�#��J�;%WGF��C% �r	���#��ߛ ��@��h,l9���9Ԥ�i�^c�m�J1�Ɓ�6{�7.Z�$��-8�	w� �>���U~@�+|�m͛�G�� sS���B��s�{5������@�A��x'}/K�.�*c�O�i�0��lP�� _8ʆ���X�3q�_�}i賯;�ԗbK��O;�99������lrB.�tN��'�8��". xwse핂�p�~c[�%P�"��/ ����w+r|6�*j4o� mZ���J��:(W����~�������K�'ư@�����y�����}a������^�x>]�#]��H���A���:?a�W��DD����^����"�1������V��>.�m ��ڴ�NP�l��o��}ʊ�����i�͜���JI�]e�-뺒�_F�cM�5d�q�uC���b���]�1#��v��*6�w�j�.�-���I;�o@8�J��1���`����g3���,1/����!Q!K�Q�#����,5>��h����J?|�l�`A�^��������*��H"��5���3���:�LvD��oc��,i[�����|�+�w���̀�Z���R�.בd��	�a���2����h��!
�|��g�[�}ĊA�ü��џ���O�=-����[�O�!�<�JT�_kh���I����|ƒ����͋�X���ף�立�é���$7ͯg�H����G�� .�@���@L� �����Ȅ}j���r/�9���Ř���#ʞD���5���u�Sy|�1�� ����C
��T���ie��W�����\��g1������r�u�G�w���x�쾿V}>����i�@Jz�k�dP�����B�����,\f.ka����Y���#	������d�俚��h<[��仗�<������ `�s�r�Y�ű}�*�&0��籉�׉�P鿙�s�}XV(���: �&%�MU39Mǘ3�"���n�Dp-D�Bo��ٖm�{,`ߠ&y7�2��'�s���&u}O>C0�m������+���5���gV��ˮ����\�\�q��[���lAw�t�):Z�A�"2P|�ʳ�}�y̽оs��P#�I�xG�Ϭ����\l6�M��^ 3�%dH
_/�:�?z�7�d���F(nn�k��.�9�ղ��%E�n�崑�~��<�40��3�զ6�k�a1-������XD����
���u��������L�'wR�`��$���H�P5��I�@�`��p������uպq7N�e�t͎-�߫2�sk����v@���0�N���	f$��I���Be9�w|�e R�/ˑ<��.:o�_�zҗ�ƒ�U���g�+cԸZzƉ�ZE[#�u��?��_�-�6�J�
��:�6$*�>���]b?���l$RU���+�8�m�N �c6E������0w����c}~I��F��Q�j]�
8�����RF���UCق�� ��3q��ڨ����k�p3�QKb�{#��溜��c��{��ѿ���W��'6��&,M��G�.��7�!�k�pM�g����)���Vg��6�����k ��'�[�W��NM�N'�҉pR��y4;�aom���xs\f){��­)RςcX��b�M���@VrkS�?^vf"���Y[s��)��:��pW�ky����#�ó�J���#����-�jJ+:��o|@��+2�ԲĢ	�U�u�נ7d�b3�!+E���/��L8�s�P.�X���6��\�Qx��>��� �����g����e�|��q�"�O��6���~Q�<���XP��F�%3��Rsk?�B����*�?�g$#pU�	8� �5�o�V�SV����Aw���`��߶.�p���SܲK��)��/	w���q��M�'��$��.$�yy�<`��Bk=��;���~�4�T�L;���[�� s��y���HF�m��t�~�+��٤��&�pGeO�u����7���է2��.ߡ���潹���d����������6s��Zbp���󙣊T$ht^�xC��=�;Җa������敾V�sCѥ���L3^�ׯ(�z��vr���M:���Ԅ	:�ٵ�sWG�5��a'��t8��g��Ojt��-��y�K�����c���,fkV���k]�H3L���GU�!~l�3��S�ޞܶ�7�X�!��m&�JoFz	��gu	��\H�US� #��,M��N�yTL��;�hYQ��Yqm~����������q(*��H�a��|�����x��q���P�ݞ�����Z�Jʛ�!(Fb��Y��Y�~4h���κך]��߇ۓ����� (5�s��� xi7�\^7/C�. �L��;'~?����˒�;!�D4u��X݇L�<;�;&&m���.mYw�I��j��c|�!�\�ؘq�h�3ѕX���:O� 2P�}��De����'�g��gct�9���F߰��,�����ON#�Ž�_S�=����٦hc�&�S^�Xt3���h��J�k���]��2�B�����R9G�K�7�f|%{X���1��{�&�A��#|:�9e�K��\�&�p��PQ�hc�9J���B���םh�������J�?U�W'{(c�A�?�.81��h�]��0II����
zǗ���{�s�z�����E�W~D���O�Ԕ;Po��s����"Xp�À,LQn&�p��H�)�������E�h���B$Jh��A�l ���X���ɷE&�e^2oy3��m���g�_(�#F����獅Ϩw��W,���S��D? ����.S}�2����Z�B`��Z�P�k�m�J2 y�*���o/l�|a������������Q1&�`�`sT�f���l��
R�����y& �hT0{����j�f3��HƗ�p���S#�Ր ���.?��Ԧ_�i�^���� |��0Z!v�$S*�g��Cm��rU菽�(�G�=ر�k����t�4x%��*�R_ɤ%7{El�3�i�a�M_q�5�4ퟤ���w���=}uߎ�=Jϰ$4�K��u7��7���'c#�x I�v�`�9�3���uJ�¿1���'�1�'�\ ~��w2|=Q�&�i����y�@�t[�Z�v����̼<Q2>�i�o�[��B�rg�r<R�����a��sqa�{�����8���kP�b,�U9�榖1m��@��,g����c��n�w���=`��nQ�fr@�)[��k#��_�>�Gmk�6u�I�Wz1��5�Ԧ���Yb��>��1�!
����V|p
JkӴ�<�A������Rz&h�W���C��uS������c�Ads�=F�ش���T${I�j.[���x�I*<�6j���vl���gƿ`qd�@<�� 0EO:��(�3Q ��E�{l�'Y��� o���]br�x��L5���K󷟂�ZI��F�F�`"^Sܸ85T��sɲJ�V�gEAh[�H:�O�k���`�J�����":B���^�Rm�&5�!g�̀��$ʄ��E����7Q�a����ܕhys[Ɗ7B�Z�R�i�����9S��B��gO��B�I��v����q}oNΥ=�r)�i}����d+S'��C�.�H�L��We-�������9fh� �F�Ms�gA�w\�ZMU��[��/��OtǢ'E3�@�g-�1A#%�sS̊���?���D[���CK�m�N���nv�X�|+�\��}�c�ҕo 
�}X�4�����w!�$�#V\3�I�������M�,�h���Ǔ��'n`�h��׷c��������W��򋳴]��>�ew��8#bcL���!^�~��;�O��h��x ��bg|. �^�A��
}A;��dP�J�Y�AH����N��hGX��˺κ�Di��|�s��!�n*n��kL�9��2�܍꩑�ÖP��iҮ�^]�v���T�� ��yç�r�4w˵՜JE��z�C	��1_�̋m��@~��#�oCR��=��*�=;��W��d5��Iv��?E�����΃�j:�2�!��D��n��g�4����DO��j�B+΄���İ*���E��4b����v�)4o"��Ȩ��.��n ^�d�!�W�7`!?�Cv��4��k_��	���	NT��Lfʧ焤�>i
p����G'�^w\���7����w:g�~:���ߠ��������%�O�޶�t� �F����Iu��D���:���z֙z�j�>�D�#j�
\�(K�f�1-�Ǉe�ǀ����ڒ��5Ϟ &p��N�1Eӯ �;��_e����G��r�JJF}T0�P��?�\� W��,���aU����U3��k�Æ�'�q��h�GBx9���}ʓ�}�#)�Q,�,��`�-ٿ��/��>�lt�Y�~.��r��ad\�,4��h��V0�ѾĤ�����91�O�f1Ɛ�]�^��}*���@��;��[EN�]o�^[. T>�HH��}E8$��i}��4�f��$�xъJ�d��F�$F�ƊW���N(LL�܃�i�@-��D��#zH��p�LR��31,��e����&&���R3�JT:�Fh.�웲�e�^����`*�6��o��v������t(#N�����a��b�/V�)	TKn�X(����?'�똌��Ď~��;����f�S_�ᭌ�6[�)̼�Hdŧ1������aŲ��� �z��V�V���I��~��e��Ю�nx
{2f�6ڋ(y !h_�~�h���t�5����8����韟ڃnTw_2.j��I�[���Z�]{Zmu]���^7Fr6�Ek�ɪ8r �'�Z�^�̳=��9G
ng8�%���WR�G��Cl"e�}6�@J�9%1W+*9]e%�7�%ő�턀�3�F���j4=�.\(���39Vas�-�P���7Mj�3(�y��0�Z�i�����n\�V�n��r�:d��I�_M�	?�����Ld�`��q�m��p�B�fq���zTii���~L�buu�}�fj��ޔfHϜ<��xL�&�Zi?F�XعCrW�T�OŃҦ\�7����D�Q���3��@xB�k��� f�c�"�AY]�qȷ���*+_r���[��^݀әBT����Y\W�/@�m�Qu%=��� �P�;���$q��p&�ڒyc3ǵ>�f�֭Q��,Ih�bqc�f�­��}X�w�w�M���&�t�VB�|�[�o�4_�T d�|l�J����-����:�v�}ȝ�\69�c���J������*BE6����3�������$v��g�pM0�����3!ώg�ռ'�*v��ƘЏ#Y�����Q�X�]B1dXp!�#<a��IB�h֎@����<"+� �߆R�䥎����be�Y\xS|�ne�ѫ/�(���b'?� ���~уy���q׍����c�Ý����Jb|�;���?�X�g�7�S*2��*iO��j��4�`���AUm���>m�"�
e�z/s� �U#��qw)�<�o ��&m3�I�y۲����Ty���&��i_�w�B�ѹ�H���B}f@卸m�ڝX��'�b����u�߷R��{�!�X��'vw�p\��	��K���}T�,��#�}���1!ϔh����>�x�M���*�q�n��3Va�qSaX��R��m}m�*5�,��֮�:+0��k���~��� -�����Bk$*����͒T\�]��L'	S�Fy�F9�~�ް���j�q{����`eu�zS�bn�����Ѵ2�Bݼ��&�W�����{��ׁX�]Qf3S��{aoG�#�Ɔ�);������>�{���#��w�����vL�\};��ܗ,mhh������� O'臤d���M7��D���F^M�:�P��䛔���'#����s����{��5�\��>g��D����kb*FU3AD�M�y4넱��s�^>��Z�۔�E@N��k�7+�{���E
�w�����p#d�r�e%�v
&�r̻h�kU�e?D:A!v�Y�ɯ�:��3�����鰚�r��P�/�\�[���+�g�z�Hg!�Q��� ǻU��A	k9s�o��w-`�D�Xj��5�2�`S^�!'|%<��p5��QH����X'Ψ�EO(w65/ԝ���͜��k>�P��V�ћ�y�٣ٌ�I����%_�X�Ȫ}{IHb�4|���Oԡ���"L���<�E\l/]��d���M��ۆ�Γ[N"��^Bp��EHE	D��].�%��_uOs�(�uP��H�i$0�$q�s�nh�]�"͇#�?_6����4Fd�/Һї��T>��W��}���a���I�4U?��^�,�,~5��cL�����c�Z� ��:�~h���J|���:Yv��xu`�y�{Æ+��:y��!R�nw�S�:�Z��\��Qw����_*-"Z<Ģ*�a������l[�XDlցvwTv�&z�?�kQ�L%B3�o�*j+�=�.\g��.;D�՜�o;�}�y�x������`�)����f�&%�u�hVA��������,��(}��zL0/��"���4kv�7���b����)���u5b�ɈN�8$�[
#��<��g�;.˖Ȅ\d��
�=�{q�l������J��*F��賄�ٯ���,,vr��s���uL��*
FVj��������E�!�.������{�"q���Hb���\�:A�lv�l�L(X��}���:���^�p����ፘ_jj/v��xa����ȶ�nG�3�1/8�ǳZiĲ�v�3���>���X��N9[�mE������!���|�z�|�H�t-���9�:W���������+���������}�<��'�o��w����d8��-��-Y��������!1�ָ���8�#v�Ky�����g���{!NGr�g)���� -��YЩ�{@���Z��"v��9٧V~=Pe�E`�����/ =��C����W�|�����o@���^�<�ă�j�Nni�� �. ��T�� g��)�*�,�FU�,�����'�g>���ّ�,��[h�]m�33�����s)��]>�,���2��ؽ�F����}��6�Un�O�����NB$��JZ�/��h�#JU���j	��1����M��[�(d�#-���e ��3އ��G���[y�Q�W	O�����Y�@��+X��s��t��
�HR�o���ՙgx�޲�]{�˶u�>�6�L���G�������4��qM~�3E�J�2A�fbQRҭ�tH�`_�.	��{c���!�66r������{�?�?>��<�9�S����q�_��uXu� �7pV����~�j�� q�|x��u�O!�VtuwP�6����g,�h@�Y:M6f.U Y1p˲�p��-���dQ��iH����G�:�?��M�������E��o'��R���A':���'�1eG"}�����Gq)B.<�4 �N;���zn�ϨU�r��M�6���i���6��j��h��lő�Is+P0E`!�{�oYh��IN!^�(���Q�
�����b	X�M��7��s�_Α�M�*�|��^3[/#��.�i���i�-�=	jAfv���ī4�FԬ������wg|������WE̖�BTFL�v�)B�J|�������E��`3��?�*��*LR�|tG!�D	�
GdE��1Lg9�\�>[%�А�i���P;/Wn��5���auQ�񆜛p�
hU6�rؘ|ǐ}6��y� �Ad��LaId������ɜU�Kp�N�@=���o�Z��}%��^5��E���O���.��u��,��"���IWMu�<f�����TR [��s<����@}�I���%�7��l-2FA�<�c2b'��7�X�cl�@5_����n�'-ϝ��U/�4��7�|�B}��Ǻ����s���Ӽ��8�2�h`�*�������H직O�M�S4ț\$��{6i����KR����2#".��x|	�	��;��2c��笚pn�١ǧF߿˓+i ���CI���`4D��×��:���!����.P����z�e��X���ZԹ��qg\$�3�{a�9���)ͯ�Ϳ~a�D�y0� �to�Uc�Dd����)�+���8�Ĭ�3�lS=�c��g%?�����Y���OΧ�`���bW���Pw&� �,0V��HXѹ��}7�J��@%�?V�/C�*Tn����L�̈́�Qq5��D��6�y4�<,u6c�u��\�c�>���<�Q&�,�g:���9�w�԰]�w�ӹ��La���O�f��N���2s���R,������{��TڒM���8���-[���	5� a%�3y�M��K��=C'�_I"��g�"�U�����{_ӱ���� z�'�z~(�������cx����tC&��Z�)��r�Qx�~Ow�K��R�wV��i�����>�h�w�^�y1�Kp��v6_w�V�T=�Cȍ`Ț+4 �5,�0�2q����#�%+!�Uwn�}��So� �(vʒ����V�����
7p��&/�Up��3s��݆�@�r�o1a�p�2r;���T�3ό���n(~	. XE)����6־G��A���o4�1���V��1K16��5��������/֞��V��ܨ��]�xnt*պȖ
��3$��D��E�[�L�NW.��
ks#4�����'K��,�n U��t����i"�DԘ���v���
@|��iѤ2�#~(۰j���#jțy���'K� �!~��% ?V(]���f��w�S+�uĽLd~ܺ��l��~�{�3��.:���IY��b�6h1���3��O���; %��F���+t�_�6>�V)�B�C�!��ܮ��d�����mw˄�����Zd�����8��i)���EV���"k��U享^J�sַ�-21n�Էϊ���d�WN�+as��G|���b��K�f'��	\��X�7'+^]�a4�K�M����mk5�R���Ox�ƣ*�� ��I�8�t���8�0��7�_�[M�� ��`�LaHj��Y�� s~�Rf�$I�5M~%���4TM��~E$.�3?tyU���In�UV��+�;��L��"��wgV�\9��om�j�v,=��� I�#m��O��b���I�����1��qI)�mP3a�m>���������FS�h�\����~��Z�2'Q:�RD�0v�淧߫^��yЅ)vy���0I<K���jG3:+��[ȎQ�Ž!��o�{���O����Ǥ��4%��?D-I���y��]yi�"��
��抛�>�v����1��,��W�j��ZYv9�댦Da�i8�N��s˟s�q��r����*�Fn�)���{�YX�p�qqq�q ����*����JFē-,�g��C���³�S�dA�J�K�IJ��O�Va�Y=��RS�x�_�����HD<"��l �������ɝ��~�h��3�fZw�آ��yccl�f#�򱏗ǻ���P%m�N>8cJ4 qz��%�1I���N����j�l�Ӆ	�*m\~�{R���S�5	�f�N��}׊����ON��)Bv�|���qW3�[�R�v凈�j�}F��n�L|�	�C����%����S�{'~��z�ډV���ç�����-�c�(�"`~#<�7���4���sO���ha�E�:t��e�ۖ�z�ɒ��k";I�QP�S஝���)p9�dq7����6�!�g���ʾ)�K�@��"k{+5��1M�2�!^�ٌc���R�[N��ɏi���\�ot^�kiv!� O�=�u�iY����B���^_?�]��]G�ډ��]��V�����=>ώ` \����L���Ͷ[��n�*��U��d���>F��7���ua+����FJ��M��VزBc��.��ކz	��[W"Ź�+�Ċ��U19���#}����4\Q�|�6\M��*�$?��@�i
,�6��5,E=�<\�Z/!ٴYm����b�Eͦ�jKl�zo�jk�pv�e��m�2L"' �dٕJf�BL�	>�J��Z�N�A%вV �h���M�'"���/3E�2?��	�E���͒��|���`�4����XBO�+J&��`ݙ9�n�>�;��N��{^��;j2Y��8!A�Z
�l���.�o�����0�
%i��I 3����k͸����Q<n��|b<x"��n&D	�"o���H(�	a��(���"��N�R��N�p�F���,��*[���^��]]�"w73��Ք6�v!�`Ō`}^��cey��|���֠�6x���~�},�������ot��՛�JJ�Ev̭<Q�p�E�_v�M�	�y�� 5˿��X_�������(]1��Ι��?�>�����j*ݼ�:(;���cC�F���7KCؑ.!����Nf]�#�v��`I�N<؁$]�5�����'5��z�Aɞ=��5��Z�;�P9��eu��d}v[�{����ʶt�j�6j�k��Y[����������Z8��\q��TnZ�_Jb>x�Zm�&&"Y04@q#7t,j3��K��A�ї�W�cF����ռ�Tw�����#�|<ܴ��.?_-�c|şW�l����u����bo�3�ӂ�|9zCԬL��qd�Foo��Q����k�1(O-���,���T�Z��|�*r�j�n�hټ�Z�0O@g\=�X��!��n�$Z+8_�2��6+|��}�R~ۍU1
1��V%F��7����v���T���<�x�G~ [�������NUv��n]�b���`<av�f��%�D��c13!���$Vp���P�"iZ�a{{q��&
���g�L���w�w� �t_��c��pC��ڀ���.�m��a^|�q��|�4T�&�'��R�ߕ�{F���;��[�m(���Pȩ��n�N��~�0ewJ����C?�)p��t��:���U,b�9��9��grY����7��6_:0���Z��� �w�.�5����L�^m�6}���sc��0�,��(��WI�<Q�8�d\N���
/R*�r@I���o��ef�UL��*�%��R��?1��Vg���������x%�<���Yx�dN��&?".�PdƝbշ\�ܙ�K�?ʵ�d �t�5e�ο�谧��Ӑ}f$���~�q�$��gOfa@z���M�0���Eڋ�Etq�*�hUo]��ՊaF)X���#o�K�=�-^��g�ykON8�8`��H��'�P�6�6�m�߈��R�<�>��jBe��Á���7NK�̬��z<�������-�K����J����'/wו�taݭ^?ϙ�sYð�Y��C$p���cI�v�ߪ��|�Tw�n.������H{�s�o�i�p�J�!�,\kp�r����&��cn�X��,#l�b�Y_��Ϝظ�6�m��n�[]�V�����铕��c7�k���7���kA[)�%�TM͵;v�%�\W�N煦�O����{y���
o�Z�-�����M
:j�H���{��`QW>�iq��l��drD�~��μ��ѝ��F��c��Js��G5r��L�\�E���&޷�G�J)A�\�	év�[6������a�2�����&�6Q��EC�s��:�q9䓱���w���H��s����<�Ʒ9N��y]TBUO�c�B�R���������p�F#���7��؞?�ys�Mдty����{��&yi�n�ʐ\#ݏ���&�JN��_�c7`�w��5{��([�%�|�a#��i�y�R1�K���$�Ps��Ϊ�df�"F��'�k���l;fZ���S�_lZ��
R�y=k�g��mNg/wd�5`>���I�R���3�Y�̓���''�x��l$j���TW�����"��9��}� k��WI��.�s-��48�8���9��`nf��1괷��c|2�>т�:,��8�����vY�q�\�κ��u4�LX�9*,�(��C�M.��t��T��������k�/�������<�	�� �C/���r� UG�vH�k����L�H,�^�R
Ddgt� �����H:	ud⋣�P�9sI63�b�/��}Vw�l_Dcc���.��y�(
�\�0])�V�99���U�l��:$�}o3z��pq��ݎ�Q.�G�g�����t�D��zy�E���dʴ/��/C�V����C`�21\��:=�p�!|u�G�������z��c�~��u���62h��������m%��Qc��㵼�	�v�]��S�"��QY/�������v���'J���֊�_�����K�o�`�5̵�v���%��%�D�Տ��>Sv�v�FT܏.���b��@���t��Pv�E�`����/����c�I��^�2�A�2Ho�DsU��6dCG$h������+>O�^�\����\ub�)@=�&'�>��2��ب-��?�����(�ؐ\ڣ9�7&�bu=�/~���4Tq��SOX���;�����C���f��L3(�K�v��'ܬ�w�L�r�n|��e�s���PY(��3c� ����DH^�ct���	eNd1s�=|���-hy����u�Ռ�G�:ww������R/|x�YE}�ަ� �':Eq��?0�D��C��T�x�ۑP^�X��±�ic�錌���ٸ�*M�~�E�Ξ����D��k0�#ih}�P�l������F��űb�É�4@��;�CL��!7��h���`%A�:�/�VȆ��g�S����&p�\��S]} �o�F�oD눖��D�޶���m
*|�R5}���>�g�s�]��|C���o���e%v-=��r*�~��9���(��_��;��o��D>�ϝa�n$����8���?Ճ�� e� -������pb�@�Fx��[��z��ї��Y�7�%�֔f5����l�kig e����c|�����_�4@�icÄ������	��D��x���Lʕ�$Q����{�ģ�1Y��Z���FH��*j*lzJ��Ǘl̤��%Tf	�r���(���+d�$�ᣱ���l�6�Z�?��MG��ev�J8>�7�r)p������!�KV	Tf�a�RLi�2�W�l��U����>u�:���|�jZխ�7�ð�[���p�e~ϓ��s�U�c��\��=���q�mZ-�ϓ��H�a(T)n'\�-����8��on�#�W�evq�U���lK,��z*�Y����Q�O���q����O ��/M�����p?�h���u�����'u��	�4��Kw]���ρuj|xe�6)�/Ҏ3��'��~�>��W�{$^�$�O�q|�;>�	�VڰCPg��#�X�L���Ħpp������_���l���qH�_/���!7 8S�K4@j��W����V�:^��ʟ���?"�i��+SC��6}(gkϢ����6O���ڄ�H�%�uݤ�Ѹ��ҧ��g:�5�>��Q���±��W�P�ã�[��ƪq��gw�'d'��K�FQ�՘~�!Ih1d^�0��J,:��Q��H�F��#w�VA�m�ݎ�6�p5��r`��Q��h�Ě1�+ ��@��o�W��X��`�IRقep��ӽL�� Ϭ�tuo���F�� �Ֆ ��;��N������e���>�3m5|���_� �2iy�����O^��F���0:I6S֌h�in(l�c�>R,�[p��T�2$f���
'Lu9������?��<^�^X�ݒ�Mُp(=�i��HE8��Ud�N8��=IuZv�H�[���mw3'�U���YoZ3=���9&�o���/#�-���$�$A��q�v ��	p2
%��E���� 5�1�M-�M����}nF��.�=�
��Y{��$�k�9e!��ߏ�o����t�c}�g���o�{䶿��'��L8]+�)^�s&����[����Vt��F\毗f���~yd�
��u���w�!V�6	�H��9�D�t���x:�ϛ�9�/�y)Į宲s�J�3�5�L�\�"]�إȤP���$A��~s1��E��2����5��t���:g���.eS���"J��(z�t�dq�ۡ��_�� =����P��)���1TG�o>'WO�;O�e�woI�>�A�I�xeu�T"S�*�޾H�_V:n�۬e1I��fjLy=�n�ӬZ���!�d �%u�Rǹ�_ m�'�(oǻ� �A�ga�zǩ~ e�3��3�nݶ'F\_Ǧ%W��'�4�+4�}|�����w�B��Z����5N M�3V*ߔff%ɇrM@T����pw� 
�t/���7r����:�׫�,I8^M4�_��d.��TB-F��n���:�*?o�A�VA���f�j~�����l4�Ǎ]�ހs^���ٻR:#��W+���]�?�sN},��� ��a,����L�Ir���R��m���.�U��!4ć���\6�v�#`���WD%g�����5S�����xE�`���C��d�X��|���� Y��x�o�V3�.�xM,'C��o�wз8\_h|T�K�%��F����xTu`V�LeZ2�d�BQ�o��Ę�
����J��|>�Ԗ����vS�4֭#��jAMQW~�\yv��o�҇��!�o�
���c�:ys%IY7$b��fn~��b�q4�Q�#��(b��K�ԓc]�n��Qm��$M��@��k�����[�h��u��@Ųd�׬�z�Z3C  �P$?�.�?ö���3me�yJ��6N���/��EOj�;�A*T��p��	O`���h��m�qˆe��r9�O�G�
ˍv;�1���AX�A�Do}s�C�I�at�׮�얙���M�u��W�G0p�������b
V%�ļ�gH�^�kC�΢�e��p/u�𮙓xa��l��@ʁ^��R�.��|i<� ND�$�j]�Ĝ�SaNo(=�8t�F�.��V�+|���|����X��-�i �&/I���Q�9م�/�[ K��`��:��#[�U�(5�ENÛ���X��-��e�{��Oxj�h�©?�֧c�No���\��7 i�ڊ�O�xETr����Z���I�M��K��(.�:�x.�t��)��j*K�u"��Pv$���z�tr� �-����3Vm��s���6h�x]S�~����9�6yy�z<A��)���5RI����_
ع�7�Ws^
�|6����ˋ�y�tx(���W���iߣ柑��x?�W$CQY��B䥒#Wi����gFV�~��K^�����~I��_h�cS�c@�{�mh�Ru�x��SA��K��D�,�U�xB�����͍4 Mq���{��^�%?�y��� ����]����g���xB)��N\�܄�A�^����~������J�F�����4<�f�h=�^�Q�B�3�� xgzRp���(����&k�8��g(��j���ʶ/�E��o��Ɠ����	7��EƓ/�I�i8����9���(�@�Ö�w&>=%���$�E���NG�h�)�� ~m#_�WP��ou�5����w�h�w�Z�r&[��b4�[Y|�;7"�,/��SUx�2�.9�T�?�G����V.��{Pop����m���_��Ȅ�-O֊֯�}�薋k��3��j�c����S2���t�1�����'��!�2N]��QYؑ^�]1�6��3�j�B,�N!�%��ET���l-<g>u�x��q��0�����v���gޘ�)��&D
ג���Hȳ�~~�0���� �1c�;�x:�����йo:�>]��o�_�f�<����]D*u},������g��[����+X*V]��?���k�vUow�X���<&xD�� ��G�" * �D	��U\*ñt�XQ��m�C��Z���YA����2\U���]T:���b�H�<���Up?�7��ė3�_�b��f�ļ��)�1M��hm �i�?��"�F]J{�X�)��)�Pt6K�P�Ŏ%�q^"�α�Jxi�0���2��R"�T*��ey��Y6!6�w� |J>?��?�#$�+��H���j�z�����¡ē$��|�S�u�z6�4Q�55�m
�MY}v�ˌ�@���yZ3Y�S����.ͦ���|��"�m���ag��;�[�"Ky�j==�������f��&(��3��蓜�aa{������5�G��&j��C>��ðU��/%=�/��+�.B��������lg-��ʇ
��H,	"x���(��9O����O�ö���ŕҏ,���r�ȿ�x����ۺzjBep�w��%��$��W'��6�	�1]�1�� ��ys��1�;�wV�������:�L�;)g ���o�Y�I@$������J�<�������ң ք�G9�O�g��
�Egњ嚭�W�o6���N�}�G;���44�<��P@������-s({ �.�U�?"i5�� *���i(QJӨ�[�V޸CMI�c�g'�g�;�_WO�#N����6���gTdY���/6g9�gi���x	��Y�]�M�!z��������Џ��(`M:��5pB	��-E��&J�g�����{
0�E��r/}�n������� �i�E��Nm��=؍�� �I[��t�&�e����� n�bN����RN܀��?W��B[K�]!�H���h���?�I��J��w�E��m��R�w��+B�5]@Û��hS�A����?c�������D,(B�Z*�ڳn��	A����h/��K���z��N0�Չ9��i�� �{�C��3�:���/��{��"��Ty���⃅�Zʱg�V4-�J��eJԱ� �˅�Ң�t#ngimmp�����x��{�_?z���Z�QS��Lg��B�o_Ŭ�F�p��p�D����Tc[�t1��.V�T�M�:� ���,�^��}�J����T5T�0;��ێ����a�>lp} o��!����_%�b
���q��0��.gd�܋?9kaǋ�,r\���;��S���U^��z����զ���E	�=�(jsv�)�o�8���/ �D^��w)Q����DmZ�U��}���']�����@�����m8ϴn����L~
���Uuݿ5�{"���������e�T���m_�XF83ӽ����F��9��L�A��j3��F� f{�ܱr>�����?��K��wK��&13���I���͡+���s�v��.�$�<̣�����+]=�?�)�*� 
,:�����&�I��a*��wߡ�o�c��nH��Y	(��Աo�#T�ԫEᕔ��M+��AS��~������36H��%�i��u�C�{_m��KdM<|�(k�r����󷨏�m�"9�x�~�����>��_|C��9���PK   NM�X�Ɍ�� �� /   images/53a6c856-3ba7-48d9-b0a2-5ca2401e7b62.png|�T\Ͳ:0�M�w�$�w�0�C�n������������s߽��^��kWW�׵�wuu՞pEyIt  �.-%� �  @i$����N�4  M�RLLQZL�L������ �
OTG�P��Ҏ�������I�+hJ�BNU�,(��D��Z㇮�A�z�ᣑ�ҩwMNNy|���z�[����!�W���fS�"_7f����*~'�L�숒9|�#�E�Ƚ����M���m}c�oc�rE��u�M_.pp��O\$cb��@�	��	 �pe��*��F8��G�G՟�C��ئp���Є���!���wb:4�ڜ�(VOj$I�@'�Q㦷aB�g�N[��O�[�	ě�;+K��g�Z��Ħr����3�6��b7:���_$G-CDD���|�"c8W��!�E��H.Lɝ�7L�k��y4���f��0��$ɠ�{#`0��EP@��P^�;�?b�����G��lƝa��!)���Cn#M�rĸ�B�7�슩AՈ�,�Bak��Ra~�B_2��'�����Dk`Q�o��u�)TF0�-�x��o0A^�D��!�Ĥ�GZ9�:�=@M��}y�U��}x��j6�2�*=,�b��)
s���D'�%5�.z���W�A���nq�8����e���T?��at$�͛�V럓_�����A��z�f�PZ��P�{
]�>�s�]�j>N���QM)�T®�?/b-ܶ���±��v?�М�ݿ�{�4���
������5ba����n4ђ DwT�l��y[�l�AV@���1��I]*h�2�y���b�-D=�q)�	�z�"qqHi�<��L���T;�|�AZC&]��'�=� �Z���-v�i�i�I���˪��𡜴t2�p*[��˒�)�+_4q?�ت����4�=����v��=�D�����Tf�7�͚���ˈ�*?!��(���c#�o0�ȝH^��C.x_�����c;;6�G;���l_I��h$��u��Mt�W�M+��@���O��#<:`��� ��?L����|�wX�w Qa�0�Ř j�k
�Y�G\�����3�� w	���}�y�{|D��cfa!wDAJ$Q�b$�i����}�xa\X~A�Rlq!&��c���C_M��J$�(冤��g��$H(ڇ������|���WB��v�M����?Rv&�
>�L�}��]	�Fd�3�MA6�fe��	/0�O�K�L4����-�������:��h�y��rˀ��pG�����@�\��=����I�`�!�`�cć�d�ލ �!�"m���s���r	�&���@��;�s�La�Kv���� \|�r9�M*�
��OUTKaE�;�.�K��G�O��x���>"'�HIt�D�ޒw#{�Y3�Z�L2�c�x�t�l��ڑ���@�/�y}J�t�!�f<�FFF
G�G�G`��G 	�t�*>�/J_T��ĕR(i�֪���$r���ǝ����(&+����IU-K1J�ղN��Q���J�燾�|�������w�y��ے�y�y����'r'\����W�I��U���3ushS{�LSk�_�Y��S�5ؙlm���+�#�M�F�gW��s�*J��3s�ZE�S\�1
�Kz��5��C&�0C(S((q���L�<�c[:Z�֕�y�!-�7G`0����9d���i�I��8{Ⴐ�cƉ���xHy���Ѐ������� ��"a����+�N-����S=�5���J9��cȑ͍60� ;|�[<F�d�����B����fh��~ϛU��98�>�<n5v�È���c�8���XW+[�c�l�l\`��@_[Z�b.WW�e�k�=b�[=\�lᴌS�R3^[Q�n�Ҽ�|ʹ�E�ӑ��H�㤰���l�T��kn`�X�X�X`���A��D����$���Y�۠E2�
�ǘ�6m�J�l}�\����O���ԋ���$�q�5�\��Quu.��
���f�4�U��5A�[燂���%A�Ѱ�@_����S|s�(!��A�B=��
=����]AA�l�l���M���1��!I��M��{�����P�\'��g2A��@�ٮ����W��|� ����Ov���:��B}�&ߤ���ZX�LI6�Tس�Sy�=�#E ��Q��HV�h#5��A}"���K�B�d9����jnlYo�6�q���Ƶ����������	�r05R�9��)�?I�+!(�������<�ӊ�YbO(�e��].Q�KgH#�"Y�[��v�S�e�;��M�B���������W��'��ؾ�ݘ�M+GNǯ��'O����js�wN��-�~NIO�N.JHNZ��{��JC(��٬bBK��"w�Rk���[���t8;fS#�wo�z!N�
�ڎ�	EHV.l�6��]ww�0�������*���D6>��L0�?�ޅ����B����y=�Պ�To�m3�8B�33����;����FF.�{x�ށ�dp:�v\/N�n��e���q0�`�U-�L�����K'Ӹ�J͘�r�~�~�>׷��zec��������*&�?��8G3G��
��ϴp*���!��C+��=Uy�39��ϑm�꜏����M���E���6U����kߚΎ���}�_����J.GU����~/s-�ܰ���Dע,9^�o9��{k����׆8����{�yO��u:��CD�W�pB�A������g�Z��xB�t�4�t�t�w�u�����$�""}{��bӭ�#����hm���D�-mg�����	�,�$�������C�	.]��#pM�z��S'��Yq�k�e�����C�`Ճ����I�թn���E�����\�n�{#��p�ǥ:q��t�y���ީ�ڵ%2O��;���J�y�V�G�4�5�9Z������[�d��|`��3u�p��#��q�:1�M���E�q�i?�������Ʌ��x����o��ӆ8���t�~x_@z#x�4��~��Sd�]�C�y?`u�8ew�p�����U��_w��	 
�̙ ,�}%�7߆�b/4M�^h6)G�>�i=���#����V����x׫�}�@�ӥm�:���OA�~�J���3ݝ��Yסm�������/��f^��9��$Si399 �_	 � ��`�� 0 �� �W���V���X  � ����-�?�߁q! Ŀ��+(���ar��E������I�C�;���:Y�9Ӷ҅�e �Ki: 8��\0��Tп�EKUg9Y^c;&C;#S&w���w��Kژ:���X�:�P�K��/�����_*�Vr�dbv��d�L,L,�(ddd��&f�������	PX8;��23���1�}f�s4gf���afacfcc�����a�l��h�D��A�kqS'cGK{gK;[���Fv.����w��!Sw���d���i�� �?fV&���li���G�o������W����ZC����R�}4A.n~��S�jN��bv6�΂��������Ӥ�����?Mj��&���������?K�fk�,������7J�催����O��Fh��������ߩ������/O`�_��o?c���	��3��N+�rZ�V ��ET�aN�-����
݌F~�T����X�N�tH���֙Ʈ������%�%z���;��:�_8�'����#"ۂ���t�Z&���Or:���S��rs�ߦ��ϟ���\]9�>^��ϫ�UUU����U��<]�=��|��k*��d���&3�)dV��4�45!N�xP/�+dW�+(�rG���'�N��@Z�T"Vm�!�+@tǜ\b*��N�?�/��c"їB0������%I�ᢽL�����;�x��	�ǽ��N�]��D	�b�`9� t�v���F���Y޲���XM���q%�	~=F�2���r�k��T�P�r�E��hݫ�_��XǇ/�O�ݖA�H�i�q�c#��Jy�X1�y*'E9������Zڗ�.���1��T�*=S�f��c�;�����lX'X��
�-k�]�\g����$�OȄ�귪��U�6���?����[�߈�j�x��,��(,�~�א��V:?���@�h@{���;~|�[0$о/�a��N������[����g㋀ռ�Z�E��~ڴ�`��a�F��(�Ǎ5�wAK��d�'sB��T��1L}n����Lci�_�a���no#o��,E�_3R�pPԵ���])��"F�q�@�B�X�,�7�Ԃ:u{��{J5�g�Ç��9R=e�WV�G��@�Ö�ٵ���lT�4�x|L��V��*�aR�F�M�{?1����<߿�b�2cqr�HyB ����"Z��jQ��xC�r���_U���CPx��i�����f2��n Sl�:�l�I�u�zb	��M)�7��:2(�B
q�4` ���1ўy-��w�
'ͦ�3i�~��ش��)
#��?�����
�Qk�|֜dw����<Z�zl~��⺡s<��r����֙����H$,���'��I^kK:�c@.����}Gmej��o4���'�r�]������ �T1%\޳�p��]���[/��d�q��]j��^W�m%Iߙ��s��~ �9�_�?I��z�Ǒ��b�������A��V1�u�>��=ʺI���*&�88t0��8Do��Q02����!�n�b�^���]ge�:�y�$�:���8O��i#�h�Y�F�wh+6u _�<�|E�;�6 ��=H��+��`p,�z�޾��%�V�x�����m gV_��/aZ�1���+���?'�o��8�+!g.�ǩ�e+xn�K��j�y؏+��G����M�[�@r��z�p��0�O
�m@'�M:�ĳ:�44��)�o�V����8wn��C�u0�c�n�L
���73�p�c�-,Vm |G[�$��
QY-���\�2�n��a��:0�*�{}y��/� #�����5����lWɾ �U�/E��|��''��ʥ|�{�\;-�7�`�;���J(R�L���WV�{��x�/�}�e�+����/U����(��#�����_�H`��:��#MM�l+�^��QȋU~��W�泒���k��P�iM��q�����%k4!�8@�㒟����(ċ8)BL��K���	t��_���I����P�|rN�+�4�4�5�۷����R��ucc��y��#��SƆW��٦1Cq�\A���#�Z�~N�Psj\*W��f�����/]����| ʽ���Y*Ы7�;�����]� B������&�1�=1�0���*�v	����O{|Ϳ��sa*������V0���nQ������3�F����q��
��5�*�R�s��)m-rX2E��eI�Oc��9�q�@a1���u@����,�ٵ�3:�T���6��&T��"�:/{م����;�2͵/K`���V�����k ���M��rT&mc3*ܸәN,��
M8ޫ�!�f�64<��g�'k�P9h���8�1�{�C%N��	���lSo4�ã�kB7EP/�E���,�-E��`"�s�.b^�ψ����u��/����[l��/&>y<���~:^����>�؍�RdX�[k���H>7�!j49Y�"�(Gw����y-5�NRk�ڮ��V��$�!^��8/1ߞ���D�W&����T�F�Q���/*|&���\kXSi�h����� �m�1a�H�sx�f�Y����f ����:��!t3T��D�Y �"���wJ�����Z���2|m������M��,��V�D�)Q��ǹjb�C6�BQ�Osj<�ǣ��%��ۗP��S�\?�0�T�4���3�n��]U�}�#�I;�7H˯+��Ir֬����ω�Q٬1b���s�m)��o�Y�#I*��'pd�.>��!tJ��;���#G��j�r51�L��`q��|}0>���v��v*R���;܀f�D8�l%zZ#7��s�O]��;e��V�ǵ�gy�zcmz�H@!ڷ��uX�=!�'�� �U�w�B�y��iy���hC����ėK
�٬��g&��<��������u��A���h�>V�3���E��.S��z`fF�d>
C�ԭu���b}��=�����^�.��T������
��|���kS%�u�CՈ�Q29��$K�X�h2�w*l���~z�������w"����S�A34��)7&�~%�1�5� ��9�2��ң�_�LH�ϓ���4=%�X���+}$��Z����
B_���3��"F�8��F=�M9�bd&1�{X�K��ȓC�Q�+�=�_��!�eΆ�6�SF��*�K��֗�|���A[�Y�-�����60��P�v�[���}��ȯ�6uG$��:��B����N�,�K��@og8]8��[�$]��w"d��_�a��+�%��&5�y��Iԗ�?��rΕ��}Lb��V�LV�X�=�xO���]���[S��qs��#�;M�(y1���y[Rgdx#��z�I}\�*�"��F:�ڧ0pζ�ۑ��(�=HY���_s�~�>힪
EMq�w!9�oLѵB�����jfSo����V��=���L{�ʞ� a5Nvk�Z��Lhcx�V+��L`�s�.�����b��������n����S�`�;��e��ΩلX~����
��{
��N�H����:�nn+�I
A{���揕��3p����񭏫J��������؇�0�Ao�wUs@H������N���	��0#�Ct�`e��볻B��I��=>��$�>=V��Ê�c�K�w�,3�����Y���QB&n�O�������p�T4�8x���:��x�]���h�i������X
��O� 3V�sy�@�W֯�#��e��EyYPB��d����y�J"���o��
�Ŕ�m�A%<��c޹�t�SXw1��l�*�߼��U1$8L��Wy�k=+M�r*�E����N���i����^��;{h����b4��U;��z�&D����V�R�n�׉\]H�S M04��C�7���Ca0I��r�k~4$�Ojc�j,|:���U��W�T�G�K&i�J��%�B��:��5���&����;��Q�
	L���������8T-��<�#6���fi�ύ�I�gI��7�ۑѰ�)����55��~����Yt���>V��ϑ(*z�Kd.�SĶ�s��,���K�'��H��^��H<	$K��P�j�6���-��p�Q�L�`���������M%����m�t�n�<Q��t7��B�f:_D�.!��r~xr�����W�1�h�F��Nzv�Y�ǭ
+��6�yB&�A���l8�8��{|�z 2Q�?S\D0쏐���w��$�\��z� ����@�(Y�9{�:K��8|�82�㗰��b����d��q�R1����~O?�N�6�]ݪF�q�� ���Z@.oA��E�=U"�K��8�Wx�X���8T)$+�r��OThE��Ɵ�'�lKE.���ġ���Ô,�sk|��+�����M��h��a�ؙ�P�G�v��| ��q��e^`��FtN8��@�]�(�S��� w���Tg,�&8��}�Z��~�H��oq����BѴM��~�E�ܡzK!��k1`�(�n�l}A}Ae�|L�1�����v)+��-qG�M}�}ae�R3j�� �H�� �r:��(Յ�a�ȱ.^�� �D�EA�r����/C��+x��7�*��뿔�j�bKѻzm�s~�����u<�
D��ufȸQ�Q�a='IQ��B|^�����3�x	�������/�RY�>Q�G��QU]�1yG�K�]rT��F$X	�Tp/��J������:6�-R{��C^�8���}^.F�8��P��R�݌��5�-����,�|�~t1P޾�
�prT8uA��Z�\��p������Zm������I��dɦ�
�)DA���1�ҁ'RB�d�b+��]������2�#�?��G��}�^���8��^�"��;[�I�>T���r�
�c|LҾ;q2�#��'��8g��[!T���Kv�����e5�r1]��~B���^������h |1�k-R��,4g铗2���DsD!}_�$!��RϷ7M��u�8��#���P���K	�p35�^�* �K�t��9��3�0����y~���<bx.����he�.�֝��z���ԧ�\\|z�w�>O����fo<��x���������t��x#]c��-���ݍ�-��~����c���h!a9��{�����q�xw�EX]4F|B�̑ob��\�~PȨ�
�F��AFjk����!=�]JCrAәw=q��~̒\����q�0�I`�>k�4"�~n8�<wص3��#��K����e��tI��@7�A'���ǜ�i]p�+���ko|��ZSEx���4 @&D�ٲw7K҈���Q:Y�����ϱ������"��%7��o��9�K�����]�?���$v?8vʓ�	s�:�������@4`��hU��@�@I��oer�Ew�<K�6C��U�P�iU�S�W ܣ`�e�(��W��l�l8�wn�M�͚�9P��ƍ88��6���U���
D�y��+��v����vy���%�g���2C���?�П�`|�c�Y���D�"�)&u}�o�8j��²�3�}l�D�h�@�������;�Q|{��zZ�����'�ڦA:0B/T�&��@��%����qWE�Ʃ9�)X{mso���B��;#�����ވn���jϵ�9�1$ME�D%b7��E �s"-/��w��4�y�D�0�J��BI�Ns'/d��PZ9�x4n��4Z��\~x��m�F?XM?� ���9h�~�;��V�Sݡՠ3[��Ck�����- )L���-���9t��ɇ�A6VQl��-#��Ul�'�"ЊJ��n�뼛G`���M�y�����RN-X���[C�l����	�+�EJ<��k��<�u
�Y�֌�r�"��V$| D�,�c�n�S`K3�#!У�Jak"��q�W��<LZ$�{D]�{�^kԙRa��gqH�HmJ�!�<���c�Sz�v��.�ul��`�8�K.1��� $����|V/���c�N���
J����X�P��^h�1��)�)�03ޒ�^�0:ϲ��Y�st�kZ+�R7{ԭ����4���� 9E򇢘��۔�@�F	��]�Ko����8	�S�o�R�6B�����_����Hw����J43'"{�io�|����?�9jä��6f����j�ɉ����G�W\^[/�v���t6e�y;����/����1�7rg�����o���_ɃqaA����L����{����PEi����ԜщgWe��)��M�u�s�)D���Kc��=Ü܍��;O4�l��8sop7[D��-������KVe���6���1����*^�����n}vW5G"�ۆ�Ԇib("��s��󁟇8�E�a�1�Cqp��\�E:v���i&BZg�a�G6:��Nn��
[�e����3z�a�c���cz�?�-ˉ Z���,Oh���i�f'6>��`~��[-�8f�?x�pQ�X:���x���hզ�r�s�3�#�W{��ex�����(m��m0�v_nrjb#q��$�r�j̊'�ĺ�ԑ�6/�=L���1}O^w��4��&���=ө�G��r%��t���o������z�4Fu����D�ޜ�a���阘��Y�x|hRx>��g����م��|A��R$Oh%����(�\���dڛ��\�������X��~��F2�o�^T�h��c�s!��m����b�8�{��bo��`�|O�s�۴�*z�)_8��q�Pd^+�
��G+u�&^;�Y�������n�.}�'�!�dG�tL_��'Ay����U��c$�_#T�����%o$�El��v��.��v)��L����hG�����xuFB.�Q�d9���\��H�q�[{}m������ʛ�g�%��t�L>Dmy�Œ3N�!ۺ���,�[Ou�V��5�2�.]�)�WؕM���d/�f��}j[�T��J�%�!q����T��i��5��P��1osO��u���x���u����I�I������G�:�47Xdĉ/��]VJ,S���N^P�¸�}���F$�v��F+DQg˄x����opN�2;3��@\0t��B]��2Śߩ7SȶM
q�Z��'�f|F%�� v�`ƲQ1����Fu%k1��2�e�c�j��6��?��M���d��i��NVy�r��\=�,�-(Y1��i�	�� �U������j���I����O��J��6va��ٖ���_���$�;��7�}����>{�ɻGBR[���G��f5���c����톏���j� #��]!��h�@ ��Ez��K˅�="P�C��|5зc
{-���W���iɬ>�$�ͱ�͋���X�v��²�j�����!����Һ���d3�谵��F�� A����},`�!Ax��\�uA�Z�
���@^e��HҀ��{�;��"�ӾȔ 	T�,#|&���֍��X˶���Z��!V�p�3��k��m�2�����|s愘�� �0��Y�S���.�]��^�sەA4��S���B#Po_����P�`�?��<�"Ъצ��[Eϲ��]�D��&u`|������"��,L�>=v$�{�1�b�N]��au �V�`r��0�T{�/���.�ރHho�N�`\g&��Ky(����V=x�h]�W��������e�C���j_���\�^�O6�%�H籄29^���̓��I
������Ao�5b������x-n�Y�6+��3θ���gz�\�>�rš����k�dQr��i��z����t���xu)�W���.���=�~�9����-����GN��e��������$���S��EԊ7g%ůY��V��5�g3l���3U���,�YmQ���]��%�� �8�?1��P��_G���(�Cv@��$k/�H��f�׭ln7YZ�e��' ��x ��9{D|��������{�~�$A��eU
�M!$���~VKb�#t�v1ZW4���g²���`��g<�)��氘��	�h��=��2Hu��ǀ�`Q%�
JD�h>�^X�d�ܤC�+�[6hLғ�H�$�xƷ�E V��F:ۤ�83��O���	N�1���n��7c��W�Q����c˻(��wv�5N�c��ȳ������N�U��&���^��Q�͘�{Uw.�5Q�Ɖ�!c�s�'^� <�v[NӘ$at��eo�銒��]�*��0�,���L��6�o�Z���G"�V^�5�rh�3c%�o��5�܅���4ND|�ũ�sa���	o�S�R��,���y�-:�r\�]Q�l�~T�wh��y�!Rp�]��t�<����$�����=�u�}�6����$��[�}F���k�L�AFu "ɿ�D!�'N!=���RH8�gFFDD�'���K������������EebҬio�Y�s��-���@�؊?�>;��8�[���)���ry�z���0l>b��{Xx�#��f���Tq'w7wqN��35f��<�F1�u͡���V�_5x��U�8��|T_���+o^��6�xo�#�`˹6\�v,�E��7���{|=Jum� #�0���g>����$��!��M�V�	��p�0%�ϱg�-��ZY��OO]���|���]#0p>�;2��$+�*�U���U�@'�y&}�cr2O=������6G?����)�oz�21\�^O�8w˞I���J)~7�8�A������m_&Mj4�Ą6�k���o��,�׍�O���L'�/�>R�N��E��Oe'"l�������9��o}����yS�������K��X[��fD�o'_`�� �_��ݜ�
.aʾC\4�tFf�z,`ح�c��O>�����Gnۜn���) b�{�4t{LZyOx�SJ��i�q(3$������i\�}i�Y'��}G�wH�41���{-gݨ;Q^��Or�\�����:�l�Z7�2V��|i$��u�u��� ��Oᶾ����a�[,*�M�]��Yg~#��[�[?���'PQ����G���Wj]�(�Z�0� �"�A#�(,�G� ,;"�����rp��y
�J�V:6�f�ǨW���f�o���'>U�e���4�I,`3v7��fJ�r��mKݐ�7���\�h�F#�<7�>�
e���̱��� 0���ę2Nt6t�H7-�_~��~K����$+?&�Z~@��SUiL����bo�0�o���@�4�3��5�zy���l\�s����Z�2�n%E�auF���~b����0��D6���l2i���tzۑ���5�`�U����2���z�=5�˜��tV��'����㰞-�;�]V.���n^[5r��Gk+:�L:�aK>�D���pxP���Do�!��� S$��U5-�H�r�����~���+��z�-����③Ф'-���?��'v��?��g���[�ٟ���l���?�kI>[����D�1ʉ?߇�`-*�T����jS�G���0[�-���%A>��܇Sqh�ZY��Z\�H����[�&-Yf�����m�l*����29+f�0Z&�OX�.�\����W��{�.��.F�Z60z��la��ɬ79��~�Qd�r����~�K}��H�����H������5J�8�o��h�3�z�3�̰��`����'�0>vA�;�s�Np򋞏�A�)�Q��`]���5����g���r���?-��1�U���+�S��`�E�+���I������[����x�x+����'��N��lφ�yc� gͰ�j�p�������.�"����6���O}2�]���rX��Z�����8??:�;/ɵ�l&[e�f�[U���f�Fͨ��?e�e��Uܜ��ap��C�;t�&�{EM4�jqn�,���3��{�/Z��4?2L6ot^
xi{8IN*���<�u�7��PW�|D��Pq�������i�:��T�	�������V�{2�i�`�'���q������]��gu���Y�qF�a_�b��Wi�����Ʀ�yU��o6l��/��Z�Z�
��E������k�$�5�]�9y�a��wc��I�VR�}�}�F��L`��Pk�I�#�mzπ�3R99�2����y�d��p�m&"��sr7H��ى]Z��ٍv����g��B�~�}r�p��&�9ӛ����*-�p�D�M���w�A����t�_B@�F}t�O\������!�_IJL�9Gd�4C,��~6ڞP-fr.Q��r�մN
3�Y�.����_7�n��.nUu��g�t��ܓ�����cÛjze��N������-br5]��$8����2��֙��H�Q��<�R�@�~.Ůk����q����E�嵦J_�Bd��C�Jꊌm���	F�(t��'��b��1cz�/ȟ�y�Nϕ�����m<.�u$��G��Q I�4}��yo�D����(eW�dأ��:�j��é���n�$�S����U�%AgĆ��)�(�)tG�{�'5�b���^:D�oP\>UaJ��AN_��iTY#��� ��z�3H�B_��$8��ͅ�!>x*��?q@/�}t�;k)Xg>
��
�
�D"ӫL�/�%3>��3�;�|7L2~n�Ez�X��ˎ��Wo�o�>25�-�x��pX�1�r��k����D���*s��~̕��mGh��n�t�HD�j��&4#�@o�]5I�l~���[�VY��UƗ������֟��!����I�M���hfT��d�SϞ4rK�Ͳ�XZ��q�=f_3 ��`#k0�1���B�d%�Ç*��E2�U� �\Fb����x�GkM㮗�o�?L����Y�Ԣ5l�v�2�A�A��:�
T�:����v��맨j�%J]R7U�L ?�����Ֆy�Ox>p.C5+����!I�rDWw��U-�:ϊ=�[�6�J+�.�M0��uܖO�y�OK�U���C��w�Ϳwt�!�	�e>�c�w,�����:N[�3x�Y���ʻ�bkJ�[NZ�NI�"��m�!��sVP�����(XQ�U4W�ȡ���F8�k��U�������@����~������N1��/t�߽Qrh7Rb��(���5�A٢8u�_��6š#(�&��;�]4��a�8w��[��B�w��s���Z�������N=�t;�W"F��~���Z'Y��@k�;c$�՘��a 
p�o�Ԡ��k�<o|u��Q��`���]���Xs�×�CC{��^i��q��w���-lĠ�Q��-k&��f������H�+�9y�=��P���$�d�Q(d~w�=�_I�����Ac����I��%!�=��;�_���F@��;���O�g �ba{R��5^ �={��-kҪ��X/R�5��""	�.IL�"�O��������$�r���+n�P��*�E��[D��܇jr=G�!ԟs����4G5��%4�w6�.�7͛Ș�����9q�y���N�h��K�U��=JP����d�z�H 	���8c΂�fG�!H�^|\$����i4�ۏw����Y<��\����'�U��2MUyn����@�]�Wk_��5\��v:�_�B��6��$�R�oqs&8��|����SV7W;Z�j:�5��;̚&��ƹ��;"�C ��Y\_ȇ��Z����d�=h��F���K��HW6F��}�2/�
�m�z�
�蛣�}� �*�bO�v7��7#}R�a�҇1�j��J���*E�l�Kv�CE<����2sK��	\?N��m�x+�O�K�#4�҆WvUk��c{������te~'�_��2�e�A�������&�2���{��\O5��Wy�6Kk����������;�UI��f��%�Z���,�-����e����d���.�F�䈡�'yduoE�(yl-̸��}��tV8�o���;�!J�Qf��M������h���a�'�Q̭��+W	����}�"-��\����b��⫼���h枀a�ڏ��z�{x�{�['��/�1նu��y_>�ׅ���F�5q7�ȋ�&1˥�8��s��,k��M�r.� bC�|��r�,�H��Z7��<�[.�n�2?��Fxn�8�P{at�_��Gx�g#׎���>��,�e�^��0(�&���1Fa��1_��/c�+� ����������h_�]k���Z�axP�I��l܆��\�D���5X��E`B�S(���ow�.*���I��ڃ������+"W˭ss��������NK�>/yPr��
��<!�"/n/��*���s����޳m�G\9�\�0C�M��/���^��v��]��305x�������z�`Um/�eW7����j����G�I���)�ઍ"ڏ.p)�{w}fM�Sa�@�2:n�R��6Ȃ���v�=(�'k��z	v��H���mJ����maE���{"�(����I@�wA� f�w�N=
�V_I�RFƑ�Y�t�I��aZb�#<]r����D�%A�����h"����'��<=�;:�e��s��ÇOv��~*��6G�֝����\����ᤐ�m����ߵdZ���hz�Zě�K�4��L�,�Ϫ���*_B(��1�����V�j� fC�E����G�)_������opDYt�^����Dl�6��r� #�KD�8�o/d�n�b?��%����"�m�Ւ��"-�	Q�7Cb�����|��w�
�"=tA1p�r9^%o�Ѕ���[�3��nL�T��.����Ib�YJqer��~��%�6'�9����Z���I8-����
���`�kIE_hNI�;[�Ĺ����O���Sм��U��R�1x�:G5�I���N��ɬWS�t,X5_MvO� ��m�=뉂��N���8-����F=.>��K�{[j��LV;֩��B��=|p<>f4O�_Lߧ0���ŧv��3�:�V~?*���R˲�<[������������
i`���9����9�"I	e���i�$��?�-��*^��c)���a��2-8�h��y&�ۚ�)�<�K7N�8�%2,�����5�-V�>�.�:#�C��$�雪Q*�g���J�"��㒏3�!���n*
Z����� *@տ֑~p�ڱ���r�K�ݔ����a�o�VÑ�e�^ou�s��;`>��y\�w�cR/��Q�vK�(�Xx��Nx��:��(@_���;l�Ei*[���S�ǩ�WU��V��s��_�5�r��0�m��Ӕ��9�u�m�n8�z/�x����]�^��������v��Anyc.�:�z�Z�����{��G�T��B2sW�<�/���w�l�v�ҀxM9��q�<Z�E�rl�%�5�m���u@r�Lj��GT�J�:HT�����L;���ٿ]�}��ɳ�^���������T�s�#���z�|�7��Z1)�7�m��t�|� ,1t�̑w 	��96�yb�{|Omk��T�������
n�[���M����2
��8c�,d��.6O�W$�>_�]�KOm,�	 �}�"�T�����s$6H�D��*<�\3e�ͿK|����p�3�:j�6XW�Vs�+��s��/�\�����ޯ�5��9�j�2vV�IoN��2F���:n6�(ӷ�]��]_����n׍�v}}�^^^�,u��ۜ�`G��Z�r�G�Ԗ0�rڜFu�@�J06y(�6��R�sFry`)�)�6���Vܮe��{+_݉��O��4�Zc�S�-Q��5B��F��K���Ё�t�$6�MN
�F��pBs� WP��Ka��	�F��'n��>����Hbf$�E��I+����]��u87/�I�#���)��C
�F�MSy;�)ۖZ���9v�{���k����V���_2f�t�u�{[:���T�����t=|��6=���g:��G���#p�_?m�����?Ƞn��sBǧSh��2��̢5)�D�>��/����<�ǋ�m����d�c�ܠqwM��d� ���b40�B߾�B�1	ɕа�
�8䍘*�L�Q�,��B'����� n�)�7�� eřS�|%,u��^H�C�N�Q��Y�$K3�a��hB2r[��f���etE�Z�~��T��)]o�l�ېk�����`�R}V�=���/k����6��|Ju�J��[}xSN���ӂ��y�n[]�a�&H~���g킝�^��F;R�\|�ķ���^5�_���d�`Q��u��8�4\x�+ߛ�zwat�x�Յ���dC�$k���Y�\y{����6�1jp�? �
S�%�{���u/a;2�sηՖ9|/~M��ui��\O%�?�ˌ&3�|��H�;�OLLS�o��E_z�خ鴈�J��Z��D@)3pȂVG2��AX3�e�
1q�j�?�,Z`����5a���$��mJ�$gM�HܛaLaI�F�|�g�r�5L9Pc:]�˺���R�7(n�;5��?S'��#��*��d��淼f� np���z�����",�
e���=0���c�9����F�{�l2���0���V�������n�����6��;6�H�'&O*#��R����:O�:r�Y�H*%Ϣ�5��E ��%q'�]q�g�F��f�����d{@m�;ЪMX�-jB�Ȗ�A���?'����������m2�'7�s��l:�<آ�j�h m*X�i�$��)��f�m�׼���k������*�r��ep��x	ǭ;]q4E�̓Z�͋�Gz�`Sg���&�9�$[���!yM��/x���rlRj���r`A]{C|]Byʝ�7� ��B��TXS d�����>���6
�h2�єG3:�AN�i{��"w���i)��5�S:_�i�x� h�Hi*b�GF�!-N#̍���$G�ڃ�6a ��+2(��
���=0K'�j���1�قі%�$������^�<���ꁇIۍ��f7��T��!oG�~�\��z2�N�E�E F�DPw�z/,&N�.%�=O\R��B$Ժ�{��r�9%M�%��NS{�X����{��^y���X��*{�̊��%])p�p�����[ᵼ�_�}d>�;����6�1U�-hk���&�Fa������hş1kh�,�-����֨6�D['�e+�_Ji5}$EEe�A� �F��Nkt�p�	>�N�74�aI1�Wv��i��M���p�k�Fz�5I����r�iļ���:Կ�##���!��#���2 Ey��=^B���,{��uJ'`��.���V��gd�U������{C=��-h:jHj�O�ؼ�c=n�Ju�bߊ���&�v*q�i�������>=���fnN��bN��}*cW���<٦�c���m�I;s�����|A�&�;�r�`�T���"�e�]��|�P7��
�lڊglx@���c�tC�_���mĲl����1]�o�ʫ�%y[it�p	A�����^ 2a�*M�a���ן6K~-Ҋ���E|R�2q`[\��Nڍ�!������P�\#�i�)�4�Ib���b���76 ��n@A�4�bf"tMf"�p̥A�(C�I=�d)���Rף]��,�2�}���#�T�#t,U�uTVܵ?C������9�J�hQ���e.�� ���}i��K��M��mI��R"�ڰ��!�t����ޒ7ȼ'��}o��l�}���y`���G* �:�H]@ �H�R����z�������3T�:I�[|����p&%��t2l,�e��A.�1��F���y����l���ܛ���v��&������}}Ip���ԗp����6������oW_<��%�<�|˱���=>��*�+u�[�*���9�8�2�r��Q��;�2��$�oa�w��5����ͰХ���(��z�N��|)nc4�0B� �O�Ȕ�N 0�q��<Q��h�z�m՘V�;���7}�hS�&)���c	��]�19X�B��l��9�V�Fڑƥ1GkR��6�d�6ep7>�L��)�k��IļJ��9.!�������U�/�I�m+�����DC���Vа�$�<��S�]���P{Wm��E��-
{,彜m�{����M���n�V5 P���X0������M�-֓�|d�w��I]�)������)�ar,�َQ�it.,�%�#�㔆6q�$9/���&~�ȗd����wM�@�qy�,�l�9�����և��ݕ�:{z��|�n��mrz��;����������E��^狋W�$�\��_ou��^_���8��f�U�7����T_�z"o�����s��<)�)' ����/�'JHʣ�*M�%��k��>�e�NG��fd3��HyKM��t6�6X��� ���}���
B�h_�'>�����&Y�)���`BNh�<]eZ�,�O�*����U��I���7�b;���>XG�4KMq�zJ,����f��A<�H@�AP��\�Y�pN����D�2�Rٕэ�d.�;��*|��^�NHս��^�C�՘%���zL��w����&�+,�]��,H�p�s�u�)z  @ IDAT�����'�F���o@2�qGz�@��Y��b~&]^mR����G�˅}\,�bosB�B�'���!YNvkU�:���L����t΁�dx��J[�.��t���o��岿*�=��k�ߤ���~��}��_�~_Y������|]�{���5�p6�/��8
��Le7
���^�ť�[��� K����.�,2���>���|]\�aDZ�o��%6o�#������Z��ă�����Wr|n�N�Y�ל�k��@#|!9��EAG4S�c�ɲuR��<)��YP=���$�I�c�Sʆ	�d �6!��tJ��4֋I7�Ѭ���>j�lo�3l�0�%��?�9g��F�s3+�+֕S��w�5� L����ld|�kY�9�O�EӮ�q�L�6R�Εt�NRG���w��'�|1�^�6�CT�ESlC�r�h �o-A3��=��N�qn���,t�A2J��`�[�
�A��;B(!)�%��T�p��I{lG�����������ɦ
RG$���j���R���?S\EZ�@7A`*I#��wz��w*N\�́5�w�LB�|�Z�q�������ip����{���;�3�<�ŧ�lC�L�uE�D���~ޕ��[5�>r�+~[��[�s���F�uT����M_�M]Ѯ{ӭ�M�J��aQ�nl��\JLS�yl�&�S���j;���.4�����]��f��<����{8�Є�V7�.y��H:�$r�Z=ۘ����QAB���h�xM;_7�O���~y�.v��Ξ�|�z,��SXJq���4�>r?�?��#��NV�(H8��ǎΑ" �2�|!/�Y�@Gڮ�Q:�YO�!�:�rdd0c]X��`�T���E6��#Q�C��aK��{�K�r��Y�@�Tm�lA�-o�٩� �5%ۜdi�v+��"�+~|�@߲�d �ƈ�@��c�lrr���'OOWO�?y�|�aG�����4��V��y�F�qܸF�H�&>��[6�N�&���t��׿ M�7,��T�f�:� �[Wv��lX��@ih��K�RJ�[�2&�j���M+r¢f�۔~� P'�ߠ���$��C�5�cg��\��	z�?<I<m{�#!�s��Q>Mq�����G��Q��T��N����+�c"�Gv���ְl��K_���������&��"b"��'w��� ��J6�OM���т�֌���O��ѿј&&l�"l�C���NV�6g;��h\�y�#O9�> �r�A%��o�P7�敮�M?劳L�s��o:rh{y��o�S��~��g�a\�nI֨)��Y���mi �?���ۻM�6�ۻ�O=�m��26T�{��4�Gsi�z�����o�s��<d���K�JUˀ��,���E�7�5O�>�5�nF��ˣ;�Q�u� hut���f������y��_ba���^�kG��?t�|��p���G�ў�$3�2XFL�d ���:�;9�qJ��T��{�呾p��ˤ�>�wϘ;�kAd���T���-s/:��r�)�*7ѭ��h��ٕb�^�>���>�`g�pc�Kݣ�ҧi���ڠ�	{SE����7�`m���H�� �����!�C�o�o�r<�t�����o~���w����͛W�gϞh�R0�~��Us���QD�Kf[���wҕ��ty���g��9M��(6:�2��ą�mT9!�EE��v\&��.���)q��<Ў����Rt�&��p�^h�-c�2`��`�$m���6����Ƭ'�t@� ����k�;9���}�v���޼	eRg�\8y��Y��=�HL��kTd+%��a�K�-uv���b���4��y�&�?C'����q�]�`���v�p�����I!*_����X�=�N`�ZB�4������Jn^iv-�r��y�w��������و��4�<�W�.�����o��?l��8�E?�`(7<J�'D�4G3��)nW�+]���4K>��hyHU�$��Z�Y�d���f$�(uM]�k�%�v62�	_E'2n�D �5�Z[`?��~�����߮~�����啂��՗�s�QZ�c'������" k�����Ni�X�	@4_^��_<&�ǐ9�bo�e�b ��ud��y>�$3���3����H�Te�̯��\8q��!���$D����#��2�#�%�? �T�Z\0�ώ-��Mij��Eò��º"��;W�RDP���� ��V�U|��5� ��A���\J�~��nיu�֫��Y���#{���ꕎ�/_d0Ƙ
�I�����:g\0���8m� �N�N(�$�Q��@����-����:��4����М���`Pс܁����9�lӲUOy_��v��LY�~���������f��oЋ�>�׭3i'Ib8sR���d4���X1���'����d!$iO�� �ic�hF &Kd
0<�?IP_���[��9	��={2����./�QfLgjG{7"ho5�OW/_<_�^w��q��>�G�Bkh�w�8�G�U�.���NѪho�\���$6�����Ǵ)|&��y�����Z�\�w�����O�[�(Wڊ��]�<��.;7�\������,��=�&�SZ�L!��`d,����2l'mٖ�_��.�K�-��G�]�|�A#�^i�p,ޱ��T2&d^��;�ҫEY�]���jZ�<�ؕ7����;C�N��ڍ��/痫�y�z��/��?�>~>����2wƢ�Z�����#햡�V|̣�<��c#c�y�v�Ju���y�tr"+��1V)��^0	ଣ�uT�4���c����>�l[��MǑnn���
G�bLA�e�x�<v��t�_rD;�$��l�|���[~(�X!!������]Ҩ.mA&q$G7�faw��?�%~e-$G*}xzz�z6߬ο\I�����"�/����Փ��VϿ�q���56~��߬���߯����F�b߬^�|��l��B2Z�U���}%�is����r7���N�9e6���RKmYr̕������Bw1�P�`�Ȕ;
�XdZ`����c�W7�1U`�q�(CmyjwEW@���ľL��1HL�:_���<~��v�R�
|)�A܈�U�R����<]@�b7�ai��::H@!�0jBD�2m����en�ҩ�+�#/�d}m��JE��@Ή ���n����9���&�~T]��XļX�\� ^j��oo�����2����~q��T���G�(��A���f�L�;TB!>���{����;5(�J��ęҧ��k�����z�3~�Ǹ�k���9�y�3�f�u��p�3�<�m|��\i�<�ɗ���eh9�����6�T�'�ͣ`��m�u��S�#w�z�y�W���8�O�i�r�k6����C���ڐ?\����o�5U� O�#a�Ac=��|
�����I��N9�&���5�\ػ��V��`���V��iM�%�ܱb^�Ӛ��:P�y�E��ϩ%�3�+@�ʆ���V+��L)ЁR��0S"#�1F@� p"=�a���-�����Ocje͆y����haR�/l��?(����sa	��A[���tCp���7����5�����bCZ 4tǚ!4m�!S 6����C��Λ�\�B�֠�bY(A_�d0w�x��K�e�e
Ԟ�}��~��ۏ���|^}�r����W����v�^�^h�����q��g�G¥���e�~�����{�6#� Bm�S��/�5�Ϻ{x����Ƿ��~��O�����<���Y�Xn���8Cs���j�L������QC��F��� �N�$r�
}G'���H��<)1�Х����X�bt���#=��7I�5@���~��Sl/c�|����px��
���S������H�$%Izq.)X*�j璱�{/_<[}����ǫ�w�uGq�����w<_��zc�N�!�1q�fp	>3b����GN�	�j�@���7�9vRG�km����R���^����1�i�Cc΍�s�s���:�v��y]��.;7�R�9���&8�u�n��8�������*����|����N�&�9����k������5��R�~J<�w��|�	������q�w+���B���m���)��f�@اO������»^,�l�>����G����̏C\�O�0�F��	r� M�{�Ad��hVTt̕�B�o�Jف ��BC�!����$�+�s?�	�`�ARDz�����ɞF��@� ڃV�	hG�������K[�}p�v��톂[�r*$���C}�������ñ���v2էײ�N�7�b�P�x� �v���b���ϫ�ߟ�~���������׫���߭�������{�,�!����/kQ�H�%�9��_�E �3��F8_Ç�|���vyQ�˗��Ǐ��N��߭���'aﴵ�^����vN�p��=� N/���#�r01�Q"�:����=JѺ�d�#� ���@�1�G��
�1XR��O���m��)Oڈ6��QN�jZ����1����<p:c�#
D��eӁ5�>��S�Sj����\�JT��\T� Hw�LxW��<_}��߮�������?�]}�r�R\꽊�ᓄP#�q��L�!���q@�K<�7#�/�_jb`�>�OL�EB���O��u9sxÜ�����M�9��߹��^� �x������r�m��fS�˯u��#���VM�T?g����:�R�#���F����>Gn��SsD��: /,:�����<��v�=�i^֊�iE�0������1�0�D��|�N��Z�x:x�ȼ��A�M_���� f3W�b�E��k�}#n�����j*���h���7�j�E;��5����e�E4�砃ڑ��D0z{�g6��=-�R%랋������3����Gc��1wÃ���R�X��G��l_�G��e� ��BY5p��)y-@�{m�ZE���(��a"a��ϻb'�ǉvC?�_��:v�x�s�5�_)��rq������
��n��Ri��;+>C�')�sU���0>��7w�ZX/Vo�h���ᇷz��N?���z����ε��L�&۹��j�����n��?<��-W��z�(��Gg��pc���luj��75����R߄�a{����Gwpq>����f��?$�0H}�,��h��c��N�l3��c�!�>R Aa���1iCD��L@�Dg(¾L�]ip���ၳ�M�� �~��ͷ���?�/���?���~�:��a���?D��V?���}>�!p���;��$dF�R�?ڗD�;g�9G)r�ʾI�K���|e�9K��ky���`���܆]��g=�eV��iz������rӳp�d��y��o�L�����g��~��;��<a:�sΕ�i����k�ql�|���o?=կ�xL���_LW��x�%�0�iSK9�N���S��ãǒ�2ë0m�+���k�ebde�#�`ΐhl����Y��z�1gHHȌ�58s/���5��#��w��k(yΣ�$0x8�/c9�EI�,� �!��ǭyu���;P�w#[C6���@��J�� ��#=၌S�	B�F�@>0�R:�G��oZd���a|��*}F�̣W���x��@��C4���H���ձ�dG��ֹ�_����Y����?���?�^+���v\%�xA��-����mA�i�C�� p�-����O�_�����?���ӟV�}�C`��|�ӧ���xq����������j��:)L:M�`M;Ơ���`W�Z� ��ДbR����v��V���$2��D�D���Ζ�=�Sy1�� 4>�c!M%>� ����6��D�.ʐ+:�	t�O��a�l65�):m�͘P��ە��m�J���+58շ��g�)���ȽQ ���m��w.�CL؆]Ͷ�&�y�F�������@G�3��j^���lJ�cp�2��驪�Z6�y�Q�4�l��|��8����Ǚf.��z��z�>��^6�ϗ��ηY�+�&9Ue�����>��D��m�,��e���.t��Kb���89�dF�Ï~��I�Յڡh'_�S��l_��@�;d���{�J�#���`C�x��ZG�	���Wtb�IaZ,��X�̍��#��"	�2�H@�x$1x!9-�o��\�x�
^��6��'�!�Lq�i�N ��j�*ic�S��%�	;�>S���2(�q9>T�H��H�N>�b/	��H)�� �J�I�C�Ru��i�d+fw�������fґ>%��	�>|� ���T��V�����7߼���%B	�4�R[�>m<ugAF���ǝ���9��\/��^�?��w�?�]������~A��볶�.x�x���ė����Tϓ��"M@F�EkӘ���T�@j�rӐtr��O��'��H�"o*
!Dm��2Y��(6�TNY���d�ak"�,_ƀ�I��ѩ��x�6�Ȥd��,
qj�j�<��Z�=l{���|��<�$M���BP�eG���Ԍ�"�W�<��/��?�X�w�{�y'��~�i�J?��w��m\�?��� .�0~k�r�$D0�5Nc�e�?���g�O�sҀ���¾F=���`}^�K|�����2=劯pp�vB��j����<x{�_�^��M�J�I�����릭z�Q��X~�8Y�s֗������7�F����N)��~�D��R��5&mD%k���|���OtN5_���������G^:j����?$#c����Z��.�fA�TV�lc�k
�|*ꡊj����%��	S�#�c}�9'�m%f䄘��� ���g4��,� }���G�-7I0	\�33�<�ҷ�8����!W�A�����s��%�4
�'e� ���6$Y��]�n��%l0JN��e��|C�$OcW�0��+<�Q����J'�X/xT}���������O�>��>U�T�
{�a��b�6�
��Ф�َ��݋���.���������w���IA�?�{^����z��7
�nl�3W*�����K�]5��y*+��'���&���yJE>�&U�i����J��=��>�a8"8t��lM�@�����3��VG�7�A��B?p8�Ę�g��T��%chtg_��lscɬ�+tʉ��l�r��W��#a��V�C�#�ȋ�o���Q3�y�����=x��	�_��W��Y��C�Nۂ���3y;�e-K9[��q��>	������f����%�P�ÍTciv-��6O�,��<'c�9�Yή|U�%�����Z�v���I���s�8e��������mm1V�
������څ'��µ��n��gzx��va7��E����5�/X���j�yVu��̀�<��k4�z�s�w���.D{)^��H_�U��D҅�_����Γ�K�	��T�YQv�]�eJ{����� �_D9y�7�+����lhS� c"Bi��B�SQ���u���ڴ7�����/���PE�N�iS�Z�i�!$�'x����0#e�sKR��f!��b���/�I�X��	ۍQ!�j�D��ػ�\kҢP=��X륟M�k=ջ���U�a���t�w��c���� �x�#لM���\2��G�iTF���z	�>~�O0��u����^����_V���;�)���F~=r�z��9~�K�u�<����.��7Z�6��K�$�h3N�Vg�y@���+[/���($}vTk�(�@�|�h'�B��;����l^�A<�=q'�̤c��W����@�iղ�����4�!O:`F� ?� �	� ��,�]I1�@��6��/�5y�Pt f���=w<;!��N�&8~U�?�y���	������
�~��	�z�\e��(cW�勧�Б}�m����/��I��	�����m���6'k;�<�}m�4�mO/k�ʠ\�s�˷>���->ʮ���1~_=��s��'�Ǯ����Gw�٥?�e�Α���4��^y$�T��:�;���pT1�����#� #봋y���/����c=��O 	��/����~	��]�c1��z��E�<_��%�ʛM-[Z�$���K۫��=_��",m��@�f�T�v����v0/'$��G�J��N���v��d�*�����Hy/m���0&Z��
�pH`'�}�TJcD��
a�H��(��@(ARM���<����_�'� 0ͤ�f���82�K����Xճ1^�Х6*�����(*
���~b�!�T���������������W����+f�6b�b�l ��1;_��������տ�=����v���|�b��vƾ���ݔ����	�b�V��eW6��/���.Hg�r��L�B9y��_v���NBj|�3�8J���X�#�l����(��9����x��%hUD��� U�C	x@�� $�Hi���Xz�8lR��v�	BK��ť�م��:��,�������� ��◈��������mA���&�&���纃|���������ۧ� t.����,����~E��9��@�X��6�m��������d��>Ñ��k�>���Z�EnO��6g�y��� �u����n�5�]�m��G������s�zY��r6ј~��p�(����m^{h��|�!�ٟH����V�����g?,�|��`+�R� ���52O�Uz��~��O���9������'O�i-[ō#߶���|^
������aM�B�B��2r�T�C��:R�b R��)�s(j�e�&�g<�k�k~f� 6�n���>H]�f=�H���ܩ�܄�Kڑ��8�����G1�g���$d$.�OL�"��X?N�B�l�&ۏL��ܴ�`�p^�ɵ%��G	��1*Ъ1�<7.(���ŐRYh^���^^�k];ү"�z�O��V�;��C
9؏��҃<.0	���g�k'�G�i?闎�߳�u��k�:��v����+��s��{��謸Qcr0��QAJ/�Tg�&��t�ʲ	��/�4mz)�Ă-��K�xV`���#����5�4��lۘ�t:���(m���[��x�O�%`J:�>��J����|�V)�R ��|�?�0x�n��m~0������W+�^z���#�)�bE��՟�q�����s���K�қ����ўT[�u�H'�6�v��QҴ�}MTь���B�/��M5'˸��!���{������_�=�<g˜����̳�������s6�.q?J�v�1����zh�@�l
`� ���q����e�ߋ�����9�j�ST(�u@�$�9F0D��׌ϟ�l0v�nӂ)�[� ^)�Rp�V%��ߢ��"g:�~�t��9v��m~#��B�6�]����ե>�ğ�c	e���4G;��n 9��k�AD�ri{��PT$K��Jb�Kc�P>�!i�d�!��x�X�XX3�(���(7�A��X���p�ǀ��X[�gL���Kak�C�:0&5������`I�B�Y,ޒl�خpX>������&"^e��ї��ߢP�3�D��&||�K9�>ѓ�՝��';�z����3�Y���?��UoVO������-�Y=��˪R�����~���G}b�Ƿ������z��\_
��9Ջ�-���e�r8�����,chǰ_�΄�MwX�2"�YcGed�}�i��(!
M�ȳ<��kP���n^��q��>T��A��n��N]�i�I[r0�3���`p�A�$4RFo����4Б�����`�BuP��� 4vA	�������Ԡ�����fd*I�)u����SC߼y�]�g�IwNfLh�;.P����n薞��R���M��&�u9 �v��s)���f�7}��f�%ے e���|ٻ�]���9�)[O�W�Kp�v���ͳ��<��Ȝ�g]Ȉ���9�^4���H��������<�k�)W8u������x��Y�a���3Y�T�8o��qB)>��=j33N�c�.(�,jaԇ1O���HA�7��D%�?>����)�s���zt��o��o �V�h�6~Qy~����K�S���~p�I?6��C`\0#bS��̎��;b��|�~J>��9&�N���G���$V�S2c�je}՝�+���m>F�	<H<��G�ݳfkֱ��Ȳ|i�ϡx��Vqd[�hc�	g#A6�A��DP =u����ǒ�f��L�G0�v����Am�Ě�P�k؋�t(�«��.�2�ԟ�~��ǻ�	��#j6x睝����������_�y���Z�BO���vM8����|���^��Q�|���^�]�+���e��k=e'N<z�G�,P�bqn��~	���� �{�3΀�ϟg���N�H��p In��>�ΡM�=���A|ȉHD"��O�焜�,�DX��_�����G^�N������$�}�#�کGw�q?鏦`2� �&9@98��H�F�0��&�^7vac\�p"<�g��F�ح4�:+��M���TUȭ~��o�U���w°����F�z����1�^h��F/�����'v�d�����+O��|";���w|�x�G+Qj��T����9�Y�sld}�X��釼��9�ek�}Vrdה>M}��l����*n��&�����Y�����/���_y{��;GW-3�d/�ٞ�.�Es�����,<��93����ڥ�\Cϴ���`t�M��4o�Oyۮ��/��z�5� ���5�y�����]��я�*����:����r�W�ޱ������a�z�GG������5�����'�����7�������߭~~�Ek[̈���oO}ԙ�)�r�a�I�]%�1�IF�C��� �b���vy�T����X����J� V� �?��@�ݴ�'�����q��f���0���Wډ�06w�0:�eC����й@�,K��G�\挅���M�lك��m��@2a�����;`�h��'�=��X�t�����9fF�����U��B!���=v;� ����\��\0$�9�j�W�̬����,�)���d��BY�X�Ѿ ����c�{[�y0�1&���1g����~�o����Ox!�/$>Jg���j�כ0��9�#;_���w�����+��]�e��a�p�TFO
��T�(_��IzU�n�٠V]3�JX?tB���3��~�*{Z��&�T�چJ�Kx҉�敻��&yU�O^��z0m�7+n>ʺ�Z(�pk1nk�Ҵ�F�T��e�>��NQ�T8�x�~�l<��2���ͭK�)��(W��#���<���F#�v,a��J&|��)�t��Cs��£!&c��Gɖ����t�� R�39jb���p����շ|��w��-��_��x���ϫ���Wg,r���~'�7�șp��7��_zO�Z��-�#����>�W�7�����L���4�m�}��������q���渥�6��Җt�
7�K�&���n3�M�7�ϸ�GՏ�fL�z#�m������i��A&<�N'o<Im�>75�6Z���}˹gƝ�-�9n��L�T���)m���G�t���R�[�El�4�ht�����c��}J!(Ӡ�Xc�/��=��$�{�O�܀�O?�(GwIw�z���d�����]���C���5�9��ѐ>�\r���v`o	�}X�p?��Owp[�����*;���3��k�plLYT��T¼a\�o��v��J��P��8V��~	c�\ë��bHTX2~��W��88����L�<�U��P��;�%���?S�7��2E�Y�V�6�E+\��� �Dy*}H��4Ko�a��,e�������I�P��pF۸@?p��_��V�'XOOVw�Y�4_��m�3�f����Ϟ�ʺ/,`?s��){n��^�Ĵ��[qY�C�5�2$c*7V@Ș��Q.H��ƛm�Dv��E���>huG �H�Z2��68��ے�'�t�p���c���4 RL�2-2���	����7�#�#�Jȡ&oʎ��8*[*]�ZȎC��r��9]���_N�l�Y�G�3o�T���/!j����@L%��9i��x�5�Gx��!�(������d��Ŧ�EWvȓ��c���M>tL*���	<�,��o�^�����oih���X����'��!�!F	sz����,��a�g���������Ro����z�G�6,��}�)����A+u?\Hv\�]���4y�;X��p���Z۞@�4n�ӂ���Ȭ�K�9,�}h���⑎�۽	��k�&���wyt�{�６���o�n�\����ؿT���<��$d`q����4o�n��~5əN��q^�)\��|��N��OĔ&|�;�KZO�Hɔ�m��[2O�����3�y�:_'B<��C3�I'f���q������g��[�m���
��O)�빀��,�?Ǌq�b���9�A�������$��X�����?V�R�sɐ
�GS\�D��=��5����0���Mـ��j�j\�م]������g��Xm����7_�#���?�p]X���� Z��α���)@�e����d�rD�RfFpeNrJU|� @ￖBD�
J��T�(���l(���G��"��с�rlNDNޅ+��-d��;��%��%�Si�<d�hɄ:�mB�$��K��g�P���!;??����~��!��ë�3��_����%�Xm��Kb|t�ǟP����5�_jq*`�*\4(�:��U�U��3!R��qSHR��"@-<���T���?���ě����0F���U�43�Y�
m&��,����D�CW�(�(��5�hU@�@���.
���.��,���xV�'�����K��Z����F9B�1�^QI*a��)n)a��#e��m(>b}7������>5�]
��� ��_t(�H I]������9�W��aR��M5���m��Y���1����������z�������]��8<���a���w1�;e��bOe�n�C��xƤ�����.�L��}�
P'|��\�����Z�B����@#��yx� �5�7�t��3�N_����םq;|���Җ4�[^�����v�x��p���{嗆6Z�u<�0����n�u�O՗��j��<�%��!��kjb������9�λ�i�iuz��5>ퟟ���i�xa6�i��kȯim
`��<��b�7yy��Z��z��w������%0� L����x�-_��8���~����>����ӟ}�,S�o߼A��\��QL�;e��.��W���`��q鵣]_4��i;�Hf��蟠T[�}2�, �����`��®ϋS�+���V�����!�=�fl�a�����"0��Y�K6��-���z몈��e�"��5CX7%���F$d��!��4R8��7�i!9paV�]�S���@	�ĩfRv�gPL25:���p�yq9�1/k�Pz�CPD�a����	�JuZ�=��}ҝ������1|ʮǿ�i����?s�S�?��̫���X|a�/���u;�˟�C�ڐYH���U���_w��Ȥ�:ȏJ�A;H��*��r��NE�HZ��X!���F=�����V���������=,u�#�C������5ӵ��o�_�\=y�lur���.�)��%e�am�t(�nK�l-�o-%E��OS�j����jl�Le�Z�!�dn�%�
��"<��B)_sHIi1N�Z��(��~�`�{ �<#���t��>@����W���ob�:�`�u��x�"����l�F!;Ps%/��9cm�1V���6�����%���KI�ߝp�F0?�Iy��wM��트�7�g�˼o#Y�ۧ��D�sh4�/Qn�j:Mw�k�/�;�ϸ���v�q�O*j���]�k�5�F�퓺C��;`��9�����-����"������<�bSZ�uZ�\�Òz��:LU~}����oDf�a�3��Ɓ2/��ު��>���d��ɓ��o~̺�+�k~��^>������S��X���ӟ��5@~����m�j/��N+l��3�O�,��D7�(���y�)\۔c!媺i8eC��>`pxp��!��ӟ9,��Z����[�{K������뗫�/�Z=����!}�����Ɛ��d�y��x�\���Z����	J `�ƙw�(W#�z�1��%�wh�)���a-UQ� ���X�!����d�NX/�H9���zS.y����K7-\~@BA��j�w3E�JE�<��s������K}�:0ۢ��� ��A@�����s���?g��S�/q�ӎ���puHy�/�Bj
K���p�B�FA��樬!�0>j*p���6LF�9�#�RQ�7�D�)�QF�
ѻZF���Vj	��!\p�p�iu��;>��6�p_�~����;����N�����)1��[ގޓ��JLY��F1
Z978������:�=
����eΆ��s|će]�Cv_�X5]��GjP��xȎ�L©�0��ޖ�~�2M�§U�����{������'�ߣx�|}��7��t"�{�rR.�[��fr���\�o=X�TI�!��*�A�����k��?���9?�<�:���!�k�����r�'���2~���ĝ�� �,�V����&�o���qMg�3�>W�6l�����q��%�e�i7|��ԝ�i��-x�iS�m�M�]<J�i���$��M�����"�Ϩ��[�9>���hى�Cgd~�Qe�(T��)�t���X��.F�v���S���\:�̝o���Z�ǟ�^�3�o�1�ȋ��M��C#Mྂ�@�T4���/��fl�q����qGy�`q��e�b͗���p�xu�Qg�1���׋�~�v�:E��s��N�	�dc���[B�Y����(h@���'�an��L*��=D�4�¨o��H����cenHgͱY�X���xj� H\�j�����-|�+�g>�r
�
���#���,ڔ9�r}�g�y��)˻��"-0\�UֲJ��3C?0_��Oo�����J�uJʉ'�z;c����l�%��^aq�|�ɠ�@�-�>
i��@B	'PJ�SM�*�����aJ $�� 7���7l^	�Aj�\D�r�$ � ��7!���͈X��x��w�)��u�蘵lc6/ץ=z�d����2�_��z��+��ybQ��!4�Eq��OU�L+)��:�Vi�M�o2���}��a��������9�:���/W��㿮����S��A߇�l���||��o�)HNz��l< ���ǫ��]����������b����[��j�2>
W�yە�L���dA�9���R&���6�[k�L���Ca��J��o����EO��yk���e|����>�S��g���-�2�v-i/������h.�ę���M��9��v������Tx�[�=}��g`�dp
��k�,3��������֡�xd~"p�c_�?����1w�[~B����7��(RX�=,��rF?;hJ���aA�ZQS.�ۣ_=��E��%Ӗ,��������3�����"y�]s�.�0��O�M�=�a�T������k�sAg�*�o��0`;�b��,�g����s�v�z��1�����.�.�cl�a�����n�Wnj}��4
pIw0���L���q)�`$���U�i�Zj�?�\�>ק��^Jy��(ʋUe�D���F�!��~$�,o�H��^��`��W��ME����!�EG���.Ey�ي���$v�������w�P�NV�O��v7����ߺz�71Kj.�re�>i��ea�yv
����Yp��G�*�6:b��]7��	���+T�LV�B�*a���"i�B�d���Q�7.���5R�7�O��F���ᓟ�.زU޻��F �{���a��b����J�l(eѼS}%4��Rf����
��7w1, �I#�V�}�o��  @ IDAT��z���������n�}�x�Sy�;��x�7{[��gsA�� [��	��抿}̩GLu>Ą�͋�~��7L=���]5ʡ����6�6��7
�8S��9�4�'�<������S�jE���X>�A���)DF��M��[�A��ԏ���U4�ם�]�K�ߕ�}�n����ʧ����a�/�w�K:��n�x����L�-���-��w=.-�zԖPӽ������v�Eh��fK�wFI"��̃�s�s����ˌ|<}~�������5&�taY�(\�iu��9N��m�v�0-,Z�vv8���Sr���N�6i����Fa��?��J�-C���@��H�h�lעRx]v�'��VEj�Ld�W>5zeq
�ʑjK���f��X�X�N��W(�=8���=�i?�9y�k�%P�+����ߟ�jūr�n���X����1D��l�( Nx�@�<�c���x���%#33�e?�[~�Ji5>�x��[��A'Ҷ�4��}�� ������f��T���"vu�nu���՛Wǫf�VW�Rv�!@5J��pگ�d{*��B��\���`���s��wiF�n�R��fh�Rl
$�.���G�X�&�k��P�5-I8�o�,��t��' h�&P�0$S�������+��~��THǄ˴&1�a8�ŉSA��e>S�z�\T���{c*4g(�*!��F� ��
.�~��&���ld1��t�̷e��0 A�?�$N^Tmp����ի���+
����y>z���C��(?|">vP
� ~N=�}���^}C�}�u͗��#�w}�Փ�o���iǯ�G���B�C}$��PIOs�o�6Z�5�S����R�Ҹ������Z=��?r��	�r����a�փ���hk���\+���� �y�� ��x/sC�E7/3��kg�����������M�4�M��v[z�t��2�K�Ҕ��-_�Sk���g��s�i����ϱ���̌g2�s9�������|���T_]Ho?dڛ7��b=���|��>���իwH��e���$��������s��p�斸t��:0�[E����{+T���U��q�B���$�׼s۷qo��Y��W�~�����9f��!_�B�%̝�҂x�ܠ%�����Z�k�3A)��c�S�P����%��9w����&��K	���R:����[Â�r�^�=�ɏ�<O���꺛sDkL��2�X
��z-=�|�CKb��Ƭ��
�ɴ��%K~4^�.h܇���O������kxz�jRǜ�GM��y�3�~ba8��!	47P��d���B��3mu�GKW4>�����\
�F� L� ��	F�fa���HJ{�b�+�A2���&N-VK��@-�Gx��G�R��+~��DV
�2g�q���4��]SZZ��ЊT��.�=,��ݡr���P�R}�iM;J��2�gq5X-��_CZ:���Nd-DiF�y�gT���`#=d��1��vv4N��i�c�Q�x�G�fS�ͱZ)YN��u��5`0I���껯_��?~�Ɇ�"iɳ��,��N<_G~�̢HKU���U �R)Ĺ�ΰ?�kC�v��\�w�a���p�<4����]��1)˄���;��w�K�%�e�S���_��.�鴎���o^�]�g�ms�V�#�2δmq���m���s�%~���-��7x���x�o�5n��t�o�6�eZ��G_jػ���������������ױ��MN-� ��A'>�d�Z���z�+�j�_���Y�ό?���A��Ґ�z���X"Y�u����BovY7�2���$�{r���Ȍ�pg��?L��r苌L�0#8��2_%�`��DO�ȅ~�	]�bo�m+�f��x|�(c���Sh.�y����3%�t�rf_.^r�L��Q#+g�KMsX��π��2�!k��X���񁏡@���B�a��Q�`��(��^��*� �����(Rk'pI�c�z�rV�ƥ�S?�$s\ŧJ��Q�_�Z���f^��Cn���R�G1�� � �]#�����د1��T�A�2�^qv��)�W�^�H�:�2�Q�4�9s������+z�s�����S�!z��R�R@
75a� F�J*�%Dq�d��WK����aH^ai�z��>V'��K�x�Z焠����8�b�(�F�2���Q����d�[�?��'_����K������Rr�no�/�Z&��
Fx��@����Y���*9���`������#�y�!TOc�K��xyM�b�
��Z�T¤�����Q��ڱ񆅀{X�S�̬'/�yWu�V��v�ս<;< �����g���������x�%�-�J��T!�6��e�z����p����ʖ�q��~�Ӡ�s݆�n��M�Xv�����_�V�Є���=Z/�0���K��F���P%yN?�E�w���o�c�ϋ�i�۱>.����Ԗ�2�S�>�7�ϕa�/���\��pX�o�g\/����]6af���n��F����LCvYG@��-�w祐>v����]�$ǒ��ǳG����zŬ��'��R	�s^5z8�WA�������`��I^��dЪ��㥀����+�M�>��?�A
S�H%��"�D�ߴ����9g�����{N���7���x���/=`�/���H*����3"�T(U꼻n��k�w�X��4�;k��!
��t]�p�|]��Ԣ����ɣ����T�P������2��b{d�l����3A^%c�v|TTh<7��w��)���7<��a��%K;���#�~���V���V:3�c��o��1�c�b��;ŪF �66M}�O_��*֯}���]1P;{A2Uu��Q�(��1�#�beT������[���aP�4H�-��7�����eA�l~�ae�g���ZP
�؝?�&p��r$>�;���]a\�Q���k��]��Iږ��!#}@��/_Z4/x�xρ���!IS	;���C�Ey%� ����i�ew�)�c���:��/�88�ٷ�$T���,�|@�T�pJvc��nG����Ό���ƾK��Ž��dS,@�d�z�8�T�=������8S��,f��j!����c�������p�\�?�V�G��]��a������%�\�� ������p�i��*��	]w�zܶ�pMs[�w_��p�ǌ;�o�_�%l�-������t��a��;�%N�7�n��q�﷝l���wJ�<���8[�ш��7�܆�<5N����p�n���c�gf��x����X�k�'@�7H��
�~n��歞�"���K�}��(�ꅱx�T�|h����ǟ/���Uv�_�%*V.59d���g��}������g֎2,Sw6�����=��m�[�7U��qV�ę��*I� m�B�qZ��*+��b{���=�U�}Y7��,���Ȯֻ9VM����w�g�`�hA!;�����t�Űz���|d�٤Z������0�r9LY�T�Tnz��Qޜ�i��Y�vkg�u]r����r 0�[A���>yW�q�mxL�ǚ��0��>8��n��9�	�/��0ֺY��u�oC����_b�z���9�E��v����v������B��#�;<�Z�а=�U��Ge�*c��4�1~��x�Zx) GR5́� �i\�w#��k]L��?5E�0�2wT�Pz\�� �� -n�C`��&���64�z� J���|���fI��3B�Pʄfn�1?⣭�>A|�S�0*�?q��?��T�)
�|��Ք+e�el\�d@�p�/Q0���i��.���@���&s�zKyOY�w�Bt��.�OY����,�%�U&��I��"lۢ��)�4���=�x�� �Vf�������u��]�eط;��.a�2 �(_Z���!�Zw&�&�_|��7d���|L���P�7y/���Zės�.� m~�k	cx����]����o�e��t_�,q�ѿO\�Ȼ���C��}]�ϧ�1f��nC|N^�k��J��>�g�����,]**T�����4?_B�v���s�ݟ�^�z� �UǹXA2�V�}/]_����쁥�t�v���9���+�Ҝ(O�l���G�bY���M�KV��߬�_�Ο�}�²�I[�Ӳ�QS����违�p*�s̴z񎎥�CZ!��^�U�kl/NSh�u���b���/2���ŋY�����4��.L`|�q�8��A��C�:`����hjȸKţXԍ�Q����]yn���۟1�V�0m3�Ln��=�`�c%Z�v���D�gL��2V"�]�2�D��������f�v�l� ?\`�c�6���4e���r`(ݑ�V�¿�ߊ���2�뭬m��U6LW�je�b���H���AU.�u%h��S�*2T�"\--*Zr�e�ƃ�I��]�N��B���A*9�"�R�0A[K���x�)[ɲ�)S��+M��C��<��.�T����Ȣ�}Ú�3 O�Z�?~r���@�sd��֡(h�dT���IZ�H�f|K��lg����-T"1�2-胲s����.����{U��9eIQ!��Go�\uv*'6*��C��j48doC�A��mY�G���p��v� �����I>�T¼�P�^�$)���K~R�V ��V�$��}\A6W�	�����|�q��O�Iﶫ���q��|�a㗸��v�6��,�0l�2~I�����^��}�g�.Gӻ��T���uz�4�︥{'��R
�q�FZ!�u�E�?�7X��Wb�YJ�z�ï��&O���I�M?�����K�4��|�6�0�����.�c�������Ef!��#��c$u��!�����M�V�-�<�G�U"E古q�|���*�:e���'0i�g�~�`�<v3�T֙Xx0 0x�g��Ll�����l�ƌ���:��S�Oɕ����TJ�֮+������(^n�����,���GߣD�i�#��ii�x���q;N+[��
�o=pY�,�i�֭c�u/��� �*g��!͌�Կ�.����:2�8�2j�alv��Ǵ]��QxA��ڤ&�ُ�b3��K�2�v�7�<�)�W�f�+����
k�ʴ;�V���!��5��>[�����7�T���t�0l�؝<�
�����D���~���d���~H�&Ӓ(c;�����\�\���T�E9��P1flyQ�E�3O�O���`��T��e��36j-N΄�G<)G�g\n~�h���F�Ez��l�y�M�}5���lV�OQĞ&��X��?e���������u��ʼ��ʥ��4ʫk�h7�]>F�K�'˔{/S��(Y?��NǗ/_Dq�`�V^�sʤ��&�~;/i������N���Y����S����&�97�]M<�<���ך����y�Ss�6g����_�b���Xl>��������K�.�2�L��ٖf��_��o������ttg��<:�>�� �k�=7S��Q� $Fg0�Q�p�k+z���P��i����1��0b�I�*��Ø��O�x��MG.��x����çh2v��<d�����e���q�Q�zk>��ȩO�`L/��n�\�?7�M^ĕA����w��c��	�J#3^b�b���!?~�ζ��Й�Z�Kߟ)41dz]�M�_�,�E�E�b�bШ�]*�N-j9�"�u�+������)��c� yx�7�=������(3��Y$�l��}��ga���Y��Å����>�-��&�dR��b��cw�g���}�M��*96��B�NK�L��"����:F�T3sj	F�{���B���˩.��V� ���P�e3��m\!.��\�Lڻ�y!��#�BP�����xLG a���M� �R���<y$��ھ&A�|��]R>Ԑ<��*{h�L�� l�h4�UoKU6{]*����_*f*-*/2b�]��@O~���T#���N��6�Y�WB�K�q��4�Fy�<�"�zM*�k��?x.M/� �,`��_�q���sq�"�V���������wH��Ŕt�.%�5���t$	9��5W��٩UC�������֎O��8>�^���-E�p~L�ī�LĮ67El!)/�$���/��4n���[f�x��/��ߖ.��mں3��_�;�g��������po�o:�JK؆���|����#���ڝӶ����Ӷ'�j�hl��an��P��-���vz����5��9mG:	M����83Z`Ƅ����Ō�ؤ��F�;�2�X9�痲�W+G�/o��#�l/K-D'��C�7,Xw��/��B��2�@N�)�U�O9�����2�w�`]���O�uh�n���,bq��8�;�,юV �g�)�`�J1r���Z!t%9���)#it>��:q�����$|�+�V%�]�(`�5����/����Qz�~!{��O>@�r*xy���#�gO���Z	cY۵���G��l��L��/��Ơz�.��z���r�T��Dp,c�rǾmK�cM�c�!_�y�,�~|�'�I:���*��Y�o����k�aeJ*��0��RA6���P����/7 *!�9l"�(,«Th�RFUw6N�4ׂ�H�AN��ҒY��£�bF�ɩ�Lm�F�Kł�[������<x����V�o �g19J�uŹg�Ei�	��+����n�qUf�)��Z�.�*e���sG�4�$Z
+��Wt�9�=��ss�?ʗm陃��v�d��2PQe��,t!eI��jy����\�}��EP˨f���'�-1:4Tl�H�Q�T������ڳƼ���ڼy�c�^����/�t���c3Tƚ��+?�H��/qE�����3��3�6���D�`�F-��p˯�?ŕƧ�\�ݖ�m4����{�WӺ��%N����VU��K�q��8w�mKo��o��6|�f��7�v\�3|�;�AiF��oOW��*zK�ꗖy5Q���;��c�8&c7!�*_~^υ�~�g�g<�m�n^�쓲��8��¾��/�Fػ������u��7_���J�/�*eY��Dq�{�0o���޲��2���K?gI���p#-A�o?e�~��mcB}t���\�
���HCh��3/�)A_̕�H��>WX��<���{� ���/U���ߵ^*`�D����~��!�ٓ��W/������*[�7v���(�OT���qYC=֗�A�DW��G+��x������F;	�*N���2f u�z�c�QY'�:��Kq�Q;d�� ����_��7DY�˚@ۉJ`e�)��-�7#Z��h�����*������O��Ib�`n������U���ǫL�**L���)��YH����[ 
Q8��xvi8*`�X�L��й��c�X$�N�3�;��3gq$y�r��]C��Q����L�w����Qf��xe�2(��9H��xՕ~R���:<,�Qn��􄻆�D)~.�>�(��ț�0p�4�7��%an�O*� ����$�>�<p�M��88ֵȞpn�>
���zw1�D���MDrG*;kp�֍\��'�U�̙Lv���/������g]�8_��&>�/m�v\mиkW���~-�s>�owY���%�ܩl�븛�:}v��eZ��y����o�}�M��|�M���M-�K��y�<5�9��� ���MZ�mB�fr4ߙF��4�5���	lK��r1vM{���Cn��6�l{��`_�$5~��%II���6�2�	μ	%\�%�[&�;-�06�,��� g�}��>�<t�����]�b�U�lPs�펛':\������[�M�/q*\�PfF@Z�/7%N|`"_��R7W��>Hi�ВFC����^�-^��6Qf�a�)_(�QX3���K���A�(_Q��ia��x�z����ųG���z���ol>}�$�!w�ʏ��}_���ZɸC���\�Gt$)��I,q�%��g�r��}�q���]���X��m���.Y[�T�k�,{�`,g:rw�#6�k<~��M��i\�B���`�}$�hP��;H*)�1�}�ͷ�������o���#!�4e�s���l|FH�H�#_���V[=:�][?ף����,�Db%��9������y(gr��l7�'>h�aT�� �O?�!qv����ߜ�����w�����lv*0%i����R�$h�h�sx;!O����l��$S�Џb0Φ�2�;��(s�b��J��╊��$����h�qU�m�� q��4C^��By	HҺ�LB(�4�Y-��ጎ��O�r�����Z<O|���]5��3�MK�	s�G��ʛ L5��J�Ûm��a[��!��4��iE3�)�z��ܭ����]E-y �+S����m�p^	��?�J���gp���7�σ��`n���	f�o~nr�]Ҽ),��}	3穿�[�w�iu�&w��y6�#�L��:}�n�_���+�Ư����u<�z��&�Q�4�ZMu��:(�զ�ަ_��_s�q�c��_�ϲ7�M�^�%��U�y
�Dot-_Y*,�V��f*
���wb{�}V���?�-h+W�� K�k�\�!yѧz��O�:e����/�c4�����/��GXsX��ұ>�������QB��a�� ���U�%F�qb�(�@Yr-��[�:N���Ҕ��h��h$�������%��u���->*���M���9Ψ�9��z�]�v����b>av���ѮJʭ���p�����կ�}�z��d����=�#gT,���$~u�Ǉ�k6/��[����k����{���[Z��Rԍˋ?ye&�2]T\�$*�.zc�m%zqo���B��1������;�'(�*���������
�I��S���М�}t�|닯V/��M���KCE�����R� �ʷ�U�R1:Uq��a�8?�i�X �w�yN����ޱKP���a]��7�(`��8%ex��U�S@#��T�NQ���q�Ï|��~Z���t�����h�.:?s������B�d��-S�60W�E�d��,�����G���I�e�@�T`M�*Ǉ�v��^i�R	��Y#�$,i��m�V5&�0�!��Px��A+���5�J$���e��4�hy �֩<�����CH�P����1[�lf1���n\�o�m˫��#<� {ῢ��7t�Xu���0]��.|��y���T�.���tg��]������G�ߔ���7\�vx����x�7�l�5n�5��<5~ô��s���i7�U�>3ŷ4g:7��fƝ�o�M�*~:��L�^���ND@�<}o�m|-C鄖�`�_�5G۫t�k��%6�h�����eW�L��[�����5y���'±(���L�F�y���;v�����|'�1�����H5�0�v�����0q���t���  I�?RS|�DK&�����/� 'C��h��_�Ex�8���#�
V\d:ю�&���������D\[��\��Z�T�vY��B{-�Z��(���hg�=�7�z����~���%q|w�q�������y�AY;������B���շ�(.���LQ�Y�m�UA+c@�OyW�I�!�M�ˆ;�O^����KS�\r{���a�`����s6 ��pt��Y�H3�T(`���[%��_�)����O���W߮�N8�E��cC��s�Q�.B��Q
���Cu�Y(�����L#E�	��ؾ�V��	��#�>�G���}^Z2�����T�0���|���P̓���ɹ��*{����c{��ˣ�����؛w����g�ʜ���l]%�]B,8�����4����C	�CATo�+���5rQ�V��;��x����h�V���8�l�
`�:�d��e���7���Ɣ���Y�դ�0�ÿ|W!�ꁿX�Hܡ�*NQ���C�/�7���.�b��L�� �m>*o*`>b1�܇�MF�\����l�k�J�iS��I�{�9����S���G����?��)3墜n�Zn���&ZMg~��G��q�/��[��'|��ov�f�k�nNk�vMۤ۾7�m�ٵ��,o�M��f����3����6��Ҥ�����g�r�w�u���[A�#�
_<~ť��D��9G�9t�|M��]��M����}�a�/�<n-�}u�tN9�|���MM�{�4����c/��G�<��������w�kH��/�x��IQj�6��b������?(Z�u�4�!%<�D�u>L�&�����
/�Ƌ�CXY���ʐ�R ����]�F8�6�`�],_A�y_N;~������������귿b��	�HL���]�zr�bR�yǸ��os�c�p�����<ɇc�u��<���t��o��-)D��˘P��!F��m���Z�ę�c�Ӡ���S�������R�1^~���[����ʣG�W�1D�.L��>k�6�2c�m��C���-?���J��	�<��a%Vc�.BwJ*q��#��aD�`��䥩RA�f����[��{#M���'�U�2�,�1���T)B�z��0���1/5�G�~������1��x���|F��/߯��}�E�����H��X�ܮ{NyT
ɣޞ�W	��FyM������O��r��iē&zH��BH^�M�c/�
緼����%���R���+�(^%k&
�`5�z��H��l���]�*i�V$�����m@��6�����-g�-�hvm6�kz�'���R�"��e��Lҿ�?�e�nw����f���?��6:7�w��nÝ�|�
�4f��i�.M ϩ��-��h�����o�k���Қi/�:�eY�psx�mt��D4�L���<i��+e0Sˌc�iO?�ڻ������8	�7����=�W���̌���4r����RrX+0�ӱ�:$�3�П��ZI3W���/4qЯr�ej��,�$R�x����Hބ�rr*� �x�p�cn������+�P���H8��y�wz���8�f�c'<�}����3<B�������~�b������g�OP��/�P/��cB�$�9$�jf��XZ�f(`��&�E�Vo@	Ңy4���X{�wr���7JaG�}�%ew&H�
a꙲�LK��m *��U.�n"B�ӍQ������#{��)a�IW(��<\=�m�S�u��3G'X�($@n`����2�1<9�d�E�|w4���+%EL�f��``�Uk�J.>�]��/����
����Ap�e$5T�� �n��}�hZ�<����:��G�&�>�����o�?��ְ=��:ek�L�N�><~��.����x�G�c�������o�BT������ ��X��%޸���C��3��tr�(�W���<@!8�2O�+�_�W�bb�G$�k:���_�+��7���J�4@FAm�L'A^��7��Y�V.��S˾�<r����?�]��J]�\��������}/y��A��m�t٤��9�;���}�1�LsN���&���7��a��/���?����j 3�/��K�M�������4a�x�_�����?[�&��������~Ɋ6�ê��4��:g��Xm��Ve���.�� �ZV��.f�Nؙ��X}��%2o���:$NX�Q�0`�s��e-���cՇ׳�(�n�S�͹�J^�g���AFR5�D	��KX_�G��WQAN�>��i'�c�p�%��G^��h��5ء�����s��0�2n����MW�o�z��_��W���7����܅B津2W��x�7|{�o�"|����٭�����X�>��J�>;N/ر�������ʘ�=y�h��D]�S\�NA.u��T�K�o ��B��86��b�Gb�?R�;�����o�^q��	e�3=�9��㜳��U��Z��S����`3�|T�s,<����p1��>h��m�Q���<�U,,E #�_��u^	�Њ��0�C�Ρ03��V7ij��qϬ��$�J�"�9WCK�B�"�Q�>a�K\]u�n�W'�a���\]�L9Y[���=���T����6$O�ϛ	<ˏe��\Bm�����W�%�S�MCb�X����+�@xJ������B��A�$P�=�_9t�@�'�|�b��{�L|�Lc�G�5���[�J\Y����6�\�h���A�ީ{��B��b���a��M����Öy��i�-�����ujplKk�/q�~ӘÝ��7�Mn�0}�k����aZ�u�ކ�q3���tt�ٖ�s���]����a��R���Fc�k�K�t�/��L���{��ݔ���z�7!���u�����Q
 ��[r��0k��~��b_#�(��ɮk��'���B�������-��ܛ~���Bq������z�M�d+��j��f�NB�i �R�0���߫c�'J䂸�V���G��A���:?�!Y ��Q�x),(\*���{ʽ��r�#G1���y�l���|����~���w/9bByyd���*��|����Y�"�v��hQ��T����1 �Bm}g,�,~�:��=~�'��-�G�+JP��
Z�[��,�%&l��ײ́�_���<˓�P��������_',�:a&��u��>��^0��(`o�.]� )@ֿω�$��y��ϫ�M�.�F��{$��\ԡpɏI������p�y�!GZɸ���@��0j�&�J�x}��uB�D�1-�&I���2xG�%8�/�1��^� <T��o^���_��Z�o��g�����.�xk�"=̹m�J�3�.9K�I���z���
�ѯ��Z?V� �����Z�X�@;�n�X+�@�7����RdL_ު���m)�
����[��мI
��Ao���U���YGM�V��Um�ځ��z|��A�l����r�{�rv�
ߑǦ�sN]�9n�ߕ>��~��k�wܧ��v?O���M����M|ܔ��K��`缶�����.Ǘ�ܞS�6���w��w�}ҥ��6-�:f���� m����5��I�'xב���=R�k�A�����n�f_�W�	����Z�;0^8�t�!Q�rVf�81"��b
Bѷ2ϱ:�~� �*~��7�3x�1��T▽L��z,O�pc���47n��k��N���$�X����jk_��h�B���uX|��G�yﳹ�S���߮����5�_;*g(1T���=F�'N/p��gϱ&��p�L�1Z^T�2!0�X�X#Jϰ���3֣;E��ͅ��7)��g�b��
�0�'ĵ�d�st�O/�k�d y8���V뛚J�7|���͆O�}B����Q����f�L;2����p"ķ��oY��{�*+`�] ��%����fM��,�R�*WV�&H�,�͞ǵ���l|Z�,A�J�j ��(9�V=��Z��A6 ��th�}��y�apw5~@!s:�>\��b���|���x��C̑�T������=����fJ���:�vw�JA�g�E�����Ѥ��T<��kۓ�~��P����%}��@�7���D؈�R�6�oAD����ð�B
�:Y�UW��M}e�����E�����`%��!���W��]��!��*eʭe�N���aJ��jM��,�hY#��#?m��+׏ddI�@kTÖk����2�T�%|ӹ)�N_��?�n��]i6헟N����g�7�e���&t��j����[�wz�3/K�%O3윶��F{��K�ͻ�k{����a�C�m	����b����L�,H+�}�p�>���z��N��(b�y��p���;�3�i�Dn�2q�2.�U!���^4c(���.\92;)HK�+C������@�?�j$�����:��&��4�ʵ�V�P�>c3�񦔜4��@�T���f��g��4�5�o�z���~���o��Xn|#ى&Ƙ�|���;�8|�{<��{���գ'/��3f``��B�c|�@U�u�Cט���j޲`���1�0�Ü�C>�Z1u�Kx�J�Tr??9:ʺ >��8?-��*�m/��fX�\����揟��a�Q!S�*�?���������n��{r����X|<�Ó�&r�p(`*MS,�f��V�(~�����d��a�$����
p&9��&�"���v�	5a-M��q��N��9��b��%~��]�o8���m�*^0�<@@�]�6hdv��8�o��B);���Y��?q���ܲf��瘬�� Gj�>Ծ�P�-E��dWqi�;����$� ���%D���&&�twd]�ɯb���ͻ<���X�+'(H��r�h'l��0��"P��딮��֑$U�q�~vA�x�L��<<�G�S���Z�C��[�W��BJ�Ed��o��L3��_�ܖ����7ћa�/�m����F��4�Ou�������)����K�1��>�f���|.�m4�r��Kǅ�<�ןX��_���s���zi�ﲯڡ��Ό7<�YB������A�e��uA��6fa�/X��~,b��2����� �����|I��\*`Π�㍙Vf�=�x�lZ�W�q�0��K�V�g5L��@�l-{�*)$.A�O����,��Ͽ�ư1����D�DT�q?+�́�0�b�8���ߡ|�������8��i���h
:Ɵlƣ��(����w_1�?"�Ml�3xN#2��a�L�`9O���r�=p�����S>��O߳����[�5��{�GΊY7��(aZдn��k��	u����ܮEs=�왵9:yGQ�<�A��I�l�����]T�� �k�; \�~��gty��7�>�p�5�yD�����o9=��W ���B��U �N�jX��*I��M! �Øʑ�-Cu��)�=-`jLNj�;F��c��8a��P̀NM:���_��5g�4�+*��iNy�q!>8���~���J?�̶Q������ϧuʻZ��s���9���i��a�?��i����#DH��3Ïh"�,zk7��2�y�������>"E[�P_�QUI!��zl-�U	��%��ж�x�'k$�d�����?J�F�%�i��.���U��t.����F|��潼;�n��a#��:�0�������r�����t��q�_�9��o��3~�M�q�t;��nә�縙�9�&x�ߙ����v���Ļyݖ�����2�S�ҽ���&w?N�{3��-T�����S;��d�)�W(-�����H��h+�j�#{�K��1P�J��5a��al��^�ą�^���0_�sn�*IՐ���"Y!�-%�&���\PH�k8�IE��h�\p#��|G�k����uK��ı�ST�<fB%L�/x�1���W_�|�j���2�Č��F+Q�3V�����3U�9���Z�b3�JP�uz�e`GS�%(�Ld� }������)G]p��3Z�Y�3�\ �4UOu�t(n�^(�փcS�>��e��ܨx����O$ez�dF��P�SIk9V*Gj�^�t��#���hCtz�F4R�yp̹Ǽ	`ir���t����L�_��n12h��4�l�a)5e%G�o (I�������i;�Ҟ0���7�+�>����=#0���J���d�K��7�9�;���,NeQ���O��5w��4;%����P��R9���oX���?oOLAZ�[�,Ѓo�T���*��+>��KO]6t�B�X�&eWiM+A�ǵ1䡵��ߐ�r=T�V\�*�±$8��OvU�Y`�m�rUI�mC$^e�:����D���pU�/8�O�6�-^�g���˳U����Muv3���繡;��:���?�]�0�e�z_�c����߇f�{��`���v�g_����6������a:|�.ޛF�m˷a�m;�t��g�����isz�-a;��K���5����75�P����y��)��`v_�,#o
��ż����5ϼ�1h�ZƯE]ˆF	g/4"$,c���BƵ�W-r�7x���cv�1o*y.����a�4�)  @ IDAT+�� ��L�p��O5�E.���㏑�@�&�A�� 	�q&������	a3W��g>E]�JY��$���W��9˖�Xh�7��[4\�s6��(_���'-���_m�bM�a�]�����p���}�}!���G!M��9�@���X,��$�~>~��q������՛ׯV?��w6r
�m�}{̈���̸����v�SZ���MQf��˴N��*�ʗ�vq��[�V��LYB�y�X`���,�]@�W0j�.���ɠ%s`<8��*I,Tw��뢠E��Z
�5�,��z���ؐ�ő49����w�b�r:�9Y�${���0��z�5
�L�^S�n�W��2'H���9��W����M��Pt�YF�Z�H�mw�LW�������_������ջ�������p-7߳R�$�M|`���!��ʤ�����5�*�^1@懣��ZIn�!m�p���E���rI�[@y�D��u�ҋLu����xD��.!oe6`�+W�#��%?ah5�:_;L���\6h!�NѸjS�_�+/�݄��N����)n��q�Ꮏ��g����wvoʿ�����L��}ݦ{��>�o��o|�Z��F|꿚��7�+߻җ�5����)~�Y�g)Ý�ęÎ�h������<���]�'_���E�����Q�1�q�1C{���	;��8��T�H�xJgi�U�����9g��V�\'��qlYsd�%=�K�Y~b!�kk�6�����B�?h���ˡ��][�q�p�5MrׯM��7 ��Л����A���s�)������4=�;���z��m�d��/J���9��=��9��Ca�|xX�]�#�N��U{p�R�������]�=;����NcUK�0������ӕ��v�?�2��QUho�S��Y�-e�I��L����F]kq�T	bKc�@>,W ��\(����z����9����]p�W��f�f{|+&4i�ry�����7 �������(L|9�+����$x��]_s�W�?��
�X��JAQ�,-��}�pp��nu��`��P��I�9��</�Xl���v�!��X�~��_��G���O�7(�>��er���w��璝_a�D	˜~�
9w���4���0�oԔP�D$2	i�)X��ښ������::���FJ��T�%�x�(<*��7o-�?7X2W���(UC"���=혃X�i����A)"/o/��*��F�q��1?Xy��5����[�t�Vg�_e�G�c++E����G�}a��������}���_?�q���S��a^�.��/�5�v���e��7����<17a_}�����u��U�yl�6�(`��} ��;_��oe��)2-� ܱg�`�ӢE��M�����ٗo�y!���Aޝr;�s<�[������YƦR��;J�cy8g��}��&?p�� v�5��<?I-�L�F���7?���g�^5<�,�1���� � �R­�nD$�Z�e�/��#<y�t��'�2�����ʏ{Q�F�>�K��m�+�8��N+Gf�c��k����l|X�:��x��R8V�`dq#Ż��W�|b
uY+Td��H*��[�)���.��<@9D�rm�
��w�B�8h�BJKW�q�R =\r.W�b3B�="�0b��L#n�RȬ�����*��p�-�Ft���7Mu(?(*W�	K��ątl��F�Dо�-��,�c�֮'O_��`�zĎ��XՌ[�*OG2�#�(��Ï��m��2u�^�b|JBs�4��<0��AR�^��oT�NW�񧿯~|c���y����i�|�b�sv���f�F6>0Up=ӥ��5���#t�֑kOŏ�A�PQ	� m��exs�	6h~H������]N�a��/���p8�j2�Gj�U4m��զyV��|4�P�������Hrr�WxL�x`�c�~�ۄFv�����ĉL(MkN���pnw�is~7�6�m�]8�|~ߴo�o��ӝ�f��������^��k�7��
�p�ϰs|�������iw��0��7�2�����i��y5���af�e�?4&wN��l��%�蟈���c�9f��-�?�f9?�'��%�+X�UKH2� �^��RʜӔ��1�%�����v�Q���@Κ���򐿜�Og���'�q��JX�f6x���JD�Fps��|���B�j#^:�N1䇜�٤x=3gt,�>
���Ϊ�@�������b*��r��ǡ闙ya<f��Ɠ�� +㑿�]_���K�C킍~R�ji�AOPOQ�v	�]
��#E�xDG] 	��j�t!�aJ��y�)�5�FP���ᝮk<O�ƀg��[�d�Ѓ��Lv���O�4�Xu=�a�O��AEX��⒦��4��"8L�;D^a&��e�{��׫G�9������|���9x�фk�-> f&^f�c�T�<n�7!ߝ���;;U��:���(m�A����������L����j��H*�Ʀi�T$�$`j<�oŭy�E�!v�j3.#&<���ʗ7�|@��K����]��x/��v�c(����c�����T�R��3�x�t=��<0Կ[��mp O4�_�\5�q�>�z���2��͙�t�Uz�O��my����N�&��J�	���O��_�7��:��z
R^���)��\��=�%t���h���u��ug���83L�lw[d4�i��w3~��8��9�pw�o�6<���]��O�v\{�<��=ä����Kj}��>�?2�?�)�"��Ͼƾ�����������qo]����q���(�����u׻�=�=F�|�"w�;��/:��2>�3(�!����=�rk���Z�c��A��B���)�)L?*�q��T��-׉U�d%!/�SK:!tH%�������c�L;p5Z`�:d��7_��꫗���r<�ؑ1]��:���,RO<���e�I���xo�a<��O���pU�RfQ�����Z�=�@k�<�g��;��@E�s?UU�X�D�Q�!��m'
�6步-���U���Wl~�@�X~�Y�)W[�$�b��L�v���۰������Z0�^s�æ����Pi��jE�滛���Q9f��L������ �*����{���C���R�J*�<H����U��')�s���=,[Y�E�q��S�W/�����|���k�hLWh�V^6`5s������7u������7m:q�G*��2�fBJ_�뺬X�o|�����T�Ƌ����mJװ����[�bs۩Xq�4���qFZӷ�U�����
�i�����j�vZ���T��YX.%�Ts�`�r�������&L�����B�уŤ�	�v�S��<>b��_6�����U��������������/��G�v|�u�����W��",+yB%�Ս؊�@�.Ü6��Jo�5��p�J_�����N�������tf�ҙo�Z�3�v=�IU���!]-�����鯉���U_��9
�M?�o�f���JC�}[fk|�9��si��sO<g�P����	a#-=�e�:{�b���X7�/�goO9U���(#�\�,�c�����1e�$�S�$ho�k��v�4��N��{$8V$�X��ї��qDP��њB C>>st�����S����o��<��%㹷/�7��PTx!�>ߝ�~�Й��,)_���闕�z�t�}�T�U1Ѕ��ϸ�@�X��WlJ"�㕂�j�E�!k��Y��ta��������Q:^�8��xфF� k�BjL�E]��l��G`���!�u���M�TJ��,�`C��s-���a+�Gフn=U9�ʁ�T�����-��"mBu'�B��G�5m�@�\Hog|���z�������>z�z��������O�����iU�`P�v(3՘���z䒼�Yq��T���1�������c�E��Z�7��bcY��r�7�~��/I����쳁Y+���*�c-��Wot*Hɞ���ھ�<@r��iG�ã5Ե]vnʿ�l���&�]kŴ��3N���V^
��,�.�g^RH��KhN�?�[7�ei#��;�)����p����m�q�M�M�݆�F�a��.��t��my4ܶ4q;�݆��
����os�t�:�3/��]k_�9R>"�y�:��G���,ϜG�Z�݄��o|�N���%͆�������-9�^�`��m�s�窠�ӿ����k�pl�g|��VE���s.$��vۿc󗧧g�/ٞAh�!��Z�.b)cg>]GS���q�?Q�l���C�y���׹�����F�k�_���O?|���(Ͽz���؞���K-}a��Q�8
�G�u���l�'���o���j�b]a3I�4��Д m# ���Q�Tt���_a�N�=}�|��%E�]���Cc��X�U(�0
#o�_��@��#~�L*G.�N����s�NM�k��b�Z�p��Zs�^��|	�Ѯ3r��v&����f��*�
�_È�|B�`��$)��x��8����!��qZу�<�5R��ִ��+\�&�X��x-�.V3����e��W����t�Hr%��m$!n)������<;,���<i�F�ǥ�8��*�Z%��0<��Wo޿��3MT�hh<���k�ۘ�����<�ZF%�Q�m&J-1����#�p�Ԁ3���jY��~W�ThH	pep�*��RB�[t-�m�ۃ[�B�J�V*)�|�7���k��Ǭ�P���E�2�?n[�T���U9 |���ۮe:��1����S}�&~�$D�˧R�jI'�O�Ձ��q�z���� ݊�iw�KZw�oKo�洙�\�f��ۖ�q�l�%�e���m�iu��6\��HX�atU��mt&��7�v�	.��;�/�:���t�;Ә��v���gܤ�v��n�mxsOt�������mC�SD,z4��%΅�XߥU�K�*`.���qg����7���2���brH kYT��IQ���%ї^_4��	]����e_��H�!�G}�r��`���7����;�c��v�� ��^+����W�;��&{.%�'�F$҄�%�����a~R���DA���&O�I�t�ڮǌ�8!~��&fU3S^���#>�S�!G�sU!*ߑA�+��LU	L�k�AF؀���%}-�&Pٱ�����pE������3jN�FqK�
k�Kps%}-��5���kAg;�&G��4n5�:	��+5�6��E�(lh��*K���` �?�-�DZu�Le�t}'��O=��C:�E��ވx�QV����j1{��I�s�[Bͬ*`�i&<��-���K�F���}þL��~ ���0w(p6pc�J��-�Q�]����xRt�-"��+,A�B�\�Y�� eQ��ĩȪ ��&o��*��T��A!$y.��Q!�g9�s�pQ��IЎS���j'��uMގ�,���̃��"Z�(�}�Uu�y�f7���	|܄�to�;�g���2�&:3�O�[��~Ӯ>�&?�7��x˲�|3�n��[���i�v�Jo8ݙ�9^�tִ�9Zě�#���LcM;U�i��FO.OF��/֯y�R�ǒ��i�[Q������ʚ֨�$�wr�����u��u��?�$n�]����y�<�Q��ʊ;#O���e���������iO�U��z�мТ^��HS>ֲE��y�I�r��FD7I8���&nUQŕ�R_A@�j��j�!Xm��B����"�cd�%���^�0��:O#w�K��7���� K����.H���p�$��ԝ� @����5:�Z�MʁR�=��0��[���u�/�M�u����ɒ���*�o`i�&=�@M�i�
�!x40�X�Д�]�� �@r��7ٍ��
��� ��}]��R͉Z�"\ߒ̛
�
��)�����~����i��� ?�z ��P�·�%�_g*�#���m�L��oh��z�
Ȧ^ء4(��MM@�8�.-y6\n��9P�7NI�:���ׄ���zI��חE(���9�����O: ('�[�X�RyN-ad�Н����W�xI��k�D+�%�2\r���5p_�F��g�����-�L[�5�g܎���Dc	{�mi3�O�k�xs^���kwN��NkW���N�0o����5����p<�� ���#�G�7GPn���Y���tc��#����Xe�����E~'����<
ʃG$��E��ٙ����x�Z.��c�s�D�]�;�0^L�+��1O��t�Y菝>T��c�1���)�{Xg\�OF��#�5�,��|�n��?�p��Hz;@R%��+��N�(0	3�����PC��Tj�M��gL�-�����O�d���D��Mb��פg`3�pl�FB�����C��!��YB��T���R�I;�W�ռ�W�6�����p����6m�^lob���a�PU�xu�O+��
$�WV�h\Q�(H&��g#V��i}�O
�@hT�`�	�:T��MaI���Ĥ�\}�_v�Y2a�G��`x�ˊ3���<�ᕩ8�[s��2�$-�FkTU�(I�˟���˭T�WE���m8s�Jl�	5.�E���1�U7�ip�*%�^��o]��u�Rv��E˩E�~Ҫ���7���c�"k귺�R�%�(i�5���#cAl�"]���W��8�0�t��0rW�-����������|n�6��J�inß����83~�iRic�W�?��9��d<���l�׸%�g�����|.y�ex�O�٬��{�f���3�
�Z���E�핅����Ur������	�9��dL�Ū���������0zzҾ�ьvg���x�yS���`�`DduO��<���`f0\� ���w�7Y;����f����+3L<f)�)�Sfr�Iꮊ0nqt�F�Wm܇��+˔�%��ӟ������p��{>:}ʆ�s�H&��?�;[s�Y;#/������f��lG���ӕ��z	l��C3qZK%M���Vz�rKh�#,ĐuI����d?\�ſt�[�.�Z,��Q
,��C���)x�K0������ Ce,�������)Dq&��oyk$�)�z�-G�k�+L��0�+c��;�y)��Ŋt]k��bu|g^��֙"IJ��j��Q@���<HgL����zX@.;Q ՙs�}�Q1v_*k��讑��\>O���s����1�c,=��6#/TN|-3Z>��Lª*r�/���J^#�RQ'������.��-��(���;��S�:�Ȋn:��=�2"��E"YG��2# XN5�gXx��*�x�*����kɪQ��ѻ�
� G�I/�-ݴR�Zө�_�wLZ�/d�M4��.�Mz����x튧��;]�;�-��6q��w�;��D�ӷ{[�M~����M�o�c3�M�7����N�7��7�M��&����9l�ͳi���ܙ�17�	�z��4���x��E����ݗw;���Θ��3"�[�5�\~�ЏW�ν�a�[�J���l�5,`��6���AVF���=�����F���}��I�N�0g�"�j�$i����S҉�`�Br	$`>��zP9^0��X������N�(�B-���Q�D���o������q��د�`e��u�݅g��0f�P��@0���^�&n�����R� ��q'�����'T��Rl�nO!�3E]�����m�5|��
�i��Ke.:U0*ށ�����C�glЅM*Aa,��O�5�����黢[�52�A�e�͚l���SS��'������6��"5i�B�bY�M#�D�e�.���-����2���?ĊS�:Ҵ^KD7H��q�MH��4�U�����ꒋ�\���L��ECUc*K���&�j��J[s;z�����␵�GO�d6-*K�� ��_���:��1D�艔C!�}���V�
ik|ˡ�^��@���~��%�:��.������_��Q��H���s��-��s�ޖ&z�"v�����T�=I��&�[�5��a���[�=���[m�I��3���þ�|�����:�a΀�g��� �/��L�����齫��ۯ]��=v�O�gL1�=xt���̶���Ov���s�8�Mgǜ9���OE��v"_qW��k�iA�O�Pɢ;�򊺆΄��$ޟ@կ7F��<�g	2�ҏ���RWM�BN��X4v�)'��o���[S�T�(��&�t��&w�u�x��!F���d��O���Yڦ�}�`ͳe�O�縂���6�H�$jIG�&�(j���)r6)�e�s�a����3����0�^(�� <�/F�[i�nc���� Ĉ����c$���Ҙg�P]�`}�'G�'�=���U�lě�(���Ě�Ȁ�}��_��&e��uQ�J��^����$�!�嚾��H�ȣt\B��Yϵ���b�i�1ˈ�Lҡ(��u}�W�'{�	'0R�߼ִ6c���0َqj���!d$?k���CW�W��m�f�j�uhs{�4�����6
��8�)�6Z3l�3�o�7�팧��Rc6��ܛ�����\W:�x�47q��7Ý����6���$��bi��uw���H������=p��r'�	��T{�y�Y.�'YglR34"�˜��@�U�ѿ���
��XuWZ�;)���Ғ��˛z����x�p?狹�x��v�2�g�I�d*�2"�[�d�����D�r)��������KL�TT`�S<%�v�f�w,w�q�4%1�Y|�����E�~toC
 �;6M;oҙ�R7\�����1`�m"�V�?dR���L��̼@�x���d����1C�݅͡S&�'`d���m���Ţ���A`%Nm0��-S�f]MK�̔:⥸!m$��$'�x6~6o�.���H��/�{E4�+��Y�,����w�#0.Ȥ4~HW�F�f
��8�o���g�P��&Χ�j4q/z��tE�O��J%
��<*�eD����{gTvR���}r���+
��锈������s�Ζ���֏p��K州(��{�cgH#�)"#�� `�kd���u%�|�N�|uk�=�#��z�>��k�-�MkӝQy�;�QB�yن/�����:/Mw�ݖ~����ߖ�����-�����8��ތ���W�~0�e����6j܌���>ڂwn�ҕ��KE ��G�⌋{P�[�!_7rٮ�g��r��Y0)�-��i�Y���M�65S��Dv6>e�ᣅo�RF��;��'�ߌ�|V�C�3����r�9��9{�N0�N0�NϘA�\7�y������͐0��W2R�$��F�B�0&��4tթ�Ò��11�M�yf�8p����ԧ��sv��\^��r�O&�1�k�(ςt����୙1u�o*9�Lm"����P�`ƮN�� ��45�.�3y�y�B>\��/�������pcW�3��wq�9	5�r��V�
[ީa�ݙ� t��*�tC.�kn����Xo)�N	Vm\��*�N1�дM�b�5���!� �D;*�^z�`���n%�{�Oj�ʮ$mi#�P��e/��JjP�o앢�*�ǙZδ2Gs8�|�)FZA,>�V=zΎ3hf�^���t#D�*��	#?wc���%��R��v���1#%�ѕ筈f`���/uo��:�����LK:McFlX����f���[ަs]��#Μ�4�Ż�Ƶq���Jp-��l}���f>f<)t��յ��N��r7�ux��w��tL�<�N�V5���.e��f{/B7���%�H���0b<����z�E�I:�jDh�d�4�� ��~�r$2��V^$��h:��'];L�I�⾤D�!�!H'�|ϑe����L�Ȝ��e����|�q����+�/�埸�H\rU$ѥ���G�v���BS�1��I���>3{������D}��۱B�e��r�̃��tQV^b��8��B�_���xGV@��ʐ���.Ks�'�*�s�<V��=�s�(`"	H�F�兓%+@�]����R~�E�
.�.h�H�D���Wh�w�T�o�S�D�o�&,S���Z~ڠr�I抄r���n��#z�1v�ia �a��5ӛ�M��*�''|�����t�Xu Fz�Zm�ȎVq���G��Ft�IR����ȸ�h�*^���h�f5�Q񷼸d���I�v�݁�*'�^�4i�9Q/y�<K���s��XFO㌲$�t����v:N��ʯ���k#E���n��۝D�����Δ���d��WwL���|����T���FS�W�s�m�s�m�s����h8������k�����t�\������/�Y5�j+W�NL�7O��&]m�*�T�6��Y�S�j�D���{����9�ڻ�b�P�+ë���/�4.jϫFY��Մ��:�����3Vgi����߆dN����E=-�D#C����ë������R�N�O�q�-�X�3����if��b,�
b��"�<�D����Ȧ����)y�`2��:�D`�{iH�a	c�H?2^ƭ���-�N��#�t:�è��.�[凰\)��l���*��]��cN}�_yS�� s�2�;4�dL����NMi�(%�cV�u���3��ֿ`;�N�k�'^+�n2��Ԓΰ�(0}7���Ӄ
_7��әIVn3(|�v�$��Xߕ+��<�2\���߯���}�n���%����E�o���"��#A�M^:�*�$|��,h��A�A�"(H�8�<G�Y���o\� ��7��>����@��d^�c�5���x��V��Ҳ�4���+�xFOW�� ��0�=��]7i�m���:����׼(Ϣ/�����k�k�+iyrg��t��8���7�mK۰�������6�<����n�w����u��Su���>yJ�yKi�o���۽	�/�m��ſ�n�k;�����	�-m-��\����,�[P6i�1��Y�n�ﭫ�}����gpd���t�C�Uт�Gi�p;�o�^ެ�`�X��R�K���8L�����s��
�1ʣ+<P֙�>ƩN(��te���c��	+7�p����a���U�U��5d�p��L�wܔ��0?\���4�|�ZÊq@6��uȋly8� �d!��~_���c^�PGW����,^�Ƴ�5�?�#ce����R���!��ȓ�[���p�y(f�>rGF�^ͥ͢~�LrWX��j��HUҍ����V~���V0��D����	��۷�F�B�G	|�!p��}�C���֫qLWr���)�*Ț�V�Pq:�|��իܧu�lmļ��Ө|��+DS���3T���,�|6�l$,�:I'm׸BR96_]�6֪`��$V��,`�?���yc���Z9=�Ɗ盐<���hD5u����N��Ȉz@yg�Q\۹˗�pr(�oZzk�*�OLvn���ӧ��N���Яt��?�_%O�TGq=~Ǌ�i�n[za3�ƹ��9r܅�_�~Ձ/+{����s.��y�2ݤ���m�w��y�q����`���]y.�6uOy���&�����ޯ��]`U�e?r�2�!�R���[��+)��_�or��~�ۇE���9S>���(3^.�G%��K�G��ر:gt��#o��n�������5�2�@���g<�����Ȅ��o�X����j�6��:!�Zʭ�~�\&E�����)P��D�q�oӡ7�O0���)�� ������<_�~���K_c2�lO9=&�=�Ya����'�$���[��-��-�H��~�F�kH���sΊNM0�5o3�IS������=���A^9F$x�\����mSSsĴ�WS�5��ւ�����(c��Z8fԌGm���aYgҤWyR)�/�k��aHx�	���>��� X��S�N��v]�rz�����%F�3`�V�KhZ�q�4����i�7c\�)��"�1VyAi�lW�
,E"
Wk"D;3&��!PU;IF* �qI�*t�+�u�y����M{�}\n6�` �U����lP~4���_::��<i�'c=S�n�c�JS��Pћ]?�����X����<�gK��;��iZn�]��v�k�wqg^M�.�g\i5��n�;nN����ޕn�&�%������NwS���["��6�� �?'ox�vX��?��R���U���_+�<�^�_(l)����M��)��_i$����}�{�.�d懲������9���iQ���g�U��Q���o���e5�'/ǲz{\e(��qA�X�����͘�$�B?o� %� .e�$Pr��bL��f��kQM"i'Q�SQ*��A.�TԲ���'����G��F�>lUC�c�<��2�`��<��0������8�����M�R�V�JG�'8y"�9r��g�1/����'���vg��l.t�8�!�p0ؔ�/d�AM|v�W��7��Ur������̬aM�]1b��g�T,k�f�B�;4,f�{�.��$F��r���-�1Vb͢X�m���n#�!2j|�6D��q��g#�//^�~y���T�*���r�Eo�j#���4d�.�f�mH�
(��T���Tl��(p�r]&� �>��$��,re�Q�׭TťhT�7I�]~������ �i�)~���C��Ӡ��P�D�tP\�;;�S��	NC������4��I�:fh�ή�'l¾+7��o�4�D���4�n�e @�NWtg�_׿.�5_a7���7��w��r����Gs�N�m|f�����Ό��:��;�_Jki~�N��M�/�-w`�(�Ն����s�e��7)���-7z��w��P���g�r�R��?���9�u��CσdIM#�fH�G^0�8^�{�~��������%�i�tQ�K�Ϸ!}߇��St�'zJeh>"��9�؝f��l�I��7�&m%�ůt�b��XKe^9�� 1�
jx~�_|��ep���t���_� �:]��Y&tA�g���5&|\�O��c�2F$��Ƹ�jv����	ċ�C
��}�>�MN����,v�v�4���kA:���s.-߬0S72uX�B%�R���G����s�_䂨 ����P�.�5�������u��oţ�����Z������@�X�-G�Kha\�v�D
>ɗ�ؒV�
_#��Nc��8j�����_/^�f�&U����>�}��a�]�Ҳ��,�K����r,�.e4V��օ^M���_�ɒ�2%d��D����Y.����ӳ���Z�P�'a�j����A;o��;�؋3��-��WY�����4?�	X#�f��{� ��..�R��䒏��.f�}�'��Te��]�K��M͟��H��.�o�3��.�q�<;�+�6�����Mw�m�w����4:�����v��a)�Mr4���4�ϴf���N��-<Ӻkڦg���n�im�k�-B wN�|u��a��Ϊ��=�:a?c��%=g�t5\7t#_���0rf��Hb����1$\�$*{�2��`�ާ̴�c`� W&��c?3.#,rH>r��*W�\�o�V�J�̨��Ûd��T0�R���� �%ird��!0�7�A&�a���z->�R�Zz�C���I���=ot2�u���Z~�Z�a\3O3���3��:���ć��7=�7��3i�4:��^l�0��s�x�؉S��&(��fT�v�!A�p����YN�dq+�c���S�d��̾��a�TT�)��1^R��p�\09	� +��5/��G���ge��}��Jt@���V�׺9mˌ'o����|�� �$� Q��6e�-*��q-�1JT�5%�7hҴ� 3oidݚ��|�Tcp��sۘ^�x���痫���{]��b?ܭ�/Q���I)��
�_�V'���΁�Q��!d���*=ĸ�Q�fџ�J9/�ڸ�	1d锥�	�oDn�X�i[�$+��C@ Wю�Ұr"D:0h��T�?��t�߷X��#�g�%����S����QxF&��}ò:2;J4s�GƑ�����Ԑ�t7莼W=�܌���7�f��Y��igՋJ�|fXӺ��Es[�m�g�L��;~3N�f\���L�M�ρ5�v��<��װv���ǩx�V�:����ٕ��m�lK���}m�5\��6ώ�.͌3�ox�M�݆�i��8�-�4�5�n��'�vX
B
�����%u���P��ҍ������0o�����P� ߐ<`,���ߧ�7�w���5�G��}@��/�џ���t�{��ط��e���C^a�1���Y�?�ԑk1��t�^%�Q���qW��_�x���FЀ�{��{�r���2�L3�u�>���h��R�i�þ]s�1J�B�7/�'����d��͇ջ�����s�I�Sq� ql�$c'����<�귫���1���Ea�M�1�*9���X�Ii�~���,w����Ty�l��Tn`�_�6�)g�!�k�s�N	9u?���C��`΄�V�����=��(����5eWn%����K�@����Q�B"���N�[s�
��b/�ae.9	��T,��|@�Ae�[X~k���_��L?��L�R#tf?B�]Qn� tz����X�QVo伤!�/I<yXA߽=^�����~��G�Pq0��k�׫��V ��R�a��~ʏ�p���5*u��f���:#��a\�B���$���!����µiz#uhq��e��C9T�a�G/T�>� ��.�z!�ӱvP6Ro~(�.}r,�&���@CL����a�)Q�6��oy5����z6�ST�ո𒶓+�k�������$����I���e>����&����3ә�)�9�o�9�M'�&L�6��Ͻ�^�7�i�v[�:��N��<�zMw��<tۿo�M&a��F���ь�� gjgx��M��p ��-���וOcJ������c�7?���g�2coכɝ���/�~�>��axI�~����E���{E�-��Ւ�2��W��y��X�s2�����d���(��6�׬��,����3���]�U�ß����(�rS��s$�o�A��u�K����b�Ӌ7����]}��U�@�>��1.���ȃ��K^��S̒�3R΄�&�����X����k<F���{"�k�q�w��{�?�L�����:`|�H	 �����
A�@���n�I�l'g���3j��ᅆ���.IC���^y՗$L�D�Cs
�%�c �>��&��՘U���ˈ��Ǹe�}^S���G��8��"'Z�'���QZ���F��'�>;
�JRr�J ����H�2�y������|�&���O�>.��/_�]��?���?��c��'��YLa3�������ʜFh�Hd�itD�p4�7���Q)?�h��bG�i��]�4���-5Aњ=�j�=B+I:D�8����-������B
Di|����	��k^f�>RG�a�2��2Ux7_*�4k:\i�ҭ%��o�ѧH��u�EDm9M D1Ӕ�
W*��<�n��Mz�(�QnM9�
�ː6��2���#�em�.�v�uG�;|�����4M�����A�B���F�]4[�}u�ɒ�6���B�z�J��!��eq�a�W�O�E��0�<ɾ�F��.u�ظ>hz+���ԧ�;�Ξo�1���35�Y2sr���v��|جqC} �i�򔫼��Ցt�,.�������wet~츊�����o :fJ�)��)���|�O�Y}JɁg��|+�đ(�2���t�G�i����y��o�7=��3�q��/VO=b����&�j��O4��>�q/K�C{�ggǫ�~�3���z�������gϾY��K�5��s�0�SG�d
:�AMX8��yo߾^�z�2{�T��4�V�l�H�bKPGS0JYZmGCXt����!@�-�K��C>1u�c��W�$�X���l����-����Ɉ�ğ%@� |A5��/Yj��r���ŝ;��u]�kP�* ��H#F�*˷T�%���OX�l�SQ�L�l6^�^�	������_�L*�
v��,�  @ IDAT1�W)+��R)�pV�w�W?��b��o\������R�`�Ƙ�>I؆U~5�� 9�FdA��4�aU&��`��P8X��:��ΐ�?3�a.iU#��Lm$���F?U�Ɗ��ǅ�?1�F�P�T~�y3���S�t���<�TH#�&}�w=���g=f}�%^嗘��<�������0�Xx���gH[�s�~��3�b�� ��/<T٧<�q�Q�����o�K��)��ބ�.�ץ7n3ݮ�utfYn�7���.~��w�Ig3<�Sw��[���w�g����_�o��p�owNk��w�v�o�v��f\Z�m�{˕�ejs�rnI��vJ�Dj��:�g��a(�[ʗ���of_�c��Z�A�n�������`�G���X��[�*fAx�wLH�e�e�4R�����G\<�K�cO��o�p}�\�l4��y[�����j�Ҙo��|q�g�8c�F�,5_*(��|(0�Py���Qw�G;�T1W>�+\����U���%R������V_�5[Pp.��6�Fg1$���1
���NL�8~8�e��q���[�\�'�<Ն��(yp��%�z���/~2�q�ٯ�w�?�(�7���S�l�y;�L�	˘�"/m��ĉ3���ʘ�a��chj�s�@wY<�nrbk\�R ��lܔ���̳~3�FPJ�Nap]��Q�Lg?nfĆU�է�m�E"5��l�NEV9?�o߯=�j��o~�zx��Լ��^�X�MbdJ�D�Q����e�:+��rg�Ύ}��8rg��'�>�p��~�e��w?�������|��|���n��"=d*�/أH6+Z������hH+�����@O a�Dԭ~,p	Qm)�C��it]�i�*�t<Q����W��|&Z*�<�k�	�@=��O$ё�0��&쟗��F���5}_J����<�z�hu�xx������M���b�{K��(�u�bc��`>��w�V�+���V�>����)�_�$w���VT��t`*�����N;�Xe�L��q3��;��g]�V>���q�t��e4�nX�\�ކ�L{�m���uE�O� ۽�Ct�M��_��I�3�F����o�~�Ʊ<�ѿ�A_J��}��=A�N�~�5������f���0��s�˙g`4�N;Vc�� �����2`�F��y�Y.� �ư(�#	�+kh:F<`���C���-{�~�����ׯ������f������g�V��11�J����%���c�@�$w�"Y���ǡC(�H,'f�D��ٽ�#D=d�8cl}�!���V����Y=}�r"�_X9=y���}�l������ϛW�˿������50l4�0,�0,]vu�����Yj��x�,���{1��0�B&�7w��?�0� +�+�)�G7���h�(g��Ch���o��_ɥHߪt�r�<D�gϿf�)�GY���%T�R��@�Kݖp�bĒ�u��?	f6&y��F,;��>�����C�R"pыԑ���T�p���0Ϊ��x3�`��ϖ�R�:p�t1Ȇ���Oj���OkY�/	��Ɨ�ﴊ3M)��H���_����W���oY��@�B9Gn���b�>K��(Ӎ���P��U^hfTV�X��V�uխ�,�b�j�m:��%�m�:�5Ӌ�s�'����k��?R��Fp�L�H^�1����^�>}���N:at�<���o����������?���T��I�S��S/\���X�Ƙ�륪a�S�J�W�Ώ�G6�D����ul�y���M�Nn峓�^m��n�gZ>�n���]���x�mt���N���ix���M���m�����G�:�3�M�M~�\����n��J�&��o>�6�M��7�m��
wz��7�·����Vc[B;�^����{Me�d�p�#���7@ '���c��y�vV&34ET�kx�ҕ����������w��o��?�g1�:�%��#����=��3�Ȩ�
'2�M�1��C�a�D��zL̙��s�7�0V.N�0B4FN�����z��S�e$d?c,�8��n�w�C�#���Iƞ����84�?/�1��a�i����|s���nkr�n�	3r��f,��$6�%�G��5(�h�,����-e7�מ�6�������×(|����?�Ѓ�܇Е	2c�_e&5����V7N<5i23
���>aS��������v&��`?b��afP�F����ۯ7	�uQ�2����N�������̀Z��k��y;D�:3�e��AЂ�� ���k�NC����z�R�;����o�z�쫼aPF�J򊰥��b����)Lg�S�4���k��l�3����u�_�]��������?�~y�t��>�9���픧��Q�I�cd�s&�ڛM�ŝ�!�b�3�	�t.�4��H\n�dZU{P˜g�?�k��E�-��9(-��'�r���+��� ����K�
��$�1�к;��\����;6H~�ݏ�o�>^���{�䧴�cf���~�R�)|@�s#�T�lL6<+�O��o�S_��/{�ȣ8>y͗z����K.�ʚ��4��T��Ӂe7��JL���"�.9z�����_"��z�u���h��}l+'1�-�ƿق�݄m�T�v�eM<��}��δ8Xr;�9�u���=>�?`v��5k�8�w�z��)����y��p@����������g儇R�h�Oʽ�Ĺ�O�k��t7P
qɹ�ط�z�	YYr��>���-���1+3h���7t��]Z�=��FV���;�?��!F�C�߳��f�'3G�r�WF�6�� A��"����&F<�E�����s	�q�=F߷?��^o�~�L�(����~�#߃t�pK���򐱀�E�7��C��ua�<F���e@',���|j\>x�^0��$���U^:�cVԱ�B-�]��4�E����1��t�v&������C'��{.s~�3}9���p��y�>3s�%�T��l�������v�wzսO~X���[�����=�=�����[0�@:��}d.9�C���\��Md ?>���Tfx���n��@��l�y,����?�~}���u_�L\j�a�f�Ac6���R߳��ǟ_����q��o^��'�K3�.v��I�<�@՚���
�OB�f}͝Kry�u)$��k���1�)h-GͨiӘ�&%���ӎ�Z�$�?OaNI��S�ӰE3y�7LI.�T��AP%R`/�s�Di$�i�
���}�K�"�>a��N�sK��z��ibg�l�p;��Sv�0^:�d=T�
��븒��,��֞�ݍΒ,J�B u�
d��o�E�S�6o�o��K�f�6��<[����m��n����_�:y7y��Su:�m�i���n�.w�Ϯ�+�����4��6����m������� �ǔΫ���˦
�&c��D�/q�b�A��D�g�oeϖ�%�h�	�V�0�q?$��8!Y�S�@���o;^�����~Y��s+��K��x��D��?�� ���Hv�Y>�;��;�����}Ɖ���2�9��8u#���Y�c�<�=0������p�Eʪn
��$ʐhxG5%��D_���c�:��x#LT_�r�Ͻ_ޭ����8��z��)
�e䛄�G�M��:���c�`䃟v��<�� �PK7�ɤ��	G[i30��-�R�[��⒬<'i�[f��L���g0��"��zfeG��p")F�xh��Hp߳2��'*0`?x�x���!�G�p�;]�����+�֜|<S�wC�;�6�����	-�K�*D�h�̡z��BSl��v#�K8��0��������k��������O"�W_}�:6���go�@��¸���\��O��ur�~"���QI'�g�?�b�����'o=����7�c|1}��{�Q��9�1�M�L3�*G6�{�G�����{�@U�)O�Q1p��5�Ϥ�[BVl��^��=z�1!;�c*!�4��D��_/�?2㪊Օ��P�#�r��F:!	�o����O�޼[��Y���_����W������M{�/h ���ﲭg帿B�ڎ1�QwЭ}��F��y�,�|��$�R��R�����G��Q���2|Rv�]��R������~�X73d]���7�nn:�l��ݒԯ&�̯e���g���t�v�0���J�ўB|l������qH}!w�6m�2#�?ni��s)��z?=盍>t:&y��Nm���z̀�ݏ/YV���V/Y5���{�}0�qeB^�[�đ��S򮫴S3<���rђ7���������5��N@H5�F�7l�q��q�+�p�3%}����c�v�@ ���8VdOu�O���U nW���Z?�btL��r����b�?������j�����_�����,<��<E�մ:�K�4l|�7��M���A�=��G���Y�L9��\b"��A4P�Ϭ�����\ї˰�,]�\̟e�MCK��3VF���p8aV�����,Q�z���߬����s
��3/��f�>8c�R���ʑ�YL�)�G���p��ުu�`�>+V�kh)[1}�[H�$Ҽ��%bc�LQ��4��i<����0�@zs?FՃ���"cΤx�K*�P�)x9$<��l�O�U���=_������Xv���O��ę5ᛎ��%4�1��mg��@�	O?��@��`]�j�n�oeڌ}�:먆W�U��c|i�b�3%{�l�)e�)dJ����Fγǜ�L9�s�Ή�e��T�)������ŭ5}�gJ92UG�T:��G���N���=��~z�
��ϩ��3d���K>����=ʞmc���VD,�Q��ǥ*)3�eh�`���\��N�yn�e��B�tֺ+W�df��`s�.��ț�mKwS�-lv���6�������ٽ��w�m�i_�OU��:<����|6iߕ�M��z��7�6e��p�o��Lwƿ���F�dO4�E��;��A����(��sӳUhC� �Ɵ��q����&���C������w���X6;�o5���A؍�n���-�?b�����+�1t��U���z�L��B�B/f��_c͞��U�F�B�F?\�N��8h���t_Ë�cw%��p8�c��ǌc��
��r��Ҧ��n�k�2T��Yv��6���2+z��D�r�욆��x��:~��p��1�m<����WWO�G����vA,�ԙZ�Ւ#�%���l	�-Ȭ�i�9])��t��X���j�L̏q�*����&���#�9y�?��w�\��//0��`���������'�����3���	�R��Cf��؇��/���S�Q$^�'r9X+�y��I�㚋fɞ4V������O�>�y!OY�w�oй������+���?�`j*��}�O[�;\fҥK׿U��?���-
�㟾[����V��߾]���kf�h<��x��%ȣG�V���=������r�?��͝�B���E��g@ix��+�� QPTZ�kŇ<���#�����9��ݻ7�?���}�yȴ���~�����V��=�S�0�ǩu�e#̆��B�솓
4�\Z0�l�yrH��y%�y�?���7L|KE��J~���5�W:������\�)�S����H���[�H8e/�TV��a* LZw�{���<}�3�N��ȝ�T�s~�Z�TG�J	�2]�[u�q��/�!���.�.���f�&Zwŗ^�i�׶�ۦ݅7˲����T�k1n��%׍	�J��/)���{���2)�ξ�G��-
�{�\i�I.>��g���1`���F���p����IѾ=cG%8���q���M�S(�f0|��5+ ?� �g��nY!�G�ԃ���̋�;�ȓ�U�&��<��8�r��N�_���Fo�ǌ�o��|@�9����+P�!�����|�z������A�����b�i�T/(���t�_�s"�=o��	�C� :�wV���.��L�� ��K���~w��ßF���_^���W������Nz8oǘ�����I
�p�U��sΜ�Q�i�ʵ�Wup�u���R��0}�%�vcrI[Ti� �hb��#�JSeLHz��\ܖ�N4�U��A�~��1A�lY�a��[�9�C�\���- �	` }π��blhCy���^���笌Ɨ�}�Q�H�E�p-���a,d2�Va���Z.*&��bGhqo]���[�'��t���f���=pɩ�c�I�j���~� ���l��3i/9>���9��_1�����'��r�=�c|��bZӷ����(�s�eOy�����-��c.R�/F@5+�Ƨl���~��a	��;=�1���M�t�3̎�q&Ʋo��Q�~�����sR�Z��BG���˪Kx�0~��P	Ё�{�ʺK���D�o���O��g�b =d�ѩ��a~��I��mVV�(ӱQ9ŉQG�牆xه7u(o�ꖀ��֝BG��
��W2JZ���p{Z&W7��;�����m���mK3�Ȁ�Jۆ|G����i�}G��n��]>C�Y'�Ϡs[�6�vgV3��7�m�7�L��~�I�nw��M��]���Qw��A�~��傆�p�I��}������?F�٧x9��_��ho�Z�����>����!�7o^��kεz���W�V�xC�e6gͲ������j_��+H� "0z��4~L@��Y�������7�/�����6?�wq�$�ӧ���X�v~�7�����X����I_�K<��U��l�A)n���#M�ˎ���<�+)����ql��[�.x��Ed��
��#�������C��֨,�*�u��qؙ3�7��o�9����=��_0��%Y�J;˲�=�.iȥ����͈�lt��˔�E�������޴Cb]�x�ю�B�<���|/T�m�������:;��Q��8�	��,����:z�x��4�0p`���G&�9�!͜�IV&�m?3i��j��[1�����>#�������?�&��#�$����iR�(SC�iO+��͆�,��L�3S��ʞ�?��[Z�#�5O2,or���}a�` (�����V�N���~�ɣ�C+��kd7�u�BM�&�.��_���D��x��#�y۳ЀN?T�a�a�|��[_=e���r��㯞�K��=
������;�D�1��ֲ�S0&��H�BK��x��'���JOI�@v��|����fߞ����߯�ӳ`I��Ӡ�۬�x�@��!���apUg,܎S�ζ�������x�����m�Jk-SB�m	n���'�Վ���_�p[��Ͳu��)�f��x�M�㮣�8���~��濂�+U�+4�1�`���4�;nB��;�٤9'���ui��-~��ou��Y�j�k��,/D�l��@z������K�f����X���3���"���F�$�_͊i�<~�$oj��xN_�j���lϡ�sx��/��������w���C�=�	������g{x��l6��gr=�]d�/fD��a���w��-E��(�]���@N�)3Y{���|����s���<�G8�Bĭ"~�H�M�ȝ[����$E�LDq�@&���
n?"A($�20����$ą7L��r���V}����_�a���0�|�����<]��맫o��;��QG�i���:������p��pD�0O�����u˓��A&r�0�X��$NeqG_I��Ё�Du�������e��^����^�x#S��+��H���/~�1��z�Y*����tg9��7*|{�a�ң�Ua�>!�*�)q4��Z�L���K�TiĘ7���!S��*(�9�h��֍�~Ux�-3��Y4T1<�K�����`ǼT��T��~��O1������O�X���M�-v�:�?d�/7��i|%�SQoƸ�h�PǸ��>/�`���j�.͘�9iA�Zajj5S��ݔ�%Jt`��Y*�A�Ȣ��
z��aV$�$����0�1R/��8���X3U%W6"O:<�M}���ᘏ�2���w���i���+������ԕ��jLn�XY-rdr�-S�i\UG���2�\�HJ�<�QG?�o�[''O�4���O�����ϸw����Z���dj�N���v���Ɯ�6�>��Z43���I�3�g'l��m��'�[X�����a�����ɯ���	���&�Lg�~����Ѿ��!l#vօ�Ԫw�M-1�HN*����M�߸�OJ<�Mn��w�A�4�|{���n�y��5�`o������Av�r}�����
���3����,���l�]bS&��U��#=`ZV�����1/�L� �yp�n�ۙ�\~���+�/��B�=C&�����]�t,�����#�x����ĭ(~����Y��91�_��	������w�O(�#����w�w��pN�/?��������yS췿y���^��#�Qu��Vw��u)Ɩ�PRxjp�Ѱ�:�5����<�1�����8t�K�K�Ɠ/�Ƀ��g����i	xff�ȶ�
d>�1V)\���%�`{zZ��̌���牮_Z8��T�~�4��ae�Jcf�7sGH�o3�6�75��I���!?|��y[Ҳ�h�]-�]�_�����G*J�:�Y
��oi4?�x��z߮���G��_2}�c�Y,��mp�ˏ�ȉ6�����GN0{�as�2�<u�#��Ve��+��q!��3].AnC;����fkk�_����4
H|��H6�S���:�㧤KuP����U�ɆKq�L�F$���7O��~��*�v4(;[�o���a�6&�cpJ�=�U��^�f���ﾣ�|�z�>5��pVH��}"S��C9�U/r�qX���:�D�)hj��.����37�\�a[Vu��?�������e�m�o�I���R�M�&���mڦ=㷿�\c|�۴6S���߸��t���&�7�M��~��s�m����ƹ�V�Ko 5ݫi�cj�I7��Ժ�&�&��2_�u����&�M�nJ� �W��MO1j��r�6	c�}���ٻ�̅�}�����@�q;�j�{�J�)�Fn�yZ���%��e�f��?n�EuIW�v��I��8�-+:�ȣ�{ -f�ػ��蒟c��U�}�Ri;&�~�g Nɓ�j�ً�������c��� �C	(rk��[�0�X���7��\��9Ap͓��,Q�1e�b� ��H�
��±V?������Rd�h3�3�]�AO��o\]}S_9�D�NT��xk�x)�?"D���PI*E�h'��䛕�c̽�΁���z�����ηi).E֖�1̷�<i��y"=�¨O�����Ͽ�������C�~�2�rG�#'*Nf�I��4����f<�i�W�PP�K$�����ҁ��c�\�Ǚo�Mg�^�Q2ط�a|y^O.4�*?���{⁥n��Рf�1�u�' *�F�Z��C�
˓Ri�h��KfGY�����D	����#��Sz�<G��;9�E���TLs+��c�g��rNE8����#����#Oa�&�b�Y��2��4�F���FI�R6&-����\&��w��I{N�<;f�'��={�^�|�S�W4 d���Q�
\#V��`���m����{��*\_f��kNqv�m	�Ғ�t��oz�'J5����Ȭ��?.KY�z���� �+R��Eh����;�v>M[*�I�dh�kWD��aa^���[g\���?E��>�U^��ȵL�ց%���Y�&_R/hw�,�<\���z��E
���Z�M�*��BE���)p��-��;�`[9�2�,��߄/Ln��p�o1�殤�g|�kƭ�==����9FFˁ~j�j���%��4�O�,����&�y۽���m�~d�������O�{���߉t`�l�$J���ޘ��T�@��^B�2�֏1��޾#����#F���c+(���8�`Y�7�{ظo��!ޱ]̱${�4����rum̀eLP�6��RO��y`�2�E��1�AU��m4]�/�p_`�j�z���זtO�������W�X��}��Oe����k�U�$�4\K��5�.~r��L8X�x�T��sMC���Y�èRkj�Y���Rj<h���uBI=PF��LX�>� �#�D�8e�ќI2xZa���W�G����������,5~�"�����"���!ӊ�b4�|��Y./��:ϣ�+��jp���P��#\�D�b�/��Z��Y���}B���0�z�[{����BYV�Sf��0ZN�3E=dVɩ�l�����,9jѐ��O��4y0���TP�L�&,�!�:_Aτ�>ň��=��c��=v�?��<���x�9bZ�����>���m�ӌ���t�Ȇ�� u���ș�҄��{�n:&DpfO!�d�����a㴡�`6>On�)��]��<��^+OG>v���'�7vt����G���	{���@֗\T�2�A����)��L��S��s]���i�џ�(?�d/����u�"PF�tQJ�v+�t�"p W~�� 5;�����u��ؕGyBm�ךj:K9��-��Kx�N����	g+��'W�3n˱�D����&����箴��JqE��O����?ߥ���Շ�z*�E���T*[�r�Q��8�(@!w�7�+m��4��$~�\���o��+N�_X4&�Hj�U����ߤg��!K��3j�ͫt�E�:/��s�WP�>Pۯ���v������f�y ��钖ˌ~���0�1Z�9��AF3�g����ݣo��/i�d u�4�Wg��C	˓UX���|��t�T��Fo\���%{],��lJ��^�Kpθ?ȏ|���I���Tngx��s�j�5(k��;b�K�T�*#+y�ڲJ�0/�{��㻳>�X�Ng�å!{έ��q�4U��qО�]flq4PE��\��X�����Fx#1x��85�QxEKK�N�B�* ~�d����~����+
D�s��a.C�c���r����H&�ۇLj=a\�goyNU��<D��#��X����]9�
~OE�x���ā������T�e��T�d��,���'ɒY��%̻��_ �rk�9@ꗶƋ��ƠƗֽ���Q7�b�ҝ�M�F�=,�}�ɭ.xū\�@ϒ(E��q-Rv�*�[丅\9�_7��R�^�;PF�z������G��+|]s@!����4�1 �߳��c:�l �r���Q=�(FN,f�8cMڧ��@��d�!�lfoe� ��',�����h�fF:�6�j������X��Y@e�%��O�~�Q::��§Lk�F�On.A���z�p���R4�G�	�^D�*,��WuDZ�3�z�7Ӽs�����a��Sy�w˶6sh<a�v�o���:n��i:���
��&ߎox�:xJ��g�S�4�W�N� L��7����o�Z`-�zg!��#Ek�4�W����Z�w�[�ft�t�l�!7��J
	q�)ma4<AiV�]#	k����'�Hq�[�R��ۯ��"��PM���C�>��7/�m߭Y�p:�>�ܣ���C�5�.0t<~(39�ul`ȉ
�霣�2� �|�R��x�l�5V�Kåt�x�8)Ғ*ᜩ�����S����@��#�}Jɘ��9����������yl��M��Ն2F��
�b�)��?�\����ffY��O}�F����c�q�9w�!���d=䭺"e�ԍq����B����
�ǀ�Y���&�%��즙.���UFO-t8F�D���_xj$[*�cl#����Ĝ�7~���Þ/z;C�Um �����f��a7�ɛ�TD)�ڵ��M��agXj�@"5U��zG�C��$���d�B.�TF�RZA��:@f(r҇��)�ٸ�m�]M��"��H�.�F�O�5$�@N	�8]rD)N�ė�{�q�>,���f���@�B� "x ��V����Ӛ�(�C��z̷5����(�Y��O�#����O'��p&Z̓�{��44�J�j$i��1�!�[(>��|��CNV\x�z��I�Pz2s�����G�A��2af��BLA0��@}�l��������_���Ȫ����>8���9b�x����S�eC�:�ȿ�z����_�}X�ζ����v����L3��ovx��\�5hlҟ�츆���ۺ�y5�-�����x���4j�]�+H7����t���D<�qWZM����o�����m(=�m�p:m5�9�u�4F�ե��u�n�U��~L����7�}�q��x���$��4,�p�Ρ��v�1q��]�l}ĵ?��(ݞK���_d��*�JP �C��X�<b:���уf����l�bV��8�Ĥ�}Ɔ�O�V����	����k�:�9S?����>�]o�;��'o�3v8C%����F\%�_Ǻ�W_m9�/����O���Ή,��-F�-Y�3Ͻbl�]U��2�|�O�����ҪP�X�h�n��V��J�^é���Qs)h~�W���Ӗ�o�S�o�ܣ�x�G�Ig����'�8V���R���!�uc_�C;��93C�D�2�A���@*�go��:nβ�`�1���A61\��<���L�g�̀��,a�@��ϗI욆�%�&��CcRc�x9ӥ���	G)~&��]ju���aqa�Ti�/țv�ˌ��{��Yt�\H�K*�_ޠ�U_9'K�<G���g�ԕ=u/:�-�g @꿩ۥÑI��>���8��VO#6j�y%-�ԭD���k�#S�72�J�h|���F}r��Ͽ~�z��*+2�!��/a�ͧB��a���_��1{�/۴����V�
��p:O3�]ɢ��&4�܆dxSw?���o-�4��hw�$;^��=�Py�qۿɯ���۸��v��eޅ3��<�p�׮�Y�]�Nk����?�'��0l	\eO��/����*���J�o�ĕ�L�n^Í6Ti|��K��T�3��������l�&Y�`/�
��"]�N��W]e�{xI�P(?��C)�{�4fz�3�S8��r�hl�Ѐ��t����3&^�~�}ǃ%�e�p�LGǌ�s�U$��a�T�3�h�6�՞7��5b�bn�'��)�Y�ꯤ<� {�Q�9`�����I?w���S�'{�9fy9 �/�7�g^E�G&%$O��(R8.8�fS:�p�p拇����烼��T�Yvd֣���*�������~�����o�@�-�Q�^�IU9#y*�昴&&β��O��|�-ѩ�v)��\��ŵC<��ذ��b&��I+�����f�|%�O� �8�zUb|0�#������*<���IQl�Q;�m��{�(K![�b�X��X�g%'C{Ս�LEP�E�*���
נ�p���?
�ؒ����T@-q�	�N@�����1]��(o�Hٔ�J�[�	p�Z��H�؄�y��-e�#�2��z�1�.#�,��ېY�G����+p�m�2&��U�K,pБ{P{Ǹ}��#���<[�'	;e��$��]6��`��B!��=sl�- �"�%�\�|Eq�a�OW���߬���忰om��߳��|{��:��[�1��m���E���ITA�#��n�W򛟰��t��7%6�8�7���Ɨ�����_ח���f\s_q���_:�F���;܀��窬�I��v�����ߕ�62�6g ꆐm���Z�C�W���L�_T>�M�/�
`���)�@�o0��t�/��l��~�\�m���-��[mn�¸�o؂���!���AƠr����m?��~��ҽ���Нx�y��?���C��|�eg��x{�����g�)y�g;wdt=�Y3�N�n*a�2�1Ҩvm��t����A���г���?bqb�����c~��}�.�BXa���S���R
nM0d�*H�E��I]��Ӂ*�8�͎�\�,�U�#�G���[���:7�;F��]C��j/l�ޗ�u����#Wʜ�*ST��k
.:
�<u	��g�+�'��?�M�6]��Kk�s��XKO8Ɨ��;c���XM��I��0�0��� ;�v#�)X�(����|�7*X�4]��Qo�2P>x.��,��aФ��ޞ�V�]����d �J�(z�������l�&��'ЊՀ2^Yn�������C�9G�+9\�U�N�FC�7\>e�,Ђ���#s�I��@H	3����<iА����9�dn�a��kaۈ�G�FX�ܺ}k�A>ƗYM��F��Ty����a+^8QS�l�'�x8o|8u�ۿ�����{:^�~�G�KC�'T����u%/x�.~�G��Xί�+߾״K/���e��toN��ӵ���k�Ǿ�Y�u��g:k�¼�t�&5?E�*n�ʹ�⧿��]����R*H��K�7ݻʵ.���Kq4A]�O+r�y	�HnM�P��Zc��ߪ��pb��W�.���M!�Z�v�隝N�+�P����"�$�5�STr�&��Ce���Kt�3�R�<���w����ܖ�>�� |��c�!��ru��F�3J������������VzUyC��7�x뒲w��ƒ�iJ����"ٳ�;d���g������4�O�{�^a����B���Z_�K�o�=g�|�
�I���S�J=�.��*�� �"����6�N����e��zB��
~�wq�T���m���=���ҩ�p�B�)���T��,��JmA�����?б�3��,N@����#>�L?{��c {X�~�2����ۀZ�g�Xм-x����f���S`�bX��=����X��W2�c��B����,zETH�S�� +( |�wW��C�����'�TX�p��ۊm��y��쬗�Ɨ�3o��(C!��B�J]�/�� �/W*Sy�C���ڿ�Ul�sw[�i�"	";^g�
_�,�2�ke�,�aV���_�Ȣ����<�����!����#qsj(+��B�N����%�z}ySF��8��p9;rf�`��S��={_�S�X����Y-�g�?���Oq�#�Ur���G��r���nA7{~s�z����V��a��2Tm^�S���s��1��v������M���m��
��y]�m2^�]���r��Ls����:Ӻ��pgZ�\��:�l��	��6Z��C�%Ө/i�����S�nݜ�p�����vB�l�m�;��;����H�._�J�%����>}�̥��#�B�i�l�S�����㍷U(�H������O�!�@E����T�9�'�����A��Xg䞲�������u����wƉ}V���� �##?G���cޖGnި�KhLx��Z�����l�rt�2+�"��Vς�ґo�2�jt�"�>��E��?�)ˠ*�+� �c9DB�]"'�5*>u�H*��U%	'�|��P��ː�J�����w��r.�h{�1iͧV=�	�Ӕ��<t���o���d0_,��ݵ�k���u*4S��v��/(x_�ͭ������Y{��#�[!�� ixE	d�Uc����Q!��E�B��t�Y@�>��RpI3(���yk��Y.���6T*���g��-���U<��-M�#-i
��4U�J*eڠa�Ium����J]�w�OM,�b��A�Dg�2��W~y�+�Ɯ�piV$K�>�AU�P���y�!k��I8т�K�:O��&b4�����#>�O\��F�'��ͮ�xSTO�������2� �
��j!
�Y�;I�/uz�a7d��S2��o���CP�o���m����3k��J���Ob�f��%nU�x������o����tQ�M	;���f���W���voC�:�]rv��g��:�u���ܙ�:��o��k۲�kL�;��@`a�7�l	�����ę��a�C��It�����m^���#���̑}�oc���!��9X�~�P�a����9��[+���)�]p�	��~8�*}d��_>x���r�/&=ee�G��	���b��JU~A�c�Hz���4`L2��r^h�1ά�(��K����|Ԙ��]v<d�1U�����[C��������iR�D  @ IDAT1j�%�/�e���5D���O��Oڊ4�o��㌭���q{�-�
����rL�+�����pm ��#_۵p���z4����}�c챘D�.X�T4�0ϰ�dɎ2:��b��>3bΎ��ռ5��%�B�T9�Qt&I�(��*L �gTT3��@�C7 �
m�&�����x�{�+ˠ^�IP��
RiCq�ͺ�/�Ũٸ����R�l!��սS��MO�BS�ʔ�j,@`��L^F�՟i�܄HNQ�Q�F��}��AC�W�1��ܕFV�F��nt"]j���������d[��Q��e��cģ�L������i������Nx�<滕��9{�r�����̻K>Z��s�7�K��g�n҅O��m���H}%r[�����ի��N����)���&9;ޤ�67�����w��rlW2s���_ͫ�,�Ͻ6�ޤk~;��6�f��\y�5����8ו��Rxǵ�6û��%\y6o���f���mmꖬ���9Y�W)@}m���'�	�.R�ikC˭*>@��V?L�A�#ު��":'zNư� ��`�eT�)�Q���u�L< �����|�O��"'�c���#�����3[Ύ�f�j���ٟ��d������=���L�h4��=�vbgpTQd��ȭ����ai���]1q�K�|��?�
Ӄ:.��D������1�ˏ�\C�ѵD�1�Kz#����4�<�mؒ�ud�b$&M�3z�(t��X�-S�Yv�������u��U�2Ts�FM$��Ơ��ʓ��c�{����3��W�����uwiL$p��>%\)Z�ΎY�%�P^����O[�/\3�Q� ]!�
R;������SL�tq#�J9Tʪ_���ZL�|Q3�T��O�%@�*��M�A)l��p�/�¼˸*Y!���F	��o�a8z\C/=f�e�1,�z�B���d;=t�0��:F2�/On��Rn�pEFX�N3�ױ�9	t?jk���6�t-���kz:o7��h�<�q����cđNͭK�d�E�H�б����ϗ���
��X�(��~g��4f>)�PY��$�r(m�^I}m`�14-��&���U�6��&�U�w	uym������x%jZ-�a�m�7�6w�&lN�<w��*iw�������ێ79^o����w��t��B)�j�?�WP��I Ɛ7������_��g��f�tP����7N��w&��+��i�Ϲ` �����K����!p�����ޤ�O4.��%��eU:�ٷ��B�K��}Y~d[���g�<i�V��E|8��
�$9�Hj�o�`�w,Ѽ�������n��4�x.�p2/�oꎕW\p��<��rM&��J����l2�z�d҈�McZ�k�+u ��x�B�k��.��p�d�a�Z�%5�#_�&D��N�{��.g��g�6\��bV*���B�|ο\:���Y%1���'�=D"4dJ����i�~t���V1���p]kƣoCM�Fb8@�a%/h��7?$p��k��E(oˍk�"f^,� �Tq.āo�ʙы�2�ruJEo`���Լ��"����7�:4(�Dξ/�!G�8��a������W��TZ���p�D��$�O:��4X���W�����.8|�#$>|��G��xNǥ!u�&>mV�3ʱ�f�"���:�g�B>�*�(	 �9��m���Ʃۿ���7��){����n�x]|����E�6iM�E�:���7iu�u�g�/�l&�?��앆��V���DfY�g�����涸m���I�ƢHc�J�4�	�	�i!&����D�NN �#��g��� ���ޚ_��������N�C�8ߣ<�T��>to��P���������lR:M�M!>h�W䓡��t�-}2�� �\����#�Dאcȹ��ՇwoW�|S�!�H���}Ȳ�����V�������+{�����g��fwO�8i�#�oD:�U�����Kȝ�5���h�8G��Qhr�c	n&WF��[4���V��;�wJ�o�w_嗳���j�PA+~Ď�7���6SD/�|V(�7��7���̹�\��r��@GELy�� �������3���a|a�G���T��?{�V��dZ7��̺ ��;�1�~�^S-k�o@y����I�$��"�e&�	��m4���2c�d���&0��ʰ�B._W���]�5V�������x�k��q�x�l,�
���G�K|B��2IE��82�U.�ֲ�k�xĄFW^>ѩk/u[���o��(ס��|����Jӕ�6O� �ҽ2�7�H	�i1�sY����6�NCꤓvdF�ڈOx�Y�<��ͰJ��čdݒ�ZWׁ]�Z��_�QSy�/�+r�w���w�����XJ3��i'(N��[�DBC�T6�6�x�i	iz���_�uS�O�x��s��_��%�]�e)]��O�Z���Q�,���:W�V��4o[܌w���XWӛ���v�z�Q�.��(�9w��Z����Յ��[��_��˒Is�rg�U����9:g�����?�nuumd��d��y��#�\��_����f���;��C�4m�������1��'W����Y�|�[6�sSBڽ��o��9ﺅ'en�>�m�e[m�O�C�'�m���a;m{���
��޹�ը��n]<�>��I�}��������y�7�"֯�K����]c,����Rv��Q`xdC��'צID�Co��6�T���$�	���d Gܵ��vˮo]�V�pP\��׋}W�;r�F� �����A~P�����iN??��+�hួ�+F��
����I��(tÃ;_��(%�#�x�m�s���2i1�ێ~?IgZ����P�����Y::�}��&���kB�A:��r�t�����bRͪ)�,OJ�唁�._-�Q�XB��Ck��7m�A1��2�)�u�RM7�.��?���$��J�AN9�Pˡ���^%�_�Q6et�B��i@�%N��X�sXo��)��,}3�4����{f�iBo���є��t�q�[��i���&L�/l�U�5X�u�\���,W�r��=�}��H���C�\s'�W�=b��ay�皰��>���e�3��W�&��1Ѵ]��\Kl+��#��l$����c���9���l�G��u�Y!�-�#	n����b�d/�,��p�"v�������%h�^~P,���Ĺ?�_���8����y��=�n'Q��s�S\�.��K�	D�ӏQ���?���Wm�mW^<i���8��睆s��+�^2���9��p)�NP[َ#i�s�<���?�����|>9t�Xy��U{���}�,�k�-A�+oi��瓧��_/�f�v>u�}� _���ۼ��l�Ok˵W2�Y(#��8�$(�{ε���ß.A��B�+q�L`A�S���.���@5��s9��̜��r8�s2��a�WR`&aÖ7p��ɴ~7�����)\�A��b�>�\�vU�Tq�'Ek\�W!��Qy�m`�Cq�F���O;�����!��N�؝��+|�e`�����*N�<�j�`�b�Ze���2��SU��yA��G���`n��K���8~ D�6�}?��p�<�H��w�X��X�N\lN1�a�#��h��S������GS�9��465��Lv��+4�J��̐��*<�=�/�"x�����}c�c���H�辛B3]�U��Q\�X�u�2c2��tH3�4|ut�ʺ�\o󳄲o�y+�R���F"��}\[7��UvN|�]��������Cx�&Ǒ�#����kt(��i\'����lm�	g�>������[.�o+ߙ~~(ˍ�7�W�w������o�Ү�E0;Kϛ��=��w)��F�F>Ǒ�No�;��:�p�T���M��;}ɿm/�m��f&��H�,+����ú�+m���ڰi+ɻ9��ӗ%b"��9�:oRb�l'��[.�L��	�U�ߎ���_��1��2��$˒��7i۽z�:Z�?3�M;:���^�m�au!D�c�ğ�@�^��V��ke�4�-йYY��!�]���<C����}��Q�'WϹl�8��ĀAo����IU/:A޲z��xWBq���L�����΄��&���12Y�.�\ք7�=o�L����	c��(�g��ͬ�G��[�"�PF�\+4�k:Z�7�x�'�$W,0M8N�y�o�CPC;��
���/���axdB��P���"�g|�S�Q�h|[q��ı��E+�'?$3K��s����워~�|u�k9Qf�ЭC���7f
=K���4$���6_����Y��#�����fɹ���v+S�$6'��c�����J�񊮕�E$Ϟ{�֓��/8��ɒ����í2�$�y�����:�zF¿&�h�T������kq��v�>��O��6\3~v�>�K�?��A~����`��U���M�\����M��e���y`�;V(��#����*������\��1����Nwڍcyq�gk�O�V����⅓ч��l��=�0��I�~�O�hOU�θ��b�eh�6r-�R��i3}���H�*cu��(Q�i��^�/�f��F,���d�8�ꔆ�2�C�(Ӗ�-B�LN�+X����ͼ��y���/�K�����$e�3�����W�}����H!��EHNC�v�M�ƃq��}�L��y�w�����Ȭ�/�C�M��J/�C��3l�dTq��)�Ц�������:�L&]B�)�;��u����S'�������J����t��Q@�4�ߵ�3,p.�(��&�<�
vJ���#�)?�i����u�"�λb�䘣��(�ؠ�B�3
Y�{�ר�s��S�����M��Ph�s�&*��GPq�tQ�CQ�%�(�b�ƀ�7��K�,��8_o�����Զ�<�/��}�e��aHo�bT�{l�O�DV��.�m\�,))�X��*��9���um!���ș�s�k1,��H�)w�.��\IG��
���8w��9���Y����N�����R���[g�ü2�0��y	���ؑ4OY�:`#{�I�d(��t&N�ù��4��/w4w�c���N������W8ʭ���.^6^����`�0�ʆ%�w��x���r�߸��uitۺ���.���an�&��ؼ\�K���W~B��4�?`/s5�p��פ���!�͏������)r'�8��uIۖ�H�p��c�
{��#�ծ��p���	�:si�,�)��^�r'��Eo����G|���i=��mI�Y��Z����m~g��✖�]k^QP,��϶��x��$��$'V�LIBg�z�ov�܆�t�i�40-l��0e.ٖ�m;�!XM�8��8)U/�l��L�6>��?i�2�~e���L���:zJ����,.����{���&YlIj��/:'��Y�]޲.	A���+�%˪����?���Zʑ�R-�a/BgkbEK��$�:�Mܰ0�����M�9����7B'���Iᗲ_'Zg��~~
)�����}(�6�DP�ebq�\W>�sΜ<�&�u�e�Dϛ8Oo�G�m��|��Mitio���0��)��l�\�<o|�X�Q��R�RTz�cu�ɹ���}ʒ<�H�	|j��.��Z�X�:7z3�����F쫏2������' �NeS�M=@O�ʯ�����Ք\ٕq�0�ǿ�AvZ#=W�a�@�m��~��D­H�9��ێ=��[��i�,?���Ç����kfB��!��9�c�Ap.��Z��_�v?�Ȳ�m8�G�WÆ9��x}�?�Vv����}�g����S�w��?o^�9�t�K?º�y���v�6�;<�J�Mw:�U�<�9�o�k^�8Or�c��4`�#�ƻy8�7?��T�����uv[�`k?s���k��l:��g ���γ�	��؋�&�Mf��]݃�/V]��+?���&�~�����7%Sߦ���݉��M�I����_���]���Q�,}�.��ŘO����R9;�E�����"J����I�l�sS&��i��a�2�M�\M�-?���N�,�J�c���'1���='�͔#[t���.�v��d��r�lܐOi�Y�h�l�4ke��������O>�sxazQ�)SW#��lr���\<a�Ld�Xz�+���jz/��0=&�X���.G��xyrc��	������F�'!H�DGq��#��ܽ.(ᝢ�x��%���}-�t]��%��jy���\�v)�x9��dVs\�\�|�w`ϕȊ�� !����4b�scٰ3_��XGl�^�?Nt��,�u�}�|��ӫV�g���4&�~(�k����	-HӤ��R|�����x��ۉ�(�c�ǹ��]4��(�8j'������u�:�DB��!��#�g�UXr�d��v����wxU�����}�?��9+�*��b��%8ALT�c95�#x�!;�>�����gS<:���f�sw�:\r�e�!m_�MU�0nʸ��}70sw]ن��e�\>����\�<?H�#6��g����ϫq;�γ��pt�SR_��ӗ3Gz�ҽl���$�	�G~��M�q��4��!S���a]7P-;X
g[w�vn��S�i�}>�����ݕ�]�ߜ�[��)���aџv��0�D4��RWF�z�(t��ȫ�uI�&у��o��<�ȄSگ�"B�ʠ��Ɲ����;����qw]�'~���mIK��̭�궖�u���fnz�o���x�kv2����]͆�8^��Ioy��cG��'��2�f.a��5:)J�p?� =�;����<��`~Ź������޵�ɔa�PD*E`��:�TF���r�����Ջ!��
~Xcx6^wCY��C�j ���̤��o-W>$��({_�S�TK�w�"�p[ `���v�)OR`��$Rs�/�w���O>
��A2�\on�i)5s�N~e\�ٌ�O	�	5���0\B�9�̙?���j�`9_�q�������:��������s�QfDl�ǣ�ѥF�Y�{�n�Ƽ�Q�k(i��f��ৱƫ�E_����+���c�x��;t����]|��W_�5�=��ؒ�J�!s�#P�e���7yjӵ'6�6O��[Y�P�R���vY��↿=�#�2_^VzI�`ܼ#T����+�{y9M`t�:���n�~�.��LB[g�׿�5����ѹ�dM�p�'{ �Y���.��s#�s*g��i��'G�v����;���Ҏq��c������M���`�-y�4��>Cq�|�8����CfT�=?��n�ɬ]��#���-N�@_��OI�V�&��g��ݣ���7>���	��S�x�v\m3��;����:=_]�v��`:%^C����/���S��[G�gv]�tc=q=��P�WdB6u��l�F���H������_���>�Z��Y�'����ԏ������H�T|I�^�Y���͡=����T��>�J�\\�s��&���	)su�4z�CbN2t[���W�#2{�"��ӑ.�J�������'?�sd
�����y��AR\�'�S|�3��ɕ�]#�ε��	�5�AФċ��?�X3����������P�u�v��}8��m�6�G L���u��}~Z��ˍ����e��o2 ��ΎW���H[�-z�b&�8�� ����^���ރ���/�%��1��͹�*�(;9�s����φ?����5#�����"=G�&��o���k}����׫4�Η�x&E�1�~�{T��2����c�ѓ�/�������Z�Paa	:�e�4�ŕsK�mhS��9�7cn����[g�@y���>�]�S�w���e^ǮӺ#C�*�i�8с\��v����c��¶�U�.���S��+Y�s�o��#��y�6YV@o�T�W�ɏ�e&�ɓ'�7�Γl9cxT���<\k$w��E���3����l�X��Ύc��yΫ�#/�m\"�ח�Vڦ�>���]�7���w���ߕ���g�]�F�;l^�,t��[�2�ԃ3(�Z�������ygS����̱�����L~4_v�a���+�pˣ�[�����2�͆� ��|�?:�c�i�
���*�.��ֽ\����B���� +�gz���"�U�ݖ��>�w�rh����Vgm�?i��n�(�8}���.98G��Ik�Ń�趲[��"���e����;����4�&^?��ɳ�<0���:�9�`���9=)��t�a*e�p�_���:a}�}&e���w�C��8G����1����;���rTx�E��Ch�0�r�܉-��f_�7��f٘'~�2ҺE(e����Xkѕ=��+M�9a�E]����}SC�4�Ix��o�@�*&���P�03�Sη���B9�h"�a+CJsɽ�S�t�D~1^)�>�4��a����Da���]��=�ԐXa_,��
&L�w�v�!]�B�+mh��D+W�T�7it9N��bϗ�|;@֞Ub3`f�|��̑�O6���<��O����q��w*W4�ʥ���ֽ��}�z�Ru�4D9аLȨ�d(�.yC����3p*G��t4�;��F�ƃ�X_����⼟��(��<�Kd}I�����!d=���!TN�u$'�P��s���Y��E��B�nG�������_��)~ݎ�y������s��>�4��q�+3'dE���2s�\�/�k�:�P�~6o[ߛ?��YIj���gq�����c8޻F�w�=^oؖȏ�����	pHذ�����<գՀHW����!}�L�5��Mf��.࡛��dG̾�?gFS~��>/�8gz}�1�[��/�{�����,Og�C��h��.܉�1���~'MO����|'�2nY���^���I�*�)�M_֥�1�u���2��˔�6ѵ��SlU���;���h���e��>�����U��~�O }�ݷ=y�<��o:U�Q���y�x���w��c5� �Њ���kQQ,<�w	ga�����6d�}��e�t\̌��-���e�r�<�dc�����!��|�2���ɞ&N��7�w��!/�F�|�%��
-7ע3C�[���t�r_��徶#v��-G�3�Œ�]�+��Y���y;ƭ�3�EK����#�w��=\S��鴾�:&1GbV�l�a�GX
�)M��"Dos��kJ$Х��h�	�� �u�?�;ﱂ`	�}>�MD~�ʑ�
~�'��q6?U[�͜�Kt>��6?5�u�*���P@6�C��9�œؤWo�o:q�q�Ӈ��|3r�|��͛�m\Өj�5�^��;V�c�=_�>�"tZIC+Pߒ/_��}��A��MÎM|o��,�u���:晊f`�2m?��e/y��5��q�����k(�l�s�Dg����!�J�D�*���NBUܪؓ.G V�fcst��'.��0������SG�~��.K�_��iogɬ
G�aT)^#I��}N���/�uv����C/�w�S^�g��|�gqG}J��a㺚�]�W�}�^��w�]�����}����1����U��x��Q�����Oթ߮�<mݰ3^��ߊ~��/R�b'tF�!0�����Y���d�7oN;}�;�������o���8g�G��N��F�s9H�-�ˉ��;��t�ctUy��
["e�Nq��#�7�f�Fߩ�i�y���ɫ;�,�zۅv6ב\�@0?m�zS�������OA哥NXy�7��m��/�DМ����z�MM���6z�e��U�X��[i����]����P~q'庝� �jJ���"D:��39J��q�
@��+糌�T��`&����3���X�`.��C��/#�\�P�j�;&=mh��o���_�5�^��u�~l�O�
IBc�Xc���ܯ�ҹ��,N �$`>����D�۹?�,�/�1��]9�z�1* 6#8��z%���&� ��X�W�	g%x��{ 'x�9�i�ྖ���^w��T���2�4��g�W:�T��������1���r��	�ǵU�k����O�����Y�������1�����Y�R�V�% ��Xq��+1ndY��_?�,Mj�|R���ދ'����S�-�ܥ����Q�:w-M�%��g�� Oc�����nj'|�?|�\�~h��.��s �1\u�����XVz�%'K��`�):��ѣ�Lmy8f�g���O㰙5���?����/���g��"�v���)������=C����KS��Ӧ��_!���@�i���v)�vqf������#͍e����:�Fe�seq��<��ę�j�k�S��Y?^�]�mf�̀n�Cǃ̊�ϊѭ��o�⟎�	�k��z���r��?��s��^����O��g�ο���9��Z��A�8�6�[���`�>���BYiO����8o�U3@�Wf��
rLt���O<�G�V�G{궚������vOG�ͻrLY�,�8�m�u�;�De�k�n
?�{��S���Ry�	WK��	�Xg͡����q¼�n����af��"[��
H����>�4�t�J�尟Hb�\��5~Rf�o8e��c(�"����R��	�o�0��ѕ��m�<WS9O�����1[��J�ī�œ<�9\e��봜�:`��-J�2t�!�H�t�7�B�X��ɹ��r>ċ0g�$�����+���q�(��A�p�ٸSld:W@͆�[z~O��m��W:e�!&В�!� ��8`f�,9��e�Wark�E9���8O3�d�+���9��4���࠳^i<4ڦ�u��7�Q���tkߨ�F�6Z���A@�{��x�l]۱���질v6�+0��o=[�2�'c�b;3xS٤�ބ�L4�B���O$��3���ލ�u\�$ ]#3�+��V��J^��(�ɑ:��Ƀ#���YlgG���v�"��I�[�dy���<	�$�}��GշG�͈�s��q�rtI{9V�����Gw�SY�ȶ���X*�{©�f���1�x�щ;����G�����u������]H6�;�n�<�nKbwDd��Yӏ@��};���W]�/N��~}�"���>ӿ}�s�ef�9o~�a>ҜWS$ݞK36]v��4x�8����l���S�����/x��5Z�w����sbq]�[����{u�-�z���K.�c٢����SF〩�S�G�*�p�l���C�r9i�.B��j�����H��u#�q���Mq�-���!����[�LT⦤z��8�LH�呈� H�"�(���vbTYf�e���9}F�8ja{9�~��Y#k�+M�2(�x!�Ŋ*T�� Sg���N � 7y�pqK#s��rU��~��T��A���T����θ��I&uvy���u؍_"��2e����x�)Q������,3тh��9��?��u#�exYd�9w����A�:��(b����f`.5[�ɻi�#���U�\e:q�6�Kc�ҿ�"��h
\��rT�|E��Wt��m�'����j�5�/��k?���~�3΍�`_U��s7O�P���U�gy}D��L#ޙ��e-�;]��J2g2�\��Og��,�H��C:����q�$��O67Ri����̃ �|����N�L�H�G�K��';?rrb*�庍z.��L�R0��%���Ύ�2������R����_|��'�Nu�:i��C��8�p�������l�o>��{���bf�����ݎ��t��������a��~Ü��������~z�w<�\��ԪC��ݪO���8�/��t�)�ѕzȱ�.�%d:���_;�50����L%�Cv�~�d����������q�?�۝�~��Sk8�c��{9������Zw��ۥhmX2W����L�^a���"�#53�ث��!�=ɤ�8�;���-�8n�,�?��<	Im�d�C��\z�U�mAS��m��0�X�7��M{g�b���f�)9�B�$:x�w�P>1'ۉ�N�
#�({QF*?h�}��]�ks�`��'�  ��1x�fd��[C.<��.͹��yL�8ǁ�a�T/$�_ډ9�B:��Ȧ���˴n��SxI��2e��m������<��&`Uj}v��̖e��p^���	}�V�i��~���=#3�ʛ[�y�G�ljV�0!�
��4v5I.{{���NE���?B�.�\��>�bp�~���ꔩ%4�8�O'�}1���n:cA28����m��}0�1̼Ӕ��4���i(v�d�|-'�3q����#�8@����{O:*T�1�O̬��!I�ȯ�⬽���}���2;�
y⚡���8���B-Ox1Z�k���Y��>��j����
��|��3�p"�����,� F��\�~yX*X�\x�IL��Fd�[g�I��jE��K<' ��"7�i8r�t�!3Ac.���!���;뜝���t��٣���!`#�����c�V�%y���ml�����6�����tl�!p-y`��9�ʹ�N?��k�A7�xwލK�w-��Dq\;�8һ���켭��S�CE���֌'G�ao���x��M��{����7閬����%[��W����M~2N6���>�b��=���?W�ym.��Kq't���}�	�W����A�wc�]Ռ��~��R���,f�,�}�'�c���?�E�e��>�M"B��k�]�y,L���𖹦vi#�=����1�� P�:��2}�8K͍����A��>p� @��(�%�����W�MJ���ƑO�>�*����+�Xe���t�J #����1�gɫ)��'��EB�O_>�Y��z@��g�#���e�ϳ����6vɎS> �+�"�ٵ_�C�����bsY]�'3;�I�I�b.��p��:wk�I��(�Q���;9g���L��
RO���ܫ��*K<+~�r;��\*������o�+��(x��q�|�А�@r����!,�N�1
!dNE�Y>�	�u�a�7�Mg�W!�3(��b�� �Ćh�)�X���i/�!<�s��g�מ�>�۴:���'�o����mt�3tt��d�Oi��:l�9OY݌As�9EFX��Z�SiG�\�vKW�:K_:��� 3p��D['��>�B���jf��ڈ��q�!���d���oǶ���Σ�S���:�;0ԥ��4��vΔZ À`kw��� �SdD���|�8�|ѥ�������¢+�r�s�S��S��u�e)��>�ْ�{O��A�3���M`qw���l��Qρ��kXU��Qb�?%��;ߎ���[�O4*���Ni W���;�����I��c�ő99�)�׽�9ظY//�5�ũ��/��(��9�kx�^-5ҝx�!1������w3`hxY�'�̐�u�Q�<<�����U����OT����ٯ�S��)�� �RR̓N����g3��ًT�bg�s6�������)N;���O����u`�	�6�I��G8K�?G��2g�C�ٶ0�mk1�8<zrSC�Yx��h��/��2j+_�?z}�:]���Wۓv�x�5`�E���z<�;���fk��hG�ąF��������y�^[?�8�کH�2����7���ak�K�\��v��+X`��gK���;�ٶ�=�/S@K㬅Hjc��i�8Pv�����Jl�ȼ��}�̃/�2G��=� 7�$	�ZM(�*&/�K\ğ��2L���T��[ل���ފ���P�㒫s,��uf]T�M;� ���+�Nw���5{�d�c�.6���k�G�k�����ZHz��t$2�F���l4be�z pu��2�dU�Ы�%Ƚ#�'��r��b$���vG�i ����ϫ��2��e����	ё޹�s*���q�T���t/;�-XlG.�"$&�l�:Ȕ��1��Cy�;�]1[��3��|�M��XC�V�Z5,]`A�wj��'�Od�tgZ����Y�i��)�9n�S7�9�횼���O��α��sGF^E �k4͔tC��Ҁ����I��c���|=|�0���|�i;�>�g�Hn�A�p/L�le���=u�l`��i��0x��S�֝3<�����C7�P=�v{ٴ�Y�} =]�3�\�����m��9�7����-GJ _N���X8�\��h��q�u��/x��3��
��?����m[Alɒ#�{a_�,��F:��+��\)�ǲ�s��ܛ������q����w�3��p�_r����_�T��mn�����8zspj�n��嶛7m��\G���тs��y���r�̒�kn;m|�u�͢��S�I+��j<	p$�ղ��w{��
?9�d ƚ���/ѝoM0�?%)t~��z�Yo���`|��j���漷��J��5��ewx�T�՝�9�)�p��9l�D���:@z�	d�W\�]y[���h��MqL>���e�Sܶs�Ŷ�͓-��F�ڙ��4�r܈cާ��7yO��4om�GG���QV�W��;��i�<��32V��!MF�<}qq73_w�|���ٚd�����w"04E9�C!�V�|荗)���k�S���$�	s=i=�R7w�'�'x�RC�g���l�6�3�c��e���8I�������5$���;^]��Gj��TұA�E�l�yp��7s�"Η���Ɩ��y]A��w��v��Q	�43ż�t�u�s����(WC�ǖ[ɿ�^��}-�e��*߷�f�xF���e�w�á<��g��A��x���x�As_�&/��[Ѕ��7I�/	g�a�a�9���Mj�E_�r�D�3�#yd�6+����sK�'�Ζ����	#8����t/]|yi<���
����4���Fq�4�,f��>�A�ݿ��<���ȷ�.�D�N�x�N��"NgM�95A�O
G�Ȱ�ﳸ���5���v�ը�4�i���z?�\��&����#��nw����AtCǖ�����p��(3��>�&���Dm�l�~KNu���~�T[��<����µM��ˋ_�����|K����O̔g���*��Q�3���J]%�����h�b�����/2�t�����_p�e4���Y+q:l��.0]h�K�i��[��q�:;�oߐ����e��܉o�ST���|���1-yE	�IJ�^ۑ�Q�������O^�R)����U���6���U]dqn��A4~j;���贅�#�,NB�5�?�l[;�D����>p���w>�SY� ����U�[��]����·�;��U�dK���$��2�����*��?�l�g<�tx�L�;��G�횝���d՝LVE-���/��دr~mO�I.��k[�L�"���i�0��A�q��F��3x����EF^7�I���������)�a��Y;��f�x����b��������*��ؼ����L����HH����g��'��E��1�P�1�vD�k�B�X�33�q��C05b�l�����|�A�\#��cFp��f�r���H�iDƉ!�n�\��3�u'N��M�Sw�%��5s��u�K9(}�XY��0L;�2Ҡ�4��K�Kw�Nا}�2m�O�����Fֈ�
��FH�m@������I?��U<����6��
DP�Bx�����������L�ͅSchK<Ǭ�xYi���,����⎼:z6�J��v�<�ݲ߲.��-}0�Y<���c��p����39�E9�k�_�s������JO>mtג_�ؒ]��H��W��O����r��1z7K�0N=��O:.z��.���������ga4�ʃ<�ų��^h_�X���+�;�4��vv�ĕ�9*|�e�6�s������#�Ϲ>�+̥��0�0�[���|��@~rV�JG�R����߾�>/!O��wa�Ӂseꀭ��7{d�����4���s��罗��n"9b�������!*�s�9��YL�]d�$��n��L�R~^�a{��U��Y�Qʕ�<��F�'L�#Ƙ#`�A�F�*v��}�I
�sVQb���gu,��䧯��x|d�L%N�C̆ ~K�=�5�����	 ����S�o�\d��|;/��ܾ*i;N  @ IDAT"�I`�gr��n�É��\�w��}�0�Ўo{;K�9��KXۯ�a N��W���<�l��(731QM:�xdϭ�U
�u�Lw��F�)�'�4����p6ř�0�r���z���b�G[ [���;@�9A���\�� �ч�fjU&��TH�/��s�R�Ǥ�F�g��ta�ܦڂ?aʘ��SDS�"d��:�'[�&x�q��Xs�:��8|�Q���s�*�h���R�v ��\p�	��|�������Ҍ@=�DGk�?���,c�D�E��Jv3F�qx�ݓ|BGc�B:�s���.O�T�7��c�����@N!N|���<�^����M�ܨߍT��*���6T�D��9������� V�}�¿X?��:b97%��!E�82���lǛӎ]~�����	�4�ޚ�O��O�4��D'(~ʋ2_��������S�!������������;~�w|y�79_JI�Op�C�#??�!��K9�>rr�6��XO'8iM��R��ѫ��kw�%/<����]NS�M�:S����#��.:�s.t>f���i۹��y��,?ŵ��S)8˟S����c�xt��l<�K~��X���ʺ�X?�v�2�~F�`����m��6��޿�)�{��?����Vӑ:fyi�ޖ}�s,NRt7�ם8]��J3}'��t��|%=yqG�w҃߉��EOR�9`�?�$�e�L|���#�f��r��d�T�;q���g�,����]y#˨���e��v��a�x�<�<��k*�&��x����^��|���{ك~��^�>kg��e�t��S1�S�3�`(x��O�3���g�r��f&2>Hց��,��q�sU��s2�r�>dlG[����>M�l��wp�v*'���𢟾�}��i/ji13`7nev���0�x�����D؛��R&��L��Kט¼�SAG0 ����s6S߿s�8�tz��̼N�/��>{܎|����9�x���Z�]8��,�N�uO�(a�;��E�*Qg& �ϠriIП�7��w�&��F��z��m�K�7�T*F�,��ݓ���鋋�2���v��~S��ռ����eX�W��7���}8�G7�F�f���1�t��)�<5�QK��'/��WE��!;O)Z���r���=���>�T�:}i���H��X�2�hh�u��9n�U��=]�4��o�Tƙ���`�cp�Zd��f3r��}^�N��:a#r�:P�� �a�b�N�x*����2Nc3v\����9L�d�b=2}���e;��7���\��I}zS؛yiH�.6`?�ӧޠoS��,IY���%ɇɗ�X�n�b8b�x��V�^\i&���~4����3�	�HG��A�cڎ�
{���B}�s�����.�.�>aF��6S?cS�=\r�k�"Y���瀙��*�D�2;|�ƻ�9:��9� �[g�����O�'�k�?��3��2���V@+�n[�U^��Y��[o��9�1�e���1�T���Nf�SO�����>�׷��m,j���ы>����'�VE%�㹨^�O[j�#���r��Y��]D2T��X03_�|�5�[�up��`c�e��o�Y�쾳����+l04���Bb��m�w�EeI5�3L��v�<�h�36�>����y�s�F�5�-Hi�k}i���䛸�K3#�6-�|���3xO��A{n�C�i��#N�8��o��������pރ��P���8��op�>M�+���4��ѿ���y(|,(��M?�0��d�ގפ?k&�
�XxT�<��o>��|�T?I��s����z�<�_�6_2�J|�2��m�����O��/��w�'#E�B��9�#)�(SD���=�`Uw�6����p�?��gU��'4b*����N_���M��T���=T0&O�r?��/ܫdU�R��L�~�Z���.�6��s��w�_��������|�o��ŋ�"��� *���&|&�mglR�/�i�@��E�����G#|7{�셲��Gǃ���=_k�Q#�!K�c���b3(Μ0�S&F��:�o�P�#�T�-����F�i���Hǡ�fê�H�C�ɡR��I��u:�i1¿}�����wOG�@�H�iD7�k,��L��!��1��V��Y�?�T�hA*+���ٿhhb oF��G�Ȣ����]��oy�='�}�#���s��멃�LX�q�!�x���m�tJ�6���?�ۻ��;��~�l��R�������6P��rAi�s�FMѯ|��'^g0MY�hي
������r9ߎ�rt��8_Ż���m��c��o����AMIic�S��!��g����'CeZ^Y�WT��K��6��	�w$��f:�^���^u~��xt�O�-�E�r� �a�ێJ���z=!��ؔ�����C���%HŇ28���p�4:������3+Em������̭v���řѲ�6��nhh��O=O�<��7e���^��-Z�x��k��Dʽ/����O�[����TԹsN�Y0����ׯ����7__<����$=�>|E��c�|�~�A�,��Ǜ�e6�F��V�0�&�2)v��Ù~̲ܴ���м��j�$��H�a�F�:Q.o=�Yތ��,�?�d���{Y����x��oE_4j�1mQ��RL��B����Vێ�����O�"�Pye��kS��8%mX��v鷂8��Y:v��e�(����0U�)�8�Ȟ��~f�o��Z�8���A�k��)����)��nmUk�����>jߗ���m�C�f��ܽ�NA�a�j_z�-�K�����=���v���.����8{6��Թ�e���`\�G'!�E�6�z;���NGoi��GH�V�`������'��ghۯ�ܙ��L+�'���U�
��Y,IakHK����I���\��OY�2ŋb�lob|��I^X����B�?�%�1 �Ǽ�4PB?g��!eo�5
f�,�հ'g2�2(Fg��a�_���vI99_�g����2$�v�L�s�� m��_,��W���F;xS��^�寔�ѽLE#�:zF1�W��K��.��H����ͣ�]&�����<�G�il�Hfj�Ȅ""*O�Ȧp��Y��U���f.�d��K�����SVN�5�?ԩ��-�O#v	~:W���O�ڭ�����1	0��X�	�� ��!�v�xu�%��5hߤ�~���F��Ӽ�����<ݻ���O�A�B�̦Y����8ʭ^%�r�&�M�z:��x���]��
��{�N�����,�wd�A�����@���χ����)B�O+�W��*�U��`��Q����5��7S����F%lk�J��L��_��]����0p�?�r�q�2%r3��;@��5���o�GgŖ���`��p��c�u��RY�И���N��'��Γj�N��F��%<�ym����=�:�k��Y��KY���T����n��J�t�Ϟ���>��櫋'�[􋖈��M�������y����m���*A�D9�.b0�ԙ~3��~)w�0�dc�WY_�NL�.�\��+>8���
�t/�$/��A��~>u7myz��5���s��d���iy�~�ѽ|�>S����p��J�8_zQ?�G>Q���hsS�\f�\?}ε�Wʡ?bϟ��J�����}�>�,�0��7��O�{1͎z�Ӛ٧�>�lR����;6������o2c:��6�Caܼ�ͧ�.�����O>��vy�!�L8�� >�gO'ɱ��w�%pD��o_�~�	���7�C��a���<ѥ��y���qN��M �������ƋG{��k*�)s��"�(�,�$=Gx�3g���D�ah��w�y��fA&8*܁c�PE��)��sY��Zzt�f\�S~3F���e�x�,%̚���ց��'v"'�b���2�c��|�,`�^��|yGG�4#?��|�S?y�K*<��4��9fϑ	�D���58׈(rz�ɇ}_�g�}��(6c���޴oie���ENl"�4�T�S��t����G���ME�>r�b��:6��.pt�,H5n����NwYvyڡF7H�C�A$_���/�@�a +�׿����AM���C�&z��ieOq��Ch�Wd4��ۥ:�붎�|�V=-��һB�vH�z�l��Dwq��� ���'e
����^�"�����t����t�?Q�!���6n���Ҿ����KG�����!%�q�����?ǎ#��3ѥ��d����y�YUѝmf�~%.B@��zW<;Ϝ�^^�Bj7_�:嘜?�h� ��X�[UT}����Hv/���r�O���"Ψ����1����-��U�q�]�#^w�Ky"����L�ʾ*ؽ������vl�|�ٯ�9^dp�](�;��lfĴ��^d�*��M�zcw!��=�d�'q��8=��-+�����\�)��֘i;jt�MN|�����G�y73y��L�꯬�hr�q��U%V���PV~i�?ͫs����ŗ��E�q����'�ҧ��<^�䄙�>���GбJD���2��>g��0��^V�>�Caw��
��&�J>�ٓ���� �X'�8���K�#/u�U�eR�|yR���G���������3���v�N�ۖ��˚�!�Wq���` ���of�;���{����W�@��Ŝ��ü>�������F��Fu��	�Lu�ي�=S�~4����T�'�a�Řb�(jw�";y���8�aR��p���tN1���8״�த�9<t`gdUK���e�sV7C)Y93��C��|�8Gn����=[q>�p��2�5�6ۛ�����a�1���>�U8IT��/3j��=wf��i�r'�=2�>5/�1o˥㸵����܈��zx6#Ff���a��.'*t8l�95�۰�F������azv��J߭�����0�#�
Z�'\��Yi���=���͸a��%u4�W:�<��A~)+���b�;���2��E�W�k&ћ�=��U:3`^G�&�t��'��k�������q�Y�U�t^l���Y=b�Fj�S����[��� �Ki#��)�������ܛ�>_��_�v�c1Gj	)٤ԣ��Ҫ�z��{�wP?[�V{GG�3p��b�W���;��!��g�%�Xڦ6�8����i1(��+:��A*��T,��A�mKx�q͏��K�d<�����̩X��'�鱬pॏl'�^�� Q�t����W;���c��LN���&��i����C{��W����Gt�-#�SgFl����_�UO/��`�:����̢{�roB��qW��.�Q�A�����������D���"(�P�;�����_ۄ�+��v�%�J�oV�\g��*@p��J]�Wn�?����O.�鷟\����8`y�(�<w���Mui<�gf�M���rı���t�}�Ed�g�l��j����0�Z���Yq�>������{�O��(:�(��տ�8_�og����w0�s
�=O{��S?����>�'�6q2>�~�V}�+C"�e�3���8O�l�nQ�B� #�*j�'�
�2F��x,Ř~��{�1ƣl&8kbS	�	nΆ+����п���QJ�`*�[���Ѐ�����<r��h4$^~��S�䍷�������n#�YBӣ�Q���K$g�j6b�xsq��	2�T'��Wh�4����a:S#�*50��i�9Op�ֻ�Z���o9P�Y�%��2�A����w��긥�ǚS�	3�|����� z��n���؇��%P��N�8��e�������8�����R�>ϋC?���:at_�G?�m��y�̢��LYɿ�6_�������K�L��t�#X����nG��I�ڔ2�~c�ǩ�����yǡ���u�Lٽe�q��-�Uf����G��˿d���[�[�w>��u�k7�ہ�C}R8|��\#��<[6��̬}W���Y
��u,0hO��	�ڑ}����K;������Nݤǆd�Ym��l����۸����]��è�Х>�����ɹmjx�֒����7�K�)��Wy�V]듑ɡ��ml�N����#@<F��+x:�p]�}�mI&�JC�&�����>V��e���n���E��}��ş��ʊ�ۃB9N:� 4����<{� �p��E�<:�+8����I�M&�q�Î�*�S�/�tq/ލYϛ7���J�8R�2�|43�]\�A�}���KL�E��n 	=��f�K]~9'
����O��	�)�6>N��+����2� ��kvW��1�q$#�L�$�~2[�n�q�s��ŗ�}t����_����&�X� �gV0��"��Wy�Bd|+�����)o�,��)��raz�$��%st���K��P,3^��n�	/t��~�(rL�����`�i{�xh�Q=|�ty_�.�3U0z� v����|������=rOZ����R��I��`,8�#��䜃�!��Uح����#�3�+�ۉO����H���( ��V#��SR�$%����(L#���s�iV����N�5����Wi�gf��L^�8�3��=�K�VR)�Õ/�m��Rډ�}��d���qh�z0�Q��!k�u�]�Ll#��xq���ց�ݡs����u�v����1
1�e֌��@W=
͌�ѻ���5���S�ޮ�63�>�N7^�L ������#/��"C�o�k���ër�D�w�Z�|p���	{�b���:|�9?ut�����V2-�W��^m^۰���]��e3�l�͒�ۙ2���p��f߰�9�8lh@*������r-/�u�+2��ڬ� sU�'9y�9��H�ԝ���4�mX����!ï��mCR�T���M���\���v�u����/�:\o�/�G[�� ��Z���۶nXj�U7K�O�>�c�?���<��Q:�s����V���WY����N�>�tٶ|�j�����-&�;6Z���-�]>�;�m�WܩlB9�'�t�-�k�L���؟u*
#ee]��丐gDg��1�)n� �Y{�'�u�{~�������
D�:`A�-���i��vE��'��Q�6zī���&?o�E�,����"�v� <�{�2����s>�0@t߲��R�7|�F�� ���s@q$-z�cǁ��w���*:ŔILh����������g���x�-���a5��Y��q�f��gg��Ͽ���������uں�����)�%{��q7N�+���!Y*Ƨ�FV�VXN����Ir���^�U�Dt�+}'٫3���8�`���'Dnҭ0X9��ǕJI}����e���Ë/ℽ2H���ؙ=}tڷylfL�S�k@����C����<
HQ
���7sߤ��j�wzh̲a��y�?��L�/�,�I�!$/��`�#�8�p��owk�p�rD%�7+��Ԡ��!�+#˕k�ҕ�W=ӎ�SEo*�j����i�(�z��ud"�"b|w��K�3��(��a�8��ˎ���z7X��>�4m4�PK|tm���Uf��m�Ӏ3Z#�����%�«|Yz</W�O�N�:Zr�����|���˔ϻ�5윯N�ǀ+?2
mNF+M���M &m`�Ľ�	���N�+��<���}�]��M9��u�Pw6â'��N�L|�O�6⥏�t�F'9����f>8�:K3)�`8��������䝇(̎=���вL�D� r��ڙr���А�/��͎h̮��G`v��a���n��G~.��"l-���P����8��2vB/�t�2�5N�Y|���%��T�e
N�;��|ʣ�E���{�:v�]Q��'i��_�z�XN:[��7�G��6����c˼��O�������KM��ՑN0� �O��fW0���������_�7/Ǻ-/��Z�1��\?�&�i�ok>I]��Y�s�U��|���\��spH�J��ϫܼ���q0��q1���~���yf��8��3����㊁}��^շtE����r�ɹ<!�x�ع�^΄�2�y���-s� !6R��&,���	RV���̆=�&�w�^��0yl�׿|y�����G3���=]�'U��c�ͦ"��#^� iC\S_V�|�O��t�)y�H?m���9\K��ڱ�P	*e�L_�[dNӮ� ;1Y���%ԗ��f�Hz��Chw�>����,>���?�1us�T9[m�$K�i�S�=��1�x0�v�DK,�MQ��9W��)7SL�\�	L�	�ŏ�\Yvpj0-vA�ntH�=�I��w:b�
����Pܹ���q(A|�P�Q@�tDȹ����A^��G~{��3%�aO61&�%%Ξ�Y�َ��ˍiԽ��g�jd^5�
g�J~�w:���I�#<w��x�%���rڔQ�.M�Bw<�h:��/B��ӏ�d�V��a�IP6��_G���&�,��`�*��Q�%k�aVp:��Xy� ��
�Q��N�_�'[��T<'��MnN9`O����S��3T��z�N��>�G��32f+�>��LmgIC�-x��I"�U|{�v�J���w#��{�4�˹���e���#�Ǒ�<E�*�ǩ��8���Y��]iW�[�Vf�?J�*����:���j�1~_�pE�Z�v�`:K]���~�����]��a�@�Ouغ��>�:_���a]u3q��p�Վ:�{{�6"���.������|�m�9�v�ey��gt=��|�T|ͼ~�pUN��}}��\��>��	x��ٵo��5��m*��ex�L2��{��=^����x�S|�'�=e��y��t��)�>��`&}��n�j�*���Wq���]P������g��T��=�Wʤm6��<��M�궽JO�Ϟ%�r3���{�%�Sw��]���_i]���rnf�Ѹ9�ໍ*󕧲��I���sF1-_��T߭}k�M�t�3~f�U�%NU^$�e���_���>����䡿Ŀ�}�QM�f�tB%���%%�W��t�lZ�:+���3z�L�I�P�g���;�gsx���mj}
�1�ȓS�ʥ?�?�4�����{�J�6k��So��HFJ�хv��f�<�~�߄���x�F�����1�TP�J*8D�3u�b 9��u�@<Y�b��H`p�9V}��!c��uނ�:[�q c��1`B@�A
`h��k_��)��Pz��]��
s�6h�����ip�0g��8P�Hz4ϙ�F�M��ڐ�)7�Cw���|Y��x�����=��x*�0oŏ�
���'��蟆V�ˉ
m�V��l��!�q��%�e|1��I>�>��"�)p�!���q�n�qߘ`*����s��̍w�(<�8 �3�
��ˌ;�_ȑk~�Ce�7��������i��?Ө������<+����/��F���	t���Ȅ��,r�Fe�=��?�hf9ʩ{:l3�ˉb�#_�2��|ٰ�����#߮/���(�#y/l�.� �@��w��Jo\����,�rӛ�^韧�C�ü��cw*DF���D����t&�:���#�}}Νv%���nYt]�FV��U�:�Z�&G3�_}�u��70m�z��}�O}����t�o��zi+l[0�q7�%�t��}t�}6@v�?m��ֹ?����5��ffI��5p�����8z��3�`�ߴ��;.�Xf����ĩ�w���s�e��~����b���cu7��2rT��]�:t���!�(��2�ǯ/���w�He@�&�C���I����A�2��z�����y�~��>����\mJ��O>�4�샋�?���Qwo�m���߾�.:��(�>��̓��si ��E{�_�9\N�w������4�>�-n�8!I��y��B�\��%!��7b��t����K�<řٮ�����*/��s{#�E��у����_^��?',O��-o_��a�'�1O��A�ض��3c?߷��$F�jR:�^�s(ƴI�˃�q~�>��y9�����s�V[�(M��S5��~��2y)��ڼ����V.�A坾��ޢ��yf4��׊DH������|FΌ��kNA��}F�N�{��z���7���#�P�lu�5�2�2D�4�s�r%�5G8a���<��b�I|`�Qz�YAT� bX��T-������2��'5>����<uQ�!����	a�a!t���f�kʖ_��;�Oy��(�{�8_�u�Z��á��b��ũ�d�dۆ7��Y�q�x�k�2�{�t���[Y�|[�G�Y�,	ϼo�p�.��v�ng�{�1�%�N��O�hu���\e�}[Ꜫ�J1��2|F]�H~��>a���g�^�a[��`�:�ɧ�hٝ�"M�ɳ�r7<]���n��,-*�\�@�v��,ܟ7��`:%O�h0Tt�r����y3`f���lҥ7��T�
;{Cj/��N���ԑ�f�إrK��e���˟���u���t�̒�t�����Q�4;�uP<)@�6Tk�S�������{��9�׻:�����S�l}^ͳ�8��m��N�0����dO^X3'��W����ƠI��0x�X}���,Iϒ2=Z[a/�o�h�Ƕ�P��X�yaV&4;�;�����j��9`x`Wcm��t��a��4�z���:�_<`�h�k�`�����~.|#��K�s��闆e�+��o���8`�iHE�٢+����;"ʹ�n��M��q�;'���J�ڞ��|���Rg�fC�ۗ�p�#��q>ݓ6�r�e�:�)'���,y~�͓�ϴ�}�~����:8�F�엺[�!� !��+G�[�>'~���)�r�Qp�@>*פ�m
�b����y��ճ�yp�����S^O�(�M��x���+�b�^=�V����*3_ڧg��L.��|�� ��TN����*v����'gv��r˝���^��)h�ͤ�������9�c���5C6���N~�7�{�Q;��s3w?{v3��G{V���\gdn�e��GG?����O?�,k��\�K%5��;s�܋�`�����[�JHZ��᪊R�d ���n���4���@�Q��L8�z�Y:�g��y��&|ީ7�Z^��a�NO<BCd*!��$M���*����,j��$���%U���ix������Ѓ�e
/��V�+�0��s0��oGh;_��`)��lc��+�;Y*���u ��2��̉�+��I��,���h���7�fd�}b�g�`i���#�n�n|�<��4�-�	�5f<e�@��Ca���T��dx�b��Î>VE�꡴Л~|��}ya��&no�\�N�y��M�-{q���?�3#a/:οq����L[�}�4O����:���|��l�9���t��� ��U����������K_��aqt��'��/N�Q��f��$i:j������Bl�j8��jگvE�t%��~/�K+����CN3Y��42�P�8u�Y=�ky�Jq�9�����0O♅q���Mޱ���Y������i�8{�r��N2n	�&]��'��r �ֶ)xw�k��N��rs�u�X� ����Ŷ҈���'�W��ˊ6$�.:ʓ��M���Z�"�v�h��ul�|x���a�f0��D>���rJ�;	���	�xn�g�&=�Ef|�}�i2��K=����t���B�b �M��<��сu����{ʥ��,Lp�|-c���B]j+���/]��-CK���#�rŜ#�ȳ3W3��}��Ye� �A�i�?�{�O_�6ˏ��|�ͳ�?�`�5������뮺��>�Y�=M��ׯ�D}�q��݋O2K�]�p���P�ք#g۩��9�O��0g�����s�[��L͵���z��{	iR��?���T���$��9X����I�Y���u;���7������r�q$3�_�-��򷿫�z?�#��0����M�Wq\�v�����k֬�֯3��t�<�r�@yU�岀����j\9s���W�;�ǀ�E�݄��mg��Fy���B������ۍ�*<!Oc�-�p���=���^��I7{��=)�l*_�'�2�T�_�Q�U�U�d�#Q�L9��w����Y�t|�1�tuJ�M���	���Nˎ���`cْ�u����:Q)E����2�-G]i\�7�{i:B���!K�:E�Yy�24g�E^(�ı�m�`2���L*����FR#�|�6���q�W;Uz�4]��C�E�q�2P�2�|s:��w㎻��!�����0:`�M�)}|���d�o���܏�7�t�:�N�/�UZG6�8��峜e���M� �[�=	�t�6qGG��hΗ�IGMh�t��B�}�Jw,k�6��Վ;����{�{��wY�Ws��O�W�p��i��]��'v�����9�W3VVt����A�K�
�a�=�S�l��A�܎�z�An� ���t7�\m�^��מ�A�o�yL[�c�_�拋�>��MbS��\��.����҆�n�q%.�^���C:9��Y=?�>6��vɣ����{�0|�^��Y�һ}��_F����g��� ֕�Ի:�-Ɣ�D��
�G�|���䎃aiў)v`���{L&��!�R��'9
��
O��.����u��R��o��搻�p�t?g�O�h��gI��-[�>�V��M�p�Kv��G��R���J�7ݿ���fo���sL_�m6̧o>��sNp���lU�苲�^���dk��<9��@�4�_�&�铼Fǫt���>P�h}��H>X?�� @�r����L�}@� ���0�
>�|չJ������ڜm�4�	/h�UD?���?���+��}`_�N��=����4ϳ���EF�q�ǽ��ӭJ�2��X;∑��*��:Z���wt�|*;�0���Mc�ͷ�z����C�{?4P�f�`����Sa��NP��'��hp����:�g�D�f*	�:f��̎�E˗��?�j��/�ٞ_<]���xEv�{�3ViT;���Tz����g*eN'9F3�՘ݪ����a��	�:|�3ˎ���5�/"_�m���[��y9l��:_1��K�1^#k��g��M�O0Z����^r7�/^<��I�<��n��sݸ�I�9�� ���$㉯�^_�dQ��ϭ�_7D�+�э<�i�lc�2�y��bw��@M#�F�������){ʟ�:b3R-���80:c�ᠹ���M�4���������Q�#�.t��-��1'��8`���i������?��b?/��K�.����ӏч|�lI�2t���m����h���<�м���\;ǻ�G���a
h�*��_c���:���`OL��)��gK���m����Ճ�'H�Yv�=~k�LGpH3�����g���l�)�U�9����ko��g3���l\���XBx�.g8����!\�tw���Cn(�{�����Wآ#un�)K~�A��jñr���9���/u;m����˽�Lf��ª��_���ʝ�θ��8�`��@�n9�y���^!��ʋ�e�.�m��
2{n��^ۻq�����2�F#���<)�0�s���;1�s��]$$'K�D��`����&I8����H��u
f���+��۷�|}v��o>�3�>�Y�-��Q7�d�)��Ϩ\�׫#^��f�,���v;�q��_f[�Gu^���_�f��;2!�i�"��a>d�4'���<Ӧ>�O�Y��5��M+X�hh;M �BŖ��Ix�k~��Υm�Yq��x�en���aZ��q;�9\����yAv���7}�����_�.����w��M�>t;Sj���)��=� �rL�8F���Q��J�:�tNJ��ˍ�$3Y��iu�s�����z���:j�Co6:� f�f��qL&S���W�9>y��,EYF���Aa$�goxO���R�����H6�D�>3��#�#�0�����t3/������,]�K�q�Ҙ���iЃW���S�FOf��H��d��:{1@��}$Ň)y_�3k�G�sO�!Y~m���˦��ԍ�1p����;��C��=j/` �Ù1����L�o��O�iW.��1�D:�tB:r؁\v �_8�+��-a��a“��'\��]I�Cp�˶���v�v�V���L���.���e��������5Ӯry��}��$9�����%kkdƍ,g��	 ��[��g��)�9]�i�u��h��W�]����y���ZD�Q�q���,k����Y��+�2�f�M^g���ی� �s;���A^H>�͏Sď�8�=^q������#";Ӎ�M���#��<���ʋ'#a�~?��{ΰ��>~�vrC��ě��	.'��}0Ȃ̻WUʀ�}�)#eF7�c-��\�ɳu�B�v|7���
i�����Ik��_�5ó� �c���+~�O��T�?5e�%�x�%���G�v ���~����Ƀ��O��L�>���9e��W
|/�
˹=@�ѱ��3�a����1����7^�K&�S]���
/��{{%�h��9f;u�S��N�����S%l7�З� ni�׹(	(��|pȁ{������ذ<���Y���)���R=�%����bc
fKX�:<x����|��nɑN1��B9�C�e;ۍ��Yi�3Gڏ~-9����q;633����ɞݮ_�<H�o~�NT�����Ŕ�7-�vsF��le�+;*�g	.�����\fu>E��D����|����!�����1�8"�j9
S��N�k/��uG�ą�>�)S%J*�z͐<�w������md��Ouq�I�!u�+ |���26F��W{�I��z�X�g���vㄨ���2r<�EҰnG�� ���Wa�1��=�hOr�5��������Hr((�uU`�I�/��Y�w�F�i�F��|�Nl�8m���L��i�A�頽mQ���(�L;��5ó�=GѦ��Y���Gܔ����wq 8_�jh ciN�1���,0%����󀑼�S<g�N�#;��C����QO^ף*�����)�G]l��Bm�'�dFp4�#���'���1�#�iK��z��ڞ<ms�,��	��$K#�<>����1[�O�8�=�_x�3|�n#$0p6m�����^��p�@u��=���%;C�+�@˦	>`���C��:���ԭ���_�`0��[2�����[�fژ��E�+���z��Z,�f�(r�S�d���޽쐾��F�7��>��r��뽽��qO�Ŀik�W��8�\`�g���Ln�8q,5��
1��*ӄ��yy�{��@{UZRZ�؍=<�џ�=7�_�.B�a�9��u�lol5�z1�k���(�����Jo?T�\�d�Bρ� �{������3��M閈�������3���� ���}QN��'�0�q�%�q��;P��'�܇�R�ރ�r�G�2/O��,հ�W����}��>g�톿J�����׼�����/��R'{�S���+Ӫ�^σ¥Y��y����ϩ�D��J'���g�~��V��U�q�.yIq����#,_���y+�3���.ʾ�eVA��m��V�����\�{�E��^�q�+��s�2A���~$=�)ծ�\F����vF8t�UD��-���0;`Ѽ�g{�:y���� 
���9�Ð�&�2��VP'�Mj�;gĐ��;���m0^ˆ�6��gy?�x�"�0:���9��&������8
�I%�h�>e',��m>����>�L�П����/��DÙQ$����yjZS�i�uvR�F6#�\OȻs�G�tx5��3�>Dt�W�3��C�iG| ��i~:���h�7�%��O���E��p��:u]�z�޷�8|q��:3����~�7��4��x o�ϐt���	��)���W��[ж+�u�0��`X�|b;��n��ե��;���H?�O��3.fh�1�Ei�
�t��F+.���r�#�dCGA}m��5#�����3�\u��$�T�㌠X|/ߦ�턎�ǂ�is���z�����z�t}�<����r������C��~�9�'l�����:ӆ39��Ȃe툇Kx/�0e  @ IDAT*�[�� �@�w�s�)G�3fa�z���/�{ε�G#h�Vց�Wv(I>������,w�c�'��(L�w8Û�;��U]��%��чh�*��uaĠ�Y�[(h�]��>��0�̚%N����|Y\�?1P����f�!O����elp��=ߒ���;V�k��O�v^d�l�#���ŉ��((�X��C�Y ��WH;�w���zW���\
�S8�:��"��FO��p�D'.������EU��M��1es����&L����һ��mM��t�Ύ�e
k�"e��ND��:W�����l��������N��?��
918�x?|�7S�q�o��F�q��ć���L}r����X��2ypԁų�G�Q�ɳ2�K\����^&Gq��7/����S��r� QO�Uɀ䤘/MB�dI�.ӎO2��u֢�r�B�̇*G�=#_Y|7�AFe��پ?%��<��h,���������?��!�-	ˣQ^�m��>�{�(E&�ѧ�ԭ�i���K�o��N��`C��յ�k�)�־k��4e�`cl5�>�v:|�d��2���!k<�;�*On1�]/��5Ζu[����Yh|�7��=����8)� __
0ږ:���������7Ů}��rOn}z�{h��,8z$߆�tk�Ǚڡ��ݓ�i�"��O�/�OPq�9�q*7����0����G]��9~�|��?Ǵ�ܫ
�u��!�O�{��=3�i�n�`
����J�Xy�M0�f�dk;�菩�FG�9D������ږ_�cj�������Jt~�-ݵ���ܮ�y_����7ҏ8���#��q�;v�}��|;����]��;��{:�q�[�$'i���<��,��o*�意�}�h��S�:ɍ#ű2R������ȥ4�/�l�[��c*���Hv;�CÙ��w8� �
�_�'^��[�]Z���/s�p ����um������~�1}H�Ŵ���5����z�W<�:��J��N.davᮭ�[�#�C&F$�z�&E�����T��#xo�N��E�i���O�׉M���8#3�`���Fdf���HN�	k��z�\?[��K����٥7�=��)��^q"�Ӕ��)&�0{���!��rl����z�@b��ᡟ�т��pM;^z{�.�+۲d�:_F��-��{�]m�W���K<ϣwIS�)���^^��#�/>ϺK/�\�i{��7�2�&���U�(�9{q/-�������w�ۑ��H��h��ʐ��u�َ7M�v��y(kJ�١� {�2��[j���{�a����������^J5�֌8�8������Н��G����(��)��1pQ�0C��F�_ޅg>�b4&oZ����'�Ԗ�A��������0*�F@�mI|*�R����D�E�s��m�y��h��5҅�il�������t��cu�i�{��Њ7��n+�����͝x�5�y1�6',0x�`s0��G�/�X/Η�����)S���s�𑣠>���u��}�
��?�C�FGT~:u+�S�	
F��*�b�� a�O:�x�$�ˁWgW��:0ZX�v��1�9ׅ/��yε��wR˟�+N�4�³�m'm�!g��{|g荂p�t������.���x�LS$��-��\yFP��|�����(���i:�Pz\.�7���&iKnh��M���}~U�cھް�y��N��ϯ�{��p�q7�7���x�Xp��|�:�An��y�
<��)�'3��(�;�k�����q��*C������;���k�6xG���o��(���7�v��'͸~ڞ���'I��Fw�oXIl�3���{��5Ӧ�up2���qb6��N���(�C��%j�o����:`�������\�<{��L���d��~�k�����9�"s�Xץ>1����e�´V�����v�K=��)��g<Alr��Y��X�q��We|�,˫@���܇�\���~{�`��ѝ�\8U6�q�L���87�q�ne2��;Փ�	ۘ��r��HjZ19���C�W9<�l����~�Ӂ%�C>C�^�_�܉=�cưs�~�oB6q�ȿ<:�uuM�GGN���S7��2O��3쳨0�*R�Hrm�Χ:���qΫ�jg��
�P^5�J@�߀��{/�4��N7Ơ��|���
ܪ�pT8Gи0�Y1
g�k�V���>��X�1Ĕc�ꌸPs�:*���)^��O�^h�F��wV;�i�F|(�~�p?�����u�}�n�f�(��r��2��E���a4\�S�〙wƘn�g훼E�\#aDȨ:�tuc�l-bt���bx�ѡ>oH*7_H��?��r0w���?��P/�Wx���yrI��{v��+u2�F�f �(�-L.N��gČ����h?���搸3��3�A`w@�<9�]ñdq�w0Qn�x�+����34�|��^+�z)��x!n�w_��aǸ+��6�x~A=p�� �.��CǮg�٦c�*�ny�?��z�F�����+������sԏ��g�=���:7M��Z1εP~x!ω�I�z�x�={�6�=g��@����y�=kmp�婭�,i;AWǰ��(���6ޮ7�M�οӑ�䖕�6t�.�c��8*^���H�wRF��� ¥�%���<��!&m��8v6��S�ScE1rbS��vK����y�:X���d��F}�����Ǆ�%Ǜ�਋��a�o��p�������x��sf��/m��yIn�˼��p>ɡ���/r����#��� ����S��K��X���9��������P^�x�YF�7�t�)=�[Y[�<��p�|��XC�v����������|����d-쯞f�w�F>�Y��{�5�Q|�=b�}VkK�Q�t�w���-{Zr��}��s�T��m������	�M�1��te�>Fw|��]�_f��
�;Z�'�
��B���it$FD��^<�{�-��Z�x���,�
�#�|Stӛ��<�.8��퍐-NJ
�P ���>��s�]��(�$g`�,R6��@u,�m`ΎbU��zƀs��[��؞:M=�F���(Tg��N�_eb@l�0#_Q���<]��QBOG�q�`�/�iǎ��N��SL���f0O1�(��(Ɔ�\?���g7��O�ث�?4ލ�D���I�p�x`tk�F/9��$yr(�;�q��5W��h��O܏'=\����ɜq�{�IK�͠D�x�G~�)#�)=͏4�1�	}�
okTS�<��|d�G�+e�Y>�xH>:O�tK<^��Ȭ�� �W;ȣN�my4��?9�D�x=mHҎ��CsO�����v�ew�/�����:o\���ew��+���w9�tCa��@v�>k�s2�I[�u�su������溒��E�����t��94�s�%a��!Ѯ��G|���o����zk��ɻÑG;n�[Ϫo����	�jltzwhl�:�Ռ�ϴ�$#�<�K_ /��������W�4��;��!���ș4��VT6-5NG�e��{�sۨ~��2 8S��S�9��J���O��!p]d�r��5�on
̳nB*Jz3��B��]y��lp:�"]\�Y2��8$ax�����K�'���%��pqh:��5UF��4�����������G��������
o���1��7_f����뷂Gڂ�m�@G$�v�T�D[�e�#Ӓ^��b|2
�2�L�t�7�w�\��cv��f�ݸ���6W��GEMI���,89'�C?�-�)"����U)��w��&� ���eq�!�"�(���b�y�nϧ!��E��S��r�v�V��=�&p3ϨR�!/ǘ"�w����:���<]t��mR��֨)C��/��X#<�)k���2y%���煌|Y��9�W����o��Z��9�v��9��k�R.�e��1����>[M�Cq|#��'����{A����ٻ�Ww<��B�)w���{���x��m�8kஞ~=y�3����B�pz`�����ROC�PvB�>B�\�;߷Fc��Pm���St"%����7����5���Ϩ���r�͔UG��7��Κ�z��O��$�4����i[0q܊,��b���栁Wg>�&�����Ai�
�lG>C�'��x�[�4�~��w��u�h��(��8���YǾ�~֡��+����LB���Z�ҩ
�⚎��u��L}�]����
q �9 (�
ꀓ��#�h��8Ϛf����!NBGs���]Z�sή�n']9�o�.�Y���5��mz��k�	^,�M�|�~R4� un��ނ��]o���S^�O�ܼ~���fT���Yô��Yե�^�N&�aJ��KB?�/�1��kKsƧ�����X�o9��TY���y����쏵e��H������E���*��H[�>����o�:e\���G�NY�،�lGݾz��fXS��]f�'+�٪���w3`]�α�Y��Q%��?08��=���ڞ�<~�͔3Rj���H�>�y�M������Ŵˎԍ_bz4�>�4В��>��>�u��A>�v��f�>K\��|�/��Y@�UW3���[���	1�3�gX���v�ٰ*�"ú��k������m�IΔ�q�?�����7���`��s�������W�z5u1E�+�K�8d���12C'0�NnGc0��4#�젷�^Q��;��r�5_��C��xS����`��	c4Jޑ�������X2�pG��`�PS�����5j�9��R֔���.�W_��:|��gH=J�����¡�5w���gX��j� �;���(�N�����Ȅx�8�T^������[��H�ҍ���|
I듬����8Ɨ\�����Cu�۱[^����t1��i�{A+'�������쮳4����ˆɟv26^�`Wr��q��q ʋ ���-�����?;���=�Q��>��x���y*��n����fǃ{���s�cG�4�=�Ӛ�|��������'uj/vD����	�uH���i����#�xe�ץ ����7Kow����CI�:��ϴ��+���'�=�5�F���J,�ǌ�"?����Z�m5w��;��!�.�^����6��Ɇ�utrIm�(Ԗ����4b�w�4�S�sr�7��5�RǞ<m4p�?G�So���Oe��`Ft9Ȓ�6�i{^��4��82�]kQ�V19��j�'��͹�!�	�v*��}=�A�����l���t�َft���/��Sq�N�^tY��
�O(��틜Uь~N�W�8�%���^��>N_�$r�kX
�vU�E���:�u��~;�C������DV���SQ��r>��w|�Q�X8��8:���惣Ϟb��A��c����U����x�Z����#BC C�l�7�|��I>C�P L`(�W}M��3bƛ���ə҈t�9��E(��eTz�=
�3h$5�=SZ���~�Ӕ����h\���#e6��"sh8A�c�<�<)�I�p{򝶋P��]8q�|F���v����C��s�4F�Ǭm�3a���,�ψٳ,�����H!ǡ�5>pCK��yk���=�t^͞��!x�X�<��'�.:?駰��ܚ~'��h�;���٤��X\4���7p�嫯|��~kx�w9.t�0Z��G�|ByY�/Jy�8`���#��@�1���h��S��ĽC�W�fgr����Fit:W��%k���@+���Nu���ӎ�yn����?7�z�9^o�G�]�1��_�i6(F�#��,�3��ʒ/�h#���J��&$e�D0�����櫼�`_�S�7���A�B��*/}e8��H��1vT�=�n���p��:y�C���-���G�)x�OYO��ݑ¿��U�O��v���U��&c�!��Z�t�n�����+�$��[ƒ�J1��(4��t���ct!�|`��é��s����G~������IHOٗ�Ъ�jCg�)݀~4wK%1k@^�5,����7��M�"�3�`m��>���G�RRW׊�.O�L����ؚw�ogW��tN����A�G͸�&�>�f=����a�ӸԼ�9η�
z{J7jS��غw��Һ�_}NMT�n^�o'�]�Kj���:P�C$�slV���0q�����c^�hf���8S��Me�D'��*l�7���k\��J���5�����k��=�A��4�3��S؂�4�~[-s@���@�9O,V��v
2'|�ä����،<;mi
���$�4��|=`>/4�x-��zE�btխ�.����֬���|lHg�pOY:�����Q�9�#���(��uڂ��Q+L:�i�I�|-oe:�?9����9/��֍��� �+_�FQ9_�?���7eu0��}>ƕ��s#C��Yy���8�=��%>e��n�;�c��S�1��wdQG1|�V��rq�#�I��a�\���1�ҳv��{�t�h᪫��<~��ޝ��O.�K?�+���_u^��TǈW\o<v]�w�Ӏ)ltOh���OؼضCq������*��'m�4�7���7;�~m٧���l�:�zI�,�ulR=�0���!bu�dJ�[tB>8?xx����m�2�*��B���cт����Z���?z�ȟ��';��nx��>���O<���'���t��\N��)|����8<�G��w�-^�0~W�O����:p9��6�X��Oۜ�{y[�A�/�@���/,�8a��-�ɕ��>�?=�~4AvH��
����Z<�S��������q��@y5������=~�/ �P�GmJ���Cg�Q �>�S��|�{~7��Kr������2�K~|�S��ח_��7�ɒG��G9_m���	�y�N~�\�;�#���,j;���?��X���|��o=EA�7��9�p��N�!��O�܏z��Y� �*��ޯ�M�,;}��MAJbZ�15��]�ȸr��)x�ΏFt���0mI>G��V��aל�`�'9Bk%��޶a���>5���O���ȗ�y��W��͏w}Z�������Q쎔�i����~w7��B>�dq*S	�3��h�5f6�����^�=z���4���D\<���_��7G�!�rZ�wmR��7e&೎��R�5�?۸k<�Dh��)YA�۸t�zU��59����ۣ��h٩^�	7��}��e_��T�;�w���<OҌ���)�^��U^��y���H�}�c�7^��_��<���Z���A:j�
��y  }��y9�����t3��;����Nۑ��C�Q�)��-���G���Yr?�!X���{gC竂�:�} 	?��q/�Vp�`���l�C�M�ɔ̻��TC.�z������ U�g�2�ӟt�EQ'ǩ�E���۽��<�ҵ�A�>���K�NC�(�-I;L�)�t��wM����u-��IO,����H�ж�t�!��i��j��?!$��W3�<�$���uq)��sm�D�������ef?#��+򕘌�$}` �O~|�)A[�p;�w��F�Ka���ns��xsZW+��o?x�oKf�(osߗ��/�)������09=���r;z��nx8�|nZ�w��P�k�S���'!f�6B�K7�N5�D-� �Y�����=���9��Bc�L:�r۫S�.]����ԝ$M� �	�).ْ)o�8�?ⵗ�2���r��i��>u)q�o�n�n���!�8!?ُ��,��S�ĆS	��/��T�$xi �j��|�i:%��(���&lU2�+��:U�v�IZ;b�0��:�36����"��Ι��Ԩ�W/��#!Z~bV���&n8�Wc��'�P�{e�1��m(�q�;��@�<J"�Z����T�F��2��m���MCe�9�,;嘧_g�*[6u��e���BϞrMc�Y}�'12�bX�li����R��7�Т��к=ρ�3wW�������)b�����u�~J@���4� 4���[��t+c{?0��X)��D5���$�"�@�� m�[k�A�(|�c��ҋLn\���ŵ��|��}L�ѣ�Ѝ�C�lp��)���������KHj�;��x��N��S��c�y_>2H�qǼ;�xV�[y���k< ?\�r�U�!k/w�7��oX=/zY��|����`�Aw8^x��bTkF6��C���%��L�$r452O�ڍ���4�QHf�<�i�Ns�YӍ��@�ΰs�W�.��#`�>�Q[?��u$�Q�8i:Wu�����--�<6���v
:�@������OiɅ3�'(��ė�i�{�8y�z�|�ܤ�ױ�ޒ3[�\��Q�nօq��X���3�:��t�isj�e��Ls�{��>f�o�	��,ݡ��M��:{��\��,+�3����� ?��ٺu�*��];���Y�d���T!Wm{��s���O?E.��C�-�B�����u�l.'Ӫ���_�}@gh�ӏ;ߜ��58,�eA��Q*�	�a���Q(Z�6O�����8u��pgd�@&ԥ
���J���s�9q���i ��(���ĳt�_��_e��|r�;��  ��2R(��|~&��;�sķ��g�^R,���3cQU��� �h)?�JF�V5���m�	��QS�.�Nk�6R���Vu�\�h�f�c�l�i]G��>�b8m��E���o����׉2��!Vʵ;
�a�]ǯ� �:��!���@R�Q:so;Z;&��H�1$v��"��3
�1"�K��?�q�L�u�M��eߑ�����T\Z��y��mF�v����pxS�Nb�۟*"x��\,����W��Ό���2E�{�����܍����S32���Om	�X�g{�_�h�������߆��#�|�ie�==����֛��F6��7TW�ꇋ�qsV��F<�VF�����k<��>:�]�yO��O�ٴ�,������㦭��/�y��u�x�#�q��l���g�(__�Ƀ���a�&���c���SQWyi�}��j]��ퟌm�褏l�;ps���gu�4������}��e鍺��6H�`�W�>�|�2�Xp�O��I�|��N�����%�~& �9�v���w�L��uYH�D<6����>ɗ%��sC���'��A5{\���c-�Q��%^X��%�������$���3<���sk<�������\���C�|ʷo;]�K�=�D�}�*�1��E��V��P��E�J&]�S��,�Ğ��Y��H�)_ +�$o|�������ک�pa SY����m������qVϘ�
�It8��Y��4���<@N�&C���;�^��r�O��m�u&O_��?�s�x����ޑG@����+H]�W\�!�Ð�@�'}��f%����ӻƝ���������]u���;z�:�S6w����He�ȵ|M��S�Ry�K%��C�ܹ�i�M.P���)��J��]k,A�@R��Q��-���Mu�88:��������R�VʈםL9�<�7��8O����y!�J8�Q~��ӝ1��<���A�ӗz}�k,#'׃Y����E��~J�C�&��!.�����*�|.����3^��#�=��Ӕ�����:�J��N�$��Ƒ��N���{_H@~��8��z뭷�XO����0M!�Gg	�Q�����qz�V��8_�:pt���,8�H�����{�A|ׁ��W:ONB(oY�
[�K#�,�����G��(��M�u��˽C��>q�c�%���\���Q~��5���g��1톣�:w��T`�V.qm���硦Ve�c���ۗ_~��/)�)D�!Agч��U�U��.]QW��\�C<�����$*�t�c��^e�){ݑ/.<�=�8�o��mf���{�kx��tL]��{DvZ;�K��mJ�<ǲN�YYv��x���T�H�y0��b�^>%#�=y��A&�f��yF�/M��Vzp����n��4��w|�0��}G|򆤼Bf7������դ�Q�D(h��,�q~ӝ��R��rr��=�O�N.\o&����%��z��+�+�$
�cSl�SN. u$��w�F��jiHҧ�yh��o��L�,���l~�ʭ�I�	�{r5k~Nu%5�l}���*|$�x��/o�Q�^�39�e��/�{��u�G�w�]��\F�>��ݖӘ�?i�c,�[�u��_��=!n���7�I���F��2���� X�sS�v|P�^��8��#s�W>*�{�Pjͪ�bl�=�X�"*9 R�����Q9,:4�a���N��t�����z	�XG�0:�@Tr~�~�N��1�4��=��8g	���RF\g��[7)3�z�k�v�Ҕe�@�C�Sq�G�Ft">=����ӡ7[�Y"J#٢u��<����3q�"<]���ȹ�H�!�[�b knv�˘�t���9�ɓ�|�����裏:U�٩I~���:K<�V�m٩8?5��py��5�ѯ1���'�t|��2S&�Ƃ��u�FF#���F�QM��CF$`u�����o~�?���q���Q�DD�_Z�3<;n�/�E�z�H�2Ń�v��Y0�r�����5~����0�Ty&?'���?�{�O:�d,���9ә=Jp��Ѥ8��|ڣ{r�s��v��>\:�=+�h���;Oҵ=#��9`']��"g��+:
����'����{�^����_�7o%�qqG���c�;�:,�@OqL�Yg�c�HM��+V�s:uݶ�I�2��5#_\�`�I6M����;yX��}6�e]�Sm0��ϡK����W���Y�4dG����oϛ���K�?ض�Y�c$�M��Nf��1�GeC����G
�=U��К�8�aq�J��5:�����10-���ɭ ��n)���M��������t�uI*��7���M���3W�6�@��Z+ܙPz�V=�$]I��u�t���tl�݃��uΎPU���n��;[����T��]��������집U���T �Ċ�������,���WK�������9D�7r�}uRbS�����K��hƩ�(Q��R�Y��}���k{̃�*���D���I�W�:F�87��_�)�'hG�o���	� �(pj�nؔ�!ݝ��g�*#0�,�)G��rCeaj@���Y�_	�4X����uf�)�dj��~��!��4O���Q|�O]�d��:��:��?� Y���N��vI��5ge&2��g�Tx�����/n��>�T�G}x��?����޿������?��ԉ�_N�>��S��Փʛޠ�1V�j rnǹ�C��J�Ξ���^0ZxR�hH>tTFɫSy�Mt����(���`p������m:�X:�:�x���lHyp�/l:w�}����;�N_5%:W�F��~T8�#�� ]��>���N�U��\�d�!wz���߿��?���oq�?����Y�2y?~=�K{�T���@�#7�������|ۆt�K�z@ޜ�EX`��Г�Sf�\M/;o�Bwi����`�#{m��(ٗ��&�w��]GǺ��ތ�n���k�v]nÿ?�Ŗb�m�:��������y���|�u��VG>�ӎF��^�!-{�W �"��=SX� ��}��w���@�^�{�2���<{4)@�G�+�\�\�g:3�=7/�)˽N��;�Q��m�I��%I�N>���i)۠�]F�Sy��u��<�΁k[�������o�Q${��5�]N_����Ë�6����CC�:g���=a^H�=�i/2����&-1�k	X����'O��Ĩa�_|:���=Ǹ��*7��r,����{�皀��q!I[WU.B������Эx��<}2�2D�;P%nC��S5�z�l�z�s=�J\0��i8���D�2R�N)V�z*��Q��kR*p����^�8%եZ��L��&e����ڝ2�����,e��اӕ��G�=��Gt������R��5���b{4�3J##g:Y��O���z}�~��w�E԰�����6x~�Qa��g�~��Q���A�~ey�)��>��|m���a�*��"���M�&��u�@���x�ì��:�G!H�:տ�������ſ��u�>����pX�k=�p?#�m��Sˤ���3|��9�C��}���|�f�ӑ��_��%�N��;�߻���[h��e�e��������H2��3��۬z����6M�������Ag��o;��ʣ�S-?M�~��q���'�$�V�I�3{*O�4��?��]�ۿ���_���zb��3Z���<��h;��tO{"{Gm_tH{�m�A'�{-]б���9R@kY��+xq����+��s7u½ԣY\���S0�}���8�q`��a�����������������Q��v�H9	F�s-t�k���������QU"��	�m��(z��{��A�E���P��T��]7�5MW��˼�o
ӄBJά���"ǭ��¦��#�O^9�c��-����<ᇩ�\&��c���ά�5��W���{Q#ˤ�;0f���5���E�RHz�`��������J���c/�%����`z���RF<;4���3�N'�>�C��-w��������3�i�@�s�?�|����r�������6�����K�#0B�8����g{
��6�^�/{�2/_D'T
]9�;��f�;5�f��	��\:Nq;�F� F!��bCG����0uD,  @߿���VS���UEN�u�sr�S�]�ĥ:C�	x�P���J젼���"e��s���<͜4��3"[��4��hR��Q��L��nS�I��~jܦ�^{��Ń��M8��/�LaX\MqV�%�4P·dOs2�Q^#^������'�-RШJר��;��k�q��y{���Q\��.I�������NY�3���	�\�`B��}��rw�>g��a�~���?���/�����_����T��Q��_Ж����,F�u`��[f�v2��u���װ����S2L�5]�d�@V5Ќ�w:/��S�z4�/0l9��;owd����]�C����V��*� �%�̄�I;�U���隶9�~j����?�m�V���s�o�=��'p,�M#�ĕu�s[�-����"�}�)G/FpN��?�t�q���LC��f��t�)}0�:�mé��n����:� �G���թ�c����t������Yu��J�@�SP.�+6ƈ��L�Nm�S� �ئ����>S��TL����5�dh����K/��ב�Yk�:� ���Ǝ�[$��y�g��O�2[��Sm�ߝ�/�0~�V÷d�ݼj_�?O3�s��ցs�B7G�N^r��Q�pb�<N_�ixe:�/���F�+W��\|��#Eܤm�ֈ['_%_i�#N9b�|�k�D�N�c�}2�M��95v�S�[���:>�⫋O?��❷��{e�j��)�����S@��
6�(������w/ߊB�И��*���k��ɽ'�=�K#v��yx�5z�-���0��2�]���m4�Z��:T�E|�\��$5d�t����f[y�Ch��������!��\�`f���멪��ʨ��t����_�eD�A���	�~J`8������J^0f��s��ɖ\�I[�dg!�$��R�-u2�;�����UXғ�`s��̓�!�.9Nj^\��z��,U7���k�2����F+�)��V�^�$���I��|eģNT�y����~Q�o����'F��G���16bv��|�Ȉ%���ѣϾ�����/>}�u#�.�y�q���E�FW�͈�ehg�Lk0|wb�.�P�~�W�C�G}�] 1j ��Iu�0.w�L�p>��N7�ǿ��⃿��{��qZy�)Y�����`�Ǟ��v����u��S�����B���mKCt��'����6:�驎��\�U��xi5����#�F�5l?����������㴙*�MO:�:r�6:�����ӝ˥���_�
�a�t����9'��L !g�s�'v�R&a���|�E/���G�X�v�H��!m;_F�����}����y��ì�"S�`�e��W�,Srlc?N99.x`n=��<\#���OoM���$��>��.�*���Ot%�7�7��ĳ��8y^�{Wi#O2��������i�8b���[���״��6���Գ[�I�s�ݿgyO���87�9��^=�*tO��S9�����ؿ�|חX҆]߻���<#��{��j�U~צ�l� �"����8���l�t��2�݋M���ڎ�ZS����Z��;m)�[����]m<��N>}c���8{��<d4���K�c�Dԍ�c˺��p�e�)8нjy���mf��?h��Ma�����D2�#ۤ��ᣯ�|�ٗ~����~�OQW���^{����/�]�yĻ
���N�_f}vz����$c�{�?c<���oB�+�H:ސx}��}���i.��ef�!��w��#�d���ׯ�dd�et��Uh�Ы���F6��a���`N6�]Z .���7���A�3�v䋀/�����S�ܭ
Ie-��?���0:�;q�t�M)7=��;	Ҏac)n�u����)|cNj��9��㠄�U�Q ����l
�F�w(YD��F.�������7�}%Sr��ƶу��17���n��K���)���1p�}FO�Z9�����-I; �#��b�(��a���P��	P���NÞD�[��[��5��,�Y��|������&����1���t��U*�Kٙ����T��t��<�v��(N�+��3P
- ��ҶTG�lG%��RS����q�>OB[������	���3����U�{��ܖ��s��I�1۝^ <�IX`�*��ܹ+�|-�|^m��C)?�h���'w�?� yЛ�֬q�U�r�4��������N�s�S�J'=3mP�8	���F�xxl�v���AԄ�D�cˡ��g0\�w�y��,�;�u��`���依��m�y���'�&"��`r7F�t4Ǥ���G�6���[��R��-���-u�)�Q��F��c�S��ƫ���<ٶ��}�w�d����ёl#;�U���o�ӟ�',[Ud��6�a�dW���D���> &G	C�:mb�?�	�|�r���L[m�i�ͽ�����=�[�����W�+��/�/)FB�6:4c/�l�����kϪP_�f�l���t�8�pi���9&h�7K�� ���7<�����Q�|��R>x�f�s�0|f-��PV�Hv�t$m�����Dg�_�m煐$<Ljt]�:`y��*e�ِ�*gg��G��<�.��>�D��[Y�o*O�=��K2�瘇����,n �naG���Lt"��$����?F���\=�ґ�޹���>�R��|�vh�8X��E�ė�s\�n�I,s���Q
��Hm��9�� ,)J2q)&�>i�JX����Q�Y�	>
T��J �0���b�N�N�0�=��>OJ3�W���粼-��L�ɵ)f~v�;Q��Q�����d�l,^Ȳ��@V�<�>�'fX��U�g��F΅��`��� ��Ay�5|��4��Ėc���y�}�z^9�F!e:j峯�����W��i��MS���N����z��?����2rf.�v��.F'�G���?5����5�6�𾎫���*HE��/0tÓ��αr7r+O�2F�TT#u�d|���,<�<�2�K�N��0:r��e]���O~N����8X.xӺ�邴�k���f�S��+�fT=Фy%l��N(�+o+P��Mw�=�)�hB�����{�M�K{����7�a��F�ΰS�^��k�&Ӿo9�
��s�l�����Xd�\E�u¿Ail�	��]h�r�8ތ#�Ck~�i������zX2z�'���)j�}��;�xGlÆ�7�?z�&ɬ���5N+Ӈ�\��~T,���lآ�U����垚 �^:0�S��Lޢ�]��  @ IDAT��/e����������|�_�O#�t�z8ve;�3��F?�w!z�����M�h��'���(v��㭝���A�i�����|=�rz<|~�5K��AwD�K�[��hb�2L"� �y�I����Y]�˹��d��^����wF9j�vG=jS"HS�1�}��|酵����{�3*l�IF�8A/2r�%\�1ps�eU/7��
v:��%�cF�9;�TήoŁn=Cu�n��tU���6*tD
;����?�:G�D���2��u�)�8\)\~�{�%4f��J��|��ڇ�_(o�[��Ŏ���w���&����W�:�ʠĕ��8`̽����ҥ:pਕK�S�{r(q¢}i/y����چQ�Pj�ڎZ|����9�(���HTT~��g���%��k��u�&~:ò;Q�pPP��C��<�p����4q��v/����n�Oʠ��
agm����]�r#7�(�8_�5~	r�0��f��^~�ϮDL�z�~����xW~�*��������'jȣI� ���`�1[�Jx�7��D��'��+�3��5_i�/�9��	�kj!�=�|y�.�]�K����������-=�1�޺�>x��A?ʎ�U�8Kz��1T�$�8��gy\����[��0��@vF/b4�d�r�SU�H��}����BVv�k��r��jt���p����&�u�^�g�(>:7��*4���$�8���3��(�Z'X��.���^�s�+��MJ�/|��{~v�fمs�a���o��S�C�f��^U����u�"�~�=xE�ʩ�īv��1��)������sHb������#.){�X�k���փ#�rd�~2��t��Y�@B��g��iI���G.�~�nw{$EY����������R�C�9�c��Qܻy#r?����5����n�&���pr��x�з��x���)�����ƜF�3���)�ϳ�̗��FƝr��8Y3�2�
/��{n�.#aY+�^�w}�O�����J\���y����ŵ�|��O�|Z��/u{>�`PÁq�S~s����۵]�3�S�r��r��+5: x���D'/�C��\ӝ�ϲV�y��ϲ��LC~��W�gj>6����,��Wܾ�89^f���Og�^F^�h��N��x@�>'���a��䘶a=t����`��9�>ӆ��~,���u��rAEs��n�.SI��+�G��"��,<s��:�F>��t�d/ )JCd�$�,C�dotSs՜���LSpJ���?'or<ʑ\�6L�������y��(�Ґ2[ǰp9!���]�,�q�h�͹�)�hŰاu�7��谿L���HM9ۿe�b�O��`��Ο��sA��WZr���>_��`L�IQVc��OV��x>Ot���t���3�>y�"�<�Ũ�r�^�c�C�q�f�~F��Y'�j2b��QdS�O�<ɓc�zq;OY�0Ӕ��i  ���R�P��r�=6���Ou�<h��촟r.�O�}�?:᭗hgG�>�t�Q0<�?G�h��/.C$�w�����v��4�v���7��0�¿3l�t����)�O����I���2p22&����xR&��ӱ0����o���CΡ�1,�UW>�c�F���p�N�I��bo��;�6�Fߓy;$[����)>�u��f�`�m�׻��jt��In�;���|�j���XѤ^��h�gz�����E$Y��z��_�X�*�rt ����ܣ#tlx$~�v��w{�x����t�5Z�_ֱ^�S2�oD�eFO���)�����m��S�p�v��kDY������.��d��,� }ֶ���o.��_�5{���m~���D�����������mr��J��њ	��+|���'Y?��7@_�n���'����	�(��(�};`/>�w�`{g���Y3+��2�E��B�,��FD�J�������{N�,�&lGj
�~�l~���z"��7����Web?_��3#������Ͽ���W��]�����k��_�.gшS�c�J�B�7��ӏ�~q7N�[��6�O֓�:n?1]�B�ɬ�� r���F���E8zO�f}�矶�G����M�,��]%O7�U�r8����Q�KtE Y^����{�!5}q�( 0�Y�h�P4{ULd�n�&��ޝ2&R<X���a���9�<E�]�5���ZZ����yu��y�)�Rj �	q�b���bQD\�#��o�O���.�.��|�z��9���^Q9�a=���<�hR�m���h��Ʒq�)��ҫ��7�����0������>1OpF�,ַ�"{o;r.�l�(���u�J���/�,2�\���13d�,��ߎ���a�ɰ%?����9�v�
o�Qpr�8ё��?��c���~Թu��u"x�Z^P�_��3�od�ǹթn��M�U�tj��\�Vz�r��Q|�_EO�g%L��[��Í�\κ�q����"?�Ӓ	��3���i��[�2FF6=�l�6~�Ӿ��_��Pc��g�8�.Y��U�W�|�0��^�瀢���en��eV� 9F<�[�#��p<�;=:�"�F�N#^-7Q_;�Նw�`�c`L�#�ԫW�p�v��\a`�>$n�*L}S��]�)��?������-U�؍ڑt���1^p����m7�#O��� �s�`�+����zC��a��Z�EP�w��Ǐ.��w�����zf��(��	����kI�����Y���z#�[�<���8'W�m]l~����7i���`�)uHs~!_�,���m��)=�h�#6Y�}�ȽrHEv����sv��@����,b�.�&Mƽ�XR�l�K�Fh<����L�X�d�(CVB�?���I���7/.�3SՏ߿x��7z��0�^�ʧ�23�e�JKa2���3ڵZ�5ݦ�"ٔ�xk0sD	�9�q=�̌����'O�������<��s~���h3B����I"G��GR4>L`�;����f��e���*��n�rP��F���qf�ʸsO�ƨ�݄�s_#�7��k,���"E������T"��Sb6��'�p�n�4�%X��F���w�
a�c��d�a����{8�7��9��,թ��D�D�7�+cQ�Q��U�l��	�F��}�)eZ뷫�:�S�m�R���Ea5|o(=��y�[_|e�U����#8�t�mw���'�N+4C�)�k�F�����5�?��Ȩ�7X5O���>��#C��:q���Q4��'�d
����j�������e�78	ŧW<�ڻf���a*^��=��"7�=�t�p]h�����v��{U8�N�kt��	�7�@��Dt����ؓd���w���t!�f���t�#=7����q�>NJ�#-�
��<<��~x�1t7�{ �ί���4=|*�r�H��.۬4�����v�J��Ψ��%PǞ�������m;��~ח��S~ip���ְh��o��rژ�9��4�̬UH�C�>T%��r�~�ܦ����xa�ۛ����=O=퓗V��Ӻf�D�_�K�$�|�x�Է���Nf���!�h����w㠽�5o�\�-_:�ӟ�v���-��������..�aF��V>u�#e���u�Az�L�y�3��<Sr�;j�ujF���.s�^����z��OQ�I�z7}��x���Ds_f���v����] O������[xXW���$2:aQ�Y":�W����!���\}���v��ރ�B�U��� ��ܹ����6X�	&V9 ������ٶ%t�����_^���?e��ϲ���޼''�Q3��~]��O��Fw=_�8�>���� Γ�=��f�L�3�v�%���ʙM<q�7�a�`�/���=����C˭8��,�G���� p!���tw���k��IC]G��G�8_��;����\��+��W��T��o���|�[�� ����"@�).(9X#C��J�A�ٯE�l|ñ�ϐ伲!�Q;�}���Z�F�=��5 .�Kq�N�tYUx��]�V�� )=�z��̹0Ro�Qk@e�6�S1i(iI�`��j>S�.:
ߑ�E��ڬ1�����`٢�8_i4ޜ�T�{��Z�ȇB�лV$X�`���Ŕ1Leн�Yg6O�ɦ�{��L�[j#����8��;-z��:��
�t^�!���#_C��_Ӧ�9ԭ��gS�~����o�T��m��ħ��rux��Q����=�z��N��=����fo�I� �N�+~�D&���\��A}pT����@gs��V�������Ĕ�aӲ��Ǵ�_p���T�!�f��K�8�����j�g�a!���Q(�m��5�������3��9��S���-#}D7rf?+�f�n�v[�z�e4����0�`ôY�N��4b��զ����&��n�' u�l�o������6�N�h�/]�ɥ�����=ȈG��ü�ə��������z9��qz��}��;9��Q�����˼%�W�֛����}2�x;o
�U��8ai��f�i�u�r��>��rџ���D4.JiP$}.��a��#�e���s��k̛�m�$�@L��DF�C�A��:��i��|���	{?k$�\��Ѱ�{���}׼�e*Vlz����2oRr^-�����Ҩ�.}Pf�Hf]���'Y&�7�=��l���;J����Хy�u-��Dآq�1�vt��Y���F�=_>�[����~"���T�:����$G+�h��04F��E0F�۷
�
g4�g�Z=� ���e
T�$�ty��4ǭ˯/��_~����.d��`ӊ�g8Iz�YѭC��;4�*A�D7�a��ly��I-Ը�M�O��Eo�m��&~�"'b��*�	R(�:z�<I�(��ki�\�'0��,ͅ6�8sfg������se���o��q�J���o��b}o�
}�ROF�(�'�����ʓR戾�)þa}*<�]〧���xANx�S�NG�۹�̟0����?�w��4#}��<dX�C�cw`�£�Q%��,N�|n��quBo`�6S~vǻ�J�7�S��z�8r���X\:����!TfF��9�W�54��zܨ6
_؋G�	j��E���q�Ǥ|�U�[}������v~e8�ih�b���x��ڱ�x�#=�V�OYF���O恴�,W}�O~4�R��+������%�����ND��5x�9�[I*8��6*N�~	M���tj�̱��~i��u�v�rMfmG�Ǒ��t�.j?�g����ͥzspv��Œ��ٜ�(ESW��K�A�VF��y7��d  �R��t�����+�T����=��׿��S�V׃}�Q�`P���H;�>lJ��	��`3���G���I3��sB��<�T����E�!��S����QK�rΨun�ƦOI��H����/m�'##g�W2������F'�G���j�C��b8�Gsd�oz�ؑ̈|���ſ��O����_���e���\�%�4����^�ּ��Y�'y��i����Çu���z��܏�LI�4{���,�w��mT�=���u�3?����D��G$ʋ�B��I���:����s���g���<뤽�f�����|�m|�C �o�����G �M��a>ӌ�����ax�F��|��ē���tu,�h=��Iw�{�0�<�Y$�(���R�>D΁�t��9�W�H�A��1�t���:RS���#\CK1��!xU08����(nι��u�
�O����3/N0С���"�gW0�U��WJP#�띮*�JiD{�]���<�o�v���l��'={�yU�����dq�b�~0_�w��Ȟ@o����?����f��}��G�w}�	'�C�`�N!t�%-=ç��)�Ϻ�p�Q��Q�۸��F�ǉ9�1<^���E����o�L�?4O]��=�/�;~�<��7��W�q�б�Lma@���A��X�-���k�w2N�qq.:;� }*�*�3H�=lb��ĕ��W�HS��)���-7%���~�p�w���h���;�=F�*����u���nTc��y����M&�at��^0�w.����X%��#����+��	N��F;i6! ��۹W�� �ڣ��]t��Eg:�/"�l���ld~�yh�ū;
o�̶�H��[�e܋(�H���g�z/���c`�	{n�P�H� �4ޏm{�q7����O�,�ľ��^_��������3&��ޑNU&���K#>�?����1������R����5������32/>�	|ݪ��]���ճ���.y8����o���p�g&���F�嫾.��e^�J��>M��8"O�V�/�08߾x3ts�^�+���
d�a*��܋<�?�ڭgYs��g�׬�đ2X�/����Tf,y�e7�����^��^��?�a�ѽؗ;tM��K��']��z�;�MF���&e^f��g�e����C;b�Y�<����yx�t��"��T%���l���d��*o.�D~e��uT�
��UB���(�X©֍��
q���ޛػ�7}���k�3��V7��ŊaO�	�Ʃ�BF�9��<�pҌ̍Sh7w��0#�"����8���|�/)M�H��'�:F�*�j��9�/n��7o�ڱ����sC<��ꘞkJW�Z:8�;�<O7S?��V�l)�I��'2ß(��,�k�'DJ={��'̚1�v��Ȃzڢ#��l���.��w�����u4���������=�y��~yk�柞�q�18{w�x�#���̐����h:�1%x�wn��B��-��@e�m�
+���o�����OƦ�x�8v8ֱ���[V�}�@���K��t��s�*�;S:�Cyj2�����=����5u�͠�+���$�H|[���u������@z��|
�i�=H�"��*�&���<�3���X?�P)��hΡ^���C�\����|g�O�鐧��tX�����G�ʷj���i�p������o� �����8X�d(	��s~V�?��q���<L�8g_�;�r�,1�a��VΔ��p,�[�{������C������G����&�n2��摮O��U`y{�v�⻛��f~�e	[�/��0t��3�S��[�gf�2�54��,���6"r�C��Q�m�3��.�0������#�s$�ȩ��U>wxW]���ڧ��HVw1H��2�vյp�U��gq�>��\��D�����w�u�7��m������w��:�|Y�s��eJ�Y����)����:/�����[o��-Eg` �J�|�ʙ����J*Y��҇yH?�ud�~s�,ui��3�I��e��^gWW�!�f��|�q*��yPz�񯺾��66��Q�;��(kC�PZr=��W�څjl'XΌ2�j1���)5.#�~C	q!�	H�l��!�n�MÏ�؍@�$m�'��}���ҩs
,��p>�)h�LM	��_�@"L��c��R-�uq`
�|����9!�u B��-UTI��4��< �������G�.<&O����I;=�:���غ�\���N��}�R�	:�r�`�&�kG��o���g�[�O1:]�ris�3*�d:��T�#�,����/i8ofh6�~�A�c���)Z����a�Kˀ:�Wi
4�.vď>/rW�ᕛ�a'������I��t4g>�|���;�&I�<�|���]���,Ƥ� (\p�����Ld�'�m��A��VA�jxhc�v�5&1 ?85�z��ħ�(t#܌9gi�]d�A)��נ\��v��n+��������|��EۖN���H�h�;�;-�	H��:�F��,���*�J� Z��m΂�Һ�ˣ��,�s�2y�a����3� ��V�S���s�AT�`����9��<:Be'ǔ����[O謋-�qд�Rw
���u��d��3��P�][:8W�{{�j���t����O2�����ST`����I�1�]�E��O��>�#�d^q������-R9�����N{�f��ζ/n��h�R��f�݇}q6�����N��Wߖ��0�l ��T�w5�0W�"�3o#Zp�e��`������8F��}N|��?���� ����^������9(�����O�e&̧�F��HK�y��ip�V�#>菼�p?;��k/d�:�:�G�}}�1Nm�638}DGO�fׂ��������ٝ\3�R#��3�`��y>�n��<�|�Q��x�_�y�6���L�3�ڑ�L7N���.l�;ľ|AQ(O�GN�2ea.BN��+��3m�e1(Q�P���|B����~��G������)�7�x#��ݝ�}0�s�)����O���@�t}�ӮQ;8�X��rKD!�E� 8�d�A�C����C�PB�=;^��A�JYno�*}��ʿ2��;Z�:��H��܀$~%R&�$0 =ڑ���7tL18OP��'�4�QM�4�=���9o��b���Z�F��=��� C��7���_~�����կ�u��`�� @c��sN�]{����$A�i+g��SNp��	�����).���t���j\2�,��t�I�v͡�Y���G��gM����nN�8��T;Q�L�TY���iZ�o�u�T5ͻ���x5? �Pn��f-�|�o�0񓇼�7��i;� �'��N��RC����J�!r�}��Z��Z����J|Ćp��RǴ��4r�V�=��O����L��L]K8�3tcd��@��D��f�L�lT9W�[:��lG��,u��"�f����o����#èҤ;%lu�p�}ۇ�+�ؐ�k��m��g_&�I�n>#j��bg�z;(ڰ�I��M�m���G����e��L�Q�$����sxZC���)�M��w�~��]�6��L���ë֯M��y��2S-Y�U{Z� @:LWw���m"��}�z.���-���J����K�����^'O�����r���lu�۬�%��k2���V����%N<�T�f��͹�&lS�?�����\MC~����߹�(�f-��z?�j��#�����?����ʖy������g�<�(���ٳ7�C�)Ǭ�|�&���~�%}"��=�|�6C�J\��n<ڴN�����pw'���d�Lq��w��q��`������}!���j#�?T�2�z�Iv��X�e�I޽)��X�,���G ���<����%�۠o��d�~R��� ���w���3|���WiE���s���p�p�4Nس���,V�#z�.�(ګlְA�SANP��Vo+�$r�(��#�k�0䚋�*��������a�z�z^�&fb���9I���qf�%]�a�� Î��� c��9����-�F�'��ů^�p��e�����|�9{o����p��m��� M�N*�q�����h�?9l�l������<��Ae��i���c܆!M��ͷ�6��WB�Q�zh9a�7G��Ox�.���2T��5B���[C 4X��On�dRS�TD%�a���
f`4@����ʜ����? �֭��c�]���|
���˟_q�}��R����\��z�����o7(�Tg`��sT�ڱ�m��EA�ϒ����S*i�����#w-�]�t�V�h��MDB��#�յ�2�x�훗�B���OQ�����c���Z���3|�x	�@N	ڸ9K3U�롬�ѫ*�����7k���t7�L��і��T]��y�����u�S��%k�L&�$�}�+bg�r����؁ ք`� �7���Bnt������@��w�j��<�qf�7���q�K]y�z�A9����jOyD�x����Q�;e�����Y{���Xu�<��zs3M�M]��0@��bI����"�֏�j��	�լ��p��U�y
6��Jzf`}<�ƳWN�6�6�n�A׺�!�S��x��!N�7���>���t�p~�m(�/�N����6��u�ì��f<�m�;��G�G���ҏrI[���S<4�px6?�y�=>��#J�T~��e��̵w��,z���"�u�$.�y�Xx�r(c:�^�偓3�0`��у������Kf�@�x}N	)������L:G�8��=��(���/����cY͑rK���ǡeP�S�{|��@����{΂�:|�ퟣx+a%ﮮ�����ӕN7�-��Өå33B��W���:u%dD^{muG�Y�8��y-#���f�0Y{c1�0©�;��6�A�)"��l��G�B�m���Aޡ�3%�z�2�5��ԟ��tpt���~=l���I%�����w�ܢ�|x��ï�#���x³�G�.}gɾ�@>�u�06q�x��w�yg�c$3�/M��C�Gϱ��/���:��y���-ؼ���c�=M�ε���wc�nڤ'y�Z�m��V�uD=䦨w|Ұ����ki8KZ[��՝��)�qi�vL�+����O��0j~k�#(�8<�H>���G�]S�~����蔇����m�7/��"y0����٦�L�_T��}����i��m[�����l<�u,��z�C�?(�2�u�!WN�Mz7�\������ʪ|���pE��o�v��5���ϐ���F�E����ђS�^��q#<��t�r�-��8��y�=O]�5� ��qo¬��,�6(����+fk���������(�!;�?d1�Kgo�:�
��2�8�.������34�}�����%�٭,�љ���E�AY태���P���;	a}��϶*�oP�;�2}��>���)	:���I���G�Q��3#D�����5}f}�� �	c��~�݄�	$W�=�r��C�Z��sV���������&���Bw9��6��__2�s�Sq6���)�<�<���)������Dk������f;l��/Z���(r-��+ɣ�<��}���t����	��|���F=�G����n�������q��=��z��T"rr����takyr������CPJ*[�7�R8-^I����RM���D9~N1��нqz3���E��<�[�٠�ׁ\E�4\SUv���6S�.�s��΢�_�}{�i�����r����@���Ό�g�t~��i�^FP���y��z
��U�9��oc���dJIo���^Sre��[E�^u���L��aڈ�e�Ԉ�d{h~N���Ǉ_�q�7bݨ�7C|�V�ũ�\���>lF�$h�o������?4�"E
�4��R��(]�tg��>l䭙�U��鵿���S�*�R�!�È��!Mu��Շw�_X�#)��p�86����X�g�a�a�h�%�Eۆ3gމ�i_���Cg�8����
��2CJ%��&��ѫ8�bX��9����˔��Ԇ�wL�mrg��q�FHsா��'��I���P{1f��+y5�6�,gz�J{d{Ýt-�_[��:�Xu��4�7���(�П�F���b񏮶�T�+�\��8}�O�?�\�s��OC벽Ug�l�\+|t�vi[�f^�E'�o}�ȵ���S�ԧ���-ƫ���c<t��wyLv���OX8�8�-e,��1��?�㖪B�X��q���̎I/�AqT�[mƒ��ugc� ��7����uތ�:�����	��9�Dv�A�I
��W���Ti����j�[�y���E(*���%�H�0����*m��	���%�O�DУ8��p�\����mf���ɧ�⌹�H5�g���)�|"��q�Ёl����`���]�d"#��CRj3�8��e ��88y§�pA�"T��Pྊܶ�|?���?�t?c�;��K=����,�>ᵫ��ub�
�o�nʵ<7�"s �N�j>�/��H���`���@HP�0͹�{�(���V^o�A���
��>W��[y�>�k��c9g!�N�3-��� "�LT��%�鐤Q�4?`���$�ɫ�4 �������q����S�6p�g&���_���h� \� �<��2�Y�+l.����)X�8�T:��3���=�D-#vi��bf��Q=w� F~줣%�nSG�~�!�DH�A���t�_�g$ﰖ�֭;AG�� �E_R�����:Au�\m'.�jz�a����Ri��!E����˸:M����k���xl0�FS��l:M�Ou�Ntt,�έ�κ�QGgtYS���-2oB����π/~;�7��t��,];m��>6 �����a��3�|p/|	'��s�Sft��t0H#z0��7Ǆ��\�9�s�gaB�����or`R��[�N�9O�AP��O��>d��6�3A��t�SN�zX�p���jQ?�ˑ�<�9>ֱ6Xl�'*��7�3�a�J=Ԇ��M�k�f5p�����Aڑ��V�֝�k�ħ]j;-rL����r��Z����#���L�_�JE!�_q�%]���8@WnW�����ik^{�?ǻ�쐧M��gϨ˫/���ۙ��M$�t~�?�n�b\�-ۮop��x�;�n��G���l8�-|h��^Y�\��_`G���M8A�n>���(��K �d].��xRAd��D����¯�\~�ۖ��Y̯� ��x�Ro.;2�O��*X(��9��@xI��2ͯ=��|�1��i���rˉ�;��c��K=#�y{���޻�xK�ç��vF>��=�u�%���މ��l#���&ބ��\��"�>:�"<[��Ҁi�\��{ׁ$X��k��V2v�n�y����߼J�tv�kt} @�r�6V��B�=ci��u��3� �.O|T�W��]�����w�����%��2�4�Vx�CgR�Yz�hO+��휼��Yu�"*�穾!�J�$��Y�%��<^o֚$��䣕#.	ֈMo�Ζ�Ge5BR7x���)i�g���!ce�0+?�,e}��ʴ��d,�XTB�����d_�Vq&��� c`�d�q�Zt�aCz��ܺ&��>�������H�v�3_��}N�ϒ:v�n��':/��?;6_A���S,i(ύ�ϑ/��O��X4$;����FO����Q����hG���k��(�1}f�L7-�KO����il��s�uѳX��A�Gu��M;B���x'��k�֙N���o.�7����|9�����{�n�u,m���]��#��^�G�R�)�i���S�as���e"d'/G�q?K�Ε%MC�V�8F���8��E�%���:�~����{���be�QW�� �q�j{�p��~���p��:�欅�4��=ge<L6�M��z��O�=�t�3xs`|����_a�s��l8����2��d\H�s�L:����/�7�!��q�����V>�s;���eE�q����T"5���0T�6��d=�� =KxBG�u#� �0���B}�c^���VG�βe,*�൚���{ۛm��>u�}���>6�TF��/hr�0��>�k97���m:`�<�r`��v#�7޶ooU�6������g,�ȓ��?�M�G,;z�}��s��>��y���M啚��m�I�V0-�ڣl�CPG����W�,�̳�5��g=T�E���n����\(;/�y�ح[g,�������������݌֗/Ə8y�ۆ����2��^��*S�p�޻�>�ɇL�2s���������4�j	�`�0j�El(�)�eԘT��Q�јe�� R�2lu�0�i��a:y�<{8i���s�JU9H�����a݄r�0OJ����z���f�N���IH��|p� ��=�{��̑I�M"A�Gv�w~ԣ�9��| �!�������T�z%��g�qa���X�Ǻ�w���������l'��
�c�|o�ׅ�w��u,'�R����af����QB�����L��_<)�ԧ����nt�Ȱ�g����es�ý�<�6ȣ0�G���>v��Ӥ��+ڃ��n�`�n���4f�j�t�t��e��P�d�61��w�����][�D�E����u�����χ���e�|���yW�lK./�G�(S�UgFbqs��r�b��_ʞ��E{F�Z�לA}����<��q�$�Y�.�pSH�<ܻw�ْ燯����i��&�t�]]O9���	�H2�{{����8?��k��~�uVy��؜70�U�hp����=v&�4Ü��ô�Lӆǎ�3�l:�Q�L���L�����<B`���7�$���=�x��|�#7|���q|��p�o�8�6�����g�ܔ�;��p4��N�*3O��:��P��[ P�i��,�g!�]vȿ��@� ���[:b�f�c���OU�c8�ӎ��2��'��?�̓.3�뼍x�/U�g���-�9��zl��!�y|h)��[\[�7�3���<�ki�KG�(��U_q�ر� �>�ͷIw�/i:�%��`!_�9׿����|���?��e}���oI�������2�����6�65�w��^ԩB��0f���8)���j�C��g�k����c�K����<�\~p������g�lOq�I's\ʄ�'/^>g��c�@y��'���	�O!*ɯ�sV�z�*X��OB2�)a<#g���[���8`P�����JS95#|i�`Gh"%��YVTV�{
]n�[x�����|�L9��k;6�l��P�ȍI�����ҘCP�"�")�|S�ⷼ�1��᠉�CKr��R���a��sL�8�P6����)��z���3���GL�x�ݻ�w���ǐ�y��9U���<��,�R�w�͵i=c:񡯋�z�|Ķ|�%�q�-.?�A���P�/��P�7RϝI��{�g(��X˷�F^�n�'���Hn��t��:�/_�y�1Ë�tm��L����i�>JQ���)S����x��)�x�W�Y8̣�;�x��~��߲���<J�4NETP��U��꿶6�������C۰G�c�n	�a��z�%��q�㴷�[�ɚ2�'��2$Skǌ���Y7~��Y�O?�$��3�/G�M�{Y/m?�[��<-�E�u.���ޙKg�W:~�1�p�*5�4����]G�Lz�8�ceW��_�kjt{���&���mz-]�o0�����̐
&���B��Ńr�YA_� �����W>�8�1@;���-D��ѯg�.� �=.-�l�W�Y���~��Q�M�����]?���6��ط�x���o�2�`S�1��1YZ:h���<�@���~�uz]v��ԟ�����[TV�ύ�r��_}1 O	%�����`�IW�*����,�V/��k�U�*����k�	��o�4[���~���]e�Ы��:oA��I��˒��q��zй�U��4jPT�Љ.I��؂�M�J#lm"6|�=)����9����>��q�E�8�\h����:�)�Q��H�qC���|��xM#{���Z~6�)׼��q轻�:��6.��ܟ	+n�T�C���1΅	[���t��AG���*fM�\��1sI
�m7�S*X+ Nn���_����`��.��k�;Tx+�����2��7�@p#H�d-�+٣ׂ� 3�=+�0�t��^ZP�+�$�Q��ja˳87���Q��6����	b`�y&��?x��>�Oِ�5��q���}��8�Bt�5a�vj�ε�(�J��X�>�	�ԥ��#�o��!��]�4d������|��G��������������`�Ҧ��+u�3���V��=+��nrp{�x2��\�S�P��-O�v����Ӱ��l��Yx?�6���G>��ׇO>�$����Hshϔ���^8��z�n�"c�V�1?�)N���	�
�I�����g$���3�o�/�#��W>�\_(����U�`���/�����o����\Bmw��k(F��}��e�Fq�r�y|�N�\ϭs��Eg�o��(WU�Oq:���zm����vb���ҷo�	�g5|�k�yNY��0�_�n`��ʚ���X�%�h�=�1��h�4ۮ��2���j��y�㭒��P  @ IDAT�����I6�7��n���u��mm_�α/ҝ���߾"4� /��ֶ��T��c�6@�O{��b�?e�&̸(�g 3�vpB�?S )PoҴj���/���}Q^ӷ܄nlM9"omKn�%���7{n���5k���Ҩ�۸��Ӣ/���^ab�ang�`;�!QmQa�q&��l��Ϝ����̣v��׊^�<�G��f�AR��Е����ȅ2�GC���#4�-�'������!�K�Q9�/��W�����ㄳ��q���ܺ��u�=t�:��ߚ�9����1_����bA=~��D%ZEc\Y$3��ICO�7(u%�	b+�
-�`��0J%kx�VA�T��Ma�e	�\�m sH߸?���IVi�>aL�R<���8'�i��Ż��ꭋ�c%���re7��� d^���lL!$���ƽ�!8�=�rL����+n���|raRx0g�+�o��޻���¼�C����;��N���y$���pq85k'"�`���� �r���O��.p&����'�o8/ݮ���1��;���[>�[�:c֑��\$�8a{#/��7���q������"g�|�1x�0�u��(#�����"���)N���)_��Q���_�������?&�]f;z�.?�=zϛ�Ge���-MT>�)@lh%����;��ܜ�;���.Ǖ�c�/����z��'�m`�3�s���8�9z��q��}�0�%�	C�L�O]�1�I�jC��q#�s�E�L�<�He��� �3�=��̆*��z����Gf���t���-bj)�pxZ�ʅ#0�B�~�e����,�#M��n�c�)�}�y��:q�^�?���nm��R�)�p�q����Wg�[/��a�@k�<{�_$��X�i7��28�Tn���V��8�i���%��A���T�[u������a-��-��tĳ�&}�mZ�gtNy���͜3^�1M�o�Dd��џê�Յx��tg���V���Dq0���u_��\���t0g8k��6c?�s��tV��a4���׈�:�"�g�r��ǿ��O]�\��j�fX���]�NX�^��Bgӗ'�^��C��p�|zQ[��@�b�xe�e�;�6��?���ᔯ��U�"Ry��O�sp������T���
0FC46 4�a�
Cǀ2�bd)��5��_��� ����s��U&DQ���3���[����-}�	�yF���y_��<���0Mwt�۪���s�]�*rly+�`�)-�9Q�*nu3�+\qu �=oC|\�0�B�-�B΂A*4�;^c��A��Ct����������-7b��F>�z����W�~���᫯����'���p�ǖ�q�p��`���#��5-ߋN�z�P��b�y����\)x���aQ�fFƲ��wԖ�0�vP�7�#�ݦ��`n����'�|Y��V��ϵq;Yub[p���k��7"��b���>&��ީ;s�az�°O�ޑ����]s���}�^�{mG-o3��g�([eT�K}��	���/�<����<ps-��͛���|ӧ�:�$���n��&� ��4���֡U����o���f�ěP>ȵ�����{��s.L�\��c�<���/i�_��|�Jz�*�8�K;�7�����a,y�s䷌�γ����d�I�d �F�'Oq�����Ų�[~��E�B��Aޕ_@�P���P����f�:̪[�qr���cZ�2�L�_Ñ�3Ao� ���_���7e��m�D��o�?�ǉ���b%aG记�?�x"��C���P�q6���ڙ�yq��8��J�K�3_:�]��)�N~�m�:�,�é���:�R��T-cb�����ܭ��Z���O�"�n)�Q쬑S���o��}�N��?'L�8ۧ�㞓R��L1�x�ڽؖ����$`�76'��=�W�F^�Lڈ�����זKE�άg_
t�=��+�(���T~�5n�����љS��wx��+7S�8�܁q_���H�%^��+±ǳ׼�pv���*��|���JL�쟇i�=+�*�EXQ6���|���D�1����8t�����i��Ŭ�~4�K�x�)�9�(�z�������ef��������6�{�N�(0�)Ж�ܦ91x��<$q��?������x��Փ86g`Bv�]�;��L�"4�.��B�x`���p%��xg��wx\u�&F��6�<�wMQV�1K� ����[�=�����g��a%���o�a]NǉY<[O]�_�6Q���`j�:���>\��T�����W|��q;@V�aO��7?��� �4�3��m���=�t�)�~�Oq���\q�\�P�Kg�N���V�:b��e�g���4�!�W-$:1^�W4��S��p�%u����I��سe��a�
�����]�[����A����?g�'�<{h�UU����q�qv��������Y�lz�}g�t����5�~q$N�g�3޾�Ŏg<�t��Z2��}��G���yMg��a���s�:Q��ZGi�M�GƑ]�yk{(L�<ˎ.,�	+k�ؖ�4.��<�n��*����F���7��.��B~�E	�mz� �X]�#yU�֥m���.3˼�J�{�c�0��:�=�)�Z'�q��RfJ<e��g:��	�����
r8��Y�їU���7�ӵ�ȱg&_��}�/6E/8������C�N��W�0g�ɩ��-����f- )h;�Dw�/Q'�t���|lӗ~^�C�:��R���ͺ1�#��̡L��I>�IR��r196�CDx��e����t�1ُ���_����_�|�Q���������+W��ZN��5�Nt��39L4spEA9������C;x��+��:���\:`����}��z�	9�~�ʿ?BxL@T.5�N�����A�&5�j�u����J��*~�����Х�-1ς����[G$.�@}7|�K�
�֯#���,�ؓ�N�rG�qpęCs��a����Q�L�|EHTY�q��K��9.d�|ĕ�bs ?�g|,��e�=�<��/�ĩ��Wg_�&���Ň~��A���C��`p���9w�?��C��o��1k�>��Ǉ�>�����Xxh���8��"�'%p@0h�(^���C���v���p�������s��+o��[��H��O�%@ʌ�e}px'���<�Ϊ>m���N�b�.�7]�#�>"tV˻Xm��]�s�����@�S;Ӂog=�X��~�̘��W���y�3� �9���:��H��2��*�Jޤ��y[��os�t�_Ə3������GE�M`u�Mj+�COå��d}�ݻ�^��>�����⠟~{�9����2K����?yL����=������r��f� �cs=�+ӴI��nϡ��ڵ*0�X>�v�+W�GK'�ʜ�~g��8�#���b�Gۢ�9�}f�D��f>�[J��@?��?�9�v�]tnuh;�����k�7;'�~��3ĎO����$T`o��u�{���/S��<Z������ҳ\�Ⱥ��u���V䱣��Hx��>6�m~+���ˬ�7Tk��`�e�N׋�]Kg�={�G��	"Oe�+r��]�2&-��y2k�\�V'�W�g�'��p�L�)����Hj�b�z�s��U9;���=��6��?t8�wd�s�(�o|۔�Ӵ�5��ȶ�D����3He�^/��8H]>�{J���R����J�/���sT��&��Y��RB���|͋<ts�o�5Sc0�uN�??��0��?b�a�N�3`�=B�4��Ҕ�2�UsN�Cj�Q�NeY	�VQ�
�K��Q�]^ P	��#�,eEKz*�
���N��W�U�L׸u�;8���B7��S�3�q�5p�<z<cF�����iEj��� o5r"W�B��Hi�cA���9�m?V��܎���5�����Eo.�����δ$��sj�+t���՟���G>��C7E|��-O���.�n߽s��7�~������߳��]�G��zgSB!R�R�������ˀ�Wǎm�4Ǻw퍶7Nձޭ������F�YXU�,r���&��g���v�YG ����������Q�g�����D�P�~�>A���Ka�L���l�x�&i3;�P��J��0{`r&A�od�^������pE
/�]��0h�9ח�r-����P�M������ȑi=�� b�<{�r��F��+i���3��93�,�k��9{���͟y���;lw�[	ݿ��ٜGy�)��g��^�^�oB����5��r:��:e|7�Nd�W�w��4yW'K!�!J䞏�����T+4F�#�N���}v#����ÿ�ۿ���o�dy�f��-��̟����+R�e���mHK]M��@&��r�b�R[����m���!+3^�"�U0��#>��o���پ�4i8�pʆ�փ�%k?ḙA�q��о/�d�|����e�	K�2dH9S	��,���3+n�y�X���i��S_��+޺��57��9�W��Wo�h�'�����N����^��1=����>���-�~sL3h����`�Q1�A��Ox,����S���ig'����wϰ�>y�㵗|��)1��_�̒�B�|u���؇��S=��po"�mI^�?GI`&��0	���Jk6��ԫU7�u���ʷ@��]���L��2̌n��/��x�7>	Q:�ũUY���Ȥ��\	r·[�,bJ	 g�^��V/:������R%L�xrM6���H/4)���y�ɔ��<[V���R���Ka��y�u��ԏ� ��^�ؔ
>�J��ⴽ�-����0�����������7iy��}6����6�{�V��{������g6矾��|���@�������]��O>v��_�#^ �ȘH�t����c��s$��[����W'�Mz��}��|;Y;��A���4�������?�?��Yԭ��Nܖ1_�mx��1��i���9��������s�H�C�!�J$a`s�s�8�,^V7�2��c��ƃy���&���oΣ�c��\C{p�YΣ7�S/�8e�1Ή��e;ܞ��6��U2��������K߲��������{�?��۝�^�ہ��w���9jE�wm�<���t��zDfP|Tg}�
�3����<����Ď�'��9w`�Ko]�K>2ˇ�MG�	�W_}u���t�����9�˷~}ܯ�O���m�y�Zw��a�s8O�v�����	�ܙm����>@%m�,, �k>�DIw�Y:��x%jK����c�|�/�W�C�|L?ԾQY���A���t�`�\��.(�WYR�[����'eem���[�����H�[�!��
�^dw- ���cf��Ι]�T�0��IfWW�5Z��U��[�[���ȑ�c?4�3 �0_X/}�ٴ��9ߟL8�S!�V���~NXRsͧ�;�S��L�Nx^ �.�'g�kzl�f拵_��p���p��^(��t�ho�^8U���&��)V2�qy�I�TO���	���
��Z##�DԎHw�R1��G�VaxP��R�b�B�d�I�ʑ�<ŋE�yuZ�8Q\�/-#MԄ� 6_�鶱��PX�z���`_Ε����gx�Q�+��������
��y8�	�1���q���.<�����w��h$t�4fMY��;��g�3`������`�����Q����8�1wV���e�n�툟�)�aT�Q=oˮ�9kࠛ
�v^�C�;��A����0lgl�K����ڐ=�E��}����/�<|�/�,;�B��~&�m��mS�78�s�w���z�J��.\�>Z�4���#C`�M�����3i�i��a�nb)o`���1��8Ѩւ�8`�oy�9��#�);:�y4[�)3�N��V7ܼ��.70�eې_��S6��sp�1���l>���q���<�$�n�Y��}̻�c���l]\3�0���o9�-�J��7"0g�\�ԓ6r�N�Q=\3�
���?e�뫯���cJ�c���u	�o��̷m�Y�萦�踓���9rJit���8F�W�c8�A� ��e4D3�d��+�2��tm�qn՟8թ�g�:yC���4xR���g�q�/��I7�aa�3c�{s���q
*NE�M�z�x�
�r�2���*��+3nQ�T������yD(2��Ϝ��ku�Y���o��u.$c���UoRr����elK��.w�?�łlT��Sfq��\�Θ���u��»�-56�����Щk�^���.V���"D
�d��8!.�{'g��8���oՕAz�5�QrR*�
�`0b�mH�����H�C�Y���� �q̛	N�(7���"�FG�S |<o��4��Hݼ1"�&�j��/���NM�����S�1�r7�)��M���`C�|�]��q��tޗ���
T�0C'�ix�2��뺇��گ[�PLg��u¼Sw�ųg�tq�)ww���_���w�?�1z��GJ���ю%W1�D�FQN��߱�����kو.���
��� �ݙ)��{�,�>�#FM����w:
��ۘ��}�A��×_~�-"�#�����L�� ��C�p�n���T�҂��r�ϔ�2��}��Cvً��ݥ|FGp���Ƕ<�~�5�9��3�"��1t����e��~ʚv!ε�9V�6a��d�)gm��
��+f<�㬊��K�p6须���Z��|��=6��=�}U����ܸ���Z�o���w���!�_ۓF7�ç���g�)��l�m�7��B|LW��F�2r������^DY>D�����=k��g����q�=z�����W����<o����g�P�m�5���r������Bnf�ݞ��������/f<�D�20�aݰuk�X��������]�P?�d��RęQ%w�N�;�&�{-jw�C�p�'IY{$���vm�>NX� o�6�F��eʻ|dV�'H��^�ؔ��-1Y7LiY�	�:R�Z�t9�&h�3�E�)Y�M\���y�^	H�(�8u�vgLR��)�5ȟa�w����`�b1h����)}8|��&iT��R
�8�:�ڃP���K%ع�b=��r`���㉿F����K�f_�F�����/�۱QT�+P֊��6$.=�P8Qd�y��7ĵ}3�R��r�?���@��PA��~	��V�� �)m���&�UD͗B�ϻ�ʻfdY��;�$e�/�ē+e��=
K��2F��1���.��~�N6�e"	�Bs �Ӽo�(��̎o��ܺ�������b_�CCk�}�G*/��� �����y��8���|:s�#(�p �ϛ�&q����r�MN�h˶�d]�,���u�ة;~��h�e�����@�ؙ�B�2�2�l|��9�(�GP*޿�+a��6P��_c���܆����$�iW^'��((|/�ٽN[#~��ƾR��!����M��R�4���|���$�����Y(Z�`�n�ƒ�ʥ L{B�/��Ke6H1�v�ޙ��3��|��o�g�Q։���5b�%�Jx�ik��S>�6��di_֝zqP������ ����2�H�&>z~�yiϤ.�b��\x��.ס������,��:�G�:`:bqb�$y�Z+wp*C؀��r7� \��N��eYK�ü\q-!�u�+*c�g��o)������o�2�D��(��8v;b���qѵ ���b���Ϙ�#�m)`����=a�0�����#�٨c�c����-k��#5�,��Fo [,��1|^�f��|1��&�?J�Q�)�b�h˗��C�-49���W�4V8�)_�c�.mj��H)~�y�$��E�n��_
|�E�L�����k��0��*w�����Ys׉��V����p)����yj �%3&��Y��\��lg��靇�k�>�s�z�
��=:YK��4�DR�y����ifFLz��B�J��0�T�p�h��K�ˡI�i����bh�R2`� �4+Պ��1�A`���--%�=S�����{x����`�������~�=���[�l����:r6�9�}��{�~?��)�{�ſ<"�3w����}<��G�Jd�n�̧�8���S:����e����M.���?�k'���PV��ؖ�c��Z/y����֗w�s8+�Z+m�@�����/9�`=�kO����沎��?�JJ�#�	��_J+��U�Ƨ�֞d�?
,�����H:/��|�s�f.iڄ9֋T�L�E�[:���s	X<֮'L��+��nfb�O{�mz�0��.Z�^�Ͱ����A�o����9��Z|�jfS���^.L���wY#��_����w�e��k.o�X̋F��m(�OE�b�q}� I	s�}[�CՁ�pY��8�Y�o�����s��d�p1�:��>WoϯN��E�;��c��!Y�ۣ�G��� �ێ~��5;���]�)>ew�C�-I��Cs^99>�SI�h����5s��3�ɡ`� QX�(�"m<��#.�-:]�/θq{�i^���?�f�F���Y1�+C����X.��Q�J�:�Є�����?c���Zt t>�F��d�!�c1ْ��O��ϛ��(��Y��
���A+G�H�������ZZՇz ��LX��"]ݏc<�,yy���ͶktO�{��ѫ8�=PȦ�P>��Z�‸�;��Uևq�#��>�7�}�3������XQ�(���y^�JJ��P����J�Z��(	��C~�!.>��tt�r��8b��j<�F1�)�!2�*�E�^�}�pô&���S7S2�)��^Y�C�%\���3Q��e#����t��n(OdF/���0�c�թ�	��s����ŝ�FJ^,� K��Db�p��\}��:��u6$��$����)�|��`;�ʋ����!��)�a��k>�k�!�P�p���5+������X	~���`ig+�77�;g;���w`�3��<��f��QQ�;m�Ψw������w�v�􄍈aø����Y����V��g�U7۵�{q���I����\��_�^hɶ�>l$�k����GG������_����gC�ڝ1�nr����aO	�lI���3?�m=���V@m�;%�/Ka��W�
v:��W���I�58�QW_�[������{8�e�6�I1~�������c����ދ�ԑ��E^j��p9G�Y�7��#��+]mRr��<�t@�m@�K'�k�,����U������O9p����M��6-�_
[����ChQ��|�f�_^m��3�4� �u���	sK"7Xu����̏p�'���r���fف�c��K^N=>���������r-��7��F�8e�_7�n�W8i��!��%Gd� ޑ��:�L�-ˁ� 6a�]\*J��/b#���Bn;�V�w��؞�R�k��B_<գԕ�<��POg�'�B�3ѷ��79���:�MH�dK*��(&%��7�Ȇ=�p>O��M���Z��t�Y�Q2��±p��� ��0��ٿ�c��̙��B��֤4I�
��39�*6)��L�����Z?:�҉��;���&����*]��,7q�[n)@���/�y2�3FI��}�2� �*���3���{�ICK×B�P��J�cnh�-�o:8�	G��������d��hE�(��(�8.�j�-6 �p=�S���|��-���;*t��d�A`t��2Õ;!v)��%S�o�\�6w�l���q���軛��8��O��0�xlխ���:4[���}OY)[g�A�A��X�A= '�~5����N�g�v�k&�A�N���lԦn{*0.�Zc�e1���.���FK�|g�|��������g.|�,�ڡIe�� ��#�D�vp�J/Y?���+U�l�H���?�{l����!�Eb���zȀ�n�9`S/�,�җT'�u��N�yCl��,f�,i�g�-e=gy�~g �`q��m�3>��L|1)~�Sԇr���l��;��-�ډ^��t^j���t�R�a��I�|��Aߘ�s�!�ļ�1����9@���㠉X�q���Z xsl/�=����?�ȷCя���F��goPҏ����?�W�
 ��#�kN.��t�^���K�k���ޭw�r9�؇��Nx����k�G�:a~�'���m���w��K��v��){�a�ru�7�иz�y�����	4	�Vv�9�$۷}�	�t����$ �O��ge��bH2iR&�}��dϲE/�O�X.�9�؅�ik���^q)�J��������"P�T�E �d��9�;/?���ų.Oɷ�Š��J�0y~�Ȥ�I�Py+�)#�m³h�M/s	�L�(��椎�/n�����B!��v�j��������O]��L�<�I�,A�I�N0P�����'�N���L��Ѹ�&�&�����tО<�,�	��cB����C�ˠP� �IY.bh��HE�Nq*����‚`�p�9��K�jي���ꀫ;�	d��A�ǲ[��$+n?jtA��|a����4��b
k�R���MZ�FL�4��67��m���ಓ�0� �t����e���우n����8�~VC��/3 �#��dߙ
�Db� �`���aY��/[B����^�뿢l�&ƙr�5wC�>~�p�|��5��y���{a)�f;Q���GK!���Y[��1���f��(Hc���5������O|�=����ҎH3{�����1ܠͶ<)�Ϫ;� S6P��>�҂E;ԁg�q6���lp	å��W����!�A3�z-δ��u��A�4$�����.��oB2S?�ɾ�E���k[k�V$��W��2>��4H�T�i��>�2:�.����(����em����i���2|�~��I|��A�5����m�˦��}|���;vMz���U.\���P=�U��CY�~�Y�bG�'ۘ��ޜ��gMf_2pf�7V�~�Ń�q��މë��f$�b�CG�#���NX1� S6,�b�/c"���b^i8�ȼ	>�-[�ͮW�\8�sa,��Ƕ�I\eq �D68S�W�6��I��WP��6ol,9cv'�=gVu�,*}�(]/m����0����R����J�Z]�c�,�� i�o�	�$��ϖa���)m��/h���vr��N=!3����N������C �ڀC<,k���� �d@(��i��^�E.�4%��N�L:@%�zA����Q�*B�h���Lҡ��t�dF4����	�)��ҹy�;�|k��f����V�:��w���R�����d���3:Qu��kg!�t��SÉ$>��#<}��;K�_��jc�VR��P[�g�4���-X�7!����gK�s)�ث�Y�7~�
#sJ��w��m,��x���$�vL�bg/��xg�\��E�OIQ�w��i�L'0���v[S�j�N�6�=,=D��%�/�T�u��\�T���gb^d�i˛~����[V]Ic�:7(��0`�#��j�3����W�~4��_�«� 8ğ|x���H����`7��L��S�:��؅�Cv�m�b5dk{�y�mM��A�x�5:�x�0#��x��b׎|�.������\\z�<���#�}�v��Çm]D�w�����nYA��8����ڥ�u@䑣�7�-�·ȥ mî�^_�u���bv�d��)��猃334��V�a`�9I�#���. 6o�U�u(�O�x�`h�틶�)���;vcf�rg����ue����*���h{�϶��S,|�T
�}l��C�gL���|�#Ã%|�/�:���M���`1~ޜ�yp�=Y� ��'�m�����>�|�K��.���c��Z�����se��o����N�5k����H=�W��|9��G�ڼ2���g����3p�K��y^H)i]�S��	����z_f�7�۬���7��o��]��!����N�`4��-��ߑSR����40��~�,���ƽ��`�� �z`{n��C�mt�W/�!��~��Ǿܪ�OJ�D�f���~��(�

����w�����\\I�H��
�7(����웽�F�V�����RN�Ȝ��K�7ٞ�sh�7߼�3��?��2�MTU�v$
.���e2�c8}ίY(�b�7��|Z�)1�S?��3u���ΩX��Sc*i�Kr&LJt������x�q䘸ס����m��ffpGS�D�![8��G�`�]t�2o�HW�k<>����̋t0:R��� �#F�����:
dC�鈩#g�<���٦,��:,Y�U"�V͘�,�zՄ8i�`�69KQ~�Wd\���r�%����\ѷ�Kw�K�>�:��deQ���'�d��җf;��S7�`G1�R�h�'sc�Z2'�)�Ǎ�IL��7es����@��P20� ߼�"�9�8PCg��>�����j̤bU����G��"7��%�_�����݋Y\���ul;t�A��Fs��c<r�ԅB]���|���1=?�^��>s`sn��V����D��{C�x�����:�)�H\ݨ���f���y@�� ��<W�C�	e��j�۹�i�XDSTKǥ�����-��)$]�o�ҷ�V��S����/\�5���co:��P�^�s�x#{��=ov���x����� @翾L��A3,�y���bFw.���P�l��b
�����3�*�g�DE?A^���E�NZ�� w9�_>?���~>�������������Q}��N_*m���52�6����o�æ4q�`DM����݌�d�Z9�R�.�@���?��a��82c�����aCNmK�A�'�>iMhܫ43`
��&��nH�g̦�O�|��k'e���,��A .è�%�"��Bb)c�Y����AފNq�Hґ��kkqŅ�qy'��<^;S��MP>�ێ��>D�gL=_=��Ɔ��䇥���#,�s�G�WYl�
<Wf��0�9w=���i�:���M�=)rZxd�<�tx��vG�lz��#�x;�{�:`}@�Y��4&f�Y>8�����]|�7@P�y�����+6�t������#:g����,j�GG�����8u�q�V/u�,K������/�I� ��@�K�=o��A�࢏��cUy�SvmH�WNgn�(��)�n�~�sn}����iZ�q83w�Y�A�x3X-�#h�6���؞��o��<�a��%4�����a(�8�ɓ'hIr��H[�	A�OxH���� !^y��Gy�\���Q��sfG[o<�eF�q9x��#%~Ë:��L�WhQƺ��6�_�pXGY#&������h�رz!OՕ\��xyJ�&����y��L�M�dL=�r�	&"�ʠ2*����֟mM#c��ҵ�N���S���E"��&�����CX�k��Aqv�'�%@�<ۏ!���kt.�I=�m�KC3AF�3k�F�x8��(;�P6ۤ�R�C~��)��S���c�
��h��\���W�$.#����~���lZ����L��$�"��[�΂������CC0"s�"JNӑ���t,����(7ٌ��2�W����ؒ6����~���6�_�W��X����E�L�ܼu����_~�����O�p�p�l�+���P���K~����Ѭ��7$�+��PO�.:2�e����Y�^�M�M�$�o�w r=B� �2���H��KFδ�7?��.�����|� ɹ���_�u�
�ۥ���tua&m)�bRT�::�:�����#�.׋��S|K3]xC�Z3I9���;�B ����ɳ,g���6�{[ ���E�D��fu�8`7X ��ͳ���O���x���� �.�;7�G����[��\릴6 }]�������W�V�3GM[�s�Z ��L[�iӹN���<������妎�Ƭԕ*��]7a���;@?`��t��7�:���8��YY�P�I�؏�>�E~����������%٢�2�$�ɕˆ9�Jcv���ͧ8d>2�?:��	J�c�Y�v)��%M��K��A�O�?e44�����2�����~�+�m�@��M���d�n`�Յ�b��q��������̓D˺S�j�,�.�
N�`���n�g���A�:D���s�s��8�jI���'Ù�:��Ua�����VL{&]>�1��Rf6�O����w�;P_BJ���S�&�_�B��~t����W�������'������ɡ�j>2��=���,%C�	c��s��)%�l���=I�)��33��*>�r�}�%�� K��ף�ԑyV����\��n �`Be���;7^�o�sh6!4l��`˳�Zo���ؕ�`��Db\ǁS?�
�g��K��Tedi���#i0צ������Ζe@wً��"���F�D�E��)�E��o�-�����l:�wz��L���+�xs�٣���?���]�#͖~R�۷W>�o<�����������/|,�Gݶ'e�E9��L���V�z��^��L9��ə+���Na�[����JY��Ӎ����Riٳ��d�~�� �(h$��9Օi�oҸ^dNl8H���"�B��R��U�!�2r�'W�Q�"FJ�I67q��%Q&�a\{b��OS-HG,e���T}�vz�u6z�O�ΞsW�������ͩ�x�����m�P�z���d�r͎�q`C��ކ����4�����H���\tY}�ӽ�������MSV.r��	o�!x��B���U���xY�nU8 ݼ�: 71d��ǂ�ܺv��'���}���s�0 �`�k��w���:��pϞ������F�ɧ���ֳ�e}ˈ����.6��?yn`�M�bGrl�N��y��������n��<��ڈҐ(��->���}�`h����"��d _�<ʵs3]����]NI6����`�&g���q�㺬�ȥ��un��e�~H���c��6̶��z��\Ϛ��+}�0�6����:�I/3�y>ϲ�������L���v��=Ǽ�!��h�؅�����"]��kSOxp���,�8�`��Ƶ�Y��r�dX�������8 7��s�δ��T�m^��Ȯ<��	7���NҚ��m4n��Χۗ���O��.4��˭z�9q�{���^^@�������U�[�ʢ#f����X�hfܮ����)p�3zQa� (�ۂ�j�꨺�V����<����/��r ��ҭ9�]:io��ggˮ�G��5u�p��b=�~gh�
��b��oM>c�i]�kL�6���&���ԃ2T��kje�.K7���]�����N\\�ؔ���l?^6�}vdkJ~8P���,��v���3�gO1q�:�#߰����g�?���������ɏ[���x^'��6D�>:�67`K)�k�X������F�^�W�㠎�s�G�\U��8.s�N�lR�(�`V�Mk��0��hzq��&�����q�5��� o_�a�71"R&��6{Ӭ��� f�E��P���Kz`V|2|�/�3�r�w��$m3��f���s7KcC(�Γ�8�v�v���J�K�t�������8��Ι��(1y�6�*z��vh�˸��0 ��4����G���QEqZiBj�r1�Va�\�W���"��{L���U1V�3��5v�X*w�:d�8q=a����e��q �	;=.�:^tHG���=���_� �8�ΕyK/al�,/�jx�e2׫�	tʯ�%��S]��G)��@��a����U[�ƕ���g8�>�2^;��<�t�����e1�&�sJ@i*ƒ�H�M�^�ҖhY��k�I��:��� �۟��XgE䜭t�֑.~�V�2���>B�6��G]؆��ѻ3��k#փ׶E呾(�.��<�^�`�-^���+|�Iy��7�Oe  @ IDATKH��O��=�MZƁ���u0��-	�tA�5���_s�lx�m:npq�˂V��s6�#Ŗ_[}�8q˫ϩ7�����_"+n���^���+ޘ��@���z���z��Z���=�K':��� ���la��r+?l-��!σ#mEFV�vbq�݈��#y`��`e,m��[&��כ�o����m��<���ZZ�!)�vHy�l���^�t������n'���"��Y#e�բi���^TEo!�D�c.���!N��� �%2�V�+�ӊp�Z��'m��M��l�ΗjV�f?��%Kt�Q�%���G�.yκ��l�q��s�M_�0��4���D!C}-�v�#�Z[����<7M������I�@�T�V����`1u�A9לc����zT�)z$���Q�i���Wq��zIm�x���N�Џ^�$A��Rs��ĔN���+0gIF8�Ij�#��"'�Yڞ!���{JKǴ�Pǥl��*��?�&��g'b䴜��q��S���<>���3�}x��	`Z��]�qGͷ��&�0�XB�:�`�M������������_x�����W	�6T�u���7���Պ�S��,��t<ʻ�	i�;�IZ�\��W>ۧS�qꄹ��t]+28���m,��Ou$�/���>wJ_��{����W�����������������"o����B�^|J��Gf����9�|��qބt�;o�:=��R�VG�����|�t8;��<���V����������[��khM�^=(/i:LFv�ڂ�
@��*�b����ё>|���=;[������-i;����3Ŭ�)��)A�:;�Km�}�[S؆6�D"=�x���MN⬳ g���m �fw�:���3i�זT0��_ꛙ.w�w_��ˁ�MM��Vo.tƲ9��]���@�y�>n�3��P�I�7�Օ��?����Y��絭u�_x�Yp��o��_u.M��I�5b������/]�q*y�eFl���ۤ�(���K���:�@�9Rq��L8��l/���>C<��Fз���3�R\��&x�
q"��M�^̯;�6z(�֍3���S������ 4�>����_m�҉�Qg��DG�8<,z�D�g]��-m N�W�h(O��x��ԣ��O��N�e�C��k����1����!���-/��(���I�F��ͪ�qX'8گ�K�2�A\;3d�Jǘ�ޥ2��?��ҧ�_	Çk�r��9:e�5��U��좑��2�A��I��[�Fw��ң����U��J�<G��_@q�]Y������́wz��o�rx��7�W�6�%9?*ܜ�`aS�)$�SZ<-�7�`�m�dv^b��R� ���
����H	ҁ�N e����g�;^��gi���Q�H+.�%����:�e�-�ܓ�Ev y�x�pa�Ȼ��0��
����#�gv$SO���Z`���M2�9�s��}�wAu�(�u�����%uLtR.�"GZb;v׀��?�#�	>5���%0�FC϶�ڦ��_�Wiʒ�NK�l}K��������t��Y���ɓ�0�����R5Ц��[Ɉat5���^~jai�3�Wa3�&���O29x���1����9�B��"V+�J�8I�u�%|����z2=w�8�q28��D���ȑ4P;#�3*v0��������#N�t�_�k+�2�A0rxm~����ЁM'�lp���c���`��,�i�F�s�b������ ��Sl�N\i^�!�ͩ	x�^�Mn0t�����7���\6 ��(_m�#�����t��uq��M7p�@��G�gڿil~I��/:֏Υ�l��E���u)Q�8t��3.a��r.��N��O�=�V���}�]�3N��r�֟~���ipHK�t����)Q�I����9.�ީ��M=��B�3j�m�߹i��r�����������gO��Q�}DE����:9�[���EQ�L���!3���3�9x��<��WҶ]sK(p�ك:+���^
�;�ltC1�^�3'-Cx%-�s�6vL42؞�;�2Ox�z����-^\�1�Kĵ�����x���1�H��+�Ll��;6=�Z���ʣ#�����k~���)�`��?�I�e���g�/%T��z�G��va]DLsl/m�B��/Qt���d�Ʊ�N_�U~ㄈYa8��o	#A=&\��M�r�h���\b��6�p������>:$<#�P��:�g̺<}Ƴl��_���Ѭ�����|Ϟ�I��v�K�Ȳ�ǝ����Vx��;|����+��K^/�b�Мs؋o�)�%P eHPf�
gH�8�-7�&�W�|��8](}����3:��w��͎�N���N�خ��Y�Iځ�E��fG���髯��+>o�5��,e�6uAߝF�A W�|��������3�'��f p�2����h�e�p�Q8@<|���q��58k�@����?2�?>�Wr�R�ʑ��{�4/��A�I�Ǵ5ڨ3j�vʣV�t8~��'f}�T��K7iu�꺖l|K�5����
�_R:(ʣy�*��A�A��r?~�8����}�n>�.���f�|�n�g����L^���R�<��>�P���I������=���:b[֑�층�8� G�d�pD�ri�LxFW�϶w�|�8�IS&٫G?�H98e���U�΁?�����h��ufT�p��ҙ�?�@�յ���uQ�u�t:�Ǵ�i��P�׏o���v^Zxg�Q�.|~��{�g�����>�C�$��i�Ge�>u0�N�vM�m�����<�PX����|�M�'ߙ'm9����f���yS�����e8^ڠv���Gan�&}�H�mX�8>n�X^���+xpv]y�'1�&���k�t�eՏfA����shi��8��ڐd��Ԡ'C�όy���m(����Pʐ�s�0��V ^���{qm���a;TJ]��d⸜qeg(4���/�C�~���.�<^CW��TK��[��û�><���Ǉ�|�֧�g���o{���	����򥍶�"i�uZvxaH�9U��©3���n���i���C�1���Sٓ�}�&��z����h�� J\>{��˜�QZ����E)��)Q�b����B�T�f�O;:_K@΂�t�))�+��rp칀�n��LD Ӌ/�a
(R�����?jW��R�I��x��]Rlh`�\_Ҡ��,F��0�gl$���H�Q^CHc����0���)�\B����G+{ׇ�Bֳ-�}��§�X�̽�S�C�?^�)7�*�������ttg~�㌎�d� [�t���*�#�z.6,ꂼ8k�k��p|4�w޻������D���^8�Y���a:��S6t;�'���ٲ�u:?��L�w�>Z{��a`=��)�G�ʠsؙ��@�o�e�J'$�C�����Ϫ�ʯ������_�5Y���t��k��R���(��P^�����[��a=� ݳ�8p�<f6�	3u :h}��'|����|P1�$��TWq�ѣ<YWʖoÑ�#iu�� F���G�D��~���K:����άWʋ�e�;a���?GIiPf�<b�Д�)�/u�@��dp��;i�5�Gu��Y\�mKzg?N�e�w�R���	4�Sg����L{v+�3fUK�Θ~	��֣���Ξu;�~uP]ȗ����L���m8��bsevS�kמq��V��� lCeEK��f.������c������d�f�>��?��UW:�����_o���_�EEˏ|*�Ε2(��m�nH�9�|݌S&��@X֙@kHGT�@�q��wXGj���?��L�6(`�q�ӎ;���]Rβ:�:�XEu&qB��$-y:[X���But53:�}/]WA�:X���t�ϯ�j?�A�m�`M��`�4[���>�!�qPgB*�m�o@����e���|�Kl8�q���{�f��9��3�Ln��ީ_}*o�˃�Y
mס�z]�Zec�h�ò]r$c)<
;u#ދ�2I�7@^YX�GaGP^W���缲3c��NHx��#}��!��8N��6m?Ѷmy6m� �MO}����:f�S����~�<���G�F#��F�Lʜ��iK��\�$Pű�.&ӎ���u���1��E8�;l��!e����؛��g��}��)����n���od��G̀�P��*Z��/i)ĥpl��W8H�rz�1]�͆Jx�{�c�:b\��6ڲ�AI�oG,��~�lZ��9ʁe�]����<^������U�V;��`݂с��W)�����A�x�*¶#��ӟ�g���޽���ϞqgN9�4J��ѻP\�汘@'��&�	{G�]�5ζ�:$��la���@��Hӌ�1��;:�릿��h��%p�H��N߁M'n������{�+N��"��<|��?��� <�A������V��fЗO۱�Ԗԗ���̀a�g�L��.v�y��7�����?�����~��@ԏ�N�Lי���:z��}m��̀A���u� �/|g	�[�B;�g���\G�N��q�ԣ�U�C��m��R���R x�{i/'=8��!��ĩ3(�::S�:Vu|+�ft���8�2�p��Hǻ]�G8\_1��5N�31�EzB?��3+������[β2����<�T�^c�f�U?��5[~P{��8_�H��Rq��u��l��ڴ�T���اN��9��)/�"���>�4ۙ��G�>ű��=�	�]����(a�Oi�8���8h�W�8GN,,g�i��4��%�����}v�,��o ��f0=I��=G/v����%�Z-)�����/�撒���)�&\FDFfem��hvt� �~F{m���"���A:��(fz��m���Foj���3Ffx'S?#��� ���O��v�:��i9o3��)C3�E�eYN\��뤭��l)�B���#��_}r2�s��g�{0X�����X��z�QǏ��v*�C)��/��x%ou�����w?:�[��v�+�����y��&�������{����nt�P-ݗ��[�.ȣ��<pt{񾂦}����b@^���_��o�_؎�̧�9��?՜κP=��?���ʛ]y[���ۢ}9-g����g0���2Q"�a�t�ņ�ʭ�c_��pX��
�`;���[?9�L~��+F=�$p��̠I�iL"5K�M2�'�<+�2J�h�9�p"]ϛ�)�&�_K�]��L�}�'�c���~�G,�*|�C�`;��Q��l���x��D{��2��1t�EhˊS"����m��g��<�y��sJs��ޜ��r\��Oחu)P�G�s\��� ����FN���ͥ���j��R�7�.�]R�ZR�*��U�L���{�U��ʗ��M�'B�rs��sF(?+�����u{����F��,|�
�:Q���+R0�'���Y9tR��|�����w8O��>ʷ2�`9�w����'��d��OM�&��mxc��p2�D��N������mc�NF~���D������d���^?|X9og�w�}ג-��<��R��L4�\�6WO)xQ��:�L���p�m����d���>c"ޑ���S��'��=�B�]g�l�rF&�<�=��5��7�wp�h#3�7���-���²�=Ï�>����/�����ar2ϩ ?z�@��w�o>���Aw��a����`=6���\�&�[�:�,�,��W&<f���������6�i2����6\{�խ#4���LO�	\i�&�r��9��1��QZm�>p��q���Κs2��=T���V�p�v1�Y���ڼ����v��9�C���9��|tpOF��g�m�����M;�&_���e�^8�������Hg�)/�:���<[\�v��~�IxY����� �9��9�t��)�>?]8�	b�oZ��6"D��H5�G��v�VC������*��n`w9��l�Ǟr�J�r�-
l�ODɵ�{S��Ũ�-�Gn��O��y�$����)�������%�'呞Ͱ�;/�gB��$��L�Û��[�������E�$6��l;��)Y]m-U�!é�����=��6�V!�;{2�O�έ�ȿ���J��x�3���<��e�FlJ����%'[z7�빡�y0�6wo�'()�v%O}}�JYB�h�5��]�l"f�q<��Pqd�I�{5u{��^��ͳq1S8wS�m˘�9����\��L���ѐ���a��\�I��nJp��\��P���գG�__��[��c��n��˼����*SuOyҔ�ף���JC	s���j�3Qo�ޮ,����--8F��"Cx�}�	�+Ļq���t",��������;x���1��A3T}�2-�� �s�Z�LDa".kp���"5������k���0�;�#�;�!���	|SPp��gC��/ؤ�{6����}e�6�����>�]Q/N�톻uF��"�|����n������J$�s+jԭ)�B>Ng`����ʕl�Jv��8� ����Z��GM�\��S�u��3����&���Ýn��g��$괃Ky�1 �0�ǽ q5G����'�d��G�|=��h&�n�x9r8�0A`(�W��C�a�=tQg�6�����s�ށ~db�/󧆷��xȥ��ku�在MeL;��"`��3�8֜-��8i��z�c���Qv�|�jqޡV�L�2t�5�.������mc�10/ܞ��~u�Et�m�C���Y�LzU�hd+����	ǫ��>��Ƌ8Nt��a�$�t��<�,h�E�*�u_���D�k��:d����J�orV�j^ys��E��'�Q���]��h�t �� v*[Y�e-K��m�������S�9�*s_uD������yr�>}Hwb��q�����柾�S.���<��ih������޾��]�c�8ŵ�Y=(�4����>�XR��n;�΃���������|���rʹ��S�캫�ɲ�Mn^���{Zw����9���oj_��b-�L�q�EH�	�kDLYY���C
<�S# H�	�a�K��>�DeM�w�*{���06�����ฉ�
a�Qc<��|�P��L��'���t@��P_N�(����qע� ,�(z����t+�m���ӵB<������LJ�J�e����^w��q����[�^e+N��4D��ئ̄_��Ba��@�ݬ�>J������N��pJ��޽��^3]�ۇ�v�.��J?�2���$���;��7���\!̽CY`f �Ygo눃���'>2�� YCwy@�z"�]��iu2���艷)_y�eX���s/�FV*#H�Y����~�����)se��3�KAh�RL@��08W�D�u`*h6t��s���{ �2�Lz,���|o��ۄj�/,�h*�÷ Չh"-�]����޼�!cpr��y;mi�IІW��Ņ�V����@U��+b����1s��Iˊ�9c�.�Zc����Wy�av�Á�,�c\)�M�u����G԰�O 1��#)���Aq/�]�,!��30ڻ+�����!;� 6�<�z:*dryʹ��C�x��:VF�z��{�7t���Y��î�'��e����Kt��wW�|��:��U�8'�h�9���I��+]�)��F9�����W�6Hn�Q݆`�e֤:�74�ިƔ���2W�S���o0�W��&� MVNWւrҩ�<Ss]��������0N��}�y�������I��l{G��'`���M�Ϊn�K���%����͍��-l�m�)�j����p��~��Ndo�ؔQh��O8W��yJo�yS-�#_�"�#<z�=zC%�dƮm�g�qy��9r���S���M3�/�{������#��NSnmcҡ��N@��}���*\������D��q�u�,��-v����w��x�����<��Ϳy�8�ӛeo�AR�|?x��Y�S ��vv���x]�I��v^)�YO�"e�w�׸�K���2��j���NgE�0��!y\�W��-
-��Ex�!����Ԙ4�u4ի�`�p����)���� ��%���`���2�d��5�� ��y��Pfs�iW���.'ϡ�?��R��3&Ӏ��=6ʁ�ĕ�s �~�ݾf�?L��3$p3<P�����{�C�p����Q�e���*^m�|��y�*�9h�P�#ogu	��.h��yP/3p?�6������$yJ7xE���,(�z47����p)W4H��zg"�3�	o�0�&/�Q�h��
��J0��۲�e�7�D���C�����j��P�>p����2���q��x���)ˎ��1�~(|������\�0�����9W����xU7gTڇ��y����!G.[��I�������0�����E"��A��ʌ�LsD���s�3���	�#�H���ۡ�}�r���r8�_~��ٽ�F�2����r��@�"����޸yT𦗔�9����ȿE%u��K��C�$�����<�CYd�~o�I�PkoNN����[�����Y�w�����L��D�f�TV��V6�q8��fC�)��Ks C��6�l+/+Wh2��t��q�Or���&���Kq(��u�+�U��h�s�4�9�O4��G�ϣ�F��Ng���6�)=�&C�jI�Lw�(m��C��V^�I�2P��Qg�G���rk���җ������M��Ћ�=h(ג[z�� ^_��'}0�V�ib0eL��]~:�j��6���������7ڿ?4qow�R~mڿ2��z�t?z��[�d�������u��!���-{��%��>���*�#���rXhG��o=���m�ՠ]��ÿ!��9:�/��*y�F�iڒ��?&J��I�l'��.Z�p�u}+���~6�v�����-}[{���lcb��������+UP��\tbǔ/"a�V)���'Q���2#�!!�dу���H\x\�g
b���>%�q�߇��(�m���xR�<ʷ��g���k��cY}����)_��JY}~�l��4�'��I��UcW��x0���̈́�
��a�8ty�<�_l=fn�C8��vB|��IQK�K����ʳ_n��6Gt���T��'M��hM@����I��l|�M
����Go��&b=��/�q�����}�kp׌��XG��g/�TJ���ޓ��}��z�x���'���}Jv��`�)X
��%J�`��y�AГ� -�+zb��|*)�����Ѓ�rE��[83�b�����|Cw��7Q=|u�����И���j�jh?xu4�f�F�.ۏ�9�$Ouv���Wẃ��q-�m�s|����f��$pN�1��ҡ=tNg��Exą��7V�+R�Qo��m��}y���0L;O�2�臏��p�{Z����菣}����ѫv�{�/9>7�k
=x02����|eAǆO"�/?�y��`�*�|��P���!��Zq6�r��Pܾ\P���;'�W]qd�m��h@�(~�?~!�����P�#M�cp����f4A���C��+g��� ��	Ku+�����.�:#ڈz[��j"�,
�>彗9��svxW�D���<�59�pG6����L��%Jf�q��i�lea��S�:����6d�:�)�ȧ=�?��!i����(0���?�ަ���-��x�'��Շ�ô#�Z�u�<Sd%��y�ew�����e2�sѯ�:�rʺz�\t��Ώ��|���~�������s������%ޓ){@��?@Z��#�Sf6{�oY.��s\'k��N�`���]�/��e��,t;Աv7σil�{48l����F��q��8�m�3�%�W'˰tM4��Ar5�;2$W�r]���^5�h�R��"a�����ɯ6)_�hv��a��8�Yt����_7Q}ވL������֗��G��l:�D� �>���qv
�ƏQ�LV��<>'rD�(d�>uy<J�@&�ܜ�� �R�qQ���:轰�ߊ�ӻ�x��O��_}�i�]g�A�$8d�.mW��)��\Ob>�AQ��N�=��b�Id�hy.��S�<a�J�~��.���� $��qS�bf?U����d��,C`�o�9?ǇǤN��V0��D$�"~��^}�*����0֚z�ZI�͗��z�.�$��n����5�􆍋���M*{nQ�����{=yܼ��H���� ](�M���>�bP� k�l����p��f�+���%�p9s��rr{�I��s�Z]��3;8Ѐ��?Y�.p��Bw.9�(w�d|7��8`�ȩcxV^΂ȃ#��}�^>�yx;�ɰ�C�>��:W>�6�`�P�1�W�9P��2�����d� ǲ,���>�e�4	�P��sB�=�������
<�׮�q����b�:�qN��O�7r��5�?[G��06�m{��Q���C�Uڡ3�����V���yz�=7?�F���Jx��3�<�-fY�H����Ï�>z0N)�R������qhԻ��&�d�.�ǉ#C6�Ï��2¼ >�)_Y��f��螣�9\<���<�������|���h�`�(eyLR�|x�����s�A���Ǫ���+��藼(�N�u8�iW'�� �e�~�&jR����0��W���T|�9b���n�ڂ]������s��}!Eg���4Q�r������� 8��r_=��۶,��N�2>ܨ|d:�r<�[.N4��͓�yW6w��b.3����:�K��?��t�Q{�uFֶx�_���&Zz	�����F�0��G�L~��q�|p��X�J����O���O�ZK��])�6.��ֽ��O%v�u�;��'�K�
 |go9�GFK1_�,A��~lKz�쀚d�h9� �izV���eao��w}��j�I�$��^O��_m�A��o:�zc�4�j��%b4d��E=�[�)E�&�z�o�>&U�4.@�H{`���3	�U��W�GAx����;6�4?9Dذ���8$x����12�0WLt��]���T�cyq��6`"��m8s/�Ml�=���u���I�<�B3�(z�H�'��:���3�繚�p�=��6������GE���ޗ������u�}�k0c�S��烲��àS��0������u(�%#��,��`���Q搘�!�l,�ZK|Xպ\�'��_�[�w�#G�3�9�/s��p����cu<`?�7B�F9���ax�������a'�p�^���e2k���3�1dw�B]�@"'�n�<o�Dv�%-?ů�:Q�� ��G��Q�F�����E��Mɩm/�8-�w�g��y4�F�a�Z?��E��1��vԵq�����5k��=��k��6�	��ce;���qU?�Aٳy��yiֹL.N�M���5������V������៞)k&�:�N��b��yy$�df���(!l%�IW��h��Y�l�S>�O��9ǆ�M���_���FVї�ٖ������򹴜���.���z��9_�ݵ}�
G�pz�q��Kx�7yT�-\K�u�+��;���:|��]���8��N<��+�Q[�V�胡+��|�]���6��Z�)c����J��l��j�����d�G=��s�]m'���2B��/��KD�vKܻ{{�fa�_��)d��0���"������$m���K���I�,��cCͥ��N�vXn�D�f�zoz��}2���Q�>�t?-~Xw*N����ɁL�\OP@ڞozݹ��l1|��v��)˴K��|5y"K����t����pq�D��4�^��q�r�+�0�!����r�z������;�  ����Q��{�[���b"�Ic�C!��h��u�=;�Cm�g>�7��ܵ���[�&� ���7º��H�*�_/s9�oH�"RJ�xC��U賔~�<Oi��F
�F�#�
��^$��C�٫<:�3ys��t�n��Pw�7Ŝ�= h���>߾2~�
���Y�G�Ƽ�x��"*��ޖ�J�h���L+�X�uM�~���1Qgp7h^�)���h��l~�`T�)oO&�e�贡������������x��Q��Y_�yea���.���M�	'O����aJ��}�{je_1uV�{���6$��!»7[?��7�r�i=�IC�?&G�`��&,��bk��P2d(}�8.&�Ǹ��Vÿ_d&Z����}����9<����f|�e��p�=��B��\���U�)�W=~�������	��oÙ�l/�1��:A&�2z"C"!�΋�yp5�u���d��`�o�E���V�o��&}.�����p2�r+Z�j/�3�`���h:/��h�%��T�)��}q���(�)Z��A ��ge��1����Ũ�uJt�N��u4�v�-��a4Y�������-�2{�=��%)�wEW9����hZ8�g�R��'c�q� �$�E|G����B�"~d���Yю�Gr�>���P�.��ݔ���|�DR_�i(^���N�􌬨�'��L�C-�y�I��G)���=�E����hk��ޙr�>=����q�[�n�G�s�u���R5�E�'ꘗj��wm�X1z}�[y�����D�7�ܡ)��o��ڔ��Ik�:{��v��)Q�[M#0��b�ى��ʡ�oyQ�ց��hM��ء������%�k��lD�m#��m�:hbj�bj�l������ӟs�t�n�#z����!�D����>�4y�����1���?|�\�sz�FY�
^���$�� @��_;#���n��lI����[e�<���'�o��e(�m�>n��ۍ��g�Y�����ҋx�Ͷ���4�a>.>j�����:`�	�=�r�����6���u�vPVd(��XVv8`�)�j:��<�#�ZPa���Q��7�fnqC�/_�;ܼ�p��Y����6Gc�ׯ>��b�SQg7���o�9�5���U��晞8�Ps�Bg!�FĜeXy���0H��Ӊu�._�Ŝ�@ϡֹ�{��h�`GP�H�r��/Q����fu*�=��m
���c��I��˫�D�E�͋�`��U�:D]�����6��?J�8~������8���.��%��p��pN���ֻ�M�Z�dv*��$���t��.��w�j���	��;}:$����Wg�[��W,�+?/�kHw�3fE�.��-�{~#':g(0�����nM�����`������;�U?��X���:Q,��V�qn��F!F{�u���4�g�0*��q��Á/�2�xC^i�;}�C�o�Cfʂ���w�y���L�&�Qd��f��9�O}����~���Hcr��B�A�Ƨh�t��[c
�d��FK�5�C��s�h?�����t�%<�ˋ��˹Q�:Jǐx�g��q����� U�D�)����s&"`g!M����5�˸��7�ՁLNԳ�<�|��#<�H�LG[�P��2�!�����g�F�"Rp��K<NGN98p��с�.C�Ƀ�O��r8_+�Y�xB��&�{;�o\���x�i��b��v�=������5�9s�DWC��I����4y~��V`�h��J�����δ�ڃv���Ĉi��~�{�k���:_�/m�ypv=x�f�Ʉg�كaҜ��6�=s�Oх�"���- ����FH�Ó���#[�v���#�`���������#|Js:tq�97�D{t��l���t�܂�H��t;��5.~h��������/n$.���&9B�m'#��B���z]`�u����`�M5�V�Ew�=Y�a��+9k���]�4�*8�p��w���)�������N@Y����Љ.sl���@ҕ�L��{�Ϸ�O!�u���P�k�c���e�YM�9Y9b��_�ݺN���"�n���-�� ȳ�-��2h�U�{}� p�jOڹ�z��Ę�Lр��-C��������)��2z:o��R^�ۺ#Zмє�g��d�s^����l���*b��z�"��O�lb5g,<>3��
�9`���Qi�����tv�p-���x@�c�X��ܵ�����nҾO���q�G����sBs�8��A��Z�S�O����i��9F�C����R��g][C�i��R��s*�_����ݩ�xc��g��(�W9f�_���&�?M������r��S��1�dً�����1|Rj��/���r-�BK�Q�u�6���折ph�4wG���qnX�a��\�:'��۹<��3Fֈ�v�m�[h����%_�W޼�9i�N�<;Y��^pp���X�E��7��uLk�v8��3�ql��9�9�)Y��9�|�Z�Y�̺Ϙe+o΃	�=?�c�N�1�qN���(>h�`H�f�+V�EA3u�sv���պ1���S&��=��_����1�2+��c,�7���s8]�y������.�A���9d�3�l�O/i�������;.��I�?UЦ�q�å��$=��2�(��*zzF�Я�9�`��{��F�~�Ӈ���s�JcV���1�i;Y�cz�����Zt�o���Жn�&ڵ�Ec�H����w��������c�g�\�=�����|d*�楌��|��휨�iy�m�ո�q
}&��IX��z؍:{�:�r�$}�������Y�R�N�%�㵶#�	(�E����"��Vﴖ�^�ww�?��r�=�����t�.���l�����b��n�s�S�@գy�g���'l��[��`�\�=<����[r��9�?���Yit�ޞݿ�����.*�0]�$!�k#t�K�NN�͢Lw�3�O:��?�Wϴ���9�=�<�l��Ej��n����8��i�C�噴v���(��N��$C��ȗ���Y.�e�r"9��z	���^R�By9`74��P�v�(�ʾ6� ��Y#�@��i�[�F�sVXVQQd6>zR�'��gz�]?O�'��9����	��#������B"v�!`�b��&��ޕ�y�Hf>����v�<�'<�]��XN��9L��}�l���+w�7I繟a���UC�j��u�I��?�+�(�89�"\�&(x���2���#��aQ��?����oI?}*�HG��PSL7n��`�6%-\�p��u�fo��z���B�9'�VU��5,�X�/?�?�a+�؜ ����_�S��⍆�^�[
b3�'��Ə�R5���ɹ�ξ���r�s�4�CbN�O� |��+�3�S���nh��fX�DQ����%����S�=���$({zG��
Wa�M�qt (uF]7�Ӽ�g�i�r�Gy7K4{p���FGǄ���D�z6Cik�]��#��c���w?�}������m+�������8*w����B�!���h{�o�P~���2������z;��K����׵��pi/��?�ē�3T\��r�_��h#C�tr(��I���}��S��?���w�3���5N�DU5F��[p�0 �J�8u�,�P�T��![�m�;����s�:R�'���F쒍�{>ϯE[Ώ�f�5s���.U����q��C�`VwP�5�k�>��FL{�1�{�
8���1ȼ�!�
���8IJ�,��_S��`�R;�ސ�;���'/~|�ݷ����}�hUY�um��}�15
d���ކTشAskƚ��w5��q��cs�*y��� z+[�ﶣ�=~X���);t�>4���a�]�3�M�O�~8���$>�9�/�V��65��>����F2#�����iLd�	Ll
5�6s�))����PY���Z����m$Y�Ar��Ұ۶���t��m�S�(��M;H��d	�Ny�w#�����f��&W�Xx�c/�5���~ε!�"��;����<&�%}E����;>�Yf#l�P�o��[�E�0���ח�7��|���8�<CX���iT�Q]ڙ��)�`l���6S�33Ɵ8&?���V�s�P������u�+;��嵉��]��W~��U�՜�����  @ IDAT��Nl��S�A�z8�B������Rα/^��+�C���sG���֐�ǽ=4�>%��r	��-�ǥ?	�<��|���'���:Gı���S���{�ƕ�s���%^��������D4sw|z�~�=jk)Q�o5\�~5|k|<�w� ޾}�t�6zѵ�{�n��uѣ�gNKÂ��6���L�7"���K�u�c�q"S�׻7x�?�W���(�բ #ot�v���2��Eo�p(g����Y�N���+G���m�*���@���z�M�Ws�D�,|�n��{���w�s�z�c���F����([/y�}J
#��8c)O8Ý=��^E ���s��G9ʭ��.-���:�F֪���K�gm�����h!SC9���u
�#C�Q�S��l�f�M�8� ʃGV�甾�Ō�.R�G�<v�N��ǝtO�&�,>�MoH��a�i/�f�Cϧ��R��grUzUЧl�"'$��X�	���8/��h�7怽(�l!S�'������r�b���"�z���Q�ᄑOt�7Ä��u�)-��cH��c$ċ�ꞁ���䏳��!�=,� �U��<h3��G.ё3Ɖ��壥ǁL>�9��]��L�Q�Q�k��彙a�������ϝE'��f���ž݉N����_$�����=�[����FE��]-[��%A#Wp��[���6wO�C�9g��Ǔ��e�����8|*���qN��~���pL�Iw�xr*a"�� ��������&>�N+������z��D�p�mO��xM{nakÐ�9dVf�����5?����'}w՜���5���>�����Ë�g<�d��q���A2b׎�{�����o*��<ӯ,&��75}�P�<�+�%�l�E6�ν��g����t����a��U�����sB(�T��w5�z����o7�'�y�ׯ�N�4tԫ�z���#4<J�*�0R)��T��<��]kP��8�qy����{ރ-{�(0���+O9�>_rSL����6�"T�;dcZ�6Gћ�:�n��_�Nn$�ބ t[�9��N1
���K�4*�Ώ*d��T}Y�$b��;��S�[��M�����8������ˬr����Z9����L���j��k���s7���j��g�aB==���խ.*��1:)G�eDE�n5�}=���Wz�6��ys�!��j0�2�<�Eq���1Ǡ���S��ٕ��d�E��|NIR�S�hSȃ�Ը?�z�Ѕ�W�J+b��~�߽����	��A8��Y�Ac,����oNFV]�%r5�P�&��%#d�2���T���c��9d�l�AVC��:%����N�=m�mtQ� �d��#5茾�~�}���2	��h��kD�1V�*;�6��0_��lGHp.C�~�8��u���R׮��(ی"�u�O���K&�;Q��h�J,�Y8���X"E
�e;��ܳ��t�� ��ÊL��<�]bc�eZ��>��=�:l�\���C�Y�I���,�"��~KgK��#��y���u��L�h9�1�5����пg�uD��a`ڍ�NٖtC���.����Mrv�r�"����u���G�B���`�ۮ7ixU���-��]J��d�0G)�M�>�P4�q�_�nsS�&�x9�7�2C�t�a��E�p��o2���ZtGZ0>$/�k:!'Y���߶+�!�i���>8Y��}������}(��Ϗ?��/? �֝O27W���ͥ$�wt\dX����N�=/,^v\��c��%_��׈Ń�s����?j1�O?~8Nף^f���C�H+�H�q��8�5����@%���o'�Cz���!���l=��oo-�?m���&ғ?����c�Y��޾�`��O�~=��i���KW�J����/��5��������a޼��>.C��m_�M����X;��U|���z��)RX�ۄN�l{K����4.�<�ʤ�V��{Y�)�(��E���K��u��?~w��^bs��䐉�\��T� �k�l��O�p�QhW���I�T���%[��ݷ/΃��4�=�z���Y	6o�`"o��e9_�;EJ|ڎ4.	�e��(=4�ri �ˋ����3^}�=�{�oP�jރ|B�aW��jg$�@o$���L�]C@�}��E�B=n1�]i��j4�)b��o���B���9�M��1qX62�k���E<	<y"��D���Ãw� �S�w�~�2�:y�A���Ǿ��0<�n��Wg?��2��k�W�7���"v��=��k�E���~O
nhJѿnAc��ɨ�(0�8h�,�T�-:��d�ܡ����99{p"�]Q9��1��U*�3���=�.J�=On�W�4��nN��[��W�p~}�m�+`��6bg��n��8���}��i�����Fn��ݝz����<pAC�)g����{9��i+��8ݫ@�t�+��u2�h�v�:�;a�߶�>ޠ�]��t��ϟ���F�N��4z�ͽYI�^���`�i�E�o����%?8�>�3�u�L,b4��/O?��F���n�I��&m|�S�a��[�HT���>�|K���u�.��K�f�e2��E�`<�otI;m�Nz����Dέ�-G<lj3��dG0>���,m1��y��Em�z���.�z޲��MG{ܬ��Q�OϿ|�ض�Z��y���z0�*��r���F�~#"��E�`淉�q�gfu1���]���땇�� 8ҕ�6��&D����y�5�bf]9[y�n�'����'��vJ:G�D{7I��ӽ?;��?{�Y����E��I����z�M��q�>���n���限���E��'^��^�p5��ș�՞Y��]���|�h��G�n���_������>���"^�;u���R3t[
���t҈qSM�Q�.3p/�\��s����1(HS������_I�Fǣ��.8ꚕ` �Y|����2�L�����y�ȇZ]5`W6�b��rHrhė	!�飏�}���X_��@p���n�Xe8�d[~��J��9�&&�Oh�:���h��C�Z�%c�8��ϥ�=���������o������<�Ue}�	!Ŗ�(����&d���<�O�_r�/?'=��-K�S�|��qh�?9�O8gG�{��A
�Pb��� � ��sLhJ�/�����4�=�����%��FJ�s�y(�����{w����04�����)��s��7| ｔ�����Uܘ�͜�+A�h���W����6)����5��s�@�Ͷ�K"U�gȀ?�����5����b��t1IinD+G.y"G��R�Lp��H����{b���(�y۰^3#"����\2'���u$Dc(�o�&8���[��)��@����.vi0�C	.����v`�<�b����{r!��0N�ln�<ʸW����]��P.Ga�Zp1����
b|�ƕC��uNt��4+Wy��e8?�!~]tϹ�:>��Q4Zgk�6�2����l��zNH�|:��S)ҩ����Q���1�
��1,�@�x!b#�EJ��ң�#Cݰɳ� ��g��K���O��	݄����`�9��E{4�i|��Efh�O0*4�:�I~��@=��X���m�v�P�/r(�����u^e�C�0iC����g:�܌��H|�q�VK��^CGg�^L�G������qoC}����_h�m_t~/��D�t�Qz��ah+'��_{�ro�������K~�_�4�@���l�<`��˗�1��{�g<����2��XtQ5�A۱I*�b��\��I�i4f=��x~���A3ul1�O��Ǔ��>���e)�_�Ա��6����qY�<8�t�!�y�'8T��> I?ʾ�k�60�YzX�L�����v`½ѵ�+�)����y��ݳ/?}t������W9`��v�?����^��铱GS�����Hnkꙍ~�t�{���16�Z�!�L�����9z&��1�����yy
l�ʈ>��׭���E��iO�A2Z���S�.8�&FipJNQ
�e��ۅ �=<{�ɗg�~�e�z'�dGaa���A�Dp�4��s�=_7�6��)Ă�"�X���WlB�⨡�7�4�A�SHh��'��������������������χ:����+�
eV�fCY	���~p����8R���X8i��I;`0vsJԶ����N=V���a���S=G�#�q�Hɉ�P�"e"L:����QJL�Ҕ���K�G�;���s4z�O��ɡ����J�I��3��b�5~���������L�gر�������18?J��e��l��5����8t!�p9������}ߞ���������'��O>9����>���q�D�^�f�F}nM�|��w�O�QU?��9�+?�EX�>}�c����V=��������^����>�t�B�ް���:83z��E>R�=���@�#��K�u�@g�e�9��ܟȎ��i#���o�iC�g�������4�>*�/?¤���I��`$["$Ώ7���NA[�5�F�����/�8����2��|���׿���5�B2r��Sx>�ᇳ����S&)2y��K�I��vJ�/Y��J�!���"�����i+�'�@��P���O?;�կ~}������EF����7<o߾������M:f#B耏ګu�8�'s��r��ߚ��Q�o�m�#���hN���/�蔈�>n��u��{T`�h���μ��7�?B�`XE�$�� ͗8������+ހ�<�q����u��볯�����n0���Z����������O>^p\|�C��ǙB^D����/|9;��e���5MgI�W�9�����Z}�0����q��}��N���ݨSdI���u�D�՚���E$�\~w�=:k�9�W���1�d����3_r�NNE�K2;�2��_���l΃�����y��%�����I~*�}!�g��v������y�(�)��=�O����O����3v�x�lBr�i9����E�q��LtW�2E��L��uŋX�Z3�����������_�����u/]`��vo��������)>`�{p�aL��i&� �a��,��R`Gϗ.����.��?�ȅ�~��.�A�x��V�l���*�m��]�����	ܦ��ӝ��xe/��xY�^]	���~v�������8B�y��PA� �!� C��(FI��?=�(�<o=.^�(�� ����y-SsoHuY~h���T�(��P�5��x�����Ĭn�۔���E��t�&f�e+OJ��p�[�Tc��NB�����g�<�����8���%~�<N%��-����K"�:[�1���Σ� ��Mù���]1��s��H;pN��ky�a���%��1�R1�Tdd��D@
̸��z�7kq>Sc8q��Ew���S�>�}��[����N��'2`��`�ې��*>���ǌ��H��N��N¯��<�x�7*9s/�{�ق��݉�޳���b����_~9J��o�=���4F�3�N��>({���|��W�W�3'L��!�z��X��q1�(����RD ����'��p�z���Y�ȝ{���C�ߖ~#_��ȳ�+��g1����Q\�~������o��)���E��Ӝ�/��b��I�]�fpiN���+��:aw2ğ�af��I�/N&�<�MFÎ����w[<����_V��qL��t��V�����������I����6�u&nO��}���+=���1�?�������}��ZF�`a��LG��`�����q�S�h��_L����������"*D �:|��I���RGF��3/��Α=�!�1�L�92|�!�o:n�s-8D��?��_%��P��S�����Gvr�M��A�Vt8�gqe���@�+Jut��	r�,����/~�n����_Oѻ:��.}������EF���گ~��������F.8a��)��W)��,���\����
7�[dK��K�4�7�8��3���;��s�]��U˔!2ף��݃�][;du
��db"2�KɊ��&
��іe�gsg�u����9�*\��g't��4���{tڶ����-d��se.4�gs�U��K�t�M��J�"�`r��o9�9�&�����$h6�X��t��}��ٯ��ٿ��_�}��'�ю�����g �����-*P�r�\��%7��td��o�&c��S��ڶA�6���\�DrW��h��r霉rI��;��O��w�i��Fv��j����.��.N&�)��!�	�W�o6Y�ν���|=x�i4��J_����N�C��g{\�� � ~��S�p0���b�C��S1V"� ��-u�ڹ� �O��S�`��n'Ȅ�?i�n=������5��o�p��?w�O���컔��(���ء�,�6�9Pf��V�zT�
�\�{=7��gh���t���*)��gwI�u�w���Qc��H��h��z�Ɓ�$h`R7o�xО�v�u~���Uz�++`�Y��n�����91E*�Z�$J�� M����zs���Ӭ�2ТC�9�����ǟ}>s/��	��>����2P�;ǣ.So[2o��y��II3��r|(cƒ����}����)��+2.5d�����O'n�#g&�-g�V�ɼN��9?���Z����G���٭����%+cDAL��=� �◿��~^��U�����k�3gB0C�`�CԁA��,O8�w7C��g���|#壿��a�>	�{9��Z()�N�!�?f�8/�%Y����f�/���������?l��@�:����a��@s���O>������~�_��g�~�M�М�:Aͻ1��� �#02�%��-%�ތ�/X�J�JT��黌�s����m�p���)�_��Wg����Da���όy�	pbo��}���~��h�w����g��u��x�,�,�rK���	�M�`�~����~��O���&�c^���4w%�|�՗��������k�6S�O�C�T)��xm�>P���~���7�u��E]��?�<��i�/F���W�o���%o㿉?x��}��D%�A�j��K�Ca����`#�t��!�I�բ�����"F�H���v��׿N�>�#����}z�漱+*e�6��?���¢��V�_�w?4�r�,YMN3^כj�.�G�/k@�\Ӭ���oG�u9Ü5C���f�L���ݹr�s�s�Q-�B�@7�>�F���(36O[���'��i��I�v��Gk��F{��y�6�wo�*еݿ�rh��=�����tՁ�I�����& �ёf��9r��d���x�w��=�)��0b) 2�+&^�zYG�Y���k�^�M��o�<)�{�������~��gg������~��/���ky3�*JQE<}Y4�~[{�צ��� �n�v����)/8��]���a������K�r�"�U�w�EA/��Wa�頋0�Ff�1�#�p#�z�~�65|If_�y>o�<nޛhу�'�[w�����>�=��5�f{���JG�	��b�ט��}��Y|{���L=��WĀ�H�y��D�_:ib�:��`��Fn��ī�7S�E̱�����o���3�ꢏd§⊎�J�]I9pt�{S�a\G��|������x:�]�&ᘧp��n+�����9�_�Ç�e�\۷�ᩮr<�<����9���y(��q����?i&�I�Q��gpfBoRѯw����2|K-]V9<7.�?gl�)ո8��� ���9u=2.oW_��ܺe9�]�N�#��/���`�`�r�[!���?�sT�g�P�"F�Sad���9s������� �y%�>o[Q�z����нh\4���{9����c!
fΖO�<�>�`�	����"��"Q����̓�/����ƿ���g7l��q��ȡ[C�����,�HqB10�k���Ù;>�n�nX}�y��&��9Y9�&rO�'�e&)�2�^8r9��g�Y���8&�?8�( G�%�q&܇��'z9��&gۮ�q��EtŇ�Mju�u
��&2�hΝ!�u(o���YT����9<g�
�t����E�}���r�Oo���Gz]wM�xC�DW/g�ss?ܟ����1�����|_� 3W���8s
8^�~b4z�κ7|�^���<c�M�o�ߪC�����3R�=�WG���p>zԔ��iO�|׽�@>sf$��1}�� ��3dkr<�j�P�i�
�>N�y2|-Z�=��O���>��Z���n���D7�d��aC�M_��?�^:�.!'cg���9^}Dn���5��!?��s�r���sD��F�pt�O������g�U�0�9Js/-��_���Z|��O� oO�q�^q�c�&E9Z��+|[��[��[����	��x���p��d;���P��Q6��>|e��>��?�O�u~��>�f������S��^�ͷ����괉�x�����������g����_���/�~}���E�M琦�ym����͝ҁ����|�hC��-gk�
���Z�<pvz�OÞ�0/M��)�.�AJ�G$�'����}u�q���?EP�ᖿ�F�'NC����Y���(��	k&�=��ӳϾ�|� (o�1���z=���ezql���n����,8j43l!��i����\�E�z=��o�6��<��@!�#����"39X%���1E�w+����+	��X�_��OS|_�[��������E�L��Twy�՝�^P{&��U��4����A�ۘ���qX7i�n͛A����Ois�FOQ�/&�=i��ќ��I�0|��g%�������qp>�&]��O�p��.�4V�3�w�4�~���jm/���
�_og�.�I���<T|�ڪ��BbO���lz�z���,P����zoj4d@C�Ƙsu�����9%�9pu�k��<���K[���?ʡ�q襐���f�{2��1B^<�r��[M����1yT��uQzW��dWQe^�,i��;^�G|
�2)3I]��:�y��L�|8N��{���ON�N �Q��4Z|�6T��Hn��M*���ȯ�Q��6���9���[�@�I���6�Ȕ�m�ء_D�V���lݞ�\M���R��Λ�z���ۅ�Z0�[?^��}��zo����i�$ZP��>Z�YgI4��Fvϗ?�KE������8��қy�pT�zބ4��$'Ut�|>]?��&���k����g4|�<𖎓�_���+|�)�O�]��C�����,�<gٰ�g�=**�}4n��v��ӈε��l(:�.w�S��7o&���/[l��F{�<�N���9L�����ȶֻ�D8W�1��aB:��	'�[N���?�P���H���e���|��h	-i�����5G��7t�n�.$�t1�E/��nQ8m�ZpsT�����
��viM;�/i�X��u�S�Zx�r��i�����݋��[)/D�9D�oDb�N|	MGEW6�Ч륃#G2��鏣��Ғ?��{�>9��Ϋ����P�z����h#Hc�=����mrC��z���*��xn8q�N��Z����Ȍ.��8�䴲,\��:ٟ���.O�F���zrhU����O���5�x���M������=���/_�lCo;޻s��_=:�?�ӿ;��������(=�Ճ��J�A�$�iW��\�j��^b:�C��q��gT���t��^ė8~:���F��[�ME�v[+�>㼟�H�L`�Ғ֚|ފ�˛	��"�7h����qC��:W�JL����G1�x�O
S���q�sB&=�#%�* I�,�����Y�o�G �8B�ƞw�g�7HR��Lp(e���kK��,��<m��a�b�e�6C�~�-�		�0˸{��F����(�xϜ�g��_��ξ}RO��մؚ�%L�JQ�2�o��S���	��R۱��k�0=�Թ���Hb�p�#�%_��i�2�=E=�n*q6�jN�-׃��=�-ᨓ8j�Q*�L�m
�k7��1���J�b��d���-%�yF�v�vk�C|�ϝ�c~��C|-�^�E=J��x�;2f&苐m�0��O�H
����|k�y��>u�,��q���*��xl/��=2�(�6�:#�z\c(��FAq@�x���9�=��(�qL���a�4�#4.re�vf���n.�����h@yVa��71E�nN�b�|`H|E_�O���i'�n��#��`�	���կ�Jg^�|&*�R^�p�``g��ߙ���5�1�<d{'[{	 ؃CĉsThx��#��h�-Z����ٗ3���#�[�k��4wM(�YJ .ё��6&t��~��E ��[ta�_�>J�#Θ���Σs��J�����]�'�����-��FہZ<��V]�je����E��9C5x$dFv�e���Z��tԹబ�ך_3���F�9G�X"-9�"�����~F����{?�!�h��F'�h�3���� m$�����������h� {KU�O{��$�Y�#�Eg��=p9ǗW��f�N�g#z���:mڣ�X�G��<�u���pXէ]��[jQ{��nў�OP�8m\=�{�e�����32�|*K辗؞��ʣ�fd���9؉d���f������VѠ�o��_����TR�ROa#q��t[l��i��q�'��O�L�szY,Y��ݞ6~�+�>���i=u��4����b�ת<��<�5�z��}Ut����g��_�}�������tt"^�0���t�n��SD����8`�~8�s|Lux��B�-7�&�Y������0Y\�����שg�믊�����n�ػ�!�բ�wr�+�4������Q]�J������7���Wф�5�F�~�y$
W3r����H�3� ��Y�|#.	`���ar�\S�~/`Or<�z܇W�o?%�E?~|j�t!w�a�\�mX�y75�K�gh��h���`��sτ��i�d�f���W�L�����o6�T�����5Ú֛|�o?J��R� ClWR���p��~��p�?~��{��%�D�L6��u�'�4N�Z�M:�N�a�_i�Z�BWW��<u�z��?�5~FO��Z\]bΊ��[�sy�fѺ���p��k��1�{w�7ѷ�e�8)R6v־�ߖ����5T���e���9h��s�9$;�����YixV���IN���q�iH����Q(��;'��"�����ab�㐬f*�,�=��%?E4�G���,w]zx�A�i�?�~l�u)z�[v}�ޚk�r���:F�AJq����̻2��X�L���.�G�]TCop=�1�n6��y7�*Qd��+Co΄��ڕ菨���)?g��u����>g��
6�\�7�u�A���>/�P`�A&��F���'H��<?6mE~�3೔@����{��=G��v(m�|"��24O(�o�yݛ \��GCs��2����8ɯz1�� _u����]Ɩ�Ckm��6�_��o��@{ZA����E��ư���g��[�#E�n�T���I��^�KyL���Q����z  ����}.�!��C{�GNѕ��fDI�������W�O��(�j	o��t��T�*������!�[p�N{e%�c�������-"oT�E��#�C�����,FOΦΌv�C_�0�
��X�H�q$��5j�L����Q��ˆ�,�9�B���`�;f���gEC���3�0W�t��}���=�P�'�`��^��ىn�l��L`��D[G.y�YaFχޮ�$=��K?�y�V��n�v=�!צ � �ҫu9�`�[�䵨,&�Z pm"�����6���ߜ����y���e�^;O�MM �r�=n��|�hU�̭��#���<x�o>��M��ݨ;z~�v�C��ؔ`V>ٳ�\��8���Cs������B|O�F����{7S�}��Ă���n�D���c�؍������O#�<�e��tzcD�y�*3��p砌SC@8R�_�znAMóvB32�h��v�14�,�:aۜ��a�7j�͸�(o��ZA[a�5J��{�Í��y>`@��1��E�(���D�?~��4�����[~9n�b��*¼�.��NP�>�t�m��tu:����e��JWC���?/����V�ݖ�mI��ß1����\�p��U��G��QC޽�����ϰ~��㳏?j(�~=n���]�[mm�w�D/��C���Z��S�b�5��ӹ�����S»-�e2#��a�W�jHֶQL�bPQ%��g];o4�������S#M`H�t	�vz�d�C��瀀ݜ����kN���G�D��Ic���T �&��g�KVEc<��YP7'k��u���ehT�h��_�����j+�9�򦏟�L2��ރ�z��HQ�x�1�zd��<�%^�����]�[��A"��+>����s�x�f3�#��a����
��&Sh�I�HnJ�4�T���:��4ʾ�<����4z�uR�u����oD���$�k��22���q��g��^���Z�`��E��6�@q4���(j��c�:h�(�Ы��q%����8n�OĲkN�ۘ����|�ax��(��#m�T���>����u�u���Ύ.B��0�'j{��}���ñ�h6�� e~�\2�*�W�[Gr������џ��Eq�n�T�L���Z��'
8�=9�+CuӲ�?<����A@>�m�wz��\9, !@޿�`VB0��D˕C�ꑝtfOx���m%��tb���f?X.o�/ˮ��?m~�O�X�`�֣\*�GUѠ�T�~K���܀��؜�Pu<ݗ�+��J��Bm:�L}{��(�n��iv2\="����騜N��g�;�l�z���go�����iώx�6�qq�q+�ů�<���������ޛ����=N)i������Q��:�H�Q��'�X��<�bl�躝n~����%U���E.a�)�t�eՍ�����@0��L:V/����(���۽�o�H/���㰭���/C����{�8P�f��#ST��Ϭ�"�d�b4a.=�R�CEY���M���t��Q%zN���^�����˔����7�p��XBfz$4"W����^y�wS���]���A
=Xâ�y�y��?����ѿy��w?6����|*᪐e�D��u�	�-O���H>2(o��\��.��>.��~\�C��3��Y���{'���c�PN�fy=�$���q�].�U�>���'�RXv��~�%��|�� O��U||^�������՞�ij�������$��h������;F{�6�ss���eab���g���yסz�l�p��?����V�7�Ѻ_��vN) ��~�e�2���` փVY�{���X8��\�i6�s܃��'��4?�eъ��C���E�z�LE#�h�h0�V�MaS��0/�aõ�:xp�-#qk���8�ᵢw��>hy	�yOS�/Ç&D�����[����>m�;�P_9�Q�r/̝Ӟz����.R7�Yޮ�v�^����z���Ѳ�:��-�Lz��zy�P�B��|�C����T2��	�T��v���;����iX�#C�&be�YF�0���(�/��ҞeJ�����L�����6���MV8�3$X����W}��ǾH��w|�(Z�����ڟU�E�-�a��͛t^��0Ò)t)��c��I�([oD��&��*��2�� ϰi��7j��D*��c������Vu8:z���~p�{cњn��G������嵎Zt�Ρo-�2߾�q�V�J>��K	���Iۍ:�s�u��ə�;������d�gMa���^����	��_��DߨH߈��k�7���[w��Κ]�_D~� �dI9of����Bw���ͼ�>��:���� ��:��̓�QeyP�{��j�t�h�D�z��Y�g�t��x�V���\.KM�!t�!k��=ن�|ܜ�'�ܵ��)�|ie������
o���a?{���d�H��ޟ��W!	�I�C�Jd�Զ5:��@S�����u䀥�;���TZ�/�)g~Y?��� [ͱ"�3:���oI[&��O����볿��>Z*��X�ˇ� 9$3��~pv�/��Ȯ�&�C�>���Ӷw�F�Z��-=OA�=��ߌ~eVƣ��4��a2��I�ڀ6a7� ���/����љ���6竓!�Ute�i:*����sc(��h�5�$,=Fm��Ÿ�8M�:��Q~�G";e =�EVAv��z By�R}�����<xԐ��1�H2�FƉ"�U��/����}�:'�U_[����� W���(*�́���o�[M�|�_楃+���f2���>�lX�X���K�
��u�ypW��_����/��r��ӱ2*Ly(�����W���4un�Jxʨ�mMS���Z�qZNһY�53��|:^u�F��L���W�oQ��c���M ����Y�e�5��l�nz	Ex# \� p�M�t΅��m|ܫ����^A�!�@��=�M�"� ?�f4E����gWf�z�7m^Z���h2���9>]�7r�s�S� i�Pu�{�ΐ�9��fF��a�i�㈝�((GKdITEٳu<zj�?Z�&��޺6�[l"`^�6T<�}�!"K����|�ܞ�� ex���Z���-��x�9V�3ê�qf^�{Ν�s�8ʥT�_����Wԃ�W�@w��4��y�[�����U�I��HY&�+�u���RP��8}"BO1�m�̲�:';�GGu��u�:���tVa��'��"݊N���Lɔ�����4D8M�F�JY�un�����	Oy�[��t"�^h�&��&W���tV�e���e�h-���Ot��Pg�u*�n��ӡFtYG��v���!�~�[=��n*�v��SF)� v;Y��Jr��^�I��0�ED�s�j3���}'%=_��W��z�V�ݢ���7x���m��T��';W���|�(Ie-��jy�Ǽ�UzQ�ig�R��Y�t�9^�hdl�����NP0��K�C�'���t�˜����|b_N�8�*���?g���KQ��X�����^�v׶9tzy��12F΂odgj@C5mmG�Qxȧ�U[m9�򼏱-�.1�O���	�ϛ�!2f�#�/�o��l��~���_��g9�ә����e,O�H�a�߼u�����UJW���3`�u��ls6�p���nt�bGr�w���sp��
`���<l2��=Nmt9��3s��sL�zQg��:,�P"���ypݓd� $h�@����CcRD� k�,���$��Ǒ%n�O5z6^vh��,$�Q�����:�SJ��c�^����;�R�6�`=+�6�`kbG����Q(G���y?|x��֮���>��AϷoV]4Y��ư9`��F�-�W��҇�(��=�]�� �89�zB�E�i��sh3e��CUp�����pH���x6��?ʎ��M�SG	��G����kR�g��� r���<���}|����)���0���h�^�ă�,�SN��`�0�����m�����o�r�ZC�w�^<�[YOϾ����V��7Zj ������%c+Z����0�����"8�<�0,K��-�	L�1^R����\Z9�<]䠉�[5���4�G����D!��c��p��{�ބ��$�J�x��ψφ ���%i�Ό��놟r���쥑�2Oi���z��������\�Z�w���@>,���1\'x�"E �]���L:��dg#)��66K#D��&�W��h.K�Ȱ��k%�
_����.8qp�� �@'��s; 8;�0�x�W<��9�߶�yս1�'�&/'�[�޾�X���y�����96��11�����L�m�Ζ<�Dƴ8��^S(B�!H�>#�E�EB�W�����n������ϓ[9�3C/��B롵4é]�չ����ɟ��  @ IDAT��^�6��,+k��^��<Ap�9e�-њ���p��� J@ε�aFx�M�s�9�"j��x�3���r�C+�Z��h1pG���{��9�	DN_v_���nB0�����{���Y���h����� 6d!�[������;E��s<;�c�C��=�萷R����7�*f�6Њf�7c^{(�e,�N���=����屷}�nu�+_=�1��?��G�$I����M������]A�
������ f�g��N����C�c�d����y�anfnfn~�g�j$���ԯ_�qqW�����A�^�O���{��2	��D��w���8A� ����#��ǢѠ"�l���k .��';YPz����5>}>�W_�:���􇶜��õ�:�z�k�:	�Z�3��wb�,��C����nc酒����Z������ݑl��$~|��t��T(��;��e�n��ZSf�l�3��5�]FeGG�d'm�w�;K����N��D|�tA�A1�"��.�����#��ł��z�s�,��َ<��h1/��g)��BQ#��R���JBb5"n�Ր._鸌\y&�fZ�%�[a�X� �/J�ҽyª��y�	x*=��u��ef�ʷm�ix��˟bj�77��*���2�P�a �����;��?�V��^�l�b�'��_�]�/Z|���,��MDTZ)��{�y�VN?�ڲ.�ɽ�£Z�zn`��5�)�dK ��J'��ӂN��������ڼ�2~B��zgM��'(�wm-���h[O`��	13gx���N��0
� {��6d5�Ќ���iB�8s�A�W5k4���x�����}'�4G�ׄv�N���j���kT+/���t�2){Q�_1��{K�1v̯�bszD�����G��Z��w��g2kq�(�9s,�zZ��E��x��54�}�%�dm��.<��VT�_=Os�V[�ZHp�3����FX���KQ���v#~��7�:�[����8Q���,ϑ) �H�|<�M^^���<��ӻV����S�
*��R_��)	�.ց\mG�H�a9g���$�exQ�y�FP �����c)84A��P�ҫ�������I�f�;1��<Ac��N|F�i�D��R�#�2����H��)L\�<�K�\2�1��C�2�!!:&O������fէ�����E�O!�X�hĨ�ghx���{M�^eAqxx���9yCc�����m�����#^ETN|�G�=�7<i�bm'd�4[J<l~�.�w��Ug�V{Ӟ-Р/"~�s:k�i)T�[�������O]�`�ho���_m�7�SO�+K�g2T�	 ��{�bgT���ͺˣ��� PBمoB�{_W����g�7�|��ʣ��}�;yη�wrj�3�:[�.\��z����c���<+�x��G�5�&�x���-T��g���t^���u�S��l6Y���d��0�tʴ}��g�,�ŏ!c�ą�{�֧?�v�xK�bL�O!�V���
�:�Z������|��i7�uc�F�$J�z��A�?�^�x~[��
}�<��.9zL9����<�����F����Ȫ�]��L���FeJ���K�V0_m�dz�В�tv-0*l��x��l�:�y���\x5��lVS�U��P*��VzUJ�3 T6�I��U��P�D3�y���}L��7_α?�x����t������Oy�k�]v�aN����7h���\�a`�q���w�w�Ň�����)���_be��č�����)h�!n8���J���u/��u�Z	�����U��KGq�{��p�ޓv�1�{��z_�zn����M0����q��͏p��x$��m��"O�w΀�i����u�fy4~�/QC���7��^�Q�Ѷ���
KN��Ǽ��\x'��h��-��+����2�����@�f:
�b�[���s<�Ќ푧ō+:!�7?kݗy�:�2!B���+������k�=X��'�׏rc��(OЛD��!ו��eg��E{F�.�V��� w�̽��ڟ��	��X}P�4��Jӓ�Ѱ)�i�*������0��+m�P�/��Ã� �3���8�ȁ!��1�)�%���M�����N�[�����hI�}����!��!��[x��?�e^����k��7��������6��:���B�ߌ4=&�xA>�#���e�^7?�<��b+�4�ʩ�+��l��զK��^����Ɉ�_n8��6#?2�^gH?k���m��&,��Ho�adz��V<��56�n<O���Z8Ѧ�я�����^��!%ޮn�g�Ԓ���*�Bu6H?���𢎐���>��d97�}N��0s.�{v��� �c8���t���G����G��)cW��������9^O�����o���r���=ѳW�{�C_�2�+q�xuV���C�<|�Hm�߆�d�����'/�t�����I*m"��N��D�����_��`��ޒOp5����ʂf��}�=���H�yߥ���ˤt���L�H[uB�E������ޯɣ`�N޹�G&k99�f�Էhޕ&�w�7�"љ��'��a2�wL_
 �Hg�~��U;/�;g���C���1���]�s���G�O�W$r�θP�xEM�޵1�M]�v���O\��i8�;�Y:�%鰂O��p��I���SvQ��i۲Z25��. �|��0���xCI>�>��z��'
/��y+u+�4*�	�z�,I^���c�oQWs18�����:,���\6 83�4D�����*�u.%�2��M�7��R��u���k�ƕ}1O@�[B������)�+��w�j�[C)ܷ�}�~�}/⊽j��~o�M��ß~O&[���F��ӈ�bxV�e��Z��G��r4ʓ�����;��N=����c\ɃuTc�R��7�8�'�|�Ĺ�����w��øФFs �߼��e��u����ѕ@��xb�"�b�sՃ�Bߵ���+I8(]Q 9��M�5�̀H\N����h2����΂��y{��܅��d��� �in��k9z�e�QW����%q	��kl�*�nQ]>��˳�0��z�j���y{7���D�U��V���v �i5�V��-/�7cD�nF�eD@2^���!�s���a��z��SN���
�c8�]˵||�o�]�Μ���c6Ǥ��c5G����x�{Μ�����@�P�����(���xo�@[���;?���g�c�xt��K��lm�0B�T�<�y�̝��Ë�f�}�W¥�ܵo�X��t;���~ojWd�H220��b��c�(�*g��c��ǈ7A~Vf���4Z��w�?�]P3��)�թ�!��jH9X�"�_Õ:�+�V����	|[��Q�� �c�.�F/
u���szA�^��9E9q}�~h���+dw�w�"��Ŀk�B�|��n��x�Sd�+��x�,�`��,�(��z�6kc�~zky�*���Q�o2`����p���Ãǭ�{À�A�Ne-e`���<�A�̏ӧ_���������~��	<��/�e�ֳm�!��)ܮ�KfU��+�����y-���_%�W1�^�V��\��1��j�/>������@?��Ȏ���Ad{�7��36��36@�v	A�:S��VH`b�c�P�~I��&�2�[�������jm��E�.��K�W�a!�Ȟ:�`Ql�g��:�7��y
��'XJ;�ɴ��a�?���UhU��� D��u%��a�&���f�z6������m�P|�V�`V!: �x�4B�4@y]�A��>�n��8�/�-�K�&��F��Q3�C��UXz��;J�F;G_L�R0\���E$K�OF%�g�UwVme�d�,j�8��o8��8�R����8D�)]�^B_~[�[�)bBחbo�x���:���}/Ҽ��z�������׽�	��쇖�$+�X�̷�}�x��iݵçp˼���I��M��k���&7�h����I��sa<�8�4�I���%����Zz��|��sTCC)\�}��U��^�<����x.��P=_T���$��O_gZ ��E
�|G�<Q�l�ק��7M�Vx��R<.Ao��z�<m��ö�{iur�2����üJ[��>.�g$�)�w��-��b�lg���г+�'~^�E�()CL�a�0*	E��->зP�2vxƀ�K`��[��� �Uq��a�
FؘOh���l��Uo�����
��;�'�frl�]��%�gy{��#N��r���E����P�A���jOC\WF{?Q��I6Pf#�F�E����o�SEVxt.�~̍�H��R��72.z[�o5���>�4 �Mm�Cr�s�v.���<�kÃHA�m<�&��y��x���%+gn�]q=�W�{|ul�3j�9s�2L�
W���*e1@f[O^:iyx����;���䩍��Ld���R}̵�O���W�5K�q�>hd����\���䐡ig�)�M8�r*��^^ v��n�Q�A�ۥ�b|�
���)4�=�G?ٗ�ܷtT]��s;��@Fgx$���P�E��7�,�ox�q^�n?8���٭��*�9O˛d��M:�Y�f�&lA˺�7�(gj������ޣ/<�@�6��xK�ש.���<��\�G�<��V?Ӟ�1;�J���-��ׁ!�^�^u}\~d�O���2���F�����7����� �`*�ksgh^O�[)��;. ��7׎������q~|m?��e�����x;���cB��7�L���O�c��#�1��xI�~@0�a��P��:����`��>�u}ؐ�Z�CU*@y��
76D	D0œ�e����fxk!	�f�3�"sDqg5מ
�(HW� ؉20ŗ��J4��<�I�����`E߮�5�����璶���D�Q�ϒ���`�I�A�[��j+����V��ޗP/��)gpN�*�=�U�8����>��"�y(o}[q�e�R���2W�{+��X$�{\��g�b�5�A�l�۷�'�nd���"E�&zk�]���w�uƃ�<�6�x�|���N� ��y�l
��EO��4$%�<�q�WWS����_�=��7tL/�������L���:��׹��})��e���<EB��Q��م�|(��"����\�#^R�=]A�rm8)��6��Y�L��f�h�!�1�\Hi�� {gD�0��g�˟��<�_��͓�m����b`�l��A��X���-�HI��ݓ��_y��ז���(���1��#H���I�'�[g��ڳi~����W���]��p-|?iޖ�<��Ù��63pj�hB��/ʋ�����%���w��-�BS���m �������w�ٳ��1\Z�_�I��ޙsX��Y��^A�����:x�)�	�z����慰*/9��f�:6��l�ݾ����ɳU�Q��HNC�nXr�-R^V����9���9�E[�]�0��wsT��x��_+���{7�։��^�b�=+��摙�V�ħ�Fs��2F��Q~��1S𧍑)��o�Ca�l#�;Җ�����9�M����e8k����U����͋�_�3�~����hʘ�|F�w��S���)ޫ}ŧE��^:�{.�uR����x���vټ�?�#�S;�A������Ow���ۇ��x��7��8�����UO�(b�`xD�X���C�%l��9�y���NN�\��������Ԇ��f�kE���Kw����L�H�Fp./���*h����V�t���x%Fm9r�Jp�|�K���y���kUi��!X���N�NnΑɤ<�ujME�*nu�/ؘ�������6���ܿ�!�cq���,Ю�a�2=�g���,�3�+���(��,��ˢŔ���E��/�Z}I_�~�V�&`|�
yj�{F��>U�ӌ�WD.9BT�î���wē�c`��A6$��h��n����	��+33�f~ΪYq���ZM9�B��l�c_az]'5\ʑ������8'rV��8c)`�L�[���U{u\�ڟ�q��K��V�ar/����j�t�k1�^��@���CC�LJT]��BJ+��=�?�NˉW�`����ؤX�ŧ����S�D2����㏷����_}��j裭NN��.�s�{�-�Ye��L���J��#4{��{�����P}���Y�w�{���=,�t ����|v�j�d}>�D^m�����9~?��c{i=������z��@ƌ^��<�-F��~���׿�]��5~�
�V�)@��Ue���e�i��o_7��j��O3L�?��~���z�D�c�S��f��k��*M�;�!�{�r�$��6���������?����(�*҆�R��mg�{�fxВ�j;t�	�G������߷BCg�����/sk�i;�	?&�7�+��!W���)�~������b)��)E�=��w�e`f8�P����6ߵ�퓩3#�I�ڽ-�ǎ�2�'���n��s4�o���f*c�.�9G�"�W�����9V�08���iRF����;C�o����w�E%/Ç#�D���țt����<6VD�흧�y�<o���&��
��e��筤���أ�my�}��E�yfv'�H�7<�������mx�zy����B�{<�C�~�i��dT��}z��{��$=��ɻ�!�cLY�y=~c(�/��~�Z���B�<=p:�rr#��gm�J�����9������w�NtȠo; �۵�Y�	+��Q֫�(��f����ܶ0�����V"���M�'Ω�}���7���s�v���މ��0*�C]{:�3�6#ۥ�`Y�B�%GJ�{�0 �ē������χ?g������m���c�2�t����ɺ?�U�^�	���í�uo��9QN�H�⋷ޅ�k�-8��eF0�tL���%��"pG�`� ?�MV�iGu��jҕ�'�iǳM���G����d7C�Q˩�Fu���|0�M������YH5�#ˠ��'z�P��+\�-���9HҐ��Ļ�G[�-���s�P���f�9������wt#�bM�4�6�]��s�pyzu�A�e����;E��oE.�=��4��{�D���(l�|��
�j>�1M��oҕC���+�Lo*��p����M#��oemW���>��1�W��Wq(��6P�K��o��ozP��p@���2��\����+������ك�g	��<��wS�-Ζ��W٫�J�w��ޟU�d��-l|x�7����Y����!���d`���/!5�_)�1�-SQ~5�R�%�s���Ǜw��^M�\JA22�6�T�K�0� �X/��I�XM�}�&���S�}u�ex�J�%?�5�<|Qv�#��he�`���v^jX��6����5;u���83��҉G��mx~�Ԭ �Y�Bz���+D~Y=6�4ρ��a��U�vg 1��c��K��yBx�8*�p	�I�SJ�v���>3��W��Qy���e"�''�I�L�4�4ˢK?£ZF�c���3����疥��C<�.xO�X]��覃��eI6ޛ�-ђG�B^;Ì%\
��a;�!�<��;*��C>V&/
o8��.��[%{�4xxn�>��7�-p0��5��i����~�$eP�o��#N��$.��r6q�v<�hx��k���V����`x;|�a���./��J�;��x�gZT��qlm�W~5H���0Ʋ#X�e��u�W����L=������$�\Lǹ2��ByP9�3�ѡI�CF��s-�����]ۧ�!#>�ε�r[μ���]���R^0k'��,�H>�K�2nyH������7|�D�xh��ŋy�����ԯ���W�c�f�>���:��jx(t>iԳ��
����fϱx�1������u<[�׽��M��yo��7��׵�۝��׿�t���;� �Y[�	OxY��a�.�.5W��_ř�+(�W���;��?\�>r8x�k|:����&r!Y����ԯ��ɞ���X�2��҈3S,��� �|7�M��d��"���Ck�Ͽ�)�1�Vf�ώ����<�q�{醮U����\��V���7����{a��ӵlx�J	H|���Ц�4�_e���@�qζ�U�s�'X?\A�!p{� X��X�`����]��� P�!�����2����5.B<�ӅA�`���+��ʚ��kr��+�<G���)x�=�A��/�BH��G���i��(����b����3_|����w�U�)T���ɫ[����<�oo��g���U������`�21���t�'���-���D�/�֕e�r=½�2Z����}����ˋ���A��;F�T���������ӝ�?��L��w���Z�p�ua�}�؞:6�#��l��x�U|�Ý�^<&Hʽ!筽Ϛ`��$�(!��Ủޏ�͠����������F���o4l������~>=�;w��4Îs�]ϵ�kQW�vi�&~����ܔ�L�vϐM8[��>�!SHW�^1c�U���rܕ�����%=��'�>����#�"C�j�"Y��C��eh��Eo����7�>o���+�ŷ�Z
�u�|�~��K��E�0^�g�0�w�W_{���~s����!O�����k͍���v|�T��4�EL��}�`�R،�o���o~����[yj(<�pb�Q�����շ�b��+̍�y�f��>������N1*�4��i|e(��<O��H��4dF�������~7Jo��<�w#Jo�q���]n��z��.��#g�v!?����ۯ��Ms�6S��FY=7�
:0����d 0��ǻ�	#7o}M��[t�Ϣ����K����=k8H'&�ؘ��]����&Z���?3�l��M�2<l_�'(>ô%4�i�m� �����:�S7�����V;6��I��Z���s-(��/D���S�5�j�.�����Ra�-��a�K�����ڃ������Ό��!�U^o_:^�}�
��e�p�9U��ny>��L�1u�f�i�1��xI��(}�90�]��]���q|Ҋ�/��nqAs%���@��#{�#��BrR�	��{��of����^�3�+��^��M�0��CF~6ɴ�����HK6��"����4<8�ON�p������
y��[�ʧ�����k����"V��O\s"�v6�ɍ��ȧ:A�:�`��x́=#\��~�F��l]���/��!�x�cz zM��w�0*��� ��b�������Υ������ս_C�2�ɘ����n({�ҏ#f��s��#�Zϧ~�&���Õ7A�����	�*��� h����s�6�������DM�+��S @B�5����7���?����?-h>K�ǚ��Ϫ�n�*���dl-�)	X�1�;A:+~@o;�w�I�!���Ut�F)� �w���뇬l{��s���Ğ��{�G�ʒ���4``p�����u�^CW|I?�7��|���znUF��`6L�������xϥx꽫��f�@*p�߯V�S����?�%�����KkWl��z�?w�L�1�������r����?�l�'�ߧ�ϧD�g�S�`Ћ�yi�K<<��z�wv��;��n�H��D!�(Ey��63�+�6,��C^��;��V�A~�dpJ�Rb��1 _ۘP��"9�d�I|���C8a�\���d�G:��x�ΜyNy����G�:��/[J�i��;jCLx�UB��͍��9�sv#q�ޝ�&��M'��fq����> ��'� �I��p�����ލ�T���f�x��JJ���'.�����m�t�4�.^g�5���_���^G��&�P���^Z�MஶC��g;���1y��7� �Y	�A�ޟ\}>�a\�� 7�����>�]�D���MSD׮��aa�o���ݟ9j��u�9�NU0'�AH��)JI�dZԭ��7&U^}�^��	�xFԅ�0������;v%�7<cҾ��-U�]o���Gᆗμ:^Q�M�
�e-�[u�#���=�x�LX��E��!�:�U�����F�{����?���ڷ��f�P�'�6i���m<ys�E��=;��s��̳ʧ�6�ng�����l<���C�(s��:"�����C�V���[y��
��H汛��#���<%I���%�%�3���'Ɍ���7�#��K���/o��$;���|1�|��K��g���lq�t?l���r�0�ǘ�ǩ�HE�?9��T�ʛ�����*��$�.�v�W�.8.�<&����?��p�g��)\�BIƑ�m��쮹���_�o�E)�9J�d��2�&��a���f���Cs�^��1��|�0>�0�2��Wz���	}]�1���N��&���~vMpOI\�0+�������(���J|�QVЄK J꩝�e�peo�"�����וh����+����l���VО�������v9���y+ă�c�A�'4	�a�_�1���ꇏȹ_B�~Z�Ɣ�q����q� o&�����γq\>&RJO�hY�1ô'�C=@C���E�@�θ�>��|�>�޿a	*cp!W�D0�R�zb^�C��+�|g$	�>p��46��"�a1B����3��쁭�%��!B���I��6�$����|&���[N��l��_ꁚ�b~уxԆ|��3/'�5p��}�^���S&.��<�����/��<��U��Kך�������< ��G��XX�f������oY�l	��1�_�s�>��N�6��4c��a��`h�
�z݆�����b�瓳;��Lަ��;gS qԖ?�^�R+�:כ�c�N�^3eD�~���V�~C<J�2<U`�6�i*�9`�U���8�6Ό~��l^BJjm��Q^)ꇏ^����$Y�-)��ӳg&�;K_0p-Bh�H�����,g�Y��|V�w<D���DXaz�cG��/g+�dU��9���Fk7A�#�Æ&��# �-��g�(�����e0���D�1���Eyu5��P%��(|������A�Z���?�T��1:laJ�1K;��Û�e���ɐ���Da���h��+�v7ĩ7֜�汼oU�q|{��w��Y�_Ƹ��e�0^�k���^^�7!���2,a&�?��v	�ߥV�k��g�?�n*6�J�ǉ�`p�L��q�9T��h%�qv�ŌC���fn/��k����ps1��A����ʄ�`	N��.�Nش�i\Յ��������W���e> ��]�;�H�-��]�oa�Aɣ���a���<c�*�3@ߍ�+����o������G�����2�r�u�z��R���<~F=�f�=�-���6�Q���N^u�1w-^w��g���P<�o�
���!L;&g�=���c���P��������2a�B���2B�;����i�7Ų�I~��P�l^jۻ�<!���
�$K|n�s����'#���0�u�b�i�>�|�w���V�����AA3��G�&�w��������y�*��߃o���ˏ���?���nzG/zr:��NK�۞�d`��{���6�
��춰�������MN�d�ߑ�އ�
�,cK?�����)tKq� ��|Zf�.�-_1ֵ�#$�Y�C؛kCؘ�U��\��F=	��ԓ�] ���������@�J��]��r�)�
?�懀y�aqda�b5x���A�-:X%İrI;�))��)��+Y1jx6��)�V6u^�&cU�Ty<ӘT�b��(r[Jo�ͤc����2ؾ��{��|�\�Z�7+��V4=z���׆~��u���I�z��~�kۄK��[���u�#��X�Fy[�d�5�ey���j>u-�x�9!W��o
������s�@j�E�>�£�H������GyF�,Q��)-��̩���^5\v-��$}��Y1��!���<@5!4Z�2�'�=Gʾ�fqy�ְ�{󄪚2��mW�ks�MBg����=+����,� ��6a�m�Q�������&�S��x�R��1���C#��x����f����91Lz���kQB�����$8T�Rp8�_U_[�G��+�~�R�,F�;U�Af5��6���Wn`d�^�i���Ņkˌ�h�������5�z�}���!���?�<c7�Z�hq�󼓭3,�M��ܚ�3�I�ʱ����`��Az#��	�ku�"(/#U��!�����O�嫃!�M�J{b��G*C˰����Ð���~�kTz���w�뷠nʋ�6��[��[C���=�2*��k����=�?��Q0�[�Cn�L%���̼P~�4-�t�o������u�����������Xp5���\<�:ZX8�$/����b�B�(���N�p|n4�t'��E=����DTv��W��[Rt�`��Xi��:\sE+'�����xD�d )aڬ���)����쟑|V�����I	�Z�Zt&?ƺ� -����o�	���-������z�>lמ�ϕ��e=�<'���E(��m�i!W`+\y�U�e�y�������h��?z��OPVY2Z��}����2�8�L?����[u��@�aƈe'�
��}z� �e����G�N�_Fa�0b�"a�.d8%"�oK�#(�w�F�;�E��}u��������{wA��X��6	���\
>P��5��,�JF5��ܼ �FR2�U���os��H��D�XI��5� ���L��;%�{ќ��9A�? @���o�~scN�Z��z��Um����H_4��O�f��_����M�=���8sC�T`�ں�in��7/�f�����"��L�~<��QG���p8�c���x�n�.䵹�H��N)0�Ëvd^��jd�tp:C��~"
���qsK�Ѥp�xM�O@���ke�^�#
��8�[�����9d��<_���7�nc��X���p�R��vګ�UV[�`�]o8n�}��<�S��O]�
���E���AQS��?1򚉇�	v�̞Z)9i����oP�+�Z�F�/���ۤ�7��e��RF���e�	#;�(lt��/[Ug���{Wu�)�Z��fֿ�Y=�����ĵ�2m5q��᨝�y���2\��_���.ϵo��}5F��Vr8Ԝ�������;=ó�#���I���i+]o�|x�駻�.�1�A�3L͝�O�L�/Ɣk�-�7��u��(��N��|�0㓌����kf���-��p.��ʖ�j-�,lH4�M�z�ǛW�J�ex���.�L���;���D����#��ms��'��=4��$s�{��0��b ����̘74��a�ވ���Ml�a�|�Oqд�7/3��<oq��餕��q�_u�᛹�y�f��ȟ������MB2n$�/���W �_y�!܎���v�wE�U��w�Lɭ`��x��R��:�:�:s�9gr��?����.��7������#�pm��LZ��`H�����}�iY-�d�90�I�*����M#0W K�q�*�f6��L����I>L����+
N�dCi���S\O�g#80 ��x�?L�e
~L���&��ׯ���9���i�2����c�l��Q�Ӡ�_d~����|܏n��D�N�/�"��J�IT|��r���F���J:E�])D蚈E]Pm��/���?��Ϫ��>l4�bKm��>����C~�/�<��ą9��M�g5�E� �:��<1����{�tVL!�ɿ�<�l���3Ê��L��T�]�d	�����)�+w�K��e�i��oF�wF�,��q)�dl�S��EԨ�4��E�B��|��{�Ќ�]�yl{	Wsq|��|�Ȁṡ-��]�@�95^�ʲ*	%(q�;�Ȩ&���N38o觞-Ϛ93c�Fυ)U�p�̶9�d�[U� ��c��U7�D�gy���ҠN���ee-(s��o�q�:K�y<�rsI;�/���!���N޹���޷��f��(�6+F|C1.#h�}��3Ų�!Zu���l<yS���o��ق��Z��ɰ�#ޭ9ʩ!D���^Z��Kby��������W�����`��Х��3B��t4O�� E�%E"����~f�Fu���(�?�����p�^c�Wf �]��b��;S���2_��fd��<�3h�~��.�˨��y�W<�S$�ȃ�`��Þ�W����i�y��Lɔ.�����%ڍq[9㙭��1�o�s_��A�'��	��D��.��ⓩ����J�S��w�om��?�a�%���E�������^� �B�p6X��ys�35y�|[r'�U��jk��v�x(�	�c�4��lƾ����lh+[=��g^p[�h�-��1�P%AS[���ؕ1d0Ad����Y�8���n��l�O:��GpT��KC1~��P��&M�������J~Ƨ�#SV�jɮ��vO'���.�y�\�)�~�=_g��&?�`hV�}����5�0Obq/d�Y�1���ˁ G�Qm �,�\��?��
	�����y���T�����g�߾�I���O�F ���\�����Zoc�H|����?b��Z�3{qV�������äH�TA���p=���I0:�{��"��/�\��*�/�b��
	���y��%Pc�>(v-}7/�j���#4�<s�j�V +z/}Z#B����UӍa+��K�4�°����&�7\��'�w�션p9�5��oa�g�&j�Y��ө�r^�9�_��S6�Qc��佰WR�n��4�}�k���\���G��������í�Әδ���%�1-��A=�W���J^1��,�[뵇�E'd�&�ϒ���bk��[0[�z�r���;�|���M��U�Zu�gk	�i(M�ڤоQ\��I����I��ma�2��R�'g�UIl��_ɺM��H��7��׭�C"��|C
�E����eH0�g����r������I݊�H88�`c�0�>i�͍�t�<�s����GL9G���#h��@�����E��r#�Ϛ�4�#8G��=���_�Qw��C��s��qr\G�W��j6{}Q�c���#��1�^�Ng!�j�x���O[qw�{N���nJ�E�xQP<0��U7D>=wHV�`���q���s2<W�V̳���x�v#��x['��(����҃y��۶����8��9�8m����;�Y�g�6�2�ު=m�s�W�0R/e�80�u�����~\�/�DB�{�U�9�Ӻ�/��?W�g:�����#�G�)g�����ly�����+�����Ջ����GT>ꏖ�(�e�Gm*���v}��^��ݜ/��[Da��U�,�w�ܔMo|yƦr�+�/�x��L:h9���a�Q^��˃ʘ$�H����!�h�w��U��rF-�9�[�.2�bF���<���H�����&ry��,�7�+���5���e�KY˸݌�`���{�-U9nu��/ނ�<�a�>��h�ۗqj_ܳ��e͛]xW{(��+���Wߙ�Ϟ� ��d��!v^*}`4E�+�П��m��>�w�}|��ζ��`�������e3Y�Y��P��i�[&��d=�^ͷ[GJ!�0J�\�#����kC�G����^["��z�4=��p�=1L�Y�P��Qp�8���b�ʑ�8�1����o���k����h ޶Ɠ�#p��qj�0w���a��O�1{Z�Z�m�ߪoY��/��K޻��SxZx|la�S��obcɤ�.8��e6{z������߆ f��zt�P�9]#D�r4<����{q�a�}t6�'Ah�c�Rfزx����	xn�ni,���=׼�+�&���lN��>�������8� @�ӈO��ፁ0��
#��fDY5�NaX�͞-*�7�<q`�X�a�s�0,��ſꈾ�n�<�,[����}��"tF��-�M��=��$a�R  @ IDAT�_cޅ`@�)C9n�%����yG�N*��S�|m����q1C�0#z�$���G%���{��2y�h���x<�alS�VZi�P�	���MΛ�e�G�f� �c��ͳ��l�S8I�2*��V{�_��V��.�iU"޵ b:q��8���WM�~�����Ma^]� ���JgsU��7p������S'����� ���M]��[yɑvVV�Z�c�+����@���GTJ�܇mF���&^�%�����CC��1�Ѽ��ţ�l<��d2.�?T���&��g�C8@+</�?H`���eU����^]K���s��;���f�yã�ۣ�o���L��V�c�&�M�W�`Hn��vA��k&;O�[�~3C�+_�U*ru\}������Y�r�/��v뽰Ֆ�6Ym��+���5e�D~k���n��YL�JJ�5,�W�7�C_��q_#+��
ڢMR]���I�޿�QlSzAᩚ�� xq�k<0�/5�<'�d��y�E7�l���!憺Ѹ+����(�,�۫��x�<(��I�w����2��c	�F�4E��c:�S��&��-��G% ��[�3�tr&T�/�Z�^q�U�)�C`Q��0�" �D���~/�	(�n�V\�>q�|D$U�H�FV�iS��+������ߏ�!L`]7�����}�p)~O��~ ���uK����a�*=_+k�^'1/\1�M|��f$xV����r�-f�>B\�$��f�t�[$p1�{P6�O�3�T�Lx���B�������{p��ҙW��LMN�w��9�p(+��\
<a�o����0M�=j���hEҕ��V�o��#3W^�O�k�	��?���ʌ���oc�sdÁ��QC<)��wU����*���}Dw�;\���I ͽ��EWl݋��U~��ad
������6�C�Ջ�&� ��[9�C�8����VVpZ��τ����.����>��Ő/f�C�G��eU��^�d��l��0�z�^0@f�#>���O��9�O9hG��#����5���_F�yN�TY���(��]��
T4~���k�#~�e�R(�0d�I<j�ޖ��k�S��+�V�1���Rγ"�����y^t�(�̚�9xg�>�(���o2�.v��P��y�3wz��8�Pg~	���v�^:�~.��w�A��PD�1��-���!��z����ˑ^e6��Q�i���D\�C��x��&�@8��Ъ��sV�GF�<��<V�pf8W��?��O�ou�xt��-��;�D�i��\��<s4YS�í���ކN�,����k2h�2]}7�d����p�Р�:�.��v�߰^ւ=ǘ�.C�>����M���o()O���b��=�_����
�䌰1�õm�f89|��!��ph�̳���U���[鵗�����嫁�:^��c��<�Y�٪}m���v���ןZ�scd���M-9x��Qe�G[�+�gi���ڊ�Ņw��5�E���"�ic��W��x9�'L�\<�-�x����N̳-T�����>���
]�����&�� L����3�1���@ܘP�ex�M�1l�i�3��U~��L�	+��W>{;����-�4��y\�5ď �+�A�w5(�oo�v�i<ðꭞJ\���q-�3����c����S�� -m�!�(4R��ַȫ��l�W��#en�O�_g�'z�SL�7^�`ã<�V���o8��E���� ����z���F7����`l0x <�Xј�f����R�I���j|gg!|�����^.��������zz�o�be�EИF�hT݃ѡ]r�
�'�\��)���C5��Ă����������;�̺�m��1^�Fp3��g��	WZ6��7+.���"XU\�z��4��߅�Q��� �f��j��M�U�~�V ����<c�׏�t������ =���4���!��c'�݉9x�al�+�aZo��憡k�6��ӌ��k�[����2�X[�8��I[Q8wr&q��US�:�i�r�|(�u���e�y����a�Ճ|��ɐ[xE��6��FUmA�M�I�s�R�0�l���*�W]����#��e���e4�&nҤ�[�,�����sc���ʼzIG�R*��~3�.�"�S��W�!��Ⱦ>T^���]l�A��k�I�3�%���j>��%8ۍn�:0�m���7�?߾�a������#�ȴ�d��y��V���<]xj~gh��8_�#��{.ޛ�D[��z஢@�t�K��w ��d�7Ͻ���Q>�.|��|� ����C뤐�0�p&�����Vi5����&���6�ڡ"�<�C��Ԟ�:qMy�/`.�xCA��
�Ư�vI_�n8>��o�S�Q~�����n]�|���[�� ��N^�_�e5�0����o�����(����W�_�9�� l� ���뚰�`���w6Gʪ�e����W?�c�V��xp�=���}���S@�@N2� �*܇U@�%M���Uˠ�䀛��bUr���n V�&��Y��#���TᩘJL~I�l-�F ̷���v��WeW�����
-AR�N`C0%cxƒc;��yg��d��e���^fL37���X���#x��ۄ�I��?��p��exDH|&��Ũ�ͪ�a�a�J^������&S�OQ=|x�E�����v��Iw��[,b(h��|�H<��ʺ��g���}��Wd n���)3X	Gƅݡ_�yդ�<Mx�d����K���(e���aE��Ro��z�v���m)����r�*1�q���(=�ҏ�� *S�v��>BCۏ3�Q���Y��3�΅B��>@I��}ql@J� Xs�ɚ�jΐ����?i����r��������ad������V����,NP�7��ᖓY����4s�+Ah����Q~�;SV��^�m��r�9�U�8����=��(&��տ��/s��I�~t�~�k��+=u�&��Q�!���<=�R[4_�UH�u����D����1f.���u���mrv�'�����Cu}`pP�#u̅9:�)��2�q{6yZh04�H�ov�Ϡ���[3lE�W^h�]��7�<�$��*���l�	��8�c�(en����C����Am��ݟ�~�V����v�/��*S�z�\����9R~m��)�o�|oy񬙿����8�P��=m��ޙ�)�<�a<kn�=�tb��-�x�!y�l�f�U�Y����ⴸ2�
sÁ�6`������>��{<y��ɉ!gx���S`_<���y�ċګ3@��7��2�ZN���y�c�]�(���k�j�ڒ�sqV��#cc:k�q���Qyx��p���ND9Ó2���4��zNǰ4�y,���)���wt������3�Pپ�7�m��>�}#c��x�LO�Vɏ��2L'����e���C���p�VVMw�1��DXO�ڂ�`n`Cї��cu0�4���{��\����7`�Z�~���w���0)���h�����+\�N��ۅW@�v��	�O�0(��&��+�n��%Z�뽽�HR��EQ�\�.V��e�>XFjQg�a}�o �� �߹X<+���;I��:���TjU��;��GC"�R<H˲�v��d=����'g� ��OC��K H6�>/��fR��}�F���&`m��@rv^�vSZ�3XL[RF�0�zM#(�4� +;`�a@�f��MRWw�;C]�cǌo�owq�/���s7&�*��]_k=}ܳFA�NV�(�R�5���0)j�S�Ձ���Wi0չ��f&�fl�:SC#V�0�Czx]��Κ�Q��%ǯ�����	�iV=�����'�"�W�T�`��5�f�Kp��8壥���P�c���p�K�-�V��^��}ޯ�橝m6�8g��� ;�I���	�%��Z�S6�/�}3��eCo�A|�D/s�B��,�:���cz�ቐeTU��SF��<O�iM>��/�]��mk��a��D���V�YY:^��;�`�盔#C�Uۅ8��ӷ;��i���?��l�j%ky0�JB��]��xB����g`��pR��~�+/���ˎT���;y>����1F�8���S�r�	.��qlR?�+�3���86�myh�'��fT��%\�ϻ6��`�$��7�L[�8��ד���'��6�_�5";8�V/��߫�Ig�^j_��ŵ�Au#��L�htZģ���Se�<�棝��ͻ�a�Ҕ��!�;׹���ރ��)|�p>k5��^s��N�!�Ȉ�0�� o�?h�������`��em�?}������Iuy��F��c.��Vޏm�q�J�[m�yۭP�:8:vp<��ܻ����Q�ԭ���NNE3؛mr�[��]�μQ�i����(OÏ� 5�Qp.��;�N�8|�7��paq�!.ʊ'���qp	�_���!(f�X�� ��>
]��Li�훜�j�.�BV���CX��/�����Dളj�x�k�}�[�B�����mF�㚎⡣���p�@}�ꍇ��Z�΢t[%{�V�`7R�Y'^�AuK{�T��F�㦖<:yy��^����V� |vK{j�H�9Y�<�a�g�J�3�O�1@ՓA�3�$��W�Ch@�_�u.��X�w��/��ͻ�na�F�.��;��3�L矼nĩ�ƨ塁��>�����o�J��s!N�){����$b�>��_o��<++Bv'��;_�FyƘ�qp�����ӗx��'�"��C<��ư`I��Az��짓v���ެy�l�\J�87#��+ɪ��p�����,%;+���}.O �Ѓ���H��'U\�����a����s���
�B�d�,Ǩ����LumJqy[L�;g>�	��5���>z�V�8w�Q0��6�8/�_��dpF��VB}�I{:��yզ�&�;O�j�b�JK(eRq3�ohT]��@!j�[E� -  ��
�J/e0��G:x���&��+��W�k��^\���*�m��Ac�(nH�Ǔ)x�"���=ǣ]�#��-�8<:��ðx�9�N��*IJ�י3ap���x]�n{8��0B"ާXxg��PJ�+c���^#��m�A�IY)Ș�&Gۡ�<�;B����g܆y�|����Z���s��<��`��L���rx������g�kM�]pO��@�3W��sy2њ��?<F�2��=XxZ�Q��/�<
�U������.��qË�3�e����7�Q8D-F�jgG)� ��=s����@����f�1�=|��aw���A���?7�z���W�O��Eeڪ`:Ax1D�iX�����V���O���
�s�ٓy��xgN�n�G���o�;�������������W���2�앵V'��ɢ�f�08�����g�Qt�8�6��Ȁ{w������)\4��ƣc�iw����_|m+�Ių`�_���<����9x�Ź��+����ߙ�����=��Y�V�V���,�c8ۇ̖(��r2�l���ŻV��ꐑQ:2��x�j\oE/�������Z��?G�#	�٪��K\�=�Ye��*�f�N��H"�|&���R���q�Ù��X8�R��ӡOX2��I;T��a�|`��8 ��f��I#|� �cr"���:�y��,���Y���}��P�m N��~Sx�;鸫3��L�Nָ���%��xa�@M�˃,�(SH����`%���v����`��vʨ|_�~R[�w��	7���&�M�Ya�n��A0(s<V�;�lFC�3ln��
��Y��.�B�~��f���&Έ%'�)�f��a�٩,+uD�U`�.#�9�M{�����yn΍�f�v���Ӕ�絧����"V�Ll[^��(�n���jcZDص�`��Ǣli�޻���8%���w8`���w!e~C������B`�C�8``�{ �H�=yL8RRӗ�	���1�i	��R��|��x��%4De�W�}�#��ؓ���-F�,��8yn�O!�Nr�ХX����L1՛����^\W���3��t�F~U�: �� ?��;Ct��s�!9{a:F%�dX<��x�(xcܓ�k��HN��>��3��w��	��C�,��DuIÁ�s���0�#! ��7�ݳ�.�<a�$� ��s&̇����4\p�}Y�3�z�V�w��7���f��X�rÝ<�y���*�����#J��.vfc=1�5�y�7���z8�v�e=�۝�w��z�t���&
�#С��g��c֑A��@UC�^���1p����aޓ���)aXo����m=����Ė�p����`�3�O;��U��r�V	�������d ��{����	#�$�����CG�u�]r�թ(� �;��B�k��ŕJǚ���$�}�C�`s�2H���d^��1��}��5Ͱ����e��&��~��Qg��6�sŇ��F]�V˙Ћ攂�wO���/��]q:���>�iX9�Vg����ރth�"9�x���:����7�����a^�R��^�=�͠��?}w����_F��?wΡ�������_�҅�x��<��0������ǳu�~�B�$x�m�Ì�����EVw�"�90���<�����:�~vk����9Fx@�KC����ɃmA���<����{yETo�����9T}�y�
�k���v���y��im�J��3�x��Z(�`��6*�|t�eE�塋������iC�d����Vg�8~2l��dc�ka)^l�0JF�Ƨ�b\�7/'��Q[�K
�%�hC��Z��.F��1�x�\Gz=���&9�/� ��ѵ��P򰕮07� :]<����l5bQyKV�������RƓ���F��4�ɳ��5�/������4_��@��n��'O��h�mΛ�u<U��� O+�*t�t�y��n���_�(�z�������W���r#,�~�S����`[�n%���пg�9���]��a���?)��.s&Ե��V��Βkt�+*'�����r������)q��Y~�Q�4���1I����۵Q���5��`�o�5-vJ�w�����X�5����zm��ł�A\ ���K��،G��=��Զ��\{Q��
��wU����V�sE¹>FZ@)�G�1�*���;���=��e5�R�w�\1Yu���~G�Z��W�s�N�1tb���ڜaV�����]��,?ƐF��m�A��GhHl/�b��O�LO-��;��2`��w���v&�p�ZOo��3�7B����I_U����]�N��1�9,G����R}�m��ͫgE訝�:z�6D}gC�!����R�J5u�A���N�u\/�ms���m{��M�KP�����j� #��:e��e�k��ɣ���������,��$)�c��	isg�C��M8@�(Z�IA0�܆�����ǟ�{����LǠT�����KCg�?y���ğ�!�hz�/�����,Bo���M)QTv��c��t��u�����u5ԗ�<������/�GJ��
�|6��2�x��)�'S��g�x��v������?�ג�}��qm�x����/\̓��+f�o�[a�mt��dL����?����N9h���� �c�"E�'���w���<D"��i�Ӌ�?��Ct~ю�&�������x��M%�E����I8sn�������.ϑ^s�5|�����3��}k�z*������a�xJ�᭤T���N_�#
~&�G�z9���?'K�-ԾO��\����+�N�v�*O��"�$3(>^V��z�a�������[y�aJ� �RȁW�V�2�O�Itʬj�Q��3�_�s����_������Ǩ$�̳�W�b	^/�ypֲ%#�0��E��9���0�d��J�x<��a�[�qt�-f�3x>�xߡ�ڙ�w�vN�}�:sת����/�jg�.C�-�B��-
1�x���霨�|��x�I������yen޼ֳ��Q
^�� ɫ�%��������*#h�0���$Z���?n�<ğ�����Q����_�x7:�rc�������:/�//��`�I��9��xb��Z#_�i�y�2jZP�AgA�N,��~��[��M���@��v�c?�s�߻tx=#������NظV���P������'��׺׋��=�J�<�H�5}}^flөo�[Dўn��՗�������Z,|�y�HJ��%z/����Z��y�W��w� b�kq����K^t
��_:�u���
)��>���=��c�zD�i����ŝь���z����^���!��%�퇧OkLh}�����w/��  R�ǋ�KE^�e�$D������{x�cƛ��x.F������ԛk�0�����GQV�=b0F��(�<���s�}d�d��w�C�T}�M��!8%� \0��+0��b��a�a��L�|RO��a���9F#���j�����S��)��5��v̇10/����we,aY���ʾ�6i��)��>���s�9�6���xk���&����#����ߴ��8o�5���J��7N�Shp� ��4���v#��F�ӋN�jDϞ��3Z(^C[3UA���)�S��3G��*��ye�3�`�a�p��0{�)=�,��s���7������o�����Iyx#v|�PVC6��f���xk�,5`��^��{TK�	�5��ջ{�0֓<`�_!�#�鄗���<L�_�ȓ�~�Q�9Lw���ؼ�c��d]3K��2��^�g^�1tM�f�y��z��V�o�B�:̀"�\�)�^�Q0�������ȶՔ���+Ζ���g�k� ?s�lҍg:E8|�9F`=m��Q�o7T�iإ��4�㵟W��yxG4�H�X��z:�g~C��a�(�_b�p����i�-��l\[>�@*b��`�駟�"�x-ym�Qi��4��P�36[f��GU���s�]^�}��e����M�� i[���	'|@�֡k���ю���3���8|L�a�����HgԽK6��0�t�&��ˊR6J/���\^�♠���qbB���I�a������1�l;Q4��;�W�$��u|`K
s�n�">/�<}pK�V��jD��=�� µ�	v��R!����*<3���74��DNk����/�v+O�'y��������u��)"���� {ӆ�OoGg�a�t�δ�S��+͋��3q��E睂6ʕ�b�3B����(���1&�7��ܥ��<<�IΜK6�<�
���>ׯ~����?�ָ>Ɨp��{���asܞ�Ԗn��=n>��臟��~-�į���1f�3�n�7}3^<�)�npYA3hg�C)����;���O�n:D�%��mp:����������et�x�=�E�NL�"�6��΃���p�N��<m�=`��������4�����|�h��ݐ��gkV�3|�頶�`��)[�X��v�ǫ2�"�'�W�MZ�<hӗ*�Kf��Vfk8�a��7�Z�[2���`̪�`�UyΆ����,���k�Ȅ��gR�a����$������gc�ػ3 �GI���?j�B͐�����	�i�ƒs8��~%@!��џ�8�ז1�)�OH� �$iQ{n�|z�zZ�{���?��_jx�ECG�0���8W�g�|5� ���"�3�J�	�k	�o���b?�'1��ë��_e�������HYt�Nޖ�������z�Je��N�?�ɻ*F�,᠁}1�r����<��6�4��W�����z6W���@�0���a����p����a�*���9&RG0j8�~"t���@�D��\z�@�u���/+�ۯ뙵�9/܋����d�a=�HHR��z㇆;��K�e������`�����!x��3���O�#T�?yb�6���=��O<�}�x����Çk�	AM��[�:���#���s����gZ%@�F��� K��PD��\�e���R���2�j�g�.e$i��/ف�%��[Ou;j�B����E�g�[Z*��<l���>������o���!ބg)|#g���z��Z�-|�h=���P����Q^Ǫ6��3�Qkj ��>L�p�̄�_�k��Go���O4���A�R��Hs`x�i<�1�ͪOi�s�_�M��xg����j��c�_�d �#�e<�z�R��;���핇�$%�.�U�jS�J�}�b6�.��t��nB��z�t(�Rqz��+ZP����	��57��� ���e'`�/�kx���,�����$���6��<�U�C��R��9|�K]�P^�S�o2��?�#W����e��	��6������w����w����婋ǂ����#�upՅG�z1,�B`�Wu��[F]َ�.�au8���P��r�H�����_|�U�-��lE�-(Wϙ����������O3��������y�~�|��o��;唈F
"��4#8�a��8�(]��<+o��`��O�1X�̄�4�>�}r��EF�W_\?|����j�-Hk7d��-<]�\yw�y-ou�Q��!�ۇy�yJG���OM����yӚ�۰kgK'��`���ߢӒ{=�����-��4����YtC����'����پ�3�.pW��鉅��,-F�i�`F~�y�;ɣ�oSL=�H����o����_^�U;\����*.�pm�ޜM;����+�?i5��ں�3�\���)�Q�F���R�u�_Se�:��=\�Dj�:�%�TF���M�㞎��}��aJ�,/Xu ��w�y��.WV��Y=^�ȅ�<���T��U�l6��k�<����k0�XɐŚ�� cx���Q��8CΜ��[�St�I_˗�V4�6/���k	P��I�$O�+�Ă���^D���b���Z����:����$��|�����/w��95=VOL��UK�QP{��?Dd.�M���r�Z��Pn��~�Ⓦ���)T.PFf�4�f�J�
�Ư�~T��F��G���Ë����=C0E<e��6VyвyT̞57�?�㷇���ׇ���j0���>��Û���Gw1��ά>��w⠿���	��ux�16��N���9\�~�Q�����_��W��S�����0�W��\��h����VG�4�khm������?����1�MC�S��Rb���u��9���Q_^�W���޿ύ�p��z�:��z^�a�h<9����ϊ�ݍ	���,!i�Xi��P�*?)v�r�9��9Ƥ��hB�<m��(/&}ʃG��T�G���2g��6Q���f�Pj�[�~�Nջ'��
Oʐ�(�Ÿd�D��Fy�0���m:��f#�#ȫ8�/�jAJtJ��ˣ��ڠ�w��� ̓!p��F����1x7z�2��F[��kU�s�޻0[6��H5Ln�%��x��N�a�s���S[�5��wʂb��y1�B�ԪE�{��ߓ!x��c8�0V�R�%,�.�L	�W��S���e~*�#��>����Jo�r��LoJ	q��(�RT�%��\~�,��T���(�1��i?��򰽌A����c|�dl�#8�\%ڗ�|T��:L�ꘌ�W�p�R{<������e0��F;C�z�e�j���*���+ۿ��T�D�ܓ��|�e�FCV�}V�� p*���M��>��{���[�g�@�z���-l0�M�+Y[&����Ƶ+#/$ �����'��8F��;\Ew��L^���C��n�Nk���ͻ����_�ld�R�Tx����n���|Ĺ�&��|zsr#y�eżm.Փ���z�O��k�!#I�s���V��?�_Gf�4���e��s�>�Ҫ���U�� e�;r���l�^��Y��� 7چ�)�~`ڳ����6��ps���U��}���͛Cɫ�^�QAFgho�����\Y�r̃�|�����%�\�7��:��_����u����I{�E����.����u�mv�F�ߓ�L�I&����J-��t?��o���Ҟ���uK*��Y�������J���<�lX�@ ��t�|��$�n��6���
;@l0o�Ie�Ϛ����@��>�4d��h���'���Qjs(���\I�TxT�lX6� ����Y�@#�P�5�ISCV�M1\;���Qؠ�=��_��*2�Ϟs9"���u҇i�<�R&�	�!�]jGSQFɦ���g�=�Uny]ܸ��εl`�&����"�`¸CZ�sW�:��2�d�8S���0#Ap��5�/.4�����\��Ձ�R��r۰��TZ�Y�Z����c|��ѣ��v�Vӣ6�n5�	xX���v%eG��1^�Q��.�x����;���?�|�%��p�fʩ|�%�x�`��+gw��������[���]����FC#F���b �d�)zw"fsв�g�nyi���mi]�9��B6L�"�A���/��3��N��>����ci����5�l�rӥ_6Z�|>�L�����cVUv�����=Pe�e<�w9�?6z|�_�%!0��YL�Si�:k/�·�XK�&+����LL�������t>�c9�5C�9ʿI�0��_Z[�(�ot���Yc<�$0�.�l�b�� ��Y�����}S��(ax�<hZ�[�QĀҁ�62"xVK������F�7i�;8ux��Q�q���+MߧAOG'�t���� @￻ �U���L�"�Fc�3���։��"|���i;/�k�:�m��O�ڹ~�f����Ӧ��~i*K=�e�C	s1�Ki����gS�e���xGm���q��jP�����6�f������$�U8� ��  �U���yVoè�>��.� ��w�V1r�Sao�f:b/W�`��[ً�	���ê�M�BF��M���{��@��5(�=�<t�s��L����MD�q�_!JO���@(��<Je�:?�����-�x�,��'��r��O�J�ӌﯳ�w�n^�o��g.�|���x�M�5P���l��;Sc��*=�7e@�4�l0u����|3�[-���s���*�A�1�>�a �ĳ�N)N�T:}��`%�y/���]���%i;�����/���Jq+ �JʣN�	���� ��ɞF�����Bm����w�~��A��ʧ��X?F�l5�c[Y��1O>3@�<@VY�-�SV��]g�j�
�Cs�:���G�6�N���f�Xm���l�	�>uh-��]������������G�n�����)W)�l��ƴ�c�gpՠ�eZ�'�Z����ԅ�F;W��*S3!	_������i̎7�}�=�~��1�\}I�Q�pT]�Qc#��%��%�/���V�i�%g#�'�=����f�L��cND�3���=Z��d�&�U@�R�e��fj�" ��X��:	LoT��S���3�Z���ڡ���/	ۈ�}ڙW1X�G*�eSf	u@o�yɍ��5ݢ�� Q�9g%fB�G�n\�TЄA\����ʄ��?���,m^�aJ)GX%��U	:G��4���Lix�bGi���{��	`g��\��>IW���5:�h*���N���jvO�=x|a�.�fz��:����~Ъ��*�C1�\�9�뇯�w��O��.�B�����f6�3���� ��6U��lNF����ب�紀�y OH�-�S#ރ�_Jp;S���^�����.���9ˤ9���hOK�1�o�����[8�����݄�i<LK�%3��8ш�_%c�۵�Z.�����k:�p
y��ם+���6��$�j~���8���i�OUZ��n�$;'�_m|�Z�}tI1,4T?��L%�<ED�C/���:��pn�	�]0#Qt#<��{������h�ה���-|�xԀ
8�O�^�v5�'ώ�.P�r��\7l�I~~T�a["�o�O�<����6�R�^F{��LNeSpB�wiL��ݜ9]}�)mЦ�0��� {����|�l]�������4"?����w�bLm�龎��)~�,Q��GG�Ҷ��D�Z�A��{�u*�l?u
;�)����/h:�;��$z��[xٹx�8�(�fR�7ә{��G挗@1�#	=����c��Y��+l'�q��	�KAP�-
,�2 �ϵw#l�Zy�4�gj��jN|�t�7[�p=l��ꘁR0�Th�Á�]i�i�W60�35�&PZb�=� �|��";�Ӆ]-B:���j��1��.����r+�^�2���o��W�"^�&dt1���d&��S<ji���\�At�V��O�.W5�a)�T�UG�۱oĻ�u�g�����ի�,D�ٷ~l1�����fh��~قi;+]��ЩË	&m���"3�L9v	`�RR�Ş!|iQ,:,^X�1OӢNW�5����
e�r���|�J]6��';].G��T+./�k��l{g�:���Bu'!Ơ�v�y�'������3Hk�^݈���/2�xwpIѢ1]�_�w�`��Y�R?+<.��]WU��E>%��n�78e�JK�р��XL�K��۶IZ\p�;esuh	z��b'#�9��sL��>*�'Z�^���ؐ-0�ʧ���X3Vy �w	�?h���\LV����5��U0��,U�l�Z�z�w�1�o���b���fC� �&T��p�{/��H-PY�"�W��G�K�FUAl�rP���rZ�xdC��0���9Æ��
����aK� ���Ǽ~��?�y�F>y>d#����#���>5gӏ#��^e������Lg*"٭J���Ng{��`��*���Yu_���;����~v�^�����O�����LO��rr�p�F~����~����1~�h�B��d���)%�Y���b���t���N�������*�o�=t}��������W�h�@Y��}u%���2Ҽ83̓|h�V��N�GP�%�/�;�Z��￞��\��/�P�q���ۊ�F�m.�ߴBm�;h�B(��!��*�ɉ�~"Z����u�B�<�z������':���	5�Mm��`^�*���M'񹁅09�m���q��	�)h��e5L�t��0cC�L�rP���X
 3���|�f���S�W�� ��>��d�W*+DW0-PzWľ���>�;��׫��n���wGLa�MX0�?ϦT��T�Ѽ�;t�:{J�����ի�ow�O3�t�3�V��t��4���xXgV��h�-)����^��6��*��~�a��������a.�@e�E�Ԫ[~�*�h̷Lws,�����Nb����֦M�:e	��Xo���х��]ո�\���*��sC����V�@-4��z��7���
����J7�y`m�t�Z:a���<�Щl~^���tt%d��}���������l���7��G�����#�>��\�l������>h/�����`7`dJ{!�V�_�Iy�>��5�i3x]W�6n����n�Wz:^�e�bP"<~�p�I� �&gw7�"ŋ�0�~����D.��)%Nv	_��ն.�#�cw�b�7	M|�X��	S��w]	u���E�x�_��ٻ��X�t&A�D���7R�iY�x]Gc���Hd�F����u�q�[6�K(5�c�v����q�CL�3�TX�_6K�m�
��ݟgPs����cZrn�����XX�{����j�f�w��+�Y���f3C��ޖ~�N����M��?�<�����w;_\:?$ԧ���b��=v��<zz�p�3��iNN@]# �C�W���:��D�:�/�0�5�����1��v�+��-G��u>������c����e�R�%WD����!�W�3�3{נּbWa9��9!Bb���)GZ�#�-l��&�O��lx�a��(�sU�VC�)�4Tu|9���7B��i�A'�*`g�DH�T5��~�%Y2�`	  @ IDATG�3�b>��:z$#���������is��P�ٔX��3��p�ڹ�HFɻ��1���
A���yԺ�_)V+g���Tu	U��aà���jg5�O�Ί0a�}�N����_2�nD�o�<��}��ȉ��;�5���4W�̖ĸaWҵ�n1���k��)|�N�1�n�1��:�{5>ӷ����U�L�^h_/�J|�����#,lG�5xZ�2�� WL�<�_���&���NN+��Q�������J���w~�ۉa"{i��PcD'c�����$И�~���E=��W��:��hnl�*Bd4�����v�*��A��h�b���sq,����ro�SYU�T�Jw��� �i�e���|��ʠÜ)jyX���uӁ�ny�+7h#���b��B��	��ٽP���:/V��[��1��܋�	&� ��	�	�\:�AøR���si���������<¸-Q�g��;�{��7!��ө'��H�ګݍ�އ�=���~���~?+�,vy� q��ɫ����;Nn�0`K�O@�?7�z���G�h�����J�g��-WaSH�?!����Vp��?��\��3�����[_��ߕv��>��^���jx�<�i��_[��Gޛ�	��4����*��K���7S`�1���{2�!e��-��K8����	�B~@P��`#�	��+̮��Z�u��A2���րu\ϟ?m��q�r"��vT`z� v:���ף��gi1���bh���v���2�:�����T�|���s|%�:���o�� ��Ȇg����_~��Yn:�a�l�L����)Be����˟����L�i���w;GС��&F��U��럋o`��ַm��w���M�?�������.����A�\Op���yB,�/����ϩ��������v����,>��ۭ���������Y<x��Mmw�A�&�?�������e��1M؇�A�Ư�kE���}��,p����ޟ)F}[���������X�&�xQ� �� 4|!�p>���>��ۣ���ܼ�2�����-�hD_�͆SZ��G�ٞ>��L��w�͓�X޶���˧C�|�h4V��}*�T��x�ƏGG�9[l��@�P��<��
�l��պ�,|�r_�N�Fǚ�;�q�nԊ8Fh(���C+�F3��h)�f��њ��u�wǈ�[~#�:��Oٹv�N�*۔�g�d��u6UN�Ҧ��!c#8�*��T3�[��/ә�ޔ���%}�a�₥x���j���6B�Ճ�[Eh)6����ۯ��t�<n+�೭	�8�h�x�\m��K�	{5���͠�H��a=j�F�l�F�id�0=��HC65J�f��MS����Ay����
��u��Νi
3�Ry�T���:��M�p�@�����Vc^�tq�g�m_���p*[-+n8U�<�����7fԂaq�������������{
�Ջ\=��}������q{NZ5�u��[Z�nk���Q���׼���1�:�A3�d�o�/�E�C�ѫ���D��{��-Oc߄��>��y�����\q�D\��E�2XYIw������{)H�3 `8MD���	��*��)��>c���wbn�'���o3P담�M�c'�m�R�⋳;?������|�ݗ���6^_�u��^'���k�fE/�Ȭ�*�N���m��ۯ�����;?|�M�������=�����wj?�+F{'�	LhD8"�����:����ˏ�w����#nV��IPVp�)���4|�9`g�+,U��S�M��U�v�����$��n	VEݼ[�����S�кI[^:<�� SCa4@H`�Kc0�.滄
����k=�}#�07�O��N.<���j7KPR��,����h�}�����GP�q�Έ������<�Y���S��5����0�Ե�7�y�H���!]Ǖ�_윻ry�d�z��T{i@�&��H3Ek�o8�,ñ4���6z�����^��{/����'6�G_f?�ӷ�?3Q�;�B`�޻�.�5�x�yƹ�g����H���X��g?�<#���F�\�|�/.e��ޕfpRv��M�r�4�8�|�5�	�S����R}� �qvR?�5�	�K��`?\����W�뷕˂�<���2�p��}D�V��N��M9�1|�ݼy#eƵ�6{(�W�ph�L>$7�,0�>>:���KΠ_�:���ә'\>��3W9ljC0}D3�b��ﶨ��	�~��>Á��˓�v�ku0S�=���&p�7G��=
�x�+�O-ebsfZ5�n�x<�3��E���޻��_|�ua�9��z�r��4a�9`l^�}�|s7bŸ�o5>��ƀ�� q��� @@g�ݖk"6�W�	V��@��D5�D!U��)��x��g��\ID���nL9Ґ,�%�H��xi�H�4_w�n�K�|��c���F�Uc��f/5_D��o�a����r."Zࣈ-Ù� dʶa��W=sbD:$���P*tZ��7o�6�c�p��+���e��q��v��sIʗ/���ND��a�hSq��:�H�
eF%�ƙ*�;�ߺy���="�q�p���
Ĵ���D��lڇo��h^5�b���\v^�Z1dz�8A�a��uz�����⨾��4b����F��#8Q#z���`4�{o��wpN6�x0LI��ߣ�Wƈ���?j{�)߽wo租~ڱX�h�u�����Mǰ�a�����$I�B�bsj�/�-C4;g�����f��
�1�sD�Ι�3\�m;H�#-j�V��8[���zY[�H�x�Y������P�z?0N�%��@������J�WY�rbn����b��i���W����6������������Mi����ڵ4֫uc�1��i������e?F��vr9zb:ap`
�=�v��o5�B'_�Mi��(�D��g�[�>zӿߔ��p:�i�1A����r9֯��/}����� {1w���!�I������6���ͷ��w�]��cr�~� =��9&��7��h�>��k^�}�8M�]u��� �����\k��o�����h������hz�S��d~q,��?��^���K�� ���6�:?q��7 &�}'�GsSƣ��w�El���)���=S|�N 4Y�_�!Դ##�f�X�R�/Gۈ��tpe����1�.c��`@^��*�6<������ʬ����X�i�P9=΁����}O�Z�e�[]l5�
V�祍O���ζ:����p�]�4wf3N�:��<H����O���
W?�[��m5S�G�����tcD'DOp}�ԧ&8��r����vfsi��D-�� �V�a���i_�"^T�qU\��.���t3/�
�f�i"��>�Az��[آw��V�v* ���,�r?����������LsZ?��Mmk�2:T���M޻�>��y}�iaS�x화,�,C�{����C��ۣ=1� xǏ]�5�KJ�����g$V�26�z  ��:�Ü4��W{��a�X�Y\T�Ujs��(�0Ԑa>�_CCl�}��,�8�iy�\K�?��H_�؛�V׵�n����?5�� ��;�ײl���6j�|x�Mʻ��N}w�I�K�^D$��k��]�ʯw�{R�!��fJiI��+\�V�����������{�_��9FigZaȎf�	ד�bT��b2�*ۗ�$��h����n��Ȩ���Pr����������`3�!���o��������11�'}Yg�6�Z�O��U���qNL��޲������?��~0�E�&������:���v4:Pj���/�?6[4r��6L��WÌ��,^4M��b���V%8ژ� ?+�̈́ys~�j��q�ss�jkug��&e6+n�y�Jݏq���jF��(��^�"��C��C��u��D�FR�u�Cǋ>���d	�q�c/Zل���Es��O1Ͻ�D�" Aw�KhLٴ�(�fǫi0ݬ�R��_�.�V;[�+<�]�ϝ.[ 6�_o����]O�{��M{K��k w:���V�����a-��kV$���3� G<����Y���G>�g`6�gҞ�6;�
���v|�f��s�r�`�HY硬`7��0�9���㳰'�� ��/�u�8l��\�QG�sDU��ZB�op D��o�I��N�m����mh��7a�_��Vz��}�	����{%���6����浟���Ү�%yhO�s����j�S����o#�L[��W	�)w4"m�Msϐ�������)�^��^��N5m���E�}tZ�<����xYխ���h��0��D�N��M��ղU�5e�>A�b���b4]�-|��R|^����|cw�Y�fE�*f��ޱ�M�3:�q뗴Ji���o����n�h�Qz��>6cc��|+O�)�x�b�3�-ڷ˳�=��3���ۥ�]C����l�.��c�����x��W��6'��}���i��A��<�N9IM���\�>�qgS�k���cS>��}�Ϩ� f@���� ���w��'�|����ϔ7�N��|U��A��^�׃[�_2�g��ܾ����v�=�j|�u�as>{&m�a���b"��"�b �}���[5�L���<��RE�
d3�@�P��}��t����d��VA������Uϴ%4��.Y���g�I�[0�`!�N��=~x7�ފ7ը3Y��û�Uf��:G�Z Z��1�*V\�g��o�2a�A.s��w���<�esn���O�� 6�!��tB�%}��7�?j�"��~�Tm��<g��k7Z�~g�Y��h+MG��QK"��Ikr�%�G��a�T�h2bF��"z0-�B,_�����8�����2��<H-�$���D�T�ĕߐ���E���T��ۘ���t���~�JǯZ9�������5����ꏝ��lec4��8d@]6��SuH'��ўe�`NB��ly]�|�w�	�	`��ch�N�p-{������~���i��r{���|gf
�1o��j4x�¥�gM�4���6{�J�$������:X�0
��h�T	��Y��xϰ:K�#$��V�F��J��C �b����0�����(�>a�2Ѭ:��5��Φ��m����3z�����7-��`�AID1�6�M�/yT6���z��D��p��n&�Ҝ{��w.�Ϧ�{��o����I����~��WN^e��� ���ò���$0Y��e~�8}�r��c�Qg�KGѴ�.��7����;=��Suj�הR6/����Ɨݟis�`���5�h����g���M��0�NA�a+�zvx(��#���F��Y(������܈�M�`�n^���n�������M���d�Uz�/S/�u}r���o�r�l ���*��ʰ�:�.���h����|���mt:�;�⩇"�L�|�qS��Yx���'�����f)����믾M;uzh�R��*���9����>�hV?�e�±��p����L�Yl` ��~��,����V�%X�|+^�/	�[�p�?#���E|��~+��O,����&�q�"w�V;�fϟ��X�Q"���Iv@	���L�^ܿo��>ŀU�M��ϣ��@���j��/K���?l��æ��rf����Ë�A�)���p���Ƨ�Dm*�ju��ؚ�pLW��ev�������1�ov��ӌ����q�a��u�O�z��]��}^Z�l���>�_�6j���6}&����l������� -�[���9FcE �����@�g�7w�����:e4�EP���������e���B;.�x�·sBڅ��R5�r��ٌ:鍣Ó�	[+!��g�VÞ��W^xb� ��Av)_d���扡in�,��)�t=�9ioa��Y0H7*a��n��al\��mI��;�G�7JyB��6h���rN⬗�:OF�{������� P����(b1T����ʅ@�RL�~�4Tv���*�Q�E�je�7ߵ�D�J��}��w�\/ʹi�0�4cȟn~�v�rܙ�4B�����;����Lit��k�׮g�����G�?�+뱏i�R'�ީm켬\w]������$r�ժ��GX�5
<�=×	jV�]�>���1�$i�~��O3����D!vY6
\�[2��)�{��6~7;3K��;
�ə���]�ʉ�O1�h��C.D^���F�{���l�!F���ojT���y�R�#{'�^xR�ǞH�_7�BK����:3�҃����u7����:�����dEh�w�\��O��йЄΨ%��������y�w��z���i���\���v)�~j�`s�z-oG�Ն6�����;�K�e��G��)M����[�+�M�A9y��t��u�c�����9���/��(��w;.�i���c�O�|��k�\݆��D�I��
�A���4� N '�+��г��k gtm۱�1y�0���L�_��N�U+~�$֧�to�<����8@f}٠k�zئ=�C_�O���Jc���^�n�l��GHp�����-\�g�tJ>�s�6Sg���+�?�Ia��2�ZXW��/~��V¨r�g�����iJ]��j(ӹ�,ad�IҌ���;��Qt�V����r���� `z@k�$�s��@|�4"�Q�>����[7wn^���K��Ƀ_���}i�u�^G`� �)'���v�5	�)/��h����_���gM����߼9Ҡ��h�][�d�{�d�6S�f��=A���
.���.������f�{?w�Z%��@���F�y|���vR����U��N�,
���Z�%d��	��i����L��zV�Ő&��?'̔�����fgw�N�C��.DՆkߥ/��~�xh]�􁤰�@n�42:�7C��	�w�k�J����K�?1����7��[��*_t4t8�
0�B��
�貹�C��ϭԫ2Ȋ��f��&�n�xo�w ���@>G���RC�tE�˗�Gچ5�~����T�E��x$H*!�6'�t��#.�����n���m۩�0j!)��vx�b����aR��z,���(A3�4bp>Ik�K�Y�޻�6�a�r[!$��an����F���Hm7���~�I
m�!�A(�*��؎�*XujN���v1 �N����5���w.\j�˹6WM;t���1�T^�?h�����{M�Y1�nfKc:��y8G(:"�'���{�&��Უy��y����Tx#�������T�@�d�����+o���8�p!��O]���8�e���Ʉ�4f�u�c �l�iM#���ރ���)mis���x)�NO�(zo��Jт%Z�Ͷb7!n7��U����~W�Sڎ���*7}<-۫�0n�!J��#$�H�ȆA-�nm(�s^֍j+�M��&�F?�}�T����chc�y�p{��
�ʀ��A��&������M���a���w�I�pe�t�v�yґ��K�`o���<�pé��ę�&s���0�Kwr[�8C�ݬ�{�����H�nJ��׉㵍kX$��0:�&���|��!:�̴�ae��r��7i�մg �N��#|-:l!G6Bgj:)u@ ���RXf�Z�;�0f	M�3eP��.lJ��G�/%V詿.p��_q����O�p���D�jK��}���&�IK�+�I��gy8�����۳��\��=�֠���`il��w����k= q�����]���j�@��f�	|)�c�o�J���K�]�?-�𮎼z��ES7pO;�]�~��l�:����pA�/�U4!�ai�6�~�Mխ��;���цt�(3�`�s�, smtS������a�so����>�Z,�H�w<Og�s���N� ?�?�,B3����iȇ��n�	KxPO&`�:�*g׹d8�O�F���-t���ǲ�f|O���~�g�����i_�XG��A�oe0�޻m��av�(�h�R���}�f$�lgɄ���hE?I6�<gO�ʳ�㪻�4}���"��w�߁�	����8�����҂��.mhϣ�g�cA l��వ��c���_�Z���j�w�'�A����?�8����,��yl�l��r���	�4��	}�Au1n���	` ��>*�΀�HF��?}R'V%%��Ϧ�*?91�"��`d�iu෍��*5h#�m�o(D}��k�g}"S�`Sy�Y�S<?���j#_[���������i_��j>�m{�}P�	����W\ڏ3g/��tٔd��W�<}��"L�!6���0�ʭ���o�~# {��R��|h������e�w<50��=ΌD����ō�˃G{�= FC�t����$?3��Q/c�TV*#��Uje�	V� �2޽�g!A�������0�b��!��MlOB˅4��[@P�o�K��-ݒ�Y`#���ҶkQ���l�O��FNP��`�:�J�Xb1X�^nG�����E���)4u�i���-:��m������Jsy�\6g�n��S��]���������� ���}��{��'�c�8vu�ix�����iQ�s��C�`�d6�E�0>Π��-HWG(�>�/��Tw�y��1�i���"!U�W�z*�X j��(���6��.6rў��l��g�S��&g�@���<W�I*"�!������������4�	����
`�~�����7�S�قa\��.M{�-!�L�9D��o�����3��t��LrQ�-͙V�i:s8^x�ױ��42U��N���'#)�n��p:��)�7=��Ʉ��+rG�Gא48���)�<����M��uՁ�����|~�/S�^�4���/��?�<��0:�-��$z����K糍c�����2��hB%�O�@�=I���(|��j��5P��*슧��&�Frux+�+�vPf��#�����$n%����>����-b�=��9���G�v�Uo�Ԭ�.N��T���c͚��F�A�ޱl��o��~���xR[ɽx~>|}Q�ga
�Vf%��-��1L@Uek:� v�.0M�޼q{�f3�:�*�T��5%Jp�f@ؚ�Ǔ�ّ*�@�@�P<���1ڝc�������efO�_a���)}�j�&!����E�(?h��/A��&}.�SC��U�h	�pG�6-#V�TKIȫw��Y_H�8�g�����i�����k�]�W��O&rτ�iw1L�����ë�sn7�>��E��޻�Vm/�g��-��cv��^�E�7�'G�i�~�g�����~<��4�+�����9�Ka��F�-���H!AjN��*vz�
�w;��:(i�Lt�	C�:�I0�����1#�*	n��'���Kg`")��U��H�
��c?��_�u��	�H�|S��^�PB3�7�>��4buڴ'�J%H���0$|�c% ���]�A5�L��֢D8U�/��8C�Q�NGLД�"N:�i� &A3�g��ҡ0i�2�69�~Z��|�T�54+����Gb�F�X	RK竱�Q��(���d+��8�-���V�,�,�W���iN>�,�H��k�g��M�L���0�xS�`e�@p�0fd�pZ˄gLdh����#iP��>>|�t�Ǵ��L+��mg��T�Z�Vs��0?���c҅O��2[����C����m뒐Ӓ^S�GL�(5����U�V����su:��tl.s3���2՜o:��0��(�Ց��rR����\��Z��h�Ы��Žr.��P�e�'wtf���oS��W�3� ��%�?�k��4�^�[g)=��Y���9k4�?ڍ��)HD:�s˨A�X���*�L�Kug�d�)��O��1h�Ľ��H�ޢ�TZP�U{�U��s)\�Vt2u7n�8�RzG8 ;&ļ�<λ�ҁ�A�
?��yBO��(_o���<������hN��1q�̣�����9]�Q�]i�����1	o�yx]1�QX�K~���-�� ��sï�3�m��~�����&��Za���T�f�A��=m�lk���p"���=&7��p}���E���V�s�
z�$�ؔA�6��ުw��؉����h��]1�W)�a��2�Mϲ�z��Ar��n�6�WM�Zɼ��!���������{�}ӳ��/�ș����:��4�϶ߛ��˴�w�Z��&��&�#x���γ�l�6x�;�i�7���� ��K8y�]��In�����k)���W�7�+�����ߡ���uёv�	��錿���p�"�A��.�v�TB(1�+�B�I��w+^w�� �DM�W��j�x]���И|JV�J _����8>ÿ�ˋy�� ���d'�y��IդШ���6A|���n���ϻ�#��O�&X}�[BX�(zL �	m�HB�������vyo����_������*�y��WI���A;#��%/��$��5��;�8���`����?�-��XL�maU>��R�e�$��Ժ	W�����u��zg���PB�~+#Z�Ƹ<Th#�ʮ3\+:4�:�vT
re�B���f��O�PA7�R޶�?����j{	�#�����MF"���7��8���-�vh�U�� ��B��-<�����7o�mJH:�&��%Α��j i�j�'�d��+{x�dS�y�B]�3e׽�݊X;<� �C?[Z���X	0�X��*S�L��
ɧ�A>�NԘǐ�fo��2�+C�4i	OʯA/�ji�d-��ԉμSex��<�_��	�G:W���~��˝��t�����ѧ�H���Ma��b��f��o2����Ke������^}�0��� �o�	��&�
1���c��}C[��Q��1�Aw�!,�W�5q���,�^o�.���ɣ;�`��oÐ|�@���-x:����T�D�b$XK�6`1 �+4F��0_�y�υ�c���1�@+�[�����p����TL�7��ͪ=�����SAp���R(#�R��$系�e}�_�
;�S��p��h�ķx*�|0�.��w|�+�,�Ƽ���s,���^ln~}[
�+%��-��Ӟ'����>)t (�6K�n��s�0k5X�~f�c�9��[͡�Uq11���a�����8'�@HYn�����^ �X|H���)���~�?����%���Q���b?ݼ�Y�ݝ_�("[�?���H\��c�H`��9S��ie�A�ì�[]1b���݂�k��n��,Pnxʟ�^�f8�����`����΃��G���[�t���rkмg��N?�������vUV�g�xxzع��--w6wvXoʞ�ӟ��!��2�TU�m?���a�R���  v�َ�5������{�~� �"�_��O	a��{�>��v����_KQp<���4UA[)o}%�������"|�o�����a�-��Q�b���EA�{4x��^�E.x�6����T]�c��P����Nh���`�Ǽ~�����
8���J�CݎMп���;iKc��
��L�F�fm�ך�`��T}�~6w����|i�H"1ɐb���>�MSh�i�Qų4F�&��H�(&	9Ң�Qw�ro� 
������.��<��gyҷ��%�Sy �JK�����k��q*�gP$B��B��g5#fQS��vQl��6�����ӏttVe�{����d�<�X�����j%-�n��Uք��v��Kc-`XZ��y��(�Nf���ǝF�����U2?Z_����#^����3	,�tF	��ͪȃ: ���Mc��1�0�X�X�{	D8�u�u\n�Tބ�$�7��1�+?�tyo���T[��Ȅ�#C�(*<�2Dm��K~�!xWNb9Te�c�:�Q�/#cZ����+�c�q��ݘ�tZ���h��?:�0VYb�hT��!�~l��˦��Sy�j�X�)4��Fe���^сŸ6
�v4##�(��b hr����L�1��f�Y���c%T#|�;d�7@���ʡJ,IV������J�2n�����T>�m�6�aj�K���3�F���~�����N��)�z���1�5�O�4z緕{�48��f�ތ��}ۖ�6��t���=-�3�~?���*�A�*�a*�A �6���򊫣7�����$C��
���rlL�+�����kp5�T�jk!�\����:����=/A��[�w����E;��M���\]���g#�o�)��(���sIi,!��u?�ػʊo����jM[V��v���c�?��i�P����oW���n	��V�rL�����7��6.���`�ƅ�43�Z�n��iWOgq�T��a�up�jũ�lꌫ�᫽�ҐNŞ�[��_e#�􄖹�x�֌�����|;�A"\�� �7��7��R.���F�'ꔣ�<��=���I�ʧ���"�6�x�v���f>e�F?�L��[x6��7�jÃ��QWd5��d+v;M� ڴ��MH�!����d������w��<��!���Gئ�U�<)
V儴�pGr<O{Y��c�-��t���B��c^�4D%�E����_0���^Ӧ���d�h������c�-9tl���!��m�D�i���� [��w��߇1@y��)��i2.�Gx�brJM��);���Kx$��1N=-�G�LR��"�̩2p\���jۜn���,���Iz׷�0w���` �\*�`�2N�u��c[Pįt�QwﻂT����$�y��t|�� r��"�*�@ND7D|��h��Z�b�T�� ^��X�����	�Fy#|i�:�)��������V�ݏFM�%��eK^-�ՠ�;�%���P��~��V�u�KN]ms���h[��u,+����`����Ν�wG�Y��������F_~̗ @�=�M �ަuZ{+v���9L���βy�Vd��W>u�,�4ϳ��j�J���ҕ7A�Ȇ �!
1I�fvh���œ��%�Y:|�p���?���ow�]�$M�}c�ې�ہ��n��mb{x�Wf�mgBRW�@��2�����<l��O��٭N���|Vbz�D	bc����!��v��SCAh��1z�y'�����RJG��Nis���T:��(0i�I������}�\�(�@��y"����s���E�	a�G��&vDF"�pg����u�\
(%N�|~�\���t=��k���>�W�x�(�U�C>}�Uoоr"?�U;+l+q��pEXmz1)g��t�X�5�B�lu�ޅ۷����v�q�Sg{�-���hk�`��Y�>j��vh+8+�.A�o�q�Q�%�S��*���u3p��\]
�Q瀵ŋ�s�eL$�昗�M�yF'�T6s
2��n����^��^&�~&̦Kۼ[q�����wHS*�{�����}��ø�w����T�9�W�n��% ���I<l���Ē��~�vU��A�F�zݔ{ם�=+��֑����m����i�W�s��lk�\�X]]/�U~��S��3}�6m=��D/�0RE�P�0����r�*���W֧o�
#�� �}�� ���.�*��yϜ�����F_>ˠ>��[� ܾqs\�}��;w�e�hh��ԥx���x��/�N�6%9B�2�7�9�+݋�B�����]�{�T�&�}�F����´Š>l���������hO{10_x*��e2��ģŏM;ÓB����Y�D��re?����0��i�= �;��'V[���ɘ�L�W�O���)�Տm(���F>q�����X���zlh�;�]qz���I?��@P�5DM��Kё�fZ��y���W��,M��$��"��&/�q)�f	�[-Cʛ���|]�%?�Pa�HB�t\@ \�:�������2�y^`NX��>kth��
�K������&�`���ԬP*c5`�{0!��So$��{��<�F%=9k�-���_F�j�&�ɻd�`'ܬ���e7�Ԃљ��4s�J��˦1����ɹ'��--���+JN����C�|�Ҩ����|�����	k	F~�%	{�U^lc�ˍ-���K��/L�hA���b�E3E0Tƀ
���ᙽ���4�W�q�t�X��8�LS:�~JKjd�d0u�X��z�mx�E�6/���!*�0�Am��$�I�3����@��1w�!���w�Bd����p6O {����.ėo̪�ܫ��Uxp�V�I��k��I�v��*��Թ�j���d��������+��j�=���`ŷ��P��v7�Տ+��	U�G�F��:w��o"L&���
^yv�N��{�ƅ�A��`�,$��g 1�K#�y7Hܼ����v�� rNٺ_�i���휐,���P|hi�څ�1�<{W�Isn�J;W6�e �5w��a�6bT��x-��)���+xfLx�1�h��}�hw��`!����d��6���{^�PV�%lՖ����h�=U��--�݂m�3����v{l���p&�@x�����s_;��n
��
?����e���@�
������Ww�}4{��X�SQdW��yL�5��,7pz�X�+�2��W�%�O��M�V	��G�S��'��ЋF�<�����%h�ʛɃN�EuG z�U�" YLt��/m�sz�����/�ն���A�Ӧ��J�c[N�8x/:lڈP�/7:����^�ҙ�ŀ�EQ~����h*�_�	%��D��[����̆ܯ�ՠ�]����:\a�e;)0��B�Bi�n����HX��	��G�Zy�v*�S����J���h��ާ5��*[;��?~�R�n��絳 �#ͮ|���+|��v� I��^����nЈ�<��غ�y^*n@��-L��w)������!Ѧ�!����A���sS:�mN�Gh-�L�N8t�(YYA3�P)ы9�<,�V5�f�Ѫ=�+�#I� YE%A�&�Z�3�%�}h��۷��fd�r
TƟ] �lr��|��nS��l������+l�v��A\�$h�B'N���K����L��4j�����y�F3� �P:n3�L����De[��ѫ�z�Mm�[9�IgK�� Q�U~<������_5zޔ���CR����_e�~�e�g��*ɀ`��MUf��&a�Aڢ[7n&@͍Å��iر���J��_���ӡ��K�������z{�ȹ��E��
0�y4����4��&��-:#�aJ��Ӝ�n�������U��tmM=�;�߹p6��i8!��!���
�G9�u2�F���d��P���]��W��E�Hɇ]���	�ƎWc�)<Y���,m���LY*�����}B�G�v�ک��M��B2k�^̕���#���"t/na��bK�`'��eE�
ӹI��ţݐYK9�LkU��Y������-&`�����,�{���ʤ��AJ@��+h�%>�.�m���^>�����/�#�Iv5�����B����p�ǁ�ɫo&��Ul!ד7ّyQ4 ��\z�[�b��7j��i�����2�=���g�ܺZ������x�C�O���ν+700��|?Զ�C�X���1��Y�[���}tԱp:���
�d�����y���w}�؍)5�)$,���X�M�lk:S��Y�#<S�C������~|�<E��Ei|�P���C�8|���W������8�����S:R5h!�׾�N�;����g� ��^���^ƙev��[EN��<�X�N�vu���3�h��ڵ]3��?�S�l���/;w~��z9J��%̃	�Y���d�<��˶c{�t����Z)� >y�kOږz��;�t�C�� �s���|�����^�y��t��j{����K>@CS��PC��
1H�>�w{�Y�[x$�3��ڴ|l�Z+_}��x����?�?bL�[�iqʱ��?5}z,;63 O�6e.���H�g�E{{�:���f0�T����B�Sx�J�*���9�!=�,%�`C��q�o�8���/�T��\®�j��H��c�-	5��k�Y�E�¯tѮ۰�#�ΙI��������t����5�)�Q����2���6��1��!�J�C[g��^��(~�  @ IDAT���1�؛��f�MF�l�c^EQ�a�!v�>�|��u{������n�o�m�M�Ib�����t��9�0�:�����aY�ƽ �F����0��
V��+�c.�ދ������?x ��4�i�� ֱ���~U�gc�"x.��FK�n]�`�-œ<�-;�>�?~Z�D@'�T}�����򬃯��6
S֓	jW.�����ۑ_.�e�#	�u`���\U�.��߹�s���ݲ����r[_|5��r>�5RZ�wo�%�gs����w��m�]�\�;S3}X�@�5n?�W�����t��y���KPv���*-���WL߽Eh8?�m��[�=�ȿ09TG=?ݬ�j��B��Z=����#��ٟт|l}�6RŚ��7�����6�%F=ږ!�o|d�aϔ@�ݭ�Kq�bĐ$lð�E/�!���t:f�Ѭp��R�4W^��W<��/1��Z�}L�ۥ�`�Fˤ`��E�'��Ar|oZ�*a���L&'
���>�i�3�?�z�W��`VÓ$�W9�y4��ٰ�a���&��_Rak�C�fp�IO���{e5}�o�UvN��ʄ��@�'<�����6�\�ݴ�nDƄA~c#�7X���$�c� ��u���e�'��,	�K���z���2��C����i�-V��'ZU����&�M"�o��I/MO%,�+��6��lwu��A2���	ϥ1�"_P�8$�0SK�v���Yp±ic҄neh�g�������!�������9-�Ր|#��	k_����|����K�ÃF�T�S�)�lڿ���WJ��h���t�@;\|��(������a�c���y�o˴�<�#�K��o�O�H�~uu�)U4z1���39�R4i�f��>��u��*��;ȩ�ү�lP|��s�b�-x��{��0�T�T�� i��)��/������}�N�45�\�=r�d��.�$��p�M��|T���������@�m&��M�@	��N9zv��iCu}BG΋��g~��]q�n�A�����+����M��0�Hc�q��=ϓ�o����>��]Oa�'�Fx���`"��d�f�V��LF"NX��U���n4c�H�ӡi�f�Q���:�*p5M�4�򎢭��ƾ�>A�R�����/� b!pPX�L-����4�ӈ�F �༼)�(-�\��|��1P��|����m�%eG���Z%J3Z�cA�JfF�!�{i1e�pp�T	K��e�D�Sv�Gt��F�4L�4@��$�����L63�]�����m���P��4J���bS;���H���K5Գ	{���<9ƫ4`�5�o��M�C��.b�i.|�$���
^�NƸ�#��WmC�����\meLG� _�2u���˂׍�^�H	|[��a�U|�l��ѾH�v�d������k�H��܎�OOXe�!�4ziҢ�cuF����Y�D�:~Z��]a��*�A燶H������1��641xC�����d�NS�� �������B�F "Pkcq�a�*�uL�ݙNc�j�I7�2� \��3�� ��V}Gyc���P/�|���u\dtu?�PWr����޴�n��j����j�PD�|�P���kK�A��bD:Zԓ�ulj��8��᧲aMxFiL��OV��͟o�Iv��'~���ay�6@`�=�a�T���+_�;ФU_���^:��n�-M8�>�l,~ <]x;�=�LVYGP�݇�h��W"SmS�����E�:�i�7�ɛ b,�NBx ��{�Β�u�+Ak�V�����'��*nZo�ڛ��Yܱ:a�>.��>�d@
���>Ԗ��J��:`Z��70�����q�Z���i+(ў2(�U�V����M��i�-��eN���!�������fl�h����fPQ��|���eM�+/%��|��#��p6Bw��̀wiS[y�"�\6�W�^7GcV"�
��u���4J 4c`���2g�n(^��҇����4Wf[��#��?�5:�=�ybC�4�g0��;�^Nş��mS!����W[	j� �گҌ $�ةhV���h�7��>y�:�yww��b?��8*OI/C��H��{!�˧h�vPQ�3���ʷ���"���c�=���^Y�[D�������C�����G�S�h����%z�M����������{��X���\��捼�-����]�SQ���uoX|��o�Ń� ��/]!��9ܯSE���"�Fw�x�rM>갚�������!�AT�<W���4����^'~��|�{^׉?� V���0��4��v��pݜ����|[��d:l!_ׁi��_��x`�c�V��r� 8>¯�0:�)X��=�a���~3�0��c���K����o/�����7�U��Cƀ^gdo�ȇMc^I(��U��6f��������)[]��:E��j �S��^n������9k����Γܹ���#4�?���i�.�m#�a�W�T��{���mB+cD_~���-&�	��IM���e[���T��c�5r�U�Z�򯢳Z8��� uP�^J �*\�a�	21�]�����	'xp�@ͫB1��d+�)�B���9*d�p,�J��3��}Ls��O��3Z������`)�_��� 7x)F�:�Jm�G�uC�b�	�G{���H��T�����w�B1:��7�it����X{��+��.sH��j�`�f��W�>����y7>-,w�~�v��箃���
�KQ�x����(�f�g��c�2j3����C�3`��19�4�iw�{G�0ڏ��Yv_ ��L4`��NxY]�&����>iDs$��C�W=�r��n�^��$4y�f�o���]ؖ��^ډAu��������`1$�yoJ��~�����2(^��yu������&<��G�@W�ܭs�@S�_z�-�x��%[/��Y)����n���e�=+hk`Gڥ#�9,2m\?P�h���{���MW�y�٪�4����aB:A���V�h�N4%y���v��8��M�+��{ �er� �"��?s�\8�6��*ky���J񱃓�G����q~������r�r�v>�NfӸ����m���Nf@�Z�h������'�
?��Ƴq~�:0@50�����w�~2[a����c8�ߘ T��](á��%~� ��M��Wn_r��5��3���T//r��$W�Z4`��W�w�ڂ3�8_�dA_�gr�vr�ԾTξ��Iy]k��Q���AȄq��և­W�n�����ލo�G�~_����M�ɠw�y=�z&0���z?e�5��{��U͵v���JpOCQ�a���L��B��z��J�轕WT�=��o2p��{�cd:��4�p���1O�S�~�WzFϛw¬�Fw��=f�i��o��w]��U�y.	�)��J�4�0`��z9�V�[����C�}�X���sȯ�kt���)<�f��0}r��d�O���w����RM9L��T�т��i�����|���i3��z�1��������{��ǐ8�a��������i9��2��	��x� �������ۍ�Ĭާ���~�����_��bf�N�^bVX�߫	[6J�5.�o�f'�i<�SL ���\޵�ӝ��O;?�n!B�V{r�&}d�QayXi365ڱ��Y�j��2��V�SG���ʹ���;z#���5vn����B���6�t����G5	'Fs����(�]�Fi'���ZaT�3�%\� NpM��Ү�#�����t*T�~g �8�A�r�7�ǎ����~S˳z-���f���?45*_]Y�η)���;��縥I���b�L#���F���Fb����ws]8�.X(�ɵ�6�r�Xm|�O�Z�1�e��.Z~�7u���ђ0��~&�b�����Q}�z�����|w����%�KS5m잆�/l�@Q�2�|�B�<ǖ���5���&m���n�A��4�Wi2�8GU���3��^�[���T�M��Y� �ޣ3����BP �Qف��O8Z�W�������+[�	
;S�-N�H�W�՛[�
��V�|�Y�8	���:WS�Z��*��!`�Yko5���Y>��J~���K��om�p{	vc�|��=~<�f����{��(@n�$(F(�'���	`K����
�޲�i�{��Fc��I�e��A 4�|���rSq��stL<��Ks�����"�L�|2>f.�/��
9�?�=��M�Z�ʂ�C��vi��wA�~8��m��Ғ�l�ӽ{/v�����u;;�������M	�_�i�Չ<!x4�]�).P���U�֝�;?ݸ�s�N��'�~��M-'�Vc�-zl���`V����M��X�����u/a��`��ŋ;'�l��<}4���3@?�e?�g��_4��,!ϬJ3��ܽW]W�m���J�}D'���t������RWS�'8�6�J�j�~:ț�Y�uL�	�}��~=��	���c��o_O>�9x���7����{��Se��ʡ|���&�T����ޅ�m:�_�Ҩ��)�V\T��3�ㅄ�3�rkD�X[bd>̼J�=@��w 9�r�̲F ̌����zNqKc��!Kg����$U�3a˯�t�ϳB�����f�᷏ �2`��f���&��� ��{��c��z�'!�C��7�斢�o���a��yʶ�HsT�bu@���T��q��H�ZW�A};��ei@F/O�F1�<iJ�0����3�ҽUay��g�jkP	����yy�<O�|�ޣ1f���QZ�׭p�/��E+o����L~w�ɗWs������Q�N���c	+�9�4��ڈ�Ȍn��,��͟w�z-��i��f���7EJs89k�VQ���n*	�z����8&�6aȶS
?�4ߥ���}��Y�x��eU��cH�T����b�c�!Y���)GP����֎����1sK�-5������;�-ӦL;
/*��;v"1�����k��D��˦$�v W��w�c�f8H�3^���Nt�h}���^�A���Ш��hߊSV��0ъfB�b4j(�u�+��6iH8�h���1o���j�<��ubR�s�`�����UL�tu`�G(���:�Y׆��G|>����	�/�\O���/�0M㪼\��M�L{1ӈSΥQ��x�t���'�M��9Npt0|fʆl���^�#����{8�I�#p�P�������lK}����!H4]�;Z� �،}Qth�"z1-�������D�J�.�Ht<+��<2\��iw��X<�
�j�P��9�XL��h��8B椸�Ug4ܦq���a�6>� n6L'p�n_W_��9�W���:h�����V7�`p��&�WQ��6�x?q��]��[��e�PXH�˩z��:�����������+ߑ4^�����p��6g����V�{�B��9hG��譶�C�$�3���ӧvay��V\�3Z/}���#�O��x"ܢ�m�h�g�۷��Q6��o�s>m�n,�X�w�o�^����f���.��9�Kh%<T�i/:��SՕ�ּ���������MX5a;s���д3��pR���\�q78>D��,'�U'�++e �g%i}J,X�^���GX��X�*pG"#.I�q��OM��3��D�c�;���ud���n��ϡ��Vf���2�gh�g�)�f��k��yl�
�=OAW=D��g����P������ԁ��uD�f�2D����f)�<*�A�!�^W�V�H�I�e^wLa��N��h�a���M���
U����S��G�6�|�GH�bA�Ŋ'�:�ݪ����D�����Fܥ�'�[QJ3E }�@s��rӻ���F%�t&�\�*<�)#+�i#Wӆ��-�6Mw���;?��Vۻ$�$\�8�eL����;�)</����|ԏ��ux�Qf��Sɋ�RN�V9�6�F�#��}�JF+�;��8F�zf̞��;�L�_�۟F�p��?w��4��P6S���u|�15SCF�����t����?�T��3�^>�v�s��kM�b���C��:����?od�Kjy�G������q�~*��Y���*��I*�O�p��[/�'Ԉ�������z$G9�s��%|KP�������:�/._�m
c���}���EX����/:�੾m`Ξ���[թe�����y.:��`w�&�!��N�w&�6�o����J*�R�c��\�:)ndo�C�ǈ�i���}�'�5_q��(�=Ѓ���� �Nb4��5��9�ƁW��~���e�0iF��L�V��Ѝ�����b��)�n���Bq�+�� ����DS;'��/�N'����j��ժ�˗���iQ��6yw.���;�L�O�o�ܹ~�f��fZ��!;����M,ە̕7��(�0}�����4h�8�%̜
.�\���ʗ9�<�9�
�h�Y���U�^g�VD�h9���.[#J�=i%��Y�w?Qwh��2�5v�O18��hy?�*�0�|��;_e����'�k|�Ց���Gi��-x*7����zֆʁPE�y�4�/���]�=������l�@a��7��/�����~��Ë�pe���ai�넚������L�?J�2��K˜U�a^	���˟���{w�/$�)�hR�/A�F�Ϩ�0\?l�拦K����3�8HV������ o�1���VD/Z������3gf��{3H<��O�"�	�f=�=������V\��5��0�>
>��0<:{д����k;�nފ�Z,�:��ڊ#��mud&�Њ,Fz�`5�c�	�'o���>�UB���T�L��sh	}��7�VzN��!���&h�><�D�B�!7����1�3-7�v%|��c�;>?�y��3��SaJ{��>+P?x����~���q���ӿ��3��k񐕾��������6��?�g����c�	��MJ��j8�sӏ����iTX@�W�
���J��A+���o8������`�ςl�1ڭ ؾ��o�y%�y�q�Q�A��@��w�&���ÿ���´��Mz�	��~௿�"v6Z�'/�5��`��B����x0H#Ne|U)F-F�Sȭ��	E����K��sک���<m?����K�4���K���a+j�d��u�y~N�|R�}f��*��	w��(�:�Y��?����ֽj�i��m�t$͝�`�t?�`y=aO�d���FOU�y��3@\���9шL�|� ��_v�����=x�|�PO�X��ڍ����?������<H�@0�|��~�?_hlh������R�J ��`Si��P�x�\l}�ؘ6.:��Ai]H��Er��坯�.���U�1�s�%2�`��k4XR�m	M�ѻ��|��L y�(�;�Aa4�6���a�}�}�ɫ��/�dגSIڋpMh��Y>O��� ���-ݾ��ت<��-�K���U0Ug�~³zU=!!́QJo�U6�*�� ��v(�a�S�_���֮N�N�W��ٓ�̷�뗇����ܝ�I6)1u���5:dOėxBX�^�ę��I�-� PXq���~:�����)Z�%�������;7�nܸ1��8��_��E�$|X� ��Y��ݛ@+�	�!-��R��	����������_�|��Ŧkh�� �Dt���wUG$/x�jg_[�B��Me��N۹���>Osh{mr��jg@	���0������v�߷�ۯ�$�4��7�2-�L��Eh�s��6����<�ax�WՑIn��g2Y�Ê6�����G�d2����=׾�a4�5���������]q@~�/`��^<���J�+T	����B�Ⱥz��fl���u��rI��� .4�I��&��G�5����q��lfzdwWW����U�>�`u� o�<'�������`\[dP�fx�g߰x@9����R�{>}�X1y&#�a�Y嗑>��D�e���yo�n �.O��ޕ��J@�2�{�4�����c<>�hJj�_�N��0�����;�a�g]�h���x��'X1Z�-2��Ϛ�eL3�e��'s�Ou������PNǶ�˶+�Dm�Ff�H.DS�|�gjvy��0����cX����׽�cr����Qmh4}1�i�OeX�W�1���0L���n�{�e�b�-O�����*@�kZ��B���5H���⏼]ۯ��]lt��]�s�?_�����Q��)�I��'�%\���'Ѷ�~Tf�4d�v��=��J/�*3���v �JT��A��nӖj���	%l�.��̓�<����gjz_q/J?�/4I(����uj��5-M�6M}s�r�8�)OFP5�!��f�y��(�?��h�Q{g�	|��(�7��9�$�ZBI��f!�gO�:�Wȹx�zJ>�w��%f���^Hී|}���F�N�?����/4ݰ;��J;����SОc�y���_�$<��Z���^7V��y�L�n����?����}ߦ��q%��<Sk�Da��BxO<J�Hy�^2Ώd�q�����ۼTo�39n�4�f���/aHQ$��p����˩��?|�
W9C!#^���9�#	��1���zc��C�)Zx��C7��o�|{���n)��~���_��|s���f+Gˍ�>�����@6> 0�4�`$WGa�`�n�Y��z��_ڌ��G ;9a���pa����'�E�w����擻է��T^ � �Љ��BmB��T���E��ݏ?�)��5c�i-RB��y��}k��zv��r������'M�����q�S�~{^:m�R�@���D7��W7�o^��&�"�1��/2G[/ߚngh���>��}�x��I�G�m��_���$��&��
`�a}'�����_��6��TL�� E,��iw������S-ӆ�x�׀O�1/��?Sg�Rl<Nz�B[|xۊ���kW�zD�ǎ�J���1z*���O���b�1�Oh+b�Q�|N3vRf<�b���ں�)Ɂ_?�k-���|r���]�ڏ^�wB��@���д�Y ;٣�C�OpM��5`V2��@�@.l���net����5ؠ��`dL�Q"OJ}@\.�TJoj�f��$��%��79�@��g	��1薞X¡��#'jd�
b'�ɷU(�F�ɗ�����H�Mm��Z�H��Ƹ���lB�Wj*x�������kx�����1�f|��m���F����߮�[z�6ӈ6�D�{,�!Z�m�<<�fޟ�߭��d�|���C���w#C�˕��ԋ�Ϡ���o[l�w1��K�L�Cm+�!`�ӷ�˖!��_�o=<X(���G�p_�����K��+!Gy�� ?�D��{td"�d/��_�B��l��;`t���T�_����H�������<{��_�hͺt���'Ճ1���-m<,}m��}ny���_��wt���K�r���F*���i�9W5�Q���GŻk2�̣%�uM����_�D/��	�pe��)㯚�#%�Z�쾗�k~Idx��;x׫�`�^O���݋@Fy#�0�y�$�C�[����z���`c�#Є7�9��2rt?7����b�Μ�4�X3��B3���mjpb44G�A���q��>#.�}�b��啣��7o��q�,%�{�l̃T@�Q��sy;x�x����LѴO�Q�Ĺ�g9x��Ff�5Z�����\ޱ�� �֌��M/���\}��Yjb�8_��ѭs��ձ�(���'I�c��%,
YH�c��!Fa�-�pq�8�*���LWax�C|�N��c�(�uie��|�;'���J�����O7_������pr���9�uB��l�\tA���Cߞ{�_�;̃���]�.%S��X�8U���T�yF���AS%�TZQJ�vm"�Me�?��fj���gI8%�8b�m�/���Π��^��vy}&Xv���Hw�aT�|y�	#��yyI�y`�OF�7� \��ݩ� ��=}t9Z��׶㰂�g���{���{����RD�{m3
_?{/n>��ZFE7�f:�6����;|�j룇7�S���}��+�9GJş腢:�-n�N�f�0��SI�u-_��L��^^^�ky�.�.��'8I�9S�&�p�g���)�J<�����?ǖ�-V�=�� 5ϩEO<Qh�w�Lër������ѣ��/YL�t�Ӕ #����Y����1j¯Xm�]�)���bLyO"�vxXL�ز�<z5�h��!��6]/���;}�=�������9��u�R����9�xPf9� �6������R��۾c��WB&�6h<��@��Ȥ��%c��A��7��������,�a�M�k�+�Y�?x�e+ؗa/qI�ՃW�}�Eg������t���ͫ�wV�EF&�$/���hچ��`f��d��t�~����́��fB��m��Gl��&?y�6�ć�uS�m���b:^���{4$D�_��t�D�pi+�ms1�'ܐ���k�e���=�}x\rG�U��ܮ�{n�}��y��A�)�_4�K})[����oa����d�-��n�h{ۚI�mbf��D�X<��I)Hv�#O\�00�, =�c��V�[��w�
�[-Kq[�*a�*o%�8�v�y��z�߯�������?]��]��w�#�EP��K��3��7O���g;�A���S� �2)�p�qO��0-�L8�y���Υ((s�fx��;�U��)�}�ݜ�>(���I�s��Ȼľ`	�<izP �8�qB�u�0a˛����7�yx�t��ɀ��w��5��@N�#!�uض��\�j��w�<���x� E:#���Օ�:�&X��|EtD�z(��(㦐��qS(�ք�({�$A}���-V�n4���,�*t�#��C;ڿk�r/�x�|#�٭��"C��\���N�*�M6�V��`Yz��ns�(A��ي���:}���gM��h��6�%�[�p}�r{�ȓ�&E&�D��o�J��F�s<P��@[F� ��q�!��`C���l�W}u�TK��~����<��,v��'��ᵸ@�Y|2��}K�-�9�4��Ϳ��7�5zV�oR��b��5���pa���O���YJɡ���Ы����\�LQX�Rg@�~�|�?WZTb*�i����"�G��}a RpM��c�~Vb��T�q1t6�w�5\������'����<�N1���y{�R�>O�$�g�Jo�����iJhV�&sC��5pp`�)Kp��}jZ����ڴ�����tH>����/�������ԷK�E�/��lq�6�OJ���j�]�p@���f����I�\�?^�� �I7m�c~�yX�E���>(n���;��yM2�3��'��o�s�U�c7�^~����|��m&����� ��{�:�&�"�h׮�d�SfC�xa�V�����B�uy�g>[��h��c���'����8W��6���b�d'�k�z�`"B�s�"m�7��2O��R61jP8f��X��Y�2nN��Ұ>�V��'��*� 6�n�6�#���4��z�gy�}�@ �|`�i�i����C�l�� #�V|Xr�LTV~�����xy���Ѣ_3b���n��9!`j:n��d�/��l�o���Eg�0v/O!~���3�M�/��W� ��#0�y��^�#\'�R�ӟ҃��L'�V5�~U��n��5?Ý*ݥ����H(ӵ�S�������k�(V��o@�ڛ��s~��/}͓d��ݴ���'j&ä�f��\�5<DCDS���{8ԴW�UXw�{w�X�� ^ߞ��nRl��T�r�M�;����:�bWf�*�k[c��<m[ul���	�׼I6m�����]���J��B�)B�Ԍ��<<=�p��FeD�x�<F�Ý�D�Uf7���o��:��x�URźp�i�O�K˖�ӀQRȘ@x�����8ϓ�P<����?� X8`�"�/�%���^��b�܄\��	�J�!8� ��n�)��:����>+�#ax:�t��@���4��,�єʤ��w�Ш��g�؈n� ����^��k{y�C2����h?#2�)�*�|u�J3�>6L醥�J�6�r�`��?�(c�J�+vN��}�9�6�DSV�
He������uv����d��'�x֞;ʰq�xBj�tD�O�{��I)>��9������L[B�6}g��{f��H3�w೪͡�V�ݹ}�i�כ{�Ӵ�	���L�&ĕv����_�C�c�WG}����8�D3���d���3|nbJx+�2�A�S�<�Ե�!F�`�m���v��
�n�9
���]>k�-�ʘ�ج������
�]�	]�#l��~x8����6U}:o ��L�G�<aSz<U�m����������:ʓr|hz*�/�����z���͟���+���i�!}3�����Fɻ |^f��P�M����>�t�݀?�fm�Y��=~�3�{|�$��̓	��6D6��cfߖN����Tޖ?l���%����V@3��>�ys���>X�¼k�Qi+^����a�8]Z}C�n��Ctb|zj*�$��Lk7	730�Ao���f�u�!���=I޸x��ج��9�f�� ��YA�S��n�䓓���/C�`#��<S��=v��z������j@;9$Gp����fO�F��M������d�l��@��Q�:�쌸!t�F'�<�_�kv���V�8�w��	��ň
ox��P�����n ���7�N�Oިd��l�O�sM#��3F+5����e]1���0;n���h�v�2�1���9���{��y�n��������� @�Ko�5E�-��M֝�ҭk.S�ht���4���ݿ�4x��+�2��iKw��ךg�{8�@��.$W�۬.��J[�AV7���=l�j��6����6�.��1�7S�?��O�}v�>"�	�����x����U��{�����_ɕХ��N�*�z�ᓈ���a�>�_�#�0��R@ҏ�/ǰ!A�R�DHX�ARc�e%O���~�h���ڌ!�RƅV����R����a� 1��J9�s������ń�e��v`����dP^��e���͹��/O6�ڦ�ε:�~.�"�� 3��Ƙ�훂S�f�^J��O�
�dȝ����֨��̀:[�"�X�;[�TzFӢ9���E#�g�adF��R����c��a���;1?�=�k�`�@#Ɣ��b���/�S�yʸ~y���_~�i���}#şf���d�¦���/B�ᴼ`���
��x#EY�(>�n�`tQ�f��:y2�~�6�!#������[�_Ʊi"�3��Ϝx�
c8�n�)���׮o�g�\�z~s�ӏS�/�'Oj���<��IFȷ焅a���ʪ�>�Zߖ���'ɃF�渲��,1mb!V�Q�OX����)D;�;�A|����3^;��2� �y���Qf6�|����:l�5��D�;b����������В�qa�q^���[{_�jY�&�p��0�=�u�zg�f�l����`_=�8�?}���f���w̶�-lx�W�8�S��u�}���ӏ������?�.��FrV�(��ۣ���\c����A��8�E��J�����a�&a*�74�%����
��m����7�Z'4���;�1�r�����Q�v7_�~+z7��!��3D[��!y<��<@�uE�2�5ݤ����c�1��X�����M=)���x�����>�p�;d_����U�)���&a}�G���M����s�^!�:#�혊\+� �2����/dș�f`0��d�b�q6��{�R�k}U7,Z�������~�:y��V4�3e�ׇ������|��|48�?H#]g��۷o�0��v��p.g��.�\izR����e��W���Ͷ������+��hς�"���/N�cM��^ܛ�0m�N�p��x˙��h�kt���(c��1\�z��g���$�=�����S!���1�כ���y.�.?��~�m[El��7���җ.���VoA���p��rx���u\�����9����T�?�5�۩o3�Tfϼ��̵Һ]���i��y��#�d�⧐mޑK��e�V2�fD1��s̲�iΔ:mG��u��P���*8Lyܳ^u�3��*�w
��(ت���s�J:���
������a�Y���	9��i3ݘa4�O,�|��b

`��)��&�b$�:�)�a�pu*�#ή>āb����h�7�l]Ye@Z���� �(�����M�8*��i'�S5�Ck<i)�Y����Q8�;�l7���Z#h���>V�P�?��%ħ���9
�38��Qp�D��2z3!S��z����Dm+�V\�-7�u^���2��Ap�~���|��������iyyK��q#c����w��>`z�������a`K�����]���N���MW�C{5Y᪓{3]Y_���N��S�c���1G�٤�uF�ǵ�â�/6u� ��Ȱ$��v��٦��l�Us�`�鳺jVnU?��Y��f*,츅��>eȣ�3� tU��Z�8�me��<�ԸiB8���ϊ:��QD�3S�`b�B�Jm��������?}���4w�����fV�x6�r��3�"� ��|��8-�d��L��~�X�� ���O�t$����}�̃�����m9���3��6E�/9�S��R�����x/g=�u�X�y��}��v��9>�yUȝ8-^M��Ҕ�L�#�U��㬭}Ტ8,��	�#q��j�Q�T֯�2�g,�o�T<Pt˒G�Q5c��+W�Qk�����?�(\f�Af��VM��{p?9z.�T�5%#�U�~�Z��- D\�ZT�𧚴�T���d{�/�-<Ss텕�kpS�08]��[|W�{|(Dƻ#��̣�-/���p�s��t�C:�*P�e�-�a%��Q4�s�脷�Wx�=ئ?�����p�AĻ�)>���䓏;���LG��D��E�1��+y�Zq}��\�����̰0ba"�vi^ؙ���]`�-y��]���3{���ihwfVJck���'e��JE[$m�v�Aк]�w���QT�������)m����>�Qjw/��2V�y<Ԩx�(����|j������z���O�f��U���DK�^5���	����a������6�lk��ߊ/�gS�	J���I���KC�y�Ub7Q��p:e}��OZ�{�ց���ɶ�u�|L�_���~bJF�ߨr�.��5*�5O��"깑������nt��M��0|U����F8���鼘܂�	�r���6R�� ka�ڟ1�eo��S)�`�o%���d0�i�V�`���Gk�{��y�b�`�鳯�,�N1���eF�	��+�x��,$��)����ťm�c�7�a�&͢TX�J!F@�����ʀˈ#��08��h�O0p�yVc��'�gy$֨�q��0��Xg[ax&�z��+�l\��u����ۿ�|Sགྷ�Ÿ9��q+G�������8��ה�1:2���4���ߵ�o�׽X1����y �j����|�a��:Σ���~�8�X2u7¶2�bCJ����M�Ψό�/>�eb���<�km�q��6^��;J%\�r���+9��ݷ_n����1�,g�m/(�X��
ǝ�|�K�����}
n��
6bd�6�8����b��_�@<O�N�IlZ�7�NYB��ቡC��y�����g�����Ym�#�J^=�G+b�E�[��r ��;fy,|ܷ8e�P?��J�m�3�$�2�M/<[���0��+O��틶�g�!����
�O�j]u���J���>���zo�d�=�K����z�{�k�\yd��6hA����)�޹��L=�+5߃e��Ë�)��}�1}�;�s<����Җ����o��� H@���*>�@�9����x�woۚ$<h q�<*��|��oݸ\Lc��N����0X�����9*�4�����h��  @ IDAT�wp�2���\�)�# ]����+�X�����C�5T�|<P��\�z'���Y�	&��G�N��j!`Tp2�fɎ�	G�l�/p?�\�4�:�զzC��͓����������ͥV�����~���o�n�;M�PGK��P/��͍A�o��"�>�|W<سd�Qq�����uͰ���~�h��q���sB���juo��>��MGY�3���
��,��J�����P׎�w�%ݽ����� {��k%T���q鶹޿�b*���D8>s/��~ɖ]�e���>�3#��ww�\'Wh�7��J�#��X�jA�U-=��*Ku��-����;i��R�k5���]���.���LY�)�*���^ݱ
W���&�v%����PM�հVy+�Jٽ6��D>�l%�w뽗��PT��Ċr(�a��v��j��ۨ�Z^HXp�8����/����Q�O[6/v���`�1N��;�(��)
E|�^���9#�	�A �0@ĂR�<�w�):ֹ�y����d��5"���tJh�oB&�m�a����#��O�&3�����
܄����w���ic�AG���Q\�@����5A�#'6F���×z��5R��wv?�yi�����b*ro:�����ƍ+�o��������YE����Dm�k#U��y�����_l���HZ���/5e\�;�����6�[9h׵�W-J��y������lA�_���������������d3[x�0^�7V��1-J�����;s�c��#�駟��ܗ�Ϯ��l8�Ԟ�Lą�%�h|����1,�C6�FJ�c|���[�P�Qb����%��L��?��`.��8�������.��g4ϖ������5�rV�:@�U��14���7��P�˛���?u5�t�yԞS��J�N�e�2`�����)C���Ws�n�n�	��AuƜ����6O��>2-g���#�wnr A.0��3��Y�{?S;�	���?�C���w�<��,u���p �E�����6�rFD�("�tӔ~k��{��h8Е;3!��q���M��3���Y��Ex=�\��A�6��i�d���$ ��\<����!��D�;������?�et\on�}�V�M�X�⪡��g�����l!Ӱ轜z���'�{��k���e����'li{hU��[������j���2�N1`ЄO�5�^�* �y�x��pc�齏7���7�����3y�l�Z�<M����'�\{nݼ���ۯCE}�����~i�m�hW�nL��{��هmڴ����ʛ�MjR8�4o�	KCo��tXߙI�;Y���e0��uy�7�w�Hm�k�4�d`���Xx_y�]Wϫk�<����Zɷ���tJ[2c���Hm�X��9� �B��'9A1�5B�q�(����Q�0z#�-+dU���� `���j�W�t���x�P�fҲ�1�Li@���;���D<[L/"�+k���yW���3�#C�S׀Lh(s�<����C�Q����#�����wM�����Yp�$�ؐ�އ�7��_�����|��,V��>�1��7�����
��K���i.Ӈ{�m�
|}��s�2��c\W�(�BD�I3�>8%��t�P��w�}��X��	�Qp�`�WR�:lj�]��Âp.���8ő��bC�H���bpu{~�6�	��U���tJ2%�&Ak
m��邴��z��6�%8F��fSz	��)�_�n����\^G���u���H*u�4�E��a�zP��/72�v�BޡK*mk��!^ǹ�V���v�̓pr�ux��i��J���"��Q<���W_5���Z8�G��{\����24�������g��l�}�����F�+8�i����Jx�u����>��+�V�ٛ	ܪB"�f@��&�1(�+m-��g�2��3��w��2:���>�1��V~�;�&[��ŗon�ꘆt�:ŧO�U�L{U�x�hN�a�/�j���Fޒ��~�]�����:�
/��(�0Ė��V��F�����ԣ8�y�Z�C9p�'�C���I�����1�2f;���N]��x�L�1��
���ƣ�6�����	#l?�s6�웊��[����lt�cS[��r�pL��{���%���j'��� ӵS����}��o�U��ڮO������A�1^�%[�h�f��d*kg��}A�V�� j\swG<LŔ�V�]�w2�g<���g�5���nS�+�UI~�j���]߾z������kM�����ͷ_��w��͵�~��׎�`�r;"	�vl�$��2�O��#~2,�U�a6��D��ePb��JrȔ8=b��X(��=U���Hl��$��n��2��-��2�����Q�ޖ����~4L���lF�{dW�����5x4�z���������2���,�{�i������ĥU�->
�����7���Ō��<��o����͛tQ��!b�@G�Ay N��\\����P�������8'$�O��o'9O�<Y!�������p�U=?Ӛ)[^�ÿ�u���<Ꙃ�oԢ��O��%o��=3�X�]�5@Q�_򳲬ܮ��UՔ�A�zyEW�-�C@LV߫�!+���Ҝ�پ�_��8�!�q;e�w�n�q*j{! ����o�秄~,���=sޓ~��^�{�X� ,c�P�W�{���AA��ގ�@�l�/a�n)�����f�.�3N�Bߔ��^�Zv>�u��?�}��?�|�ɭ��c���2_�h�p.�w��X�a�����`���/t�⢲�"�� �w׷�<�rz���QA�)3#�D�[�<�H�Ry�r֏�ň�zG�T��x4�x��ƪ�2r�3�����d�Z�F�LգogS|/K�R1J6�n+�l�*H���ʹr��"pהe�ᇏ�4�-(8#d 0䢰�*�����hJ�����pJ��k�v�
��4��<{ګ�����IF e�m�
�]�ڃ�H��4I�_������ǈb$�i���ە�~J�*���}�1t�cȦ)� h�(�1@޴��/3%�b�b����\��0mA���!�zAށ{x[���wS��
��~g�:�]��h<8x�~���ٛ˹�V�	��Q�2b0hP��l9,��cd|�ñ�)m4��2E���ġ��FD�%��ffL���G������Yjm�Ϫ�bF�������"$o� �Մ�$�`�Z[�>M�;���<�;��b�r���k ��#�;eo�����};�@?��>���"{T�P�j��ch��⁤�M��ys6��c�y�\�;�a��B�2�.ğw2Vx4�wv���2�+����Ȟ��0�����V-�p���T}���Pn�~����P�NV�U�Qz�ut
�P��y�F[=m���Z�w!ژ��㷣�������7����?�3�����|�uq�7���U��R�k�+�8W����<ԝ���ǳG�(ӆ�du0�/f����	1S��ٙ Co���@)e�P�oMw�Z�Y���a�f��4%Rn ����c�u/��b�&�yT�ض�����w�������_�������N�����Xp ��\<�'*y��q�V"���|��Y�h�a����"��Q�~F������f�E���� �U��eQAy��|h��g����Ȇ��Wt��lM�+cʩO8�7k�R�k�9�y����=������U���p��zhk�[i�<|VfY���x�Y����x
i�`��=�Ap����)���Iӈ2NfH���}L��C��(�Rla�v����'`��^T�2�3��ۻ>Sn���&Yo��`H�f˲ʑ��tҮ��=���M!��u�{ɶ�D�)<�k�U���*@W�p#pAܽʆ���xc��X�ը�)���\��ۿ�zs/ϗ3�޾zMaz�T�1�'o����73j�|��w?X;�W�@H���ft!�7Bw4Ќ6�Fѩ�H��j'�H1ȵ���PWރeġ�[�92i;���:0��>��7u��Π1����|=�����07�E�������hۊY& �!m�Ja}��������{��4�U�y�]��M�7mLi%�KlӋW�n~����������0%_kAn�� /֩�W�-`��7B�C�֭mꙷ���u	he ��?f3�`����)�?�����݌�k�������N��;6�*�<���P�ESź�ze1E���/ރ��uG�����y��]-I�3�?�8���|o[%����p|*#�F�]�M|�ݟ��&��X7ĭ�8��l� k0�Ś>	�- ����n��G־a���)5�7c�9�U;Ű��EC��,�'�њK�u�N��V=����l	;��dʸ�3��r�G�6�1���'O���Z�b�DK�w�o�Ih�V0�֪Rm��+���x��I���f���V�b�3A��2��<#�El��c��jO�0�#�}
e���(ka#���JU�~��x/�'���6�~5[�<����%F|+����_���͗_|ٖ�R�y{k��~�fxI^%��>�j��t?�ё=p0ӊ�|�Mx��pj�n\K�SdeQ�Ξ�K��FC�A��F�����s
o^�1l����.��M���_6=������K0�'�~����ӧ�O�9M!9u-ϐ){�|���^kSj�ઘ~��ۊ8�{}f�-��	��$4z�ZE�Ó�����@�:f�r�tM�i��ƀ�Ry�����7��^�=�%�Y[���d�����gj��;>���曯�<���&��ԬZ�:���~�ϟ�����#:r?��&�n60�&��W�|P��ڦ"+�Ľ������y�� 
�����[��~�k���݉��-m��'��5����5�W�����De��]�����e��/�Oրs�|����iɖz���g�����0�꜑qhx Qg��7�����lpjէ�@?8 �*�D���j*Z�����d���R������2���z�S�zX]S�*l=[�laX�U\X��V�JYC1ǖd���L�2���²m㶘�����)�G��j���b��:��8�0�*��D���ʒ��|z�N�v�o��T�s1��Ò7���2�]7�b:Ҫ�_�W�{��ۺ.�؁��`$azj�"\mDp&���Վ�
	.OB(���<yK�`9L�0���q��t�p���6Ÿ����o�X}�	����O^n��3�~���:��c��j�H#Ճ���HxW&��3p�Q����ʦDv�����⥃�u�Z̝���Fj��(��� d���2��wc׾y���Ӈ�����P<F�W2�o4}ȳt�vQ��2��T?���X"�bђ�/X�.�N�9����Z�C"��?�p����:8��Qe���=���jcu�#A���2�V�LKJ�J��0[�w�d��AA�?���l�� c��F-�_����3�O����.��vS!�I�7����q���9酲)S�<���wS�ԃf��5�W���{�N:�f�r���=R�Lx�*R��n��z
���U��>fإ4?.C�e�q���w��D��_�g�մ[c�l�W�7_���f�0zy�{�]+0�b1+]{�/�1�s5�c�_j����/��n�����>��(�{�L�>[G��	���^�E�̨y�&��A)I�e�Ҭ)T}a ����B#f_�0F�v36�0�w�I�gd��;�6.M�D׻>c������<__3(�ЄO����AN�mۄ������F�,>:���b��-��������T���`��˟a��������2r#Z������6j�\�ĵ���a��s�����%_O�q�T�{0���=T�c�����VE+w�����/g@ipe:X�����p��6����F�m>aС=�~��_��b����x.�O��O�32���.��KC���>[��,���3��=s�V��	j\~�l!�vU6���Xhp�Z8\i�w�Өwh�7�\F�ރ�/����I���O���J_�;g�^�9�\=&>��~��څo�$m�fl!<��M�G0�%��Xl��Y���m��Qgi� �~����2v����<�v��Q_*^� ����<5~�8o�.��1o9R��_%��qی+żU���ӏ	
�{�%�;� ��S嶮)Ӏm�)�2g1}���S$9Bv��u��b�~g$�ه	�<(�����/����2�UEÖ��F��7�kJ�����[����7��ß6Oۥ~�ciN]��MP�"<j�U�ʔen�=ӦV���W��4j�1����L�:�� a� n;7�>0Zt���l,�vB5��+:@iwL�@f�:����?����լ���:H����^7gv�f�Ssc}��r��&e���ި������'�q�f�b+���~ؿ�Y�y�}���Q�h�Bt^�1�D��]��"��?LL�XuEIR<sďX��A�2���;eP]����k�xc�V4>�ɔH=�?�V��OE;�Z�^x�^����R_n)R������EƋ��J�wF��fu�>�J���" �1[mԿ㍁�-o����f`����p��B.�r�7�0���qG�[Z;?�-�U��^���m����qe���*��mh�i<ʳ5�sX��GGFO��҇7�[��O�֦s�.���|q�_��~d���gq��j���g�߾}g�>i�ͻ�0�j��k��o���8}�z��b������?�����Hn3��b��8��N�yt�69��Y���a��;�qZ�1��7ښ�z^��;m������-{�Q~C��M}���O1[�mU�K<!/��b�ӣ���@e�d����J܂�������bag����ǧ��Z�y�f�6m�ѦȂ��d� �W��l3ݛ!l�,����֤,y"����7_[��Rl�yX`�l��F�V�̫߯T��B&2v�%�Ԋ��e�ch:�F����4�\����]�ȭW�?D;IЁ�v?��6ɠ�o}�v��3��#�>��ng�~4�C�+ӡ�>4��(,^ߑ��1��^�M0��s$Ѡ�Tog����Ykc���ywӿ��g�9uM���4�#�Wm�<���Dr&Z���][��<33�}`�N;�F�;�w&��cm`���Z}C��f��P�?b�e�����^8���ɱ�0��)[��=1`��7�$�[{Է`��q��w��5 ��;�Jhy��juN��� ʬ�X�K�s�cr�s�ͤY��~���"<%�j��A�\*y��m���G`Wxy�)
�G��g���b�y�b��ۣ�p���K`��
������h���J�=b��S��1��.u����	�ۭ���2*n������B���x�Y��W�J���l���f��U��m�Q�q;��օ1�"4�S(K G��럒�߿w�Eq�+⍹	MH��s_���+��9Ic��b��2�7�%�wG��b�$�v�{�0��m�z����*79Ak�ϯ[6�E��Θ3ʿ�a�6| ~�q�e� cц�Gee|9ļ�;��A�Iަ9������D
�iӍ�`�T�r��a���[��ՆQ�1|h��HQ�3��i%���\K�`K<��&C~x�%d��l�XA{1�'e.��R�傅�bQq�`s��y���d�1XP+oݪ�P|�gd¢{};���ti��U&<�D-C���k�(ǵ*�Qk�A]c��^��z}1Z�2(������NT��Ag�mh���,�ģ��B0�����R9p�m` ߬��=7�������9�Ǵ��N>`@O�1�iQv�_lct5��������X�7���ڹhe�)��_�����~\l�s�)��9�<�3�?�{���O7�m꘷�⃷)��l�|\��Zɻ���%�E
�f�F����[PP����/�Q�"3�#��q'5������ϳ�"ȯ$:�h�J�^�j?��$۬�.��b�v�Z������C��U�V�j��A��T�����/-/���J/7H�{���>��|�AĠx����f�np�yG�B���E�e�j����ә��g��Vd��G��M>i��׈�f��xn�S!�Kكx����w?�+]w�6������Aw�I����H���S]ޓ�g�fVu��bY�G����{�̩\;c�	G#w��h4�X��6���Qd�����2��]c���������⹶��홫+M	)�򐯮�U9�_�#�a�&��Pe�4���8*�:�+�����_N9��4@` �p7�;�qig�A�`�����4�+�_�1�"��O8��{)�r�H8���~�M�na�MY�,��`�Q2�����F�,��^����,N�G�����oa���Z@���������e�+�Bt�|�!�F`�Qh��R��1Ų;o�i(�YҊC�B�XHB�3���Z������p{-b
~�:����3:���
g��F�r�i���/�}�}k��X�Եh:`/F#�W	:�?7�����]i���3Fas��/|���s��r�F�E^���$Fc��*I�m&&��oNw8khC2ީ��]bP#���Hކ��pKɜ?f��:��_��L�d�� �At�=!Bƚ���ښ������?��4�� ~3�΍��_�èUL������	�#E�`8�@�O@X�5�)���~��"qW��m����=��������� ���%�a
my����ٯ�	#��A�̈́3�͵�E�?_�#=�|��E2kЀ���;���a�Eo`Z����n0՟�N��(h�MO+�Vw���C`���r�+p�
��iW��S�ј���Mig(y�����b����R��>s�O�2<g �W�����iK�F��������f��(}���fqk_~i���]HF�.��&�P�0^g@<}�x��O?o���?�G����bp�}V�Q�bD���uJ<}���y�o��>������ߏѳ����^l�ʛ`�x��o��ߖM���j�(��=2�)W���'kWr[��	+�Ō�j�������E�Y�tnI�����tcH�{	�Mݔ��.��)y�n޸:<TW�0�/T��&�x���7CN#�޴@�E�%��"������ڔ��b��皭O�wz��^��773�����<�l����I�=����&/�s].m��O�M:��@��D����W3���Z|����1����_��y�1�AM�������i�=��S�$��?.���$#����	֯��S�ItKH����b�a}M@?�(k���r@�,�����q:s@���&��4]��h`bd�44!��Ķ����2l������kc�=����bPO�0��@�tt���	qyE�b���QZ
Rm���xFv�������8�|�v��C��N������"'�M֋�N�L�h*2�W[�f�O�u��Z&E�����x=�vS9�g�l#�{W���1����l'$8�}�Te������DFyƛW�!�Je�L����׌�/q6:i�qt����[��i�T��ݯ�`+�}{�ӨՈEX��"�!�R���Z�aP`ϧ�J�Q<w<�Ǡ��稜� J�=�!��Oi �a5B�7����m/���������JC$6_�`�e�I�r�"�C���ѯ\�*%���j��6����4A�+�(�%���)��s�|�K��;�ol����X��?8~ޑ9	�\a�9k�� �⤳7f��yԣ��u�a�J�Ι����3��p��q�CF�sCT̘ ��v�#bt>�B�+�npg:���-���cϭ�+&�x��-ϖ�R�+1sb`xg��VOZ�>�*�׃Q�w)qt��ӌ��}([te�5a��^LX�n�)���~F�0,�	N�Դ�[��R�hp��m<C���M�7���U���[�F8w���<�@�l���`z��l��w����(�����[w6�4�Ȟ�Pb �z��X�]=ک|m�����[�[�I�5�����nf$}��m{��W3Y��́��V���\���q#�m��6L�{c���w����p}��'��λ wSIy�W�ow|{��(~�'�����a��ַ>	��~ݟ��L_}������j�{�8�'O;�+Z�y�m ��/a+]���xq2~��q���٫��Τ��{γ����j<��KM�\,<�
O�(#���.�m2k�%�I��kx��2A�d�
���5pX��š�[�=�����S��^�˸~����x�9�'Zz,�6�"�w�
'�MǾ�䈧Of�}� ���=�F/��x���F����"�F,C��q^��`
�7����3ui��h�y��{8�)v�݀}�t����z�\���S_T�(�`_�\UR�1ps�3y_�ã��`�X���!V������Sϼ�^r��SFT��,Y�k�խK�3����4`K��5)>�ڞ�Z��L=��n�@_�<��*�o���㡯��߇�G���F=���A_��n>��vΓ1vz3�����dP�2a��~�\��it���YHI���E����� �Tn��~j0�g&,��^+� O�]�z'���rOgX��?4=�EO�ܻ>�?����fh���y����;Y�$HӶ��Mg���n�0ft���:��c����	��aiT����K^=I��C}j�ி;Ɯ^�R�Ww��=�c�o=WR�cdH_s��'d���g��PTfOeD�DBj���q{-�>��Q"#,t�!�c��wXI�w��\�����C���JTj�u��J��&�3ju��ٸ�\B��9��1�U'ehؽ���g��~���сq)�:�������wrb�\~�\L��ö[���oǅĦ�[�wԴ�Ayr��©F���GB#���픊~��5k�ڥ�W���`���q��N��5�a$�s�$�<�c��ٌ4�������)�ZV���hƈ��;��F�:`%�*�J�� �m �Ӆ�^�$728n$�g�� #ǹ������p6��'��n�&N�:�n/�J=*�LY�j�Q*��UhA�{�.#�U������<��]�,��o��a�8��F�/�C��|���w��Cyc�����4���LJ�t��_�>3�ǲ�"R<�?�Zu��+4n�Ji͎�^$c�p� ��r���>W���*�����6c$3���d�Z���Q�{�����K��Ű�c�����O�N�~��zqC/_ݮ[y<AuO ~}F�(��g�2��⍑=�A>�e
�!M���aft|�0���!xә��Z,"���'el�&��Aw��x~���cz�:�:��B���M����A�6×��8�5<O̊.�q������~�=�.��v���ί|����K�C��j(k|�sƤ��v�����0!ؗ*��G��!�s�&�a�',��n�p��f=���9V��z��E3�U�\�Vn��ⳏ;B�����
0=j�� gT�	ߏ=���K���ӧ5/�8̸�`���ن1�z��n��ڣ-���������S���,yp����-} 񰯯�:��W��]��ɒ��>��Ҍ�Q\��Y�5��}��i��H�-�&�0l��cD�7��iΓ9�C� 9�ԩgm35_>�M��:�x<q��?2-��t�v�wv����A}}�eh��e萝QH� &�� bx߻�c즳�'��t�+P��NXr�cT�Yڐ��׏�E��N�0-���������6�S_;/9{�U��u���iv3P�q��P[����9��o��W��O���~�N���@�ϲ�lG�|4�Vr잘��7�ŵmZ��.9�L�)єLJ����2���a�1|x]ۃ����:�l�^	�5J��U8��$( �zX/�\���qO����������ژ!��!�F��~���Mͮr��oD�+��m����<�l� 6
����=�A�X�X�#�QR�_�D�H���>��۸��mA��͎|)l�v�PLc*�T%a%&�-�0SB�pS#�a�� �s� �3�#���?��\W�uؕ�&��G{N%�Q�R��1�0iJ���.�ј�<�	GF�k��k��[�-��5�� .w�@)����A��C(��kD��~F��#8*@�B#�K�>o)z]8�`b�8�l6���V,b���}4K�����=@���u�iD��gmZ���\p�n�?{1�����eFy�%��B����P[������X�(��o*���M# p  ��W|Tѧ��-�T�J��=���/"�ĴcTq���4U;ޤL����)��r���9cK;�;�c�i�L��M����T̸��O�ݝ��zyyLA��z��.���]n�����o<:���.=�>��^꧋s���f�^l[�� L�<q�Q&���(.]�\]�9���:
�3ؙ����RTr����cM�c��s c����&����{g����+[JT^��]�h�����ߴڡ�V�kc��il��=ܢ+�Jٌ"��޳x}�/�vz�&�pb�|.F�póe��M�}����t}w��=�1�sEk��+x���Ll1��>�����%Nep�c����,��Q4�s� s$��
.��o3������d���΢x��
d����=H�|�=�0\����zs�g��k�ȸ	3I����m�V��J�P�l�\t#X��1m��}�g�\=D����	u�e�!�$O}�S��b�c�y��g��p��%����O�C�pm#e�39��2F'56ŷ��?�+�m����l��2� C)Át���Es@3�/8�FT	 @连� U:<ֳ�q�������ս#�F��=�M���m�Q�����wo+��x4{�R5>��y���W�pӋ�bv�͑+u���b�����T���]}�����gl�s�Ѻ�`+�@!�Gw���s����RD�ds�Rf���3T<�м_y�l��b<̨8S��j�^Dz�D�N��">�Q4hY#G���_�d)��b�*�|���c�;�!�vC��Mbt?FXߘpV7D����:�}E�ǀ�]1��3�2*��T�dl1�����腓��O��l����h�'x"���,x�/<���"ң�#�\�'�k�UH��u��g��lZ�Uj�p��c^�e0(&�w���R�T�CL�Z'bMR�#�����P.�s���,�F&I��E����+Y$��K%��+�P��e��VJE��=�Ẑ�u��x	��q�jv�'|��j�x��	ϋŵ1���m9�'vn���_�����ϴk��v5-{��O�/�����mmA�	E������[��ٳ'y�ڊ"�>��y���22N�0�"YSY�~̓�Cz�èu�7f�l���ڙ���K���u����Fsk�0<D��0Y�)Z�$>�"��?)��"&\�d �׷|���G���r�խ V�MH�k����X$�c��2zϢ��K�&$_tΝs&�\��W�0^+��0Cz��tZeuۙ���#"V���ų1h�����3h�!/O ��է��Q~��+'Ė��e��B�Sdz��d�ve�`�	������pxԿ��
��ӻ2��2P��2��K��@�]\�W�WJ�L�W�ų%؟�O<�.��w�+f���:**�2����:�9x�	�⊟;��;he�����_v�w1�[yԊ��;�}d����LY�W��5�Z���J,����<�%|� x1��ZX0'1���o�5;Z������^s��ap��ݻwG])�GA�Ds���X聁f�~���
�G�g�k;��I�56�gbB1|S�2��D�c4�|��ړY=�h�|c�����{��@.�Ģ1��"��F�A�x���pM�:o��=���`�
z#\���k<�A�\��Q�N����S�g�>C<>ݏa�2~���</>i���wM�h�'��tfP[=}a��(�.:�>y	�S��o\��I
f�������l�Nm���'��`��'���w��M��c���4
;�';��t�w����c�B�W[0�K�ϥ�H�9���H���>~�y��B:�8_q�-�8_<�s��o_��������5�y�܅�M�F�k�����x;�x�%�Ϻ�C����/��}�{hL��[�򒋻g����t�Vh�����"h�m�	3��uX`���(#/�i2��-���	^� p?������ә�����P��;�Է{�"���� �k�E<;U�	�È$�ȢFm2B:bx*��!����*�z��g�!���є�B�Jz�;0�:�;A�c�י'�l�<��x7#�����vg	�m���oM�=o��#mX���?���G��d�ix��t���eb��>�ѱ�H8��~8�6�#x�1ɧ1����n�$,5�ֽ6I���9N8$�������7�v	���0c(�iX�	�ک���O���� BOj��A����x��w�Ey!�/5�p� `#P�.Rt~_o�uZ=%���͒sK��g%.d������=��џ��lL�FP��ay���9mCq]���髌��}7�t���v�8�\����N�����c���U�n��;��a�i������J(���/S����u���m��.��/lap�R��F旯<w���`��=|2F�`�=蜻��`� oj|�.4rb���eLw��3SR^��|�/��%��t�:a�`�fq5�S��GAV7�u��g�F����YY)Q�%!Vy���w���U�g��?*�D�㍔6d�҂�D�΄�L��sp���
�"��<JH� �K;%�,R�����=��V
��g�N�Qt��և�X�h��_F+�?}�����kZ5��y��9�}��3����c�8&��89={#^�S��"#������������)���	ς͖%`tX5�!�Dgz4����M�����~Sx��OӔa���|�T�f���V[���_�@L�S¶C*k?�C"�P����?����x����o�DSɺ�7<=�*��Og��`�	��ωz�V<���<:�����.tݠ���-M��V�:K��ㅓ����9��$'EY�Cvf��5Pmx���{��w]R��_�>�(_O���U_���i#�o2=�V�SI�6>�OWZ�jk� K����j����!�?�^!0`	�x�Dc쪫<�r��*�S=,T� �M��Dd�&�Λ<�����5Y���r�:�O�o�'X$_�G6�3<�5'�G���ni`1Ӡ/�w���МD���;6.��ٌ�W��c4���}�z��d���"^���v�wA>���c�������~x|��}�j#����	Mc���J�s�2�jh�s����ms&���w�x� #�H***%b��wZ�c����^�S1���-5w�_��-�C�/"�l�|�L�u�v�����i
ď�{|��o�0Gk����>ވ� C섄b�T�qS`X���:b%�TS�D�Je�)���mt�Ë��>����ھ}�Z��F�=g�ɯ.��b���~����c5�� �X��q�kgx�����:c��`O��T������w��~s��OU��A�(�~*�����t�ѩ�^4��;���>=�9l������~��8��O�Av}�q�&h��Z?#����|6�cdo��U��}����^� {^$��?˕<��ǔAy�4z"Nׯ�"xވ�aA����<�"$h(a��p��m���.j���?U=�����(���??l��������S�bHfˁ�@SA˘�q+��<#b)^��;S�M�`:���	eP>��'N��i��)>t�3���n4�*�B�[�s�
OQ/� �/σʥP{�yqY;)8�qW�}��V�ğ�fo&t�B�XجxJ�,�iZH;R�=���@�k�gd8HXȌ��Of�qou�Nr@�,OUJ;�`0�ᾛ�#�K8� #���BH�ߥ�BQ��i�L����?E֪*i�ȶm�6�%  @ IDAT��â�B���I|�)����:�3�W�z�A_�)�t���SߚB+·��Yy�l<�O�x�7����m��A�;b�`�x!�U��O?=��h<M��ã_<�8/g�Woj���{�m�,�)[��m������qs?���(h�`Ĵ��Ĩ��A+�E{ћo�S��$�����_f����8t���o����޽�ɬN�EĪ�G���h��I�1
m)A��Fb�&�񚼨�X��0:I��3n���tr�\�^�)������@�96DΒ��|3m��q����������o�g��|d���$�+o<O6I�6C�2�NZY�R��#�d���`���&ތ�����U���@�>�� ��Q_�3F�c�xrdse�E9*���hǆ���;wnvR�W�v{�{�����N_�0�C��`M�^�����ǨP9�d���<���ŋ����o�>M�=x��sxw������HV������L}.R��9��ỗ�qO�9o�4�Iw%2��<��.S�>d&��@�������fQ.o��jh���fgޭvN`�crC]��`\1�`�1F��_kʱ��S��_�;exW���#�\2Q\��6=v��:�]��^�;�,^Cj�����(��!F����5��
@���Cp�,e�����r����V�#���Y���c����wUM9ʢ<���~L.�9cۄ��e�-���27"{�,9�.g�N��yĬd#�"2g
��~�}�#^�]�-B��챋�yb�+�`��1 A`�k�LP8ؙ\��`����Aڸ�։F0�F�g��
Sխ�1@9ᤏ����X���>8v�~�"	#\iT<%�S�����1�0��$�Ā�Za�aT��Q6�u�W��M�H	mp�f��߆�s�H@�������)m��M,�@g�b90��������V�v3C^��.����S���	5f����v�ה��6^���cl�xA�e ��pe$΋e
�����
��N6S�4�7�dJ記����X��ݶ�jV����Ԭ����Q&�;�׽�2�2�ԧ�5@��Ν����_�?�zyY�M�[�m�oz4�7�'��ד��t��l�)�~#��\8PƓB����8xƨ
f��������/�{�_4��i�)��������g`� u^���3xX�{���o�__����m����"�]�e����x��/�]A�A9�R�q�kSx~}�7�a
��������^�i:<z4����8n�y8�����lp����
�o�O��y����yM���΄�7����Q�˳Muo )���ށ}�1����:6�a�\���>��x�3m�IuA �c����-�*����b�R�#[�#wUO_)�!i0�pӅpnq���gy��C�M��О� sJ/��L�g�U�ܦ��"��9�HV�?<�P�	;R��gz���v�rh�3�! �}�9��J��3h�x����~��^��6�^�d&��NV�d8\�"�ꓒҮ���N����I�������#�)7x?��/�#�t�����ʮ��)��VSG4�?Gy�b����4��~/c��#E�gm���虾M)2@l�d��`@����p
o��pv?O���xkj��{�:~�������.m��@�{4$H�+o�rp�| �Jw�?R߶rr>�Bz>Lg��Xͺ �<�����m�<Q��'Oҍ�A�C� �z��v6z�k� K���\p����d����=��[rqktW�¶(?�I~Р._4�q�����c4�Z����ސ�zVV�"�f�T`vz�S����m{)e�&!@��ح��@��W���M �z]��j�� W~U�Ӑ0���%�d�)��	b��^ֱ3��t���Զ�Uz)���*��L����.n�QMI8���'��7)�>"�[��A��8w;��N��݈�/��t�,7�O`���[�Y�5�v%d����}@�	)U�q��52���i+�)Sy�2���d
��8��b�,zx)͌?����`<aZ�F��X�a��b2A<A���x���`��ʰ�~`
W;#���3JM�G�Vb�'%2<������Z�_IA���H�j�ia}�c)
�>�d1W~=��o)i1�0fe��#��~�o�V�ѷ[��|�'|j���V�ӟ�'g�_�أ+Ckv���[�*��N0�x����s{���.>6�\�OwA�a���ٖ �R�Ѻ�̖PG�p��!�*�Z���� �5�0}����߂�P���Y]\��Ҏ� �$��3���)'�#X�a�Hax��~���t?B*�F��q��]�'=#��W�Nù��L���~Wⴝ��n����W���|�|]hb�j�<��!:U��2#/*���H���;m�'Huj;�ªVqH���Xr����������U�D��tes�Sntw��'����y�s�Gd�����@�w��î<���?ˠ	�b�G/vh7+ѣ�aeA�0���>��kOy��GN:9�-�5X�0O|Z4qx�����U��ř�m�i ������[p�	;�â�X��b�g��w�3\�'dPBx��x�3Tj�s�G�X�i����U�7Z+,�NG}�m��A(�>?I������.����4[}�� �Ed�F1&ч~��bߞ�j��g�J��&ܛ�e|0<Є��1�����pI�����{dUx�́���0df�$
�z�Ȉ�|Sy�&��@�]����@k�t�_}�����b�1��$�1���Vn������ýR������~|G�R��5�*��jZ����|{�����i�����%�} E%�K#�}<Y��F^�0������B�˺d���t���RN�~|;ߝ�5Kk�RxOl}}#��G�|�&����[x�T8�~w�����F�I�P5k�f��d��t&�G�SF��à�X�]�m�J�fV�oȆ}�l���8�hzw��|JkFZ����������(�f(~�j:�έQ��|��H�E4�«���C�-ZS�B�'=\����̳�~з�0�g�_��[`��^.ä�!�x�鴦X��o��.~�$E�ْf��;���ԙ,e���_��j���cs�富/��u�yv�IvZ#��Nap�	.FF��sm�N�C4:�$32�	J����	���"ɝ�k����'���S��3ȁ��T�b��h	p
0���bӯS)"բ*z_�g������IÅ׭pb�1��y��2�Eg�`{��8�&�w\��|�:����W��M�
�&؜�y�7w�W
�?����[�P%�rG�L{���ڮ�x�������T�^c��/R[��M�={Z�1#��^y���Ǚ�y�!5��ʟ%�nJ�������.�Kf���׬�]%��Z0p���X������Oy-[}����@]���0��#��?�4��,�v�g�F�]��	��@�_�^Y�Ͽ�N��Q�w����w�&��y�口K/�@����׮�yԟ�ˇn��8t Ô�`��L)ۮ�&�KZ��7ܡ���I1u���.^X���4/�޿�������B�mp���yO�67:Jx?-��껐�{:�U��$��~�>oޞ�]�b1��m6���O�� �=2�h�����㖂ON��>e6�^�����H~��9|�f�M['�mq�QF�Ŷ� ���%������-Ph����_L
��}=��61�^��uo*��VZ�)C����޽�����O)�8��6���F�6�!\�M[�WC��go�^G��gb� ��d.UYY������߂=����U�{��������gnq Y]�ĉ_������ͷVl�3Ƿ�"{딋el�tB�-�Z�ͻ�c�s�3ᜄNJ�~ �r��6���e(ѲϺbB��$h��d�%�ж���t�ݸ�G�3fe��c�&kJ�c�r�M.�J!�İ���v�����~u���«�|Z���?W�]��f.H�y�q����*.gtH��!�g��(�iP�O���ͦ-��m��c��2Z�|���?Ŧ��(�(a�9d��:�x�5�m�L�N�ɛ(�~[g�o�{/;�^�u������o8����*��g+`��&e�ɴ��C)�ii4�*q*�v�	��o�e��{kTmc��lQ�C] ,h����GOS��:GG�!������$<W3Q�R!�0�O[���r,�J<zPӦ��P��a>������	F?�1Q2�S�D1I���!���w�+�ql�&�C���x���R��u�`"��:c��0(m��Z��?eN���B����O��o��g�Y�ϊw<g�O�=Z-jж��w
��̷���a�3�u�0���N��	����&+�
o{Q~���;�C�e���Tx���O7����|B�'> ��-�v����G*4�������^�Pj�爵�l9��c��uT&a�/)�Xp�'��¬�U|=҉.�� M���o�Ɋ�յ�ŷ��®��}��d��EB|�2�ɛoi�^Ӡ���U(e��_f�$w������>o������:J�C.
t���/�;���9���<G(82BG/u$�H�'���<��2q�ef��l��8����94(6�_!�a�>j�r7z���U���'�Z@��5=9��N�6����w���a^v��x�ᰐ�/�����m�^��԰�^��Kܤ��
3)����7�=i�γAʓ8��M��*O��!�����A�/.�9 �������ΐJvw�"�­�RΨHhe���s�A�������C�G(�gX��X�w�̋�}��.-2w%���iZ�]D��iա�<'��C�����|�x��.����f��O��M�xޫ�w6a����~��X��8:Q{�Ne06����𸕲��'�|WZx��*UUFl�T�^Sgޢ8޼y�����?��Zt% ���J���Ac�������?�������/WN�x�Z�C\���x%K�~ji�a"�@P뽞q@���7���"/ʪ᷼��}�'�N<���^���{��oQiw��d+����0g>k.")�આ\eiG�t�L~xvx�6��i����y�	\���ۏj�FZ ��������+m�0�ϔ�����@	�Fc��q_3~L�vĬ��p��BFu;f���1S6�_.von����|E{��}V;�Y���S�I#ʳtԩ��c�2��I�S�+�ՙ䓴��s�ܢbI7�C�Y�n�Q�m���|b�M�F���Hy�!�w(��� ���#8��Y�v\n�{��o'dut��� � ���4m�Ԃ��~��������bV�aȤ�;\�F�:z5p'���Ap���ɳ|�l�b.Z�#|��Mf� i�dñ���PX��(,-*`�����<cr67���/�,h㇠@@�3�m�	�DA�@�uŞ��:����!�m�����d���_0�x;�e�Z!J����{5�׻M�>���Yq����N]gR���޵�i<���U��>2��!)��r�=��2�?�,u�`��`|O��#N�(.�6t��I�RO]�FƪJ� i0�p�h5��ʸ��`c�٥�9~!q�����q�Ϋ��PP����-��~�8��MxR
s_��/�a�[��
,,�K�pQṁI��16ƚޟ��e7����P����&|-��LV���d���ǋ�=^<{��I�5�Ǟ�
|{���g/���(_�Ǎ}]mkz�^�C��4��*���D�PKuf�_���CӼG�8��Rz�|�g��}����k��0B���FT������R@P�͓f�k�+{�*Z�ꢜCK�z	�|[F*7���E8�?�!��eo#U<>H��J1o�%������P��=- ]歒�'����ю�/p,�-یw�6<a��L��M�o-���º�!{�03)��\'O�)�Ic��x���M]]��**"6Z�v��f�cz�3l��\R{˦��[�8��yb���e�C�$bB^��q<�]��5�]���OQ�>A~9�w�a����z)a����-��2 ��q���{��`���)��x�6B��ޞ���y.EbCu�����]��7���X��޾���j��o���/;��i9��ʠֵQ��OY���Ҿxǧ_���KGy��rT��\��Uxr�4��fBᮬ7�q���k?��$$d��)G^�5s��~V�SG_y�ߟ���ה#�R��r�*��B"�x]����{T/�U�҃�	��+�!)%i�y��C�c�����;���#�F,|�������&<��~���ho�̆�k��b$YF`�Kht�z���p!>�D�*��%�i�P$ 3�>�3��Sh����5�CB�Ќ�Z��ᆛDQ&H+a��#o�CZ>w��޽�jsFB�1`)��1�B�`hѝ�M*��c�^aۉUz/���`o�{�V�/L@�fNf�_f��e������
/��(�12�Uw$d�x�c�T»/�y��lID��Eʆ��4$Z	4����|�D�_X���o\|ϲ�x�d�s
�\e,@������`���&�}�i�S��� X6�U`
#�&�UP櫮~���:n\�&o��f������-�6�R�I|`��\q�>�}�W�ȓ�՘��G^:|?M�J�����.��Tn��[��?�m~�XA��vO����	<Q�yFH�G6�*_~�y����o�9�q�[	����w�Ç����p6%փ���ܽw�Ɣ�F>�O8:������/"�H6v�{f�u@tp������ַ�/6�����q��S¸��b���L�;G���9b
�6���̳�����o9�	��4�*�v�\�� �/���4��K�������8��0���Ӽ(�D�A�B+��DV�����Z�˚�� I_�׷x(���2�Sˢ
J�4˼@��&p6j��1?>�6<x�C�&�?uD+�J�e��|���Iᤒ
|�k�N�r(�� ;�(�Y�b�4m̗�ĵ�l3�|�h=WyU�߆�ᒛXU�����7�ŝ[�.q)�w(����!�P��;�ȹ^(觘��;�q��m�y�n>�m�~m���)z�����)�
O9/���'�����Ҡ1Iy���y'�M��������r��tU�QY����������p�)��PsA�
�Jq�m3�����x��4I�]:�{p�H�	�{XvP#�I�33��ĸ�_���(��]t����ӝ��̆�.q�;n���T�*�k�,��]_W��e��k|:Vȹ�x�Mx}�y9���ǁ0���s�+i*/���L�>O�#��Àȱ��	��0����y����5)��V���X?�_$S�n#O�b��/�3��3�X�6]�����<E~#?j�k�!����H�U� v��,[r�J����
�!\��+��A(K�uH���^宲�8#��[TK����s��[�o,��q�V�"����صw���4Pwd�U69��q��#�������<�D���l�̳�@�\��-�&��μ:*J~�)�y��@Gːp����G� C �
<�[͟�������8o���4nZ�v�N$�y�g���|�$Z@�,q߰5�&- w$^��)auK�D�!���+�xW�E��z�N����qT\u3<��%�Lp�z�i�=`KC`�W�y�*���g�����E��8!N��#���>Z�a��	��շ�Vf�Xv��4�z��*v��חz����w��В�ʞ�2Bj�<�b�8���חV���`R&p$w�$�*y�UlT&N{�[}�5���9��s$ﻴ;� ��
�y��������l�ʐ�
+i�Xmyv�VW"�?����[�8p7������M~�e���#��(�n��
8��\�B,ޥw��t�>.L;Ҥ�:E=�+eK�K%�F�mL�F|B $��]x,?漕�.��Pײ��"���(0��R�Q
A�����LJ�Y�����4)&|��&���#*.�)K*��bXa%�����I�8�����Q�
�(ٖ��a6{�Z���k8�Ҳ���O�Ļ)3�1�4g�e����*�[ޜ��@l0�
T�8����D%k�6��7ن%�����&�Y����yB�g;�g�au�<���z����
�t�ʗ���¹�8I�Q�(`�pF�-�7B���|�ܚZ�hY:��$'kر}a'�e��@Og9$D�]�s#��ȃ�s�+-.�i���,/>�2�.�Z�J�U%����
�@Xi;�/_�}*���H��rŪ�3��B��,���弔'#إ�K��[�J�]z,�=oE��)!^�I���@M���M���Ͼy�R��x0Eg���C��r���4�I����w��3&��V��"��w�×�/�c��l |��c���6�mdR'��>�ty�}V;�!Ƥ ����Hk�m�ت�̶�9���F���-fdR��k��_$C�i���N�v����TV9댱��eU��<����Fg]Ep��چK�]��K�b�q�;�|��a��Bp�5-|��N"��%�
yQ LJV�����iŊ�>�� v�,�A��'?�#��6^ߌ"C��vN%M�,�!�)����Z���?�7��o��w���O�s���l~H�̞�gN��9��N�x�|9�U���� y,pm5[sZ��-������k�d`D�-�p�69�-T�'y��tX\�
k�G;�)����(P	6K����K;|�	�D1'x��;wz<�2� ��k�B���
�]�,�4��e�������A��ٻ��k6�!��2� q%�gR:9ڭ9~�Z�^b&v��V�è��*kgC!���E�R�b^x*���EC}���״�`�~̞N�,�u4�%*��@���0~ʾ>���O�?���s6Z�c���3L)���Ќ�MVh�$��2"�a>�t�0�ݿ�y`��L�u��!"�Nߡ����H�h=s��7�������7���@p���L��Ǭ�;�I�^��A !�e-�(��F�"���]��C��%oI!�H�⩢q��f�@�+��+vA���&�<dnTP�Z��䰚����wc���_dڂ�':�����}�\���A��
��sr	���(�L
t�
����0S"���-��?	o�O9_S"�!g�`�Wу%3���L_��V54f9��_(����E�"$I���9��=�2B%�V��dG��$r1v.�ۛ�?�^���c�l6_�%��;7�,Pi���n�c[�J7e���Z�i�!`���vº3�"e�Ow�͸���F�y5#�W9�[ʽM�#R��O/�͗�Y��x\e� �O�s%�
�o^	�J����?j�Ԗ���0W#�r�VV:���+��׈3�����g�q��%^hA]�x�XY�S������v;�vfܞ�c�.�*c����{�������'��Ғ���1�
�{>?�pwNBA9�)[�P��P"��P�XT2;�N��oO�����<ڋ���l��"���s>��=�,m�C6�+��7)Kp�p+��e�N���W%NO�w$dc��z�����FGގ����m���̬�I{�N�ݦ�Z0���J�f�f����w�8��;���2e�ᒍ��5�"5��[=�*�ʙn�?��s̲���K�<�W��uN�Cltz��R�r�!���`��C�����s�#̥�S&[��w0��g��=�-��"���Sm*�A-~�$�yN#P�2���;�5^/�pm5焳�-�~$|�:��iz	���������"���o��n�g5bSO<�4�ʯ�GtҘv��<+�D�>KQe:��#��1�����P��p�?T�\���Iϵ�E*�a(Hf�m��>��s_���j'��bU
�c���<����c� ��dC�e�X²��8'k�[6�<��(hΕ�`��U�\ ��׿Y|��/7�IX�v��s�n��Q|D���IB(��� 8Si����g�e� wDWʮ���7ro�nC�17��U }fn�A��@Js�S2�O9�,q�\���?�h=Qq�!��s���+�*F�}�{YiJ�������(�)�xL�(#�������r��
8�I~�=�(g98��&�*`�������!6�9�n���X�m疔R)��\�N�P�Dߎ�e�!֙6�ކ~��]s�ا��a>��7�-;ծ����� �(@,f�i�r���S%��Պ/Bt��f�R�T����������KY-^6��FWlD��Ҕ�3(a���3�:H��3�C�RҭG���c������>�Q�z�%H�yJ}��ez�K]��~�C��x�Yƺ�J�K�s���K��O\$Tt�F.�Ot ��;P2d�V�ʿ�}�;��w0e�'��
+@W=Qw� ���3���One���~�9+m��'Ȅu��n���K�[��SZ��pO��X��1�����+{�iNop�>�x�V��n���"��
ڀȈHL��a)T�ڴҽ���o޾S?�QH�c���\��X1Nu_U��B\u��6+��C��ڃ/~�	��9ɀ�"�:��b���_9����h�6N�����������ɢ�(s��*�`N�'��o,Բ�5ː˂�U��HL�V)ʤML��!��!R$�?�VL�J��;LR��A�/�	T������3OTG�t����Z���sOY�a�I��a"'��e�`î'�bO}i�"�*y� �B,f�g\UH�0l��W�+ƫ�g6�:<O_�2������]0�p?<(wX��F�bj�n�6�60��a�|w~�A��<�^*W�ˊ�/nZq��"l�H;�������� *�S�`�m*��O���!��ơ�t�����a�t5֦c/��;�$iӴG��*�o�c���e���4\Oݴ��Ĝ+�Ex��y<ZI6�l3�Cga�㙮s܆���u��A��Ϟ"�%�fH妆�{�[g��p����/qs����#o^�Wv���ܹ�I�Χs��Xm��0��E4i�ͻ"��a�`��W���nO���u6��� �"�R�i�4 ���K� �[��#)�Q<����E>��S��=����F5O���W���l�r�>X��7mo�=�^�OZU�޽Ê��q�G�����d��RlI�������E3��^�e�3�(��M��5��W�Ħ��_�dՠ2ʽ��-H*=��!�y#7�Av��u�<�dG3�����>ԑ��צ�|m�]e��z]����?d5��NX�6*�n.��՟�(h�P�T�܂�z�b�|K!�*�8*���_�o	c9�� U".u�7��2 �]v:��5ʻ>>��?��U�����}��O�f�W���;|?gA.9�>��������ac�o^˸E����g>�:|S�T�O�:$y�Uj��������\�g�������9ּ.;�*d�p������N�s�ӪJ�V �P��}�%�����l�U�?�]�to�(y�U����)h'�#�@cTb|ĝ��2Ԩr�N�[pt��Z�o#G�A�w+�U�q�v��|��p.���m�wq �k��QH�|G�|��)U��-dLd�
F
�����0�;�ӧ!\��0^�T���T~��D��k(��U���A����R�*<�	*� L�u�/�+~��LA����#q\�F��<�������=<�98�%�i������ ��L�Ù�T�✰>/_�"�,
ڕ�������<~*�>����n�п���Ϧ{����s���>����"��[�;�Ǒߙ�q�|��B*ƥ@R�R�3�*iYH�{��)JX��@g�Z���榌_>���^(@LzV����`���pV���BpٱL��<fsU��%�k�r!ȏ?����?/���=aN�U+������ K���	�
��36�VTii}3�ڎC,�IyE���Ug�t�-0�R��`��g��$��tţ0����g����0���8�֍��b� 	��P����Fx�#��$�=˲�_&Z�����8��q2��x� �%��og��_p�'�PWC1.�aD��OJ~��OOp����_�WsIϙ��^�����ա����/J��2>3��~�#y��/�fcV�n㣀���u�j[X�6�\c�S/\}�����S~*�A��=袼l9g�F���)_3ԘMJ��i��Y��F�p�at±t��U�?psũ�+o�ϛ&o�b���*�%�H5�g��GG���߯<u¨�)�yha⣗�1�ĝ���
]�������2l���?����&y-��t���p1|��S�^p:��/���8ᦜͼ[��:�B�j��i�)�'��}��M_��Վ_��s�:C�iC�c�� �֢�f��"��v��=v� v#mQ�"y0w)avh�j����=��MX=cX=��Uh	��Z�&@G�tJ��#N�F��@�~X'\�ș�qn0���qU�Zw������M�皻[QTk֙��M _��K�]���c!�kK�
��܄�ɠ�^1?���o-4M3k���F�L�����y��V��<�=6�Ԍ'rJ:�ƕ�<��������8O��G�؁X{�s�g�${��1�z�g�����}q����ٳ�`X�,D�����7H��W2���"��ɟ?Vocz�U�an_Gȗ�%¥��������G:�0�,6��W�]��q���K�#�pm�K�)������/E~�C&����.��CdP7/�_Q�HR�;�_cB�fm����$}�D�ߠ��Dq��p�ں��*t�9x^�r+�N�Hi}��5,6�ԗWXG>|�����s8�s���]f�ȳL�a{���Uȉ� @�PS�8<�j/^��q��U1�HbD�#=�Y*QP%���p��gg����t�" MT�S���aH�3{tn�ꕧ!��$X��2OUf�3�7Qo�L���$�J�ܬ�Oo{��:�g��N�|���2VR�W?VI�g�gW�@�����.K�he�e楃9)�۽jd�0x'gxj	�^��(}��q&ki
?��fȻVb9�톦��,s{��r��S� $�{d��' �b"�W_|���
�=�@���7nj�"d7-�陉XM�A���9������L��h���L^X&��bP+Q){���Ooݾ���n�Xm�L11�a�o�{a�$��Ն�ZԄH�ã<m4+a-��.H�@�Y���;��r�2�y�_B�L-0�]�W<١����>��_�Xz��1
nd���2a(��q�P��p���E�\�n��S��s�>�q�g�7N�e��ɆKX�h*u�S��?Zڳ_�s&�X������{���e~䗬z�,;��e>�s�冪�7?���M�^����p�Ll2�/�x�?�O��4u�圳S`i�z�B������mW�ɢ�FY,9^�gi
X
�W0���&ݹ�Z�8}K��zL
����6$fT]�mbV�4<�� �~5g��U��.���| ��$�d3/�$��j��^1D�D�"�"mW�8Y�=�l�l�2�ɍ�T��53�#&̉ŵ��dd��-���K��ŮV5Q�5A!�a�0C���^bO�>&������HXď7b���n0���]E	*���%Q�zK����7*f�)J�?t�Q:��[��_M�R0fH_/�w�>s[R_G�M��.�rm��aG|��8��P?��4��2V�����(ԙ� u"7��vO#��D:{�X9�7Tn�Rd6�Y�2t��9=�c6�<d��|e�I�c���&�vNNU�H�U�>���eGCK�[���&_yN�[:���bt������� F��p�V����s�7�QD�)�NL,��iU��_�F^6?�Er�c�wQl\ �Ɔn���<�3���5�/{�N$WI(��J&�����b|�mK�[�t��³�����R��Ms���yJθ�o���0 M���ߊ㯁�_���
8�������4D�_ߤ�4T)���<e7o0WZ�_k����a�ٴ�:��&��u�cˁ�)'�B_�����Q!Q�⎂��o>������s�C�m;dC�41'��3e�y�.�wk��sW���p�<��o��`rVy2?b �f�%m�)�~h/�<�_8\��Q�5�T<>�x�2z ��~�]�=;�G��������p�&�byx���L�R�y�]�&�C�\��2�SZ�`8|8X,)�B�­�u�JI7��W�믊��2D�w��{�j��O��bT�xu��[<��}��K�~���J�0S&���7dT)�f��R\5�ȑ��Qt\%y��]��pq�Òvj�}�{�R�܌x+��c|Q��:5ni0eڴ�7�h�$��u(W*]�mie?��r��T�;�x+1�4��d*���_���z�,U�ۙ�\apݿu�:��+�y�lVQ�������<�F(����Ҥ�ɚ��߸po*ܴ
9<��q�}E��
fEz���>��D��I1�K�텊P����N��9�ᮣteO(��(�v��L�L�F�o��S��z�D�7oviD^�4Rı�W![Il�b�'���?���4d����=O'��D��2��/m�H���H�w���"Rp��h
�*ax��w�-��oJŐu]�tD�,A���]z-a��t���U������2�Y�����A�&��Kn_�ef�LK(��6���rU��<�9��#:O˚q��?��x��-7�� ZS�w<�H%�-�7���B�'�F��F�p���h�z�uW������&M��B�S��Z�Q�tٴ���mq��§)��,e�9����-0��=����/��{ Os����؛�X�W9ңC\Y�P�C�'�7#/�|���d~��B�$��4dڭʧ�[��u�x���+��S�BҼ4\kk]U�G�ñ�_�%�u����p�G�:�UeJ	������[>�H����W�p��[�}�ٹ����a����p(�ɹ���LC��.�IY9�X�{�R�����U䟛�~����-���z�P���9�ȕ���X53	>֪�C��a㉃vT��f�vӫ��Jn��r6b,�>���a�;'�͝ǋ�W���ll�)'v�=[�[������왜Z���I�g�)�7s��VJ�D=�,�4\��i�2�%@��gr���4�},�U��6��~����y^^��gA�ݗ�?��w��a�4��}��S���Ê]=+�a�w�H��2��;$-��v���� =
��ݛtX��W��n�z��Z�ϯmɷ̑�ڻ�u~�M�a*`#
���B��U�l��*�� n��b��Cr�=�Թ�d:T�X,k�E��Z�d��������t�6�̮��X_�.���'ቐ�� �皚�9�̐L���٘��L"C��\�,+B��1�U�/��w�T@�&�Tv3@���nA� �B����q�g~ݠ ̔?AB����I[I�db2�W1�3�᱊�\G��As��zm>�Ma(\����Y?eb�C��n��n��l�SBf"d�������v�<��LC�У���AD(���z�W��.��E^�[ȕ� �P�U��Z!;VA���1w���������Nhr�� �q͡vP�t��u
G<����� �y���Y��tw���)��!��bo`%p���R�@a{ű)>���P�w��EU�\������e)���|:��<3'L~���'C��0�>g�^��2O���<�5��P�ޱ8�]��Qݹ��.᦮9��	��TȠ�ֽT|�W	�C��a��%=N&�2�^�f��Bj^��;�?{����ˍ�[Y~��U��5V�O�y�Rp�u2��O����꥜���-ΕG볽�ethŌD򮰵nw�G�d$�T
އ��*ԄWBV�Bw�$��:ր-�{B,4(	�Lke�"kP�����]සu��{�,>{����G�S��!K��0a��;6�E��R�F�9�2�|�X8\��b���5��P3���v&�g����['��sV-��1�ˆD9�c��?�z�0��Jw,��'9��Fzfۡ�>,X�
����4e���  @ IDAT6��x��\<t�U]�t(�����Т�l0	��j��I���g�L���a��k�cY��L)��o�-���c������e��g����T�d#��Ki�;�^�3s�yM��%��c �����k�Ҩ�^����y���x����0+l�#ec�r�7
���w�̢�u�6=N�����\QgxGgRe����YFS�q�\�P�偺�'޿*ߕ}�B\;w�ju��3�*�yb=A~��)��&���������A⪧ ÎX���*HK<��𪒙h�
�	`vu�������ҁy	re��uzł��A@�hz�yhXOϽ�RA���eHS�En�Oƍ3��,�i��S!Ķ�/
�����|M�I Zii���#��+�}�|0@�'M��;���aήr��4F���KM��LX��N�*{.?�lAK���t�� ��7t%Kg�$��U��_��wA�[U�~�V�������j��vyt꺵��	6�����_��F��x�m�jm�������˿Ӭg����oP�D��ա�<�*3X��l*[4dQT�k��ɓt�B�q�6"<K����6υt��T�}�>���q�|�q�F���4U�ܕ={�Q�6�*礼� ho]�O���Ж9���w�×�7��N�zE�h��rrƍbf��}�ȇʝ��N�}��Q��6n��18���-{<�ǥ�	uHQ&�u�Or{�ױk�z��yp��sv5�]�������m�	EbQ:J���Q6Y%�zg&�G	�*e�Y��H	d�A��|�թWm1�7B��΀�HS,�+�i�v�9^�8��4;h�S���pb��ӟrn�-��qޓs ���/�������*\��g$2��	�0��!h:�(`[#�}�GI}�駋?����M��(��� ~{GY�!fNq<�[_<d���y�z7 f^�rq�,��#Z��4d%9�у[�R{��پ���\��*b�en��ŷc:
�[���\�繥���P��q��;�TŒ2(	�̱�苷�%��>�&��o��sqD�EW��L��r�%�J�Z�e$s���.����n�WyTn�_���=����<���*</�e��;���~��G?��]^-��:��O��,���3yr�nm
�fD�<u��:�$��ZPŞ}m˕�2�irܹ:MQi�<�_E��z,,�2��|l��^j<���iSN�p��5�O]���G�j"�z��e_%Q�eY����1j�}�3Q)�&W��T�#��` ���@�� �`2+n��$�=c�N�bO��R��ͨ����d� ��k��������L#�{2>��c�L��I���P����@0$�����)�Ril��`i�T������jR7��b����T���`��R!�m��i ]ӿ ɛP�A�����~�[��o�\���o�gm*�����XZ�%�M���u�D�$��t��ׄG}~�!`v�J<]/�L�y�6�%P:���"��� �Z&fTU������tX>�R�Y�p n�H���`�t9!�����WWT4E�sq��
�ok��Z����KxP]�9�\��^*u�\!S��O�N&�R�)�XN��S�"����T�����"F�km!�e+2�Ok���O��i�%{DA���K�=��35��՜���2�7��GI���ᆯ"\�{գ�dxl�E�):�w2�R-���d]������U߫��U� '񕕽xO�	Z���"p��4����6J�;��9+h9�����t 9t������O�����?�e���3q���%N����㝃K�(�/�)�*΃u�Sk�u�����,��`o��l�o�uO٘ȗ���q��_�����g����%+]M+��\[@??����s��w�dU��1/wP�\Ei���N�Zf��_�8 �}#m�,�^5/�'��4��l@]��P�Ky֟Ԗ�va��R�ߗ:�x����?�E@�6 V�
�1
�n�^Q���(���t�9�v��i�/�x'��3;SA!|	-�o䮎�5c&N�-�*���P���@�$�i���>��*=6 ����^�*ܨo�t�/�]M�)Z[�%c�ڹ��I��HX�x�>�����:<k�E��Y�9g�b-u�^b���1˓m��dC3��JB:6�?d���d�5��
? t�W�U��̭b��H�����Z���І0K���<̐B��d�btA�S��inx�LH�3��U��5�y$oe� �[�G��m�q����{���GL��R��Mh3�a�T1��[;�T@W�Q�Vj�>��Ik��x;Ds���ISK�|.��y�1b1�p����$Ӎ���!#��c��=��E9�k��K�j�]WU�(�
A-Z���Hp�i%�F}Ĵ,�1T���9�-i�QV�k���$G�黗8z52�,��V���2t��t��姫Jl����J�=�ȏ+�lD�87F˦���>*���KN��%�������7t��Z::o+�:�8�SL���a�/����#;�SZ��@��^�uJ�\�\�~҉�N��w�Wyb?�P��-����|��S�me���a��zF� n�4뭼b^��0Z~4�
�P���O�+��.�4������0�+�Q�D�Ǉ��]��_���<��μG!u�H01�y�w�yF��`��2��)��F:�ΐ���R�p�AQQ�.����u�Ղ.E7-�����0��-H���{,`O�z�h���ᒡ(%h�745?)#��)�˹�nu��h�9g/Xuyz|>�Փ��S�,�x������/��������i�H�[n��9&��M�,�����^g��<|���7_q��7i8�O���#��Dξt�\,�����;�4_ ��t:�V���(�2�P?�2 � \wHޥ��|S׼̆�����_�/�}�]��n�~�8�#��(?������)P�kn�n��I�&^�"_���
eXW��K�l���~)� '�xG��2�0_�]�A��E/��ϕu��L�\��s�p��`��C^Z7�E��)�����\���ov2���}����g,�v�۫1�;���0z�=C{����X]�';�kL���t��+|
"y<ʆQ����uMk]�b�v�`r��P<^>�V�f�-1M&�&��r�b��J�ӌa�{�k��/9[���0 ��2�̀�K����ҥ2����r�� M|�$N��g`\��c<x��8U^V>�* +�W`<��\�Ɛ��ʜ ��l��k+�| �T*���\
�NY\RH���-(�9P���]�F�5]Tb����piLm F���;o� �J�]12�D���yA�i��\-ʾ,%X[Ζ��>c*��j�v4j�69����O�ɔ�쩛��G���D�c�_��a�ӏ���20��� 9��U �O���\+�UA,��s��(;�k��K�b\L���ݟ��s�қ[�+�V��I�$���|9��'�B�нp.�;�'�P�[?X�7���F���$�y�{�xL�8h���ȏ��]bsAv�ʐ�s~f$"}�"k3B˿�i��-4�BA��ȃ43�	Jĉm�O��Q��/)=#�����4����)f=�a]�0�ࠜ9cj$&��һ�7��8��l6�p%̕U>��d�i�-L&o(�t��H~�斧v(�]����5���Ȟg�اWl�`���AK�s��WNDP.�
�;�1`h�t��+��9c�?r�PU���~@����ª۟P���;�)�����	M��c�/ߝ2iQv�F�VW�$6#�6�*��
aû8*�T�jx�W��AF����|j�;��_�p��4�]�{�sR�o��6���`�_ϊU�fD�#��<�A��������]u�2�<\��1�]:�<���QB�_���#�ڶ��}V&T�r�썌E�R.��14ilw�¨�%0<	��9
-g���	o"�w�Y���1���*��=�
�Q����u�,q:�6���@\��&{��skX�9�� �Z��?A��n�Zb4�x([������&���9��g'�'�\�Gh)G��_�C˂:�](�l�by�#t���}.�1���8�����x.1�����ߞ~�N"f�yTlh��-��p�L�S')1-(MtfV^k׺�2���3d�9T��#�ze��v�a�j�6L��[�#��}��	�!M��O����C�dAxd���
*�:?#'IJ��M"��WR�.�Q����&/^�M�5U�]�`��������G�b��c��l[���s�-x���d��N���b�킁�id}�B�R�b`őa]��ńnW�n2,r͕+���P5����[�R��^é��_Zt��2�0�0\aY���u	]�\�[<��E!�A�?CW�خ(<����o���Q�+���+c�?
<�o�'��$a�:=y	��L|�C1M��R镯2�eͣ}�3{&9,�^�g'lZx���pX��U���1����_��A������ǿ.~��{��%������;{{y>��=]��?�3e��<�u\m��:��� �B3�'�CIo�H�Q$�q���Pn�R�a��T�(��M�Jη���uUy|~,�� �'�?��)؀��x�e�}�<4�:ZG��^�e�QIp3�s�\ccR�N���KhĿ�?lʏ�$�WD%I>">?6�Q��w֦��+})_�����][Pݰ�9X�o�Z���r�.?(`QB^�/�BsK������j��,��� ���@/k�{���_��!�vW����U�!छ�.
�� ���/a��}5�X�X٩��Mh�S{z����&����x-������\���
�͌��nܢ"�+�"R�?���u�-��="�&>��K��T�:���CZ��n�^p>^�8�7����K!N�UIt��Q�Y�S��[���<Q���,��\`�TڨN�$��J��G��H���<�\M-�nq�������'�#����l�Q`�q!\
�-G���\�V%LZ�%�X�ۂ�Q�J[]VoЃ�*H�m��#�pr�h^qE�m���z���u�ѭ�g�ѣ�����c�aZ�-��)��a�}"!�
�ƪ��������B�01��4��/��1�Z���e�"��̈́yU ��@*�+���^���U��2�iZ@��/��+�u�j�ߟ8�^"�\������`fxJ4�wf�èT:Vq)D�"j����kf�D5�E��ʒ5-�;@�J��ΟX��Q�t?F���	��a �=�����Pf�pC�M�p३1fa�-�%��Aw���P>�!-��J�v-��- t%=�*,�m1�p,% ����F�[�K��[�/����s�*�_��암M?�0����w�`���P���`�S6n�*U�g�fo '����K��I�.�h� ��d޴���dD*��_}zY�,�/�
*��l𝸺�C�7$��?�U(}��ɏ
|���S���W��Bd#�<����Fx���ʊ{-m,������Uh����
nm�;P���̧9�(�A�&}�ǩ� J�kl�	����-V����r8���nOIC��ζ�j`�`R�-6ۼ����g4��l�qȐ!�d.�����I�C������ �Z�Q&\������A�z�*6bU*���cWJ*�L*����-�ȗ�:��t������F�wc�?*Xg����G���&h�a(���T?+m��h��!"8�a�鰾��$z�0�ZQ��7��*���^*�|'��9{�g5�V���y�ٶ%�w�8���lrN��
�6߭R�2��)�t� �|�L_�j���qaXo�uvHѠ����8'�Й�ҳ�E�S:u.ࠞ��V�ꉝ��V��!V������r%d�a�P �|�\x��6]���替�X)���}��z]���q�VF�[���+d9�]�&�M�����+O�vp�޹��:�uS��C쐙��_��|%]1�?ū.eM�^�^�W����1�o�����<@i���m/Q��EChK>U�;�_��V�#1����w����C�����.C竑����|%-=�Oa'��S#L�J����A�CZ��X�F���{`X��g%e����D��w�#D\�L ��q�,v*A����HC�=L�L9Vs�u<�x�[Y��BI�5.)�mJv�S�v���ZM�d(�A�-��4?�𹎤�E�u�{1���;13�%�7��:U���H.�AQ[$�"�:=�4A#&_��z3;a�Y����ѻzr�D�j�$�ƣ��ߒ���iNȖ��R��5�h�F0�-g̽|�!�/�$�9:X�\����p*X����i^V��[����!Q	�o�Vެ��'�JXS� �a�#z�kϞeW�٣"�pp����< �U��C�q��_}����]w��/!������G��CO����F�F�3E�6`6hN��	���ְ�yE()�m���ս�6����f�{lv����◟~X�z�A��tY�-��{�ك�7������~e?/������&򌳞C�f�Ф%�^b��RŎ�{���wX�Mo��>VF,h�m��n����;ٳQ'�����H���b���<l�g�Sw:_�eyXF�S��I�Y�H��(4���i��5^r�Y,y��*��� ��$������21x���������2\����lv�;y�o���j)g�+���d�ql�����ϓ`��id]1�+��^�΍��g�&��nw���Zv�^�D�t,��<�HG�ź&uL_%{��j�sfM3�,���(ʯ:n��rp���e�w��5�v�܃���D)qt4�%B>��a�}�8g�,�Ж��&]��R�*t���K\i�e��M+����2�'���R>���=�n��p��(/��D�\n?�싎W/��z閲m(��Hc[�$�qGx:,�ޅ��v�"� 8$�&���~L�Iޫ��esћt̤K�WRa�����L���>�Dy9t�<���|�p�C��p���9����z.��4�ٲ݁����yfy$��I��%hũ�R�������#X��P�$w#�*L�uQ�47W�w+(O�Ȧ��H�ņK?��YR+�>�TA���'^�����?"yխ�F<�o}��˖e`>���^�^�#T�۶9����:-���G�y_q;rG� 3�·^��Y�#C�9G�����)�������#H��ne�Td���Y�'�n�Px�]2�>Y �\dP�6,"�b+př�P�y'� ��zR�'��Y�_�s�(�u���]�l R)�UE�A�,!p�ƙo^�x.^=e��9C`���+ĥ�=%'9�kr�$B�t�w�<)��5��4�G�����u-An��2����k���`�����ryW����"�1����7���ob}��~/S�.�/><܆;��s����%P�ܢTQ.*�
���qk ��b���C!H��Sz+8|Wzk1��!w9����D�)����Z"��q�x��}��^��������X��P}�8|f��s�)
�������^9�o���Ӎ�@�z~�z��6�*!N�6_�	���}�A��*��������2|�Hy[\
�p�;�����(���s�&��#��Oty%/~�D��~, Ì��S��7N�Iю��m8�K���:���v.�(c2��-��C%Gb͢ᯎG-��ׁH��y8��P�ni�|b^��"ȽB焓�P��-�6�f�bk����v��+���xU:ƭ�T��U�U��U~R�J%=�^U Y��Z�Js����[n���q�,#s�K3B�`�Ѱsx�.�C��idxn�Ky>���I�'�����{��c?�{�| Y�H[����w�`�$��W�������iǫ�}��r�,1=QVt�N��e�έw�l#�uJ�갠ʅs���MhCc�~���h�%(�^,�<�� �);B_]}����3'��V;'�훷l z�Dr���L�ϼB]]A>P)3���:�+��׷��T3�'J;�&���҅���	<'+�`���SOOk�xz˓��3�1mA�o$(�\�]8����{�!OS�DZ�M���O!��z8t ��su�V]�S	L��#*��h*_��"t��͟+W����W�f���A���x��W� -�A�4J�9C��Dw�!�2 �����(ad^Š��+��"��bYi����],�U(AK�z��u\�ܽ�`��l#S���)��JQ�r�Z�F4��,%bB`i2���³�a�K��l�Ji^��Z��=y�8⸤�G���\ ��=q�2w ��cK�7h[%��L.m-�VtI�h%�V������Xb�$A{���,��e�l8�7�>�����R�8��Ǯ�f���!�/�h3��	�BJ�H?ũh�KR/z�\�/�]egpq�_R5@�`���G3��~ϣ��p��a{��j�|I�'DS+%L��`��[�|�7�"����'���»�w�}n���l�y�3����������m��`�B[e�-yE���^�����
�v��}[Ň�8P��1Wloo���]�]�ܽs7���nk���u��@��&�#V�)�z~�iT�J[�T�alT�Q{�Qo��y��QXwP,{e��,�t�W_����S�K9U�
��;N���W���v�X�E���o�i��C�����ź<��T��Ȥ�Q/�tC�Hov]�t��U�N)���{~�Ë�7�P�);�7L^�z���]��a$q��Hi���`�[���<O��}�,#�/��_q.˵�Rʙ�7XUƂ�q#�������i��R�����F�����(���W��s��-'`����(��y�
�����َKM��J�5�m<"���Ѱu���KP�d�%3��/�����K��*>�K��R�G��By�7�8�	R�w�Q�sAs,S:�z)ە�5c�V�E�W�PV�/�e�fc=2?�I��ռ��|�_�CtX7��b�nr�UY�<��M��X�yxzxOK�޺����8�����OG*���':�|�"d�����MAҐ�[;L`/ͬ��P�AY[�VRo�0���̓���0��Wb� /0���HE\���FXϫ��߿@u@�
�t��G_���|\������QJ�So�w:��������?K�}T&���4����E�gWkr6A		bV$�L�Uf�g�¤xF�r�Lk�;T�7Y����,�7rhIMW�m�������
p�*�L¯cQ��2��
37j��wZr�D��(c�{yiLl��.��E1�4�&�����Mb@K1�C҇p�ojz~D�c"���c����ԑP��Ps$
���Wo�/'�ۘ�\*(RAR6�W} r����@ ��,&�����µE÷��ޠ�NO�F���o�.!{Ea�8c�'#�9~%̍u� *�L�(t�2��RCq�S��g��i���0���h7Yi��P�@�� i5p�˭f����^�T�@,�q��u���0'�>s蕹V�;,a��4߅�*@?�B ���䜳�d�i����GS7����2i;Dd#VB�s�(2,�(���@�u���Č�qY�I��+������(t�K�ep�(
_�TI�~Iy�tR�ư���uﮆM�ɾΑ���/��(�*/�����ϳ���+WXn��r
y���UO�V��=`w�)�u[�ȚUN�XǺ�S�ɽz���v$�U$; �G���2�iz�V|��"��%����ڪ�@e^I|�,�(���9�(S
�<J�trx1t�⥂�I��:<U+��3?ţ�,cᩀY��b+!�]��4�"�ż�{7�?�K���+н�����uZ�\e]�&��ʘ�_eJ����V0���Y�$�HS�RSK�1|�[���?�h��ћ൏ҵ��֧y���bQ������e��?�e�P���z�U�mbW����( �[��[�e��Jn�];Zo�d�Rf^�-pt^�{E�kSڢ$��S<ʭ,��;�q�ߌ	�ۄ�Ǜ|P�ⲵ�"���tW�SZ�T��Y��o;�;�,b��ְl� �HW�j�)��;CXz�Ѡ�ڳQB��H�+�uD�O�RT\�/�']��:�N�:|$�JX"��#0r�M��{8�=CSv�����?��ߺ��E(餈���Cg/Ӻ� e���7�ô�f�_�<7�N���k$W��*!>p]��ܭ�U����0Cd&��w��Q���R0VL��ـ���#��/�@�=+��H��o�zv�e��p@��`�WXCHhb�r.�-Z:!�Ϸq%n�4���O��D�'�rSx�1�q3��/����"ߥ�B
:?酽bu���3z��W/v ?�7F#�⥐���
���x)4�j��M_���?�����u�Qb��
T�7OU���q���-v�FP� �o0��a�*1J�[�>�"���W̗�{�wp{����X�hj%����E!W8M�����D՟��Wk��������4D1�g ܭ<Z����[�^+���1�~}�$�����t��;CC$l�أ�~��G��wDA�ՈBt�K˓y[&Z1�O�k�҈R, /9DDcf#9j�,k�z��S8�̷�ʜ?���%�
� I��K�({8�r�!1y ܡ�~�g��í;H�������*~x��e�Ӿ�ܔ2$��^��Y`�`}�?�]��fQ3�K�������ڰ�q�*d ����L� 4 ��(p�I�K_˩px|l B/��BO:�ཥ�2º��"�<;�p�{��*Tt��v������~ܻ���,�����}��V�%���(���t7��Eٲ?q�"�s���ݻ���[|�����#'�`=Ŕ�̡�5&�on`�b��+�׷�ٶ���.?J�B�~�`eU9�4������Yc�WdA��u�\��ꭵ��RxXE����mO�*��F�Ӣ���l�P~R�U*�r�p�?y��O�"�u����G~�/�l�v�$���~�|��Rv�#t!����nr��>��,����V���^���_(S܀����<$Ģ�H�pDH�2�q���J��E9��f��M;����)Ǉ9Ty��{��@�h1ߧ㷿ئ�܈�/�����4*�X��0w����R�-O�"x��2�w�T�E���Z�Ko����ޠ����2\��BU���D�(��x4"�^1;��~1eF9���S�UŴ�HNBH�H'�LW����}�M�~��t�G����>�4ؿ��)�B��!D�Z���(a�crD�Xˤ%�� L��+�=�^���#�'
@�puL+f�:j�3"#e ����1���k��������q�xN임�Y*�*6X�^3�K�ׯ��	�����V���R�R覷��B�VZ�lޛn|\����61������8��I�7����}�"�C�r�aI���Y:f��׻g����0X�z-�Ml �Z� vʮ&Ū!X<�/�y�,n��(Ȕ��$=�
k���~����(�n�Z�r�2��XbM�Rq~����N�2�k��J{4���s@�����C>H�4�EV\fn�{'�;	�td��ru���1ʷsB�UR�#���)�/< 	𖞱���0n2����΅x�$U���Q�ax��&U��/���S!3�\�򡫼�KP�R�\#��[?瞦eyT�<1�m"�D�(F*�\	��	���y�	lD�`J�\����G�x��O��M�x6�Qb	UJ[geH v:NT��*�($������.�6���J���p�|���/��a(E�E!��zï��5i�U ��tn�c~,6����0e�xm��߄�]h���%K��C�d0֠tNIO�F��]�ֺ$?�麈�M���ƫxر�ئ:�'���X���VC�X�,�����
�I34�fj�u��L *�����ʗV�3�\S�~*�vD�[�W��c���I,ᓰ�Rx���ܑ��3<W�Hy#X S?��{BT���Y�H����Ͷ�\��JT�H�p�B��(�nUS<���<x��6��� 108w|؀�(`j���
�7�͈�!d�@�Q%����|���>A�c�N�kC��rע��i�z$U�/�J�g�V��-���，�Ui��L��=�	l�O��S�7��!��|!:���Lu~�#
X����{j�
��v�t����h�����۹��:�;{2�A}���k2B(iآ=^}�
�8�6Jw&��S�hx|�6=�"�a��=4S�B\q5♮�����^��p!Wj��T���R�=y����G�r���IO_��MΫ���D�-��CF����0l"�6���x�A\f�yL�����1�x�Q�D	@HyL��G)�:��5.q����7*�� R)�ͽ���``= �B�"�zȧ��8MW�Oq�䖠U�%�jKKx���ϴ���p�|I����Dju�dix���@�.�;7��lX��r&��7�{�V�D@����q*q'[�c2/g.*�����(�X:���v8��٘1w	���2dc�d�1������D�A��B�ɟV�chy3�+G�
U紹�{+i6��p���to�W�����cn����)��ż�0����"hea{�w��fL!~o�^�0L���5��S�Pg_�i�����eڦ�γ��t�b*\��#�Z�T8|�c�/�䗆�zg��rV1����ʒʌ�ڇ�����/�+�Z^,/�����ݕu�5<C��u�����4�����2:[��
��M�-��+�b��?�j���:�[�1O��Z̥��m���o�	�����{��S6 ��F~�N@뻊�~�$� �R#5 @�z��0]�XY�-ԇ^�К�s�Tj=]@�m;z��a�q�C=�mEvJ��%^;j�6���zn����^nr�y��`�a~e�
�J�|`�� ��ʏ@���^�u���r����F�Gʪ�1^�:�����5t��Tn@;��^a�v8�U�'�L��N�����T�@�֍�B�HK�vpw�p!��V�����Z���mL���x6��&=�{"�,���@.�|C�0�-L���(R��F&�.�����U�y�w�� 
�ֵ(�ni�6����j"���
3�-��d�
2���?���i�!�Ay�v��<' +���r���)�)�D/�'��S�ˀ7�D�R(PF�$R�s��F���Ty4i��U
��) d��Ir���I���;P���0�.fy?u�a�0��=R'Կyu�8z�h����ų�ӳ�7��^Ea��*`;Y`yQ�ۨ�Л�Q)�,'�P�2
sϼ��k�V�Y ������([�]N
P���\~ʼ���h �xv����]�Bfؙ��{��,-h\x��A����H�R�0V�J�J˲�@R(����h��Yxg9��lр�p#��4z�Ғݫ�qp�}�@Z�R�J�{%���_�t����V���V��b5�
���ʍC�*U�URny����4��U��%�ҽ��;X3T���A�L�?<�~��p��+�28xu����fCb���e�+~l�c}��L��,{V�sr~�bx*Ч�mBM��Ͼ��{9�yn��RJ͘;�=u������W�G���Z)jh	��S
${�QG䳺R���sj�M�x�DE�2q2z)
�B�5�I[��{�����oW�Z/8��#`)O��B{� CdB�V.�,7޵��r2x����Q�TĜ�@�8(�\��L�=N��+D_bA{�Ͱ��6I�h��ˣ�<�{�=G!S��"_HHy@e|�1��ӑ�O�J~"Ky-
J�8'WDȃZijEa)�b�&�*˩l�3M��Z.��3��/>�B3S�C���[b��:5�V�jX��
��W�_(^Z�H�vH��F��Z�2>�~m�V'��i�I����F:�r�}�:
f�,]+�?��I˖������)%Gk�
�uF#�/��������>��QI��[iF	K�d����̛�gĬ~5J0'_c�F6�㥄��N�Ys�����r��~���s2F��p�D?'��^W��v37_G�0���S�.ϩ�{+��OX���n<�o�
S�k�U��z��/�������S������<v�0)���@̸��[�m<�jdt���Mʆ�{��~�K���w�S#/�����n�VȜ 0��r�w��|�{nS���߸]���1q�ͫ�lQ�+{K����=fe����k'y�)�:B�]�ex/U7im��7�4��Lz��'N�wl��<;��N�,U;iJ��_O�VW<��&�[I/����=a'�G��f{VZa��ۿ�XAaKZ��@�i��5p0/� �Dީ�q��4�_ e�F0�0巚�E	�Զ1��*/��c�Ѱ�:',a��B�x&L�_|���NQ�n�`��� ��pEʼ��i;:z��6�[���X�`����;�5��orf��?���d����q�u)f���W:{�Z<��rr�/-�)0�E���X��3ZHܲ ��w���7���^����*N@v8̡n'�7���,���r��%D�����~ژ�i����74�𳊍�߭4�]f^L�\��_V��eZ+]�`o��a����0Pv'�6$�2��މu�**�ӱ~��C�e%���R�.������\���s�\H��J�����
�<d~��8n�b�L���,��EV���Õ��b���ca�Ppr���sx��F����]K���tM�:�ę�)��h;��SJ����ʛ�8N^�]g�'w�Î}��W�d�
k���7��B�J|m�cu�,�O_s��K.�ِ�v�A+w��p8�oRJyf�,����d� &�����k��%�����6-&W�*���W+� Iz-�F$��5�H/\�OqݡS� �[�q�s��=?�t��ǁO�Y�a�V� +L�W�eˏ�2L%#x@?��ϱh�a~����!�u�(G��3I��r�"df�W�(L��*�N�����2��IJΜ.�K���!�ӥ���W��mf���8�L�t\���J��{�ip+������s��7�^گD�)��ʃ�Z9��B�eDT`:/¥�6x~{u�Z��c�$���#�� � X���xjP�9�xh���RyQ	𛻘�O% ��l�~>��U���x��+J>e�!F-_�X��K}��/X9^Gp.���n�x0�y*6p;&쪐���m)L�Jg�K���#�1F�nV�ѯ�+	�$-���0b���i��"�Dm��ـ���r��`��˦Ũ�e���u�VOCT*p��'<�L�/s�VTo_��2}g`��P4ƊA!�z�2���dg�V�p�p��[>��Q`\�<]�P͡��"x
�|�X�d>�J����al-~����/�<�qs�����<pVZ_�����^lv���ߞ������`�U,��s�l�]�����̄|�;4i�k#~q��;�=�$U��O8�
��R��D!�J���`gi� MD7C����C�Y�(V�����rR��j��*�������V��=:}N.��+�0��A��0�Pj)�=���x��J�� �R���5�R��j���V�H���ل�a��Ⱟy;a��<eX� (t����וz6zu>��U�5�;�k%u����i�Lw�wU�:/9��mM<�*�;0����q\�����[��d�|O��y⎸ �XN�G�y�]%L�߼dr?���c��nr��%�S p��2��Yo`v��'ߗ���rV%NE�f3W
~V	�ᷜ3l��(�0܄fz�M���WC�����X-�6A�q+:T���D��T��D�C8�໼m�؁�E"!��Cx�����F�񤻂,��[��Ǥ�w̔�x���������;�Hr$�&ɤV�R]�fG��[�������nDO�L��,��*j�{��I��������p8T
�}H	�E�=��<\����;��%�ն^���8����s���m�Be�ނ�a��7���W�*O��f�y��U�&͖6�f'�	�H]P_M�ti�s-�k  @ IDAT�VK��+5&W�c�Γ������&ao���N@C��J�)���)�&�;ڀ�<I��ݍ7�6�@��Ԥ���ڤ)�u���W`镈R>xû�U�à�
=��Z�,L��:B��^�|��{�Ya�b����[���Ϟf�*'�ګ�`v�5ad]�p����sh���^$`R5�46�$�����&P���A��ʧǻʨW� �B����bpr�p�NF��oP\lp�YΐG��;����!� 40s	?�pٛ�t�E�$�T%
���-ҫ�o�*�����0��;�(̜�p��A:��s3/��·p�$�x4^��wp���E�2D�|kXִT�c�_�eN
���<FޅAY91�_��w$���BY=fחlƺ�\��bs�mM��׻�����+�Sz���Ѹ�����˹-��4��K��yh]y�����U����D��Cm���<#HC�P�����}>�F�P�ӡ,����)�-P�RT6>��O�^�e^�K�V�P�$� -��#��$ �^��H�Ǐ8L߆����̙ʟ�i�xz�
�J�t�K��~��_�~���E��(KK��:f�8>~?z�f{�˖*�L�G0y:�ֲ�X�\�;^(:CԖ�J|Z
��A����!��q+����"�s�N�����D~��F���L��pIG���-HPǧ��%4��w,�~"��s~KRq.��WI�+� ��翞(��J�ܔ���:d���w�����0q���w�l˗�۷P^Q�L�\X�{f�� �#NZ�m������5�v��BT��%/�&�1��"�t��^���Fx����~1j`��ya�f'ĩ�����٣L��M
50�N���3��^�a��n� �0�_*�$*=�vR�߲�~�S.VR���
�(���� /��� �9ù��'�v�&ca q�K�yUڷ��q�O��1	�k�>��w��z�vBP����M���k��{��G�π<��zu��UO��P���tv;�
P�R�_���,���נ���+<��bL�C�6�aJ�,�Z��(ǂcoc�?��w���4���o5Z�B�O�`0��ן������S���/�M��b�@{��� Q���\�ko�#��Z�T�r��3ٲ��
Ga%�-�$W�̋�P��0�� ����EP�����|�<�4��[ܸ��,hSa�C�*T�<��z>3�Ω;@0�}�2Ddc��C0<1 p{6�.�W�{���]}*<��� ��������%7-x�97�9򦖊%0����� �EE��1��D����
�y8o���Jc�ΰ8��a�3���C�����(��a��%���uy���m�u�����ڃ��X�h<���l�Y�Ó�uiS	3뮂s��l)aM�rqHj��\�X� �7�̪=��J��T�����U{�O���n��`��]Xw�[0�)��k��D�\	���)Vy�	�@�'�*��W��~{O�X8��}Wf��M4�����к[7��]@k��Z�ww9��r�p6[6X�;�}m=�*ڀg�/So���=��و�;��-le/��bgO�4b�tK��@���I WK?A��3�߽� ���YQYC�CI��o��(�_OO+��F�a�[d����<y�����h�bQ�ٸ����Y޻B�|���j��/34�V�S��HR+���d�M��q/��|s��v���jճ��/�R��Q� �9D��̏o�OO.�ۥ_9�[�Qs)Y+��R��'�(� ��܄����7��f}-'-1�]d(���V���ʨE�-�,x�b�.���.����	{��th��c�\y6V!�$o:U��E+��X�?�v�8ٹH��c�,�Xq	?�L��QІL�OC3o��ӥ��t�[�L�I;O�N�	窫D_��ղ�QD�"m�y��.@ed2�kJ(9�<�f�a:]at�]H�,)6�0�2�T����P���Q�u�p*��(P)(a�k�٣'W�Ex���X������2dl��n��߅��R�U��n!DZ�~��k��E40�{����!_2o��`��;�b��b���#V�z��&�`vd_���C���}����kx��QZ�
 ��;t�K:����b�Q4|<;VQ@tO��}�+.��W�'427ѽ��攡��6�E|�Z�⣅��:,(����%�F٤q�!Z$��Ji�aV��\Ű�{�췮��ȓ����0nP���H<9yP��9��!Ģs����l��{����6b�B#��^�8!h�wd�Nh����a�K�fGs��,��v��"�����U�D��Ao�����4�|K�T�EAҢ�C��h99��!ʻgt>z�(yQ��§R�&���m�0;���q��U��n±��GS	sXҡ��no�O���~n�E���v���y�?��ϔ���%��D����!���tX�[���㗜�%B9�ox��������c�ݸTژnV*:���qˈݝ��Ϛ��B���{}�
��V���2�Z~���C}*�G?���|;a�>}��Ud�{��li1�Q�E��A��w�'�G�Z������/>��͹�p����3�*ܗ��|��F?̼L��E�S.f�����*�<���O]=�3
P�7t�G�V[4pLr�i�4�K�6�}����)��#�o^)�2:��{9Ɓ�}�N�J�q���v�c��T�9�N~�D/e����b��~Y�r�?;��TZyi��{{�I�:��}V}#d�SդMLܴM�cG�+铿 �*{�+s57�h�(W��n4�6�ۯG�-��'��{���~�O�?abn8J_�<q$N�)��"5��!n��'�!K�P�߽�b.�SO�p���x{�sE��h�L��L�����/�U�Sn{��e�p�CҐ!8D�]��Y�F������f������Q��(�*��o�*�b"�qh�/&��>8�L1F���!a�kz�e�lC{P��*��ƣr8�t<�2��4V�O���a3�<ͳ;��
����/q(g��-!�����(��!�0a�v�Ɗ7�$聑���d_�����/Fq`A�U��s���X.j��}C��*��k�o�Ǻ����ɳ'(_��^_2���g��w�����t��t��g%��7�˔gAnA|�8f��x�S��i��=	I����+��Sm��b��r�K�~D�wF��y�
��ʨb!ݵl��{U*�[y��!��8�p�����>wI��֗�Y/+#�|(`	��ևX"�P&X��|�����:$�moО�P"r[ �-����D�r3�kzM�4tE$�b�Rjdޣ��@/�o���9N��n�(��/O��H5��S�ڈkaq��'O9S��ߵ#?	G!�ܨ��QH��Γ��J�W���D������M<m���mK��?�a*8��e��n�^�F�+���ͅ��V�' _���&qpk���-z��r:�Q���T�ޢ�5���bn/Y�z\��(���ƺr��$_�2��g�cZyh�Pj��WI���r�:>�b���շ��2���/��Ob�RN>��v����X�]�<U�ɨ��_~�����nkc'���*c���z4��m���
�8���.��c'��!88f�C��8��H�$�#�R|[>�q�B��U�%u��-�+���r[ƉD-��<4-.���C�ݮ$���1�I������+��'<���
?mN�7�M/	�W��YwR�ɷ�^=���u��=Hhb�ĭ�����S��Y��I=���j��u�ƭ�ƣ# ?�PV]��V�;r�\[RS���#H�M�xc��Iò0���O��о��y����C�U�^�c����ʢ�W>�6�\S��x�)�؃�������c�M����@\��ǟ�l:U�%;K7(`4L�����a��9�K��]eP�+�V]�l�.b�$�
��x_h���)�?��]\+`��N>+��#b ̟sWLI3oV�x�ڥ��X�T�'�D�+C�<5;���`N��ysfB�!V0��Z^�z�N̯i9I�b\+\Q�o{* �@��_�/'hf�
��qLCIK-^4T&jɉ�q�]��G�D��i���*`�g,�����w{��7z����ٯ>�D]�{�!�,����������4e�I��2A��H����¥�[���OÆ�)��\��0* �Ex�.CS���kl���g?&��_|������;�c	�qR`g����;o�J6̌o���2V�{:�fp���g��\�T�TV���4�+
q흹{���^��Tr�MeQf���e��{*6�(,�1	���2y�����
�?���y'��sN�֫�$�����՗_|���l_��ʒ���1$� t�59!������	�n���u���	��W��(��RK�"So�Q
��6�Z����{�����	�S��?�Y�s�So/i$�ĿdD�;�Y<U!�ʖc
(�*��N�'��sH����Q��|P<��W��S�hk����;���w�}���D>8�K,��,�b�L���ЅKXc�BA�o��h��y�ܔ)�*�N���|���i��&��Ã�4�h]��;��ݕ��|[�9"Ӏ���ʾ|I���Ip!�sN�F٦��d1q�	�lZ)bY�O�s��m�}���M�w�|���]Tg����❖��ȗU�qDn�a�Ph'��UEѻ�@�E�Rʋr��y��P�%P���u��!�>�G}~om��GVZ�TzsLy�HF���&�O����ϐ[�%m�������wB��]�)ؖQD.�bs˟����c�7��w��x��+U]��:�J��Y�+�����-8%y��W\����R7�u.˸]�2�3��W�u��@ѳF?<������l�b;��`�N>uu�,�
��摗���I�4��n��h���U�R�A��m�c��M+';H er.��Ѭ5 �g<��sN1 g]Aì�N���V2]W�1��<ixW��r�c�Ԙ)����fh�*��T�p}7�$�I�Yx
+A�D�WĨ�6!�H�xs��Y	�T�Dgx}t�Qqv\p�$N��č�%� T���{���!f�!�WX�-�x�����Gޭ�=�;)������#~2<�8�	���7�>����\���	�XZ�j����G��K�� !��g�M&.w~ZТ��7d���la�*p�@��� �$�5	�Π��h��wH��ݷ����C�� �?��dVᤂw�&�T��n9M�jB�ʩQO�-my	��U�� J�,Ow�Uɹ_�X�<�u�E��J�J��#_)��6@Yv�R	���ws����/hT�FWX/$��/8��dc\���������š�������K��"�H�̒}7Ѵ��5�52⑹;Tp��T �ʳ
����a�kZ��ȴ[�T�|'D�T����QQ0�Q�'����S�O,�!��O�;|���pQ%�{�1@�U��&o
;��ҙ�S1Ml�`���a"z�-��5�qغ��exW��iJSi�oY�E�xO�cͅ����R6v>3�C$ R�;dN��+\����K6\�XT�/�?Np��an���B�]x���5Z����m>�|���@�h�+�]����-V��e?�����4[��4��S���d��C���c�~�5�{��)�q���P���V~�H�]Eٔ%O��y����{������/T{T���@;#��6�2+���L�έ��˸&U�y�? q��/|$/7�w�&����V��X�&��`ʤE��U��4y��R-G�1�]����I��3,ݭ��'�3W7/e��e��N�S��]�[��b4��,��O&�|��N��h��K�WV��1� �gȌ��Rߨ��Mnd�O!U2GH8�݌Xb*^(��q_���r.�>iS�$Z��I,񒎱m��S�)��M\-]7�-�3�ϔ�t���*�u	_\�����}P�R�:�5T �����G��P�ڛ*�]q,�܆7L�+�����0��Ȓ�4jFBsW�[��`�p�jÚN2NfN܌��BT%C�Cѝ\hc|����sr�'�zz��K�� ^:����5AZ���[�cV��;��Î��:e�b���T���<=v�ˮ�688�w!p���LO�̙����G��7q2�>��(c �Q��_�"I�F�Y�a�(\�黣طfw��W$m<x��O�In�I����:4��c��f^��[6t^��QT а�p:����\�^����
�0��<�!�'9�ט9[��K�}�g��Z�@\�����G�(l�q㬽����]V��O��!_Ή���U��xx���C�������#�.�7�1B,�P`��Z�����{��c!�͜��3'ڻ����FS�{2���<�M���j�����`�D�u��b( 1��*��@9�w��t�ot���Q�~ww����$��ߔE�x���s_4V�aq�d7���jd8��ݪh���+�C��G&s�Pf�Q5gثO:��Ƴd,�ye�~��G��?7�`�蜆K��9<Zg���%)i���;H��	�m����O�J�K�s�lΦ-�Z��'tİ�N�X���t���3�eg�X��B��k���Ͱ��:ZD)Q�y�������W�/��� ��O"�c�	�c�H�G��!*�B�� ���O9j��s��D�DZk��L�`>�&O�*h�����%���$�(�։�-��<�ܶ8wS�!C�Yt��ޜMz��E8Kv֐CZ-{.?d���4���oxϕ�_��X�\!����s���'bI��<];�.,*����M�j��P�����0\T(W�ʼ������*���� ���<�=X��Bn��O��p;��)p1{ݴ�øЙq�ˤ���p���:ǷIf�M�1(f�f��p3ޱ�EĮ%�V V
5d[����WL\랸�3S�p@���@2)�@��:�E�����"&���d� �".v
C��H��>j~fU���Z�6�Υx����d��"VJ�4���T�V�{�,�~u�Z��I�k�{�����O���!s��u��C6�t������.Hl��"��z��^n�����ŭx�d_F�ݜz���4�^D0�la�&'�;ܻ��d��a²���=�¨�C7�-솏J#	�qhec,�')�G�\��xXARpF�ߎ�
�/2l���1*m�Ţ��pw#��]��3w��3�q��z�}����=&T_d�Fk�5�2���t�A>ج-1$m���Y}�����J_۩4O%@̤���������E��8�@� � �yV��
�`Y#�⥢f���,�$� ��-.�����vv?�.��XwA�����(�O�T]�8vpݥ������q�&�\",��J9�+�Eⅆ��8@�?�[�Vv�o��i�.�B(�;Z|T����9%*Ȉ�P)0��S�6n��Z]QN$�J~����AX^���iq7}f\3�tt��˽�*�� 0�8V�]���M��y%-�d]�g[~���g~͵rNi��'i��b}�rh*[�0�*=����#��e�zj��2�h/ߔs�4���&r��24��i�m���+���%|+}����7^=��&UJ�ބ�yWy~�C���+trϳ�?{�1y�n���B�je�r�Όf �=�D��������������(���pI/������e�R|��SN#a�� �\He�LYj]�t3�0*nnp-�X��m#R��-*��x;}B�S+~���T#�"���ٰ٩.ų�/�ݙD�<E*�b(O�w�	�m=�}�Td�p�8tK�m�"8�o���.�ER㪄|o�~�$���ɜ��2������n��^��N����Ѝ�t��f�/���Z���b2"X�юA��,	^t��:4&���d@_����G�"䚲��݂�������^�|M���?���"��S۷�j����g��������z����m'����{FL�g�/�~-�|�� %J���P�晼7��t�iz^�Y_�ې�v����xj�+���((��(F�;N��g�x�r�:c���=���抽���sh'��~*�ɳ|�|OJ�!~`�`U�U����l�+��y"]���nЁ� �����0�ß��E�a��n��q���y�`�s��i��UҤ1�̑��3s�I��M#�s�kk�������Gs����ba���<?���b�B��)i�K��'�/�^6z{:9�ygZz�@��@�D� ������P��
b��иh��y���l��#.d��
?�V����C�?����E/�޵��+?�g#����B_%J%UeL����?��%��,WA�AsyH��*a<i��u��#����9w�$af8�@V)�L���%�M5]�RX�����qq�c6�W��g�T��QЛE�4���U��5�4�\�{�PK��`~�se���4�zR��F�x��de9�!�CSӆ�ؿ�r� jŽa^�4��L@�M�.մ �H72��0�L�t�O� 9'͕��e�<��Ţ�U
OP&��L��������+b�\��ԓ��5�ʯ�<}iKטΠ�
Z��ECo��y�^�2�hY���ӄ�/"�>x���4@��hΌ�\y������ud���1�8m1uJ�<#Ȭ*�I�NC���Swp��mtbiS�Q�:��,#�<�,��7�E?�ҋu!^���/J_z��.�dȭ��I�F���H�j=pچ������V�1G��JY��&ə���6Xn�b�&�dL�������G�rH��}G��1��8�f��:T���F�	�J�thNZ�A�eI3�%ڼK�y_�xZ2ٔ�]�I���b�$@���<�T-5��#�
��൶eW^R�r��s.��_�a)?Ky��0K"L�JǼ�*��
@�
�ִj�s0��D2����á�-,A�@s���]�S�ZU�=�O��LZ�������K(�,<��\�g�K/�k���e�~;�y����昸i�'����?�̝a�#ă-��ɸ����y/W�)�����k*����.�Y���� K/� Ҹ*d��;�-���P���{�����Ɛ����99_�����p�bw�R~�o ����#W�Q�\���L?1��"l(��U�&+[[�n�� ��5�f�p�aL�g�
-��䨙X��W�T��� �1�6��W�B����	/��5�' �b{��aă�� �3��"��^���y�=y�cR�����Oڟ-���on��!o� ��ʷ�6d�<�o� �?�a)����n�NZ�UN~�y��P�K��r�kG��i�K���5
7�1���A�q�z�ՖQ>@�PJ��ﮬ�I���*�0��H�:`��*a*�I����*��&�J�ݥu�NA��`���P��������'������	�O��80f�'��yX�ώ��|��1�/�ۘ�(RQ�|r��d�>�l��4:.�UK�����(@�:�օ+��p� ntJ�si��ᑴ?�Y�3~S��=�*� /V�@w<;	y���ȥL����:�����=�1�+�F�z�1Z�|+�W����2�KC�內tpb�e�]i)ϵzyڂSJ�T)�r�	���g�	�x��j�������U��!��u!��U����d<[@愩��͜RGQ����cat{�=��r;�OׄD�Z%� ����P����&���rYs�/� *L��i��;���M
�:�5�3���R��������X�,��o�ïfT5^� $�R�ˆ'<�����55����C���MK�����^F�2O��Ȼ{��?������'�1����P�F�ppO�G搝dH{��\�[�g��fz*�Q�:dY�!���A˃�~�L܉�Y�g��B"� /��0�(�5��3~�$-ٟ��^�<�}��W��~%嗞�ow�J��r�=�����ٳ0��쐏�pr���6v+#a��Z�S�_֣�/�M_
�Rj2��k�YZ�k�V@9�Ɖ��^f&G�9��b~Eo=�r�Jb�o|xX�W8�?34dZ�����S��������^Uh��҈�S�眰�b��K�(΍��)�h��_���O�|G��dʡ�ț�Z����'�G��(��!/�7[a8W�Mt$�rou��$@�~�ޯ�w�&�TEX�6���Z�2>����L���
��L���'>�P��&�p���Xn,�B&�/�2����Cna]*� Ro)����m��9EA�ky �.)WKA�H�����l��z�A$�d}�ғ���d (�U�S�8�����"{��;�p��!e��M�C����GW-����o��re�<0{�4��#v��*�.��w���a����7�$~�r������Z�\i���a�R��c��.�*�u���8�TYk�N�+]t�ca�<�۠D0�F�`�W���`<o_�7v|���%b(��C!ʷt�/^f�AWGopV�[D9Ԍ�rN;ky�}���:\(@ g�sh)ϖ)}&���/ݬ?�I��O[�3T�1����x���������	����?��_GK�iY�@�Jyj�E�΢$�!��j���7VN��v]��=4'�}����<3�Š$�r+�����[�𰹢�#-��w�i��!�ᮨK7�c� ,>w��*f
�*_��f1P)[�}|N�g퍖g+��*��.�� M3��+�Q��Kًd�k��/`i���b
C��2%��fF�z<'!M�,~'Tp�ך��F����C�- �s5�J�8�p��u�R^��а*}9P�e��_�}��s����1��DƨX%B^	M�)d|�.x&2�44�����Z9���u��?W&�\���s�֨���8�|�*/�+��D��a�7���S�V��K4��à�]X�^E�4�=�×N1ݹ	ce�g���!�n"��|�=��׶�[(P�UEp�ȭ[��`��.����xL �Y��TW朳ב�r5���^W_@8��+��+�e+���~4#���4X��S�s�nG��Ҫ'Xyl�p>=�(��X&;�Tx�B���0NGk��� �����x#|���[,S�U�:���:e��>�"M+�5L��:��Շ�,��E��HC��-e
��w�yB������׭[�`��<�烴��o���^w���¨|-�$C'e`����;۫��b52��R��Jyѵ��C���
��Z֌UF����yʏ�ՠ�ʪ��S6-�Q*�B<�rt�
�C˦UP#��N{�V����u��-�����P�5����H�i05T	}�*�%����d\KO 
�8�jG[�Ͻ�\�i�x[��*y�*����W����i�H� ) ���u�J�$��?m��i���{��_t��ex)���=�eGuV֘�QC>��h�	�֭��0q�e&����$#���~w�-�Z~ܝqz ��?; ��NXN�tp�9r��˷�5��!��ڃe�5�ж��Wy2;)g��P�Yը��6�o�tr*�r��'��&�E/�� ���$q�	�ϼ�Y�%��e􁇜z����!~P~�JlG�N��8^��L�r뭱KR����J�JD@���jN�Q��<� b�TH�>���$�]������cD��]���S����஄S{���f�0\琝qc�l�ާ��Dm��Y�{����8���_L�T�`h��Ĺ�{0���ߌ��毣�ovYb���9	��F�zC#{�F��a+�xz�bO�H���;O�g#FW͹��cV=>z
�.6o�MӠJ�VʇpI[��2KaӞzT8���״_w�ϭ�������S��<�@u���;D5�5���t%���>����[/w�vʇ�>a�x��"W�1:�_��<o_S�G���;�'4�����s�{Qd���~J�k˜�ʃ򛛲Z/RW �7|�p�Yn�{rr�������<�[7��T�����=��@bJ�8(b0��������W���,0Q�9D�p�,��E´I8�"��^�B)�/�ym0�peu�e�X�T �1�Բf����-��peȞ<�h[��vCk�<Z���o�Q�M���e	N]�|ѝ�߽��8�f��އOw��D �q�s���ȫJ�C�Z}7-�Ix$����h���ƅ��f�|�u�Q�f�e�"+=�<� x��E�o:���H���(���CfYaIPӲ!S�1��>Hj�,[��[Qāc'�9�<�R��3.�*o�\5�MZ��v�mhL�4(W�)�\H`��f�0��I>�������;�&tҒfC�B��<*����[�^�涽WyI����+g�z^<�V/ e1��� Y��tB�*�����KKS���u����*6\�r����\#�EG�`����/a�Z^rE���x�痮r�+� 
���We�l���
��-��tu�*�����#� ����iW=Ί���e�.ۚ�z�Kҿ�����w�}��1+�Rn}Ρ�1؄-�A�V__/�Lߴ��R�*b&�X���P���%��~��7�L\i���E�oX5t���V���H �%7=�`f���lo�N���9��h2̙Һ�T �3?�
�reM��t�N��
a@8�Z�
��r�d�)�4V~h�i ·B_��޼g�g���) �l��W#\����5�3����=��=|( z��sK�����_��k��X���"ܵ\c)�/���%`�O���y'-r�I�� �5�\+���[\<�|�F�`
w�'SP`�>��'~P��D�
oӨ�;�-_�2@���Wҙvh�{+d�D
t�V~��ɛ-�����C�|2%�}�(�����e�p�>��DY��<�u�ZpHH� 5��$P�o��8 �B_��ݙ�h���yD�g������Ջ������-�~ @�Z�`�+_b���4����!�G�����f�Q�J���&��!�X��G;�=�{dӋ��~�E�F�$6��)T'1%���R���bA+87��zFn�+�� Y(�݉�o��M�.�x�L=+�H�Y�P6�'*�7ZK��7h�����%񈳥�s�~�[?�9�i�J�D*��}Z|��(�x&����^�A�{sO�F&m飌�ܣ+y�4	�ÒZس�'���V*M�Q�]����O�q�kE$����".:���2�,v�t�:
�7yˎ���ʏ�9뢸Ha߮������Hbõ�/����7i�F�ʶ6�Xf�L�[^T�t�Q�JWAt8�tEDk���i��M��)']VK;�*����!�탑��*^�� \�Ϳu�.˧�ށp¿4�#��#�[f��:�� q��v������������2�"[*&���6tK��#�����y�����Z��;�[g?�)G˼h[BF!B����e�I��tQe�m�"EX����8�=��ܿ�t��W(�l��H=EN~���
p�̓�Y=�=H����7�p��'\ɱ�@>�l�7��#I��}����|�o��7q�]�Ɲx>e)[{ㄽ|3���4�+�j�R��p�q<�y�$����S��H���n����f~�}��4���(U�U�8*Q��ef�o��WF	!�
��B�ޕ1ϭ�Z���U�@�%��E���(\V:�Q���$Z�C�nR�{�|���o2���}p2�V��y�U`X*0�����lU�M�c�����LE�)(a~�u�*�k�u��f�zK+��z��n�@�(�	�$�@���D��/��_��-
� �K9�Kݽ�}JvX�i�K6|�R�TB0�Ok����)�M��%*a�Vޫ�É�M#3�,��M���]ivJU�+O7V�G�� �3:l��R��U8*^�����/^�^ms,��F�&��:W!+�H5[�a�ې�D�=崢]�8���dç]I��|O/�g�.�C��w�=�z�"̻֯�T>��@�'}�{�
�4����!C�ۻ�Ի;�l�X�ĝޤ�f�n��bp��r?��$N�bL��1,~ֳS���S���)CU�J��x�i�|�}��x�I�-R������L��f*��I�6�LK�
��.'4�o����������vYᵆR:�����`���>�V~�E�ݻ�A��Rhd��"�1vr=��uz�+l]����ÃR>\)��lˇ�������)��K��t�13�t�}v`�E��?��-����9>=��3B��	�+y`�"S����5�m:����e/;)+�i�u^�J������ MƮV[r�~�����a~�gʔt�@:����c7��i��]����z-��e|��2�Ľ|����~���{���hm�t4<ncڳ5F�ֱ�#�.����{�t��|:��8F�}��V�,� N�d$�PA4�P{��OǇ?�/m|���i/;�4c��%J�1� ��~�z�/���ѯ��<��W٦��Q޴��Qހ��N�����-0C��]�f��0�x�N��r!<�Jgl���ER�U�p'�!����g�����C?�e�3��������dqW���EӰ��e���n�JŰ�LJ�a��*���8�����;.>���|���%&�~Sy*2L��͐�.f5�+��Wq���x�p��Q�HLah�P����n҇X"��`ٯ��+Dy��sh&�1�"�jP�"u�d�g+\c��/��|�5)ZѫR�a������y�� �}-1&�0w�$U�ϟ+�d��.s��i�IZ�`�?�� �
�"��_0:�z�c�q|�pSi�ԋ�H7�'�;���ʐ[CA�e��(�h�T��u��i���o�ij30�!=-`I[ɪ7N�E匣�������G�4�GX�\�c�9-�T��t�:��!(Z�E�.�E��E�(�}�h�,}v
@�%�(A�p(�j��g��k��]��s��e�0=ARP�JZ�O��G(�[�QA`ݴa#d3A;J�N=�8��m]��Q�ꢑ�i�I t4}�����(�O�
#n����$Jkӱ~�&�*_s"��L��6r58� &h^K�>�o�8�]|��E���� N<%�y
�}��������ha�8�62g9sF��&Y��N��~�iΔ\el�&T�0�tT�r@���Qv��$ ���#�>c��&�Ĺ��V�ݝ��ﻗ��u���l��>r�	�v&��������1������(U���O��b�6����O�Wa�U��mvv��\��P�zE��CG~�Z0����/�������	���q�i�]��� ��.����FM��A� �X�p\@F��x��E ���Rגps����L���~��n��?�=�Nڄ��X����-߶�^��x�[*R��x\bN�ְ��)��k����t"�/"�dU�^
̴*'�:qM$W��rh2!s�(��8�-�`�k�� �V�#�8���i�Je�ۗ��6�[8�U���E�pN���'u�̅������s2�X���7Q&O�����;O��L�C9�pL�澒W%/Eu�8y7n� O]��Y��y�Ŗ�m�4�~���#��0�E�;�*J�CvНeB���
u�LO^)����04 �P�%I3�
�3Fd���m���B�D
5�,	o�:�[����A�L(N��.�Y�أ��=<�x6�gM��_������wX��!�34��s��3��ظ*tm���ڠ�0����M;?<��R^1Y��8)��!��L8��	����-�W�2Qv�69�Axa�zJ���%�$�|%�/����c1�c���N0�S����^�;��:�����k1���bp�n���a�z��Ui,�2�~-��;A�g#��m �47�>�2Vc�<q��
����2t���@ ���5�ʞg���P���?�tF���^��T���f^���� z��
���zXs�D���sb��t��� ̓�pI�򺊟�Ϫ�.i��s���!̣��X9��[vT�2�Z|f��1U�F�ɠf7��~u�x6+X&��|���M`��^�������Aw2�g����c�#	lx�(pt�N�S�5�"y����t͓�˕Ӭ�c.��̏Sv+�G)��C�	  @ IDAT<�������g,�+9K���6[�`u-K�ꡂ�:������eY��)��w��Ho��;K�����׿������㇡�~���/_����y���S�����P��$����Zg������a~~e����S�U��VZ�r�X>}�p���<�2�S�(����bE9��<Gvy����c��Ő8��i8�B��Iq��!��N1��s�|\�7��Z8�bꈕG�H#hӋ1|R%����#��>�K;��	���՝7�~u&�[�H�.N�
��	;	:��o~Lc���wW���R�&���+��l?拓�~�s�]�{Ϻu��&�	��.9��T��=��
1�C�o�֢Z��bf[L��>���rչ@'-�c��2v�z�J�|��h����k��&g�>x����ӧO�I���<2$r����D��*��O��2�������xW���:��lKQ�$D����U��P�U�+� �������K.�s>���r������a���(�A�瘫�Ɨ�����gG݈ w�;�^�h�]LOE����P*\���",:f��f1�=��W��%���\܆Qrs~�vA;�z΁�6>��Y����^2��}&E{��V�*�J�L�j1�
l�P�2�t���9������~�w�Ӛ�#0A^"��o�T�X��.&�+`T�[�0G�#���P�O�\t��V�{K� R�Zt
|��&�C�X�����<C�a�u���帹��9�ö�.�y�3�'?&_>&�\��4�ho)�.�����.���gh_���3��9�������L5�|�"��Ĵ_Ӑg7s�
��S�/����%��\a�Cr��%"-��3��T]L=��J��=���eM�!H���!{�kz\Ē�^�iCZ!�"XȜy�p����y�a��!���)@s��������jA�G��)oX��Z�Lg)��c�o�E^��|C�L�����\X���V�4�
�P�|����M:؛UIU�WKUmX!+U�>��3�5�K�È���c�(��{ד�US�g���Iў�1C��54����>�=~�š�OG�<�x�2W!�j����QW_:�̣h\��C�*��T�:�"�vcsHY?�
_qvύ���hk��j�{��'�,�NЀ����1��G�����#�|��F���
Rk],�22�h���B��֗�2�J˧u����I�B���
���(�em�C݀.�U����t8�ő�=T}���~�s:��͆��R� ������l����aS���`G©�u�Bfh���n�̴�[����>Ci]�I�3�����"b</�R,�ks�#g�矋���0��������Q:"�Y���<��E�3����	���c����l-��HW�LS<�¿aa!�y3O|��P~Z�)�.j�A���]�o��P�m�ܲ��P�*c�lرA��)zQ��PR��\�Wwi.;!c�r��N߼;\�݌�i�n�d�I���n� DL�c�M\�:��)'�t�a;��d�ૂT�z4]`QT|�������Z�4��Qp��wW~5zE��-���cX�0b�ӎ hV0� ]�w��ez	�Q>�A�8w�'��8���*/���.G�[ˌ���XT²�u�$�D`H-�&J�K�dP��\&1�=��o~��U�A��
��!����(���9�P�6�*�68*�N�?b�d����\��ByN����>�"�,�W����U!�B����r�ڡ"�u�w+M6�L��
��,CL(�(#)�.��U|��b��4U��J/�FNk���$�9�]���!u�	�k�z��5zӃMHUM����y�k�X�i��?�ՎcGX⭻yrBwP�>i>y�9LZis��u!ʗ�%x�-�l�TL��){�9g�f>�1@��@Zu��	Ap�LI���.]�A�w�Q0+��:��uV8|3��W��t'�U`W�L�������+�l��"H?Y�6��!;�T���y��RVq_R^��5WM�~�:��\�*aUlVQ����0��)'=��8��;�g���ڦe�'� LG�_�:�(ǽŨ8:�F�'(Æ�--�t�鈪�9wm��~zư$Ï�?�����9=f;�S�� �}�9:`J�×����x�]�1����*�'^�NɄy��F̹9ީG�\�	+M�e���tN�e��E�,8��K��*8�q�Ԧ�����w	�>��[h���g2�`^�6�y�%��)��{*�j��rV�^�;
c�G9wX\�b\��2)�Y�-��w������D_|�#��1�'�����Nt���[����!�""�J����%�F����O����𼷰�Y)<�3)fQo�&���l�bE�vb���Q�)��$�b%�Ғ#}�%iTu׊W#��]���=yDE̅���N7���<�u�k �8Y}e�m�m*�Ѳ�@A
�R�Q��J��_��S"2
�X�@*DIHIP�NL2'5F/W#��DmU�)�����I���3�)B�	�ni��s�s��[�VP��&��kCaf�8f��"fMh����Ƃ��$#b�`1_�7~�q�8�H��zƥ����KD��Yr%n�&��G���{O&i�ܭ8=�����������j�EZ%p$.���U��-��d�Fd7�u勓�ܰ�}�ΨO\����i�%��w]z�
�z�!S�kY�/gy����x1�NX'���w[
����b��bv�<�xše��I?���n��UP
���Q.�4i�ŭ��W��w�l�^�[8�y��������9'�%��6.�^�Q^�*ssۄ�J���̈́yE�VmJp�N��z�?�V���d#H0��l��wd�q�zQ��� ,�#����3m�r����0Oϗ�0���EFp[�آ�9f~+=Y'���'����/�l]�8G�#/�A�$hZ�Wq��3}�c��/�Z��%�I�**X�Q���'�;\��Gly��K��YU��h k�S�N��}�E���r�7�Qْ��S��9:5O�xX��f�{df�k��|�����cM��Փ�ig�0r�_���F�O��nZ��%�KgY1���t
��	;�ge7��E�1Ws�]!O�𥝓K���@3�Gd|.�-8���N�f���\:�rNY�{:Q��&�g�x`���i��ƏVN�2��KK�<'�*�?\bJ�lX�#F��8�����9\�]���M�'xqjmr�-�e*|%���L��z5\�M��"eĔ�8܆S(�X�o3��Fe���ֈ�LӸ�
�4p���o2��z3�[4��G���㌕��U�I۲�U�⛄h��U��������/M>�˦������w8W؝*lv�K��GV���~�)���c�Wo��y����{3bx򌥓h�N ��I���$*��^T*�ĶBH����LU�"D���k	`�̔�2F�N̒�������s�q�p7���,�jP��� &/�wނ�4��3!~�M2M�U �����"c�2�%��V���gኈĝ<��A&�P(���c!渭^��n�^L���-]�)*�1��(�����C�7���}0R2�Ҟ>l�!Q.�MhT���a���O.r�['p���Q�Ί{e
(��A�d�P��˔�VU�$*E���:��*]z7�F�Z�j�2fe ��Zuo�z@c���[�����������6?�����ZD�>Û,f��v9���p똂H��#)f�vl�.����/m�>u���OG_|�	<:7z���4�@>�<y4z�Dl�����!��X�qϱ�����������ҥ5:����Y][!I�C6v���=��I��4OZLdmu%�ZJ9QH�\p� W�!r�Z�K����c	 q��
���}�݂�-G�;�+��Z(q(�x����E��'��'t˺�_��
GH	�,�¤e�2�~Z��]^�K��
֟+�]f^ز�C�SxI�Hl{�5qbvx~�6�R9N�>�F S��;�X\��D@��g+���4c8���[\P�'𖊯��i������L=Fa�����&�)w�����[��G�Oe?(�龅Z����9_o^�ʞfN�  [C�8fu��I�"O=�_�hص �|iͮ����*�6Ş����u�Q!�-�l���	-X����ॷ�_-{�c�q�r��X��'���-Z��G=�k�Ja���kczz	���r�uU�[N����zgR5��o�ߍfI#xZ����tΰl�?���"��3'X2)����h��p�Y '��htK�M�_��>P��/�R��#l�����k��"w�2'B,��d̼�uŜs״t*O��<��^����U��"Pf�o����/�+D�tSo��(�'WDL6>�T#��D��H�Um�w�=�{_�E�'y�D���N0Sy��R�������h���G8���DY�4�Z,B�0�b����oÕ��X]�&�O\>JP���-&MAH0~�bg{�V
�8A˼�0-xfT��M#�۹Fj�N�u��#c�t�N�g�3�i��lq*0o�
?�vf�9c�V8��?h��R�����W3��`]K|C2�ҀO��{�k���3�ӻB;W�Ѿ�����p<~�3��E5XZ�N>��)+e�6D\�Q��ZrK�Syi��f�n��{ϭϡL�Y���
!��Ve�	�0�����W���m��;�'�]�fc�p��2GIq����=��L^����ȡT��{��}ˤR����mh�]�<�)a;�a�Z����+����ѯ�l��y>
�Y��8���W��3lysΩ
�b}�:Z�w��0[G�y����C�aK88��ˈ*����8��I����0uΞ�8Rn��{���\���CfdH��^���B�`�u��X�ģs��R��AE��^�� !��I��N��R�G��=�?r����#�����]����(8/qqޕ��T��S˖�"
�|���S	�Z���9��}�a�����
U�$qRΙS5{��Q�+G�c8ǻ�=6�̈���UA��rK�v��&�./9+
���~S �`�)��O�X"��t�z��e�P�MCK��{;ƒ�<��G�̑T��#m:���Q1ss�O?I�Y�'�1�c�(y�Cؤi���U���݋�n9��uGG�-� �
o D8hW��A�X���Y�zm��0�t�NZ��g0 n�۳#X�+Ͽ���,���@Z�$%?���;N�?��Iٺ��JEY����iJl��O����bM�itkI��|,?+cfi�ń�΃�-��.�pջܑ�@X4a�/��ʁi���UgJ�6BL�*��aZ9L�.�|x'p�o7iIG��g�z�ş�P �#;�s��Ӵ�#W�38��B��"��H��Jd*G�����y�U���bf�Ƈ�
N�	���{V*���"�|rWa��W��8IB\C��B)3�DJp������ѿ�Ht�֍RH�(�vo̼� dF����U�ăg�;��h�C�Ŭ�"�$��o$�^���&����t��@
`��P�U�!��#�!�P��+o�]R1A���7�ׯΨ����|S){�$SUv�������_�PvZ�WP�4��⌛���ZA����$�'`C���Q&���*A��8-<V-WǬ1��&￧�X�=7�ɜ�0b���kVm^��1���'���3V�=���ѧ�}�5�X�s��Wf�;�t�d�$�����������F����6��o�隓!�x����P�z��R����Ŝ��T� ~6Yt��c���mg��`Jr�-6t�5��5A�m<��pX�Fv�g�l�e%{LQ��sz��s�B�1V���|��P�|f���4�|G� �+����/ӻ���Ď��=V<{�I���9���;K=�U8Z��@�4-/� 8oK��p�T�d��"hI :2 ��#h<"<�òt�]�'hC�Ρ�9KIS�+ݲ�=C�*MIj!�V�:L����_1�=-l(�����U�G��0BN�p���š��RI��R�w����y�|ߺXr@��t'�K�����_�\�	Ƀy�r'�dI����u"�ə�Wu�q�ۭY��]`���";5�K�\	�a��R��7%,o���Gv�W�P���/�����=��C`���4���k@��0��O������4��
��3��
M�I��v>���ڎt�����8�l<*��r�I��T���Quj�2w�(��	���|���%��"Y�h�/4�Po#��ٕ�/D��w��m;�m�>���]��M���5n��I�l߾�/
o<g�����2#[X)������;�}��"q�5�TÏJ��/�CtTAaR&�����R�";��~!׸Y)�P|��-�~�)Z��n�s���հ"��⭗�����h���U���;� d�J��T�6�9_/�-Z�0��-��p�E�/�N�`��k̗�Gu�ZB6T�]Dy~s�hx�0]|+D���2ż5�~u*�ݭ��F�ig��7][��^�-x�7zt��� ����s�n�͵He~���!�1�/��`�n�����n��|	���/q���,?���h����I������y�-{�����A�Z2<��YW��N�]%���Z��8����g[~�!�1���_}��m�_�b�ڛI�d�ek\�(�Q�Q]u��!C�Ϟ2��$B��Is����p���`�s{-D������C��|g�I�=Jߪ��0��)/��$O��S�ɡ2O��8F4�FS��J�d�r�ޫ�K^5ꭸ�@W}��tKX�q w	n�u�$;T�Maw3�q�A�(�6m0�
�[�d��fcN�_� �,��,1<�B6X�Lw�"N�Y˷
��[���z��K�2��V^p�?7��X��-,4�$�ȇ��In���k�=�J~ĊE���W�:Qe���F7�-����G��Cn;}�Un]9)^�8$�t(�}����`�y/-3�B���7.�0۰�	*z*c�_7��T���q�v���c
r�̑j�z�����uZk���l���EVNn��J_����A����"L�Cw�)��/�U����k���쎼w珁ji�N�T���$����ݹ�����;�^�!
��L���׊å8/%���C�a7z��^��#/;]=/>�*���W�(S
�uY��M��!l�'%gy7q_���&��~ϋ1�{��x�I�z4�ɏ�n��e8�M��7�3s�PҲ�
�=�)��,s�ފu���/�����3��NQ@���I��r��;���%������z�x��2���E�dG���څ<O+@�_B�mn�k�F��FA1�������a�#B�q�+8�V.2�2�9f�qn�%���*��L�ЄY,`�[�U:�U~��&<|m���6�^6䮂HO=.��|����ܥI��q���}۷3����u7���ۡ���r1��z9�r�G�'��VPT���K�TB�(4`s���>�����/�oJZ˨?�5��6av�lfP�M׆v�)�br���U�S��w���7V3���+L�ײ�0l�����8����x�Q'C>��Rxi�1}���ĺ�𫍺Ã�Pm\�H��
�G6	�ߘZx��"s� α)�C���a� ��PVǔD�
������<Je��蜠K�;�����A��Xj�p������(��vn,����3N��ED�Y%@7U�`��t��j��N��x�(:�&�������@�UiގJX6vl�[��U��_�f��{&�GX�R�L��J��-��76S�(s���"O�s�crw��{ǔ�1Ri�#
�
�d���3���<TȴD�ܤq�"�Ȫjy����y�e�ZΞ>y:z�VXOc���T��E۽��r���QkH�9:��n�c��R�JYY����^d�]T�6�s,�.n�����cxm�|�G1�ꫂw��z-9��n0vV�k��sq���+s��rʅ�v�J�u8����ȑK�a8Q��(��r.��^���`�����4K���ds�m�/\����3�����v��W�;q���S�ihtߕ2�ν-��I�R��<��"C����{p�]�zZϝ#���ey;�?�Yv��2��bqQ�[X�9{����Goa-I�F�%nB�L�*K�{^�/�
W���_*_��l攑G�e��4�?	�hɴ ��B%��3
7�ޢv<����ė��7���!��DV��
f9�u���_����˹��b!r~�)����� l�D��On���F�5�J.��lȖ)_�Ջ'�+��3��:�j�f��C[�*{@�FH�[i%�+/~�h��a��V3�v�w��B� �j�N��.�z��MО	=�7C�O/���#������}Ѥ��XC����~���B�~��[\}����S�Flh/�vƤ������4��.���w��ET�h�G���ִ��B#d��ңEC{���#��.�_3�����WvZ���q�&WUڨfxJؤ眘U`��։�b�`��o���Ӌ2}"��X����E��J��uIEjJ 1���Ma(�)��݉����2U�֕ޱiÅ���'��\ƪ� ��e��]�[ښ��U�qr�CoZ;l��E��Js�&�U��R���������Ai3v�*ʸ᭵�+9�?*3o92j�{��v��r�L��z)r΢x�S�$	�4�0��<���l�������B��7��\�@�x��w���ٞ�y�|��LR9���M�������J��"J�
�:s厗L~�$x{��D椩 ڸ�n�"���ʣ�BEʺw��=-���JV{����!V{���8����ڲ�E�W���������a�W��JeW\ݪ#��1<%��2�"�>�\���#n�3/B�������O{X�qǃ0���O���!�ƭ��G���[x׽��§����*�=!��qO�r�x�U>큄P�m@�W�Mz+�����Bw�9�Hݸ
W��Λ8Z7oڐ�r,�#q�%�QnK'��*+�KuU�i���pMֿ��x����?��Q�_���8�^��Ɉ	U9M�J��Q߁��@@e����M]�J�\��E�`�Sc6�:�fn����O�W���/Qb\-(�/9ت{J�����{Ĝ����i�p�)�Z�z�;a$Se�0E4�A�r�g�Tx���	�@�b���k�ڙ4��)<b�9<W݌�*��)�n�x����2&�A�a
�����N~� ����d��7n5���{�	�{+0�
�tϜ��c�?��!����꠻9V���C���i5�5�Tx����ع50���z�]b��Z�����d���	E�F�%�d�0��v�EũJ��}>��������6�n��q0�T4+���+�P�2g>���!� \��Fy�P3_%����!e��bxR˖�}�{�/�0Fc8�����=���նK�����]^ƛK�+���k�l����E,~6�*K~;�f��� F���FE�׏��Q��9�1mw�I�X���uRZi�����:�n�"Lc�E+Op8K�`���b�q3$ʇ)�c�o��֯mҫn��.��n�r����r�������f9�p�H	\+�����y{_}�U�qX�����Όx@��\<�G�]�,��&��Z���g���!V�2,���ZOQ�aY;��c,R�"-X���ꐡJ�C���uL���ZF͏��rq�ۡU���d�<.�>4]h�W�L)����)�>�O%���C,bnY�Lw1���(�P�<`^��"im�?]<�̆x�0g�vã����m0T�s�xd�e�|��G�\ }�1�)�<eA^��´~pM�Sw����[~�&������\?3��)�~��G��j���8O�=�׍,��,N()��0	X�0�Ϡ��Ʒ��o<�OK�s����x�g��f�#�ұ���0�2:2U���:�s�%�P:	*c��i\�PB�}��(JU���(�(�Z8�=��4>??n�HBʜ��z�¥���u5�)�s%���w�[�̀��X�T���fs��Œtɸ�%C��'��
�G4��!᜼*0� E�2F�U���Jh6��$[��q��a|�u��%ါ�ˀś�B�T^2_�X
5ܢ|�s��q�C@8A�PM��Y5*�1ްY�Lǌ��+2��������K�����:��>>.'�|?q�b/�e�ƿu�����ʵ`�����H׺�b��{���S��?<�^��y��wOa*(N<�]��R��R���c��;g��y�~c��ٴZU�����^���ߜ;cn/��?r�=����X��L)X��t[*��g1����|l��<�H�|F7�]��k��c�����z�d���� �*PX�b�w���0筩 F+��ʃyQ�9������q��Y��Uw{(]�ws��[�0�d�
�JzQ�+4�[( 漀���� \Co'�GY#X���D�!�g��-��^k�sM��_��}�6&-�Q6yz���������kaW	u�O�,�)7h�"~�vږ��� ?�RCJ�o�
��7����y����!AP��6F_|�eVQ����_��mV���������&�o�2�,���
X:�
z���)>%�e��.�5>|?�<Q��ێwyM�t�ʛ<��G�����wD\�#�*\�_�,ӱ�Qquޚ��8�G�`%nǈe�Z���C��i��[i��XC�6Ɲ�аk�d�e�,rIyI^Oߒ{qK�R��O|yN_ݭ=��ם�w�ƻ0�eq+H�(���Sߺ�t�=�[P?�)����Qh*���%��B�mh��X��7qr�(*`�<eG�z2\��em�O���T��o�_��YzC:�$����B�<ʰ)0e����Q�R��˻��T�I����D�#fӗ��mrKG����U9@Z���s�<�(��)yx#��}�����H������!�����f��?��y���њ���;Z��ū�p���
�~$￱�Y#� <��3�
�ʌ�[6���V		^VPw��Ԑ#���e"��/�!���M��A���k�ořh�� )$�5�?r��>�
��%7�kx�����?}��\MG�w+h�!�|n�ƹ���Cp���O�:D�JE��d/iŕrh�oU�u��������⶧}�*�����2���>�>�~q�er����@) dZ�W�\,.��W�T��T
 ���s�JH�6�<�e��0�%�۩�ĸ	��܇�4nZĚ�E��ə����m=8e����\�!-��X ��� K��1�FP�	�w���pс�����R�V�D&���z��˾h(;*����aGt��R	�r��ƣoQ��V��*�z�:;]�M��x���-
�>��@Y닖�(�H[砪�ZԖyd��m?�H��y�Ù��_�x9�
���+Kq�n�0���$��a�G�Xy� -<���&�V2�$5�(ʔ�V�t�:_Z��G�(��#�����
�
�_~�0��>xo̠0��0�8�T�ʒJ�2�-�X�D"�3��$D���S ;*/�>O�o�tu8TE�y�%�Re�vC*U�[~���?`���h� �;��a%頕0�i;d�6%9��=�C�`�?8����b���8����rX��k�bQd:��!yZ7ml�4XU�{}��D��<������ýWB�S�Mwrߍ�c��%�?��u9E��*����{�����=�I�n�������y�� ���y� ���H�����&,놊�7�`Qx�p�h.����I?��≿B�����P?�-
������L��t�t�I�l+C��F	ғ�8yU84u8�P�������Pf�_�ބ�����&�ZJRI����zf��y���>�����V���M")�~�@�M^Q*Uwό��̛�@  �@`[�B���C�T}�޸O�ENk dC%�4��jM����P[k�cX�TH֨k��7�([����`�Y�U��4�+(ꃘP�$N63��w��tX�-���"�D␫���L C T^D)��N$X��Vh`��#l��RL��-=�L�K� n�If.�ڣ��~��w1x�|��t-�No�i|��$�q����MJ����k��?礟���NKR|��6ïO8�ރfݽLsx��e�qhǣ�d�7Cz�	bѯ��7�Nx��U�K`�?6���訴�yiup�A�'����H-�m8h�_�p�V˲���m�{_�]�07	v���pV�Q&?�g�(����O�c�p�iq���n�z�~�D�ȹycA����6�7#~�!⏰�<��c�۹Hz�B�匴:J�Qnғ�>�WlӪ�ee�!y�e������?܂��([O�R��ÇXi��@Qʜ��աXP��G�^�0`\�B���G��P91>CR�,��d�L���e�Vh�q�8��+�~i�q��]����О��"�_������ИuQE�"�&�k̡�~�����G�vJ x�w�N��,�d�:�W��[�Kˮ�lr���cd�nv�=)Ak�:�;�/~'�{\�gCZ6/��@áa紒��il���D�s���g*��x�%o?ePe�C���?�40�E�lܿ����}1�^����E�r��ʺ
��.y#.�W�����{@��<�/e5�Z/���WƓ$\���4�겔��~Z���w8�	��.������ʿ݅\�(��n��Q!NÞLF�W�i��n�6�U�V��-�I������N�f�zaS�'��4�ַ��y©���L� c���H<��d�&o��=xB��Y����7V���<.Y�jZ @�js������-lp�Seh�-�� �?.^�ֳ�4?��д�� ".)�=_D�|Q	sZ��Nb��棢���i)B�Ըk+}-lS����J�L��y&�;��JzfT4���H��:
�-�4���4.�Œһ�O���|4��4�O�8��jC�R���pf��x�Z ͥ<� I�',T��K�|7T�9Ay����3h4X#I��hK�tx���R������2�%�"%��G���8���`���(N���aa��i>
�wi _��|�*�'p����(�@U���L��l��� � �A��E����Z'�8{q6�/j�B����Vmi���FNE�<����b�2�{�QX�X9r�;��C+��\̿���h�t�����_�e�7V�V7��e"�CC*~�����]"��y�Z�Fc���(jwƪ�UW�h���e��J�su\�����|8�����(_(#�+F���]z��{����������Z�����#k�UH�`��@�Ų፲�����0��!
��:��ۙd��M�C�. �aL8���e�1Q$�W�rHԸU��d�qF�^Z�����,e�8-	C�U:�g�$e�<�l�lo��>%�SB\� �O(P	��OQ����[(QQVwsF�{hş�졸܅ZJ���o�5�4��{w�w����/�0jQ$��I���%�V-X}��6_������8?͉�7aw�����/�ۆ�tA�)Q��̈́��
�~�tOZ)d�9Ԩ��9lX�\uk��`���y�p	��5�w�W΃Tv{���Ǭ¼��IVc]�ynLL��G�<4���o���S�n�-x������D��A��^ᛙ|���(��=�u��c��uft+�|�K�||����@��q$�Oma��n<R��Ye!�,���=�򵼚&� n�_,�K�7݅���*;U�*=�v,��2��ÐD	Ǻ�+5�N�t\�b�gT����qgVn�f��vg%�\6Hd����90,�9&�5掹9��Fk7j���^B*Aw�C,��ӈ/I��x.�!�)<t�������e����WD,i�Y>%�XZ�DW背XG$Gz}�Ϗ�*���'�1��,���yDI� \�h��t����䪸 �ѵ�w��
n+x볉9Ư)��^��1Ij��>�fI`�=�rU���������˥~qOE	*�!���H��0��l@]���ee�%���!�]�Y�m�z|��������������qC��@Ėg���
w������x��PE�>�;�H��]���]g;���,�p��6{���1�	6����l�n������Y�#NSoi���%\�A��02G%�9���~*)9
k�gɩ,(�T�乊��Jў��@�;�P-iZM<�С�7����i�6��Ul��H7��ѐ~H�ߔ���PN��=���Yҫ�ʉ��O��EY��N���Q����)��i�H�K{Y�k�CY��Ή��Se�H������6���nݺ�4h�{���S9d)O\�bYQ>�~-�Nܵbޙ��[>����X�\!j>	�,��`�T�a�zDZ�P�%�eS�t �+��B�-�H��Gn(|��6��-��ӑq(Z:Q(Q��n 4�0j�d�Ľ�Ol�J!uk�"��k��.H���<
��q��Ni�|�p����K�~?'GW�W��6���쯉�vx+���;��6�R$xJ�|�	����/}��,>i�T���`���S���ԣV#����Px��I��I��׋8*��}:��=u:�'aD����&Xx���d��)*���t���?n�ފ�'.�&Q��뭺�D{������jt?�0;��Z{�8�`�V��4#���E�)&���J�PL1���̏0���	d��(��Vڦ�T�DW�|欱��B5(O��N�Y���sq!$x�����?�&m�����І��T`�^�E�I�Y� ��o�G���^�&_����]4�p�a(�%�!�����3@sG��g�^���S�^�˼Q�P	P�p���cn��^{rm�J>ʼs���0���B9�F넸����?��0��ǹ4/�9��������5Y�1�dk��Xe^�a(���+�����qe�o�D�������[��^e2�CAY�}���٘�Zo�mT
�N*��l�L����k�{ŘсCG</^�j�`��>�t�	���**6��g�SQ�a(�ź��̂��!/�rh�\�h����9�빕���!	O>����R�͛�k��|	� �B�C�>��W��D��)�
I)��c�U´�E�D~9Q>�λ���/#9��r�����ý������a�W��¿������2h����ȅkl����A����-��%ʞ�\Vؓ����ĭC�
�N�Se���-�l�*Hy��eYq��Û>���٧�r�(a7�&�,]3���V��P;.�m2�h ز|`O}��ҵu�}�vXA��������#/��C��O�_����n3�G�֛�����^	8��p��~�i��7����w]	��T�	?�}5���^� �5��%6ߪ%�a��-�'LQ�O���7:�qt�<��JO���]�X�b����2�� z��zY.qUX��]��	��4���! �*�
~tz�-��
Gu�s�c��-�<�������9A�������鯛�a���(��h���ʙO	�5g����2οAe�ت"���@������z���p7WcУ���J��d���-�{�����:��d
z��+e�G�e8�
.1���W��,��`^I	� ��eP��H)rW<�?	p�������~�)=��"6>���k����3�3��
��$IK�Ǭ��⶟�R�� 6������6��a��4�P��s��<��7of��74</-��^��*⇖ z-5Mjٰ���9���Jm�b�C�1�ĩRᐟ�6}�
WR�Ӹk5r�����?*d7�ب����v���b "tb�:�h�Kο��yb�Җ,6�.m��C<�L��%ånș���8'Z���̕2}�ByUDeb6����J�O�d0�
N�94��k-8�O��2�UC�:~�)Y�/�|�'�G� p�k�.L�8�12y���Y�ě�L0��X��F�  @ IDAT�p�~:'L��ʀx��a��>e�C����l��ql΃sQ�s�]�qa��(�*�Z�\�aNO�8:�9e��r|iϮ�(<��e�T���I��3��������믿�*u-J�yh�P�����?�����t�j-�������Y>��/{�1�/'ؗB��1Z_P�?!Ml�A6tx�֝{�WvHp�Z�e�Xo�_���g~�k�=��+��Kl'B��I�)���^`�o>�[+�)�M��2�:��o]s��� �p��3@�B�W8��^K�|���`��)�鉯����SѢ;��B��\�����4�^᭏*�N��n|��AU�w�ѝ�޺ǕG���-Q pR$��Q�	R.#r���;��M�
�������@:�4��N 1����2WÏ�B'�{9]��\U�0Ь|S�s��o�`~�G�˩�|g��<鑃%g*��d�0l ��V9�ŕ�~ES<MV祙�W�Ya�X�.�2�\�P�z�S��NO�L;g�E ���KJ�]t����Ygn"6�Q0߁��%��i�B�#��p6v�n	��8����u�w��g���8�_g�?�R����e��lX>���N�`����u��Bm��Zb�F�ñ���6�
?w���ok��ȹ4L��6�&�U�f�T� ��а:��I�{Z P�ldP��@KT=s�"և(_4H6�$��ĖW.�0G��C*$�(��}���)P �<�G[��Q�Tشܹ������-~��"�����S���~O�K�!Á�X=�4���,����ů�{���gX��CT���c�Sx�Z�vݎ�D~���2��f�W���>gx�%s�ܴUE�kQ78D���9{�<wR�
��^K�a������w���Z��H-x�\���7�8�&�.p�SEˡ6-3*�Γ2�zB���V��R�Ѫ��'77H�a
v(V>��m�}/0��ϰN2'�2�6�s��Z�,'ZA]P�Z������&��Z�� �O��	��~����������/P�v���ǜ���%��8ܭ�s���������_����r�	7:gO넖2Onp����l��T���Z���]���ˬ{�����������?��Ń'ϣ|�cΰ
���.w$��L���|Ew�_[c51�We�֩/�2�%�wv@��M����(.�\}�����}�����3B�ZTe����"4����\?+#&Q ���/p�.e��i/E�8"������;ﶼ�q����<ʂ����z[��^#�U9�o\}�+q��{��,���FU$���?��H�x������
ݍF�b��B��+ɦڎ��K�Q����F��g���I����~����{�j~��4�TztY^�w������	7 ��m��$p!I� ��46.��^�P�����Q�w^�b�o��yq�E��La�XH��ӿb0�x�p���?���!;��o������/�׻���-���#Ԓ�UI?�)_��t>���HT0�Q��Q��Ň|I<z�G�f����D��ү.��2��㐏�'�Լ({m�q�l��|��k,�?`Ɂ�Q/�2	Z��J�b�),Y����zw��h�T�T�T�ܨ�vHwWq6(�|���똰/c��쓛l����L��}�F���o��%Ò�Cl14���O+8�$2���K�k�`�I���t�eycC�&���<���.2č��3��3W�V�ܼB#|��)]�)_�@��� 7_1Dec��\����NW�,~��obIy����Ⱖ8��x���<�Z��a8��?��b-����<7#�ƺ�^\n��*W�^c�O�H�6�1Qn(���'7� ����wc�R	T�VqR�<&N-x������4�U�TԜ|�b"���p��WV��_?���bW����fn�&G��×���@�HD0kY����6J.�dx�->�6�����YA�Rm��r������*�*��X-i/�!�^uk�o��k(sW��᧿�aU�kc�s����@��;�x���.z��O�Ҷ���ᖢ'���I����C��_�7��x��(%<����i�Î�����8�iy��y�˧�ے��K8+�����l~Tv+x:�z�|�	���оB􍷡F����<#�>$`��DV�D���L<�ҡ�Cs"�Z��,���Dk^�Y�ŋ��:ܒ����)��M�5\:��6m�'Y�xq�򦿰�4���'���YXe�P�/��{ß
����#i�'���b��x �?!+;)��k�
����f`O�1V%�M��6��Sq�\�Ξ^'ZȪ�Iذ���(k"���*Lpb��a#)|]���*8��%��
tk��T�B��J���)\ϸIIe���{��	Y1��q����-f�P�|�a�'ĉ����J<N��F,�n�	�̭����0�|܇��G���?�Gz��w���aG�t��Ӕ����'�u3KN]#_T>:��*	!%�*=�H{˟HP�h\y�@�a#~5� Z��w�n�>���˘T:�6>-`���QӒ�'�����i�n/�PD�*Yc�hy�v����]�0J{�[���ܛ������r������ɷ߁�'�&���A��x���x�d����(^5g�yKXa�֒g�v?�pk���{�^aZ��|�c|l���E}wz��),�C:f���kve>f��!�p�m*`Mr�l���mP��ˡ��M��Z���9W�P��4��\�M{Ncm������&��6�Zh�`*���w,��ʯ�T�`S�Q�se�e�<}��Y�t~X��s�9,�0do��<e8�yx*xʉ�u�V����;w��{�p\�]�8�{�^^W�S�V��D�G��Dy6��~G�ց�ۉ�
�CޗQvM�!�S-�wYT��l߉�(��g��y��V87|u���;L|���Xl8ja"P�gEK���<e8��Т앇�3
��<8w���m������Owa��\Tj��6�l�0q5.�S���EڴcA="�'�j<�.}I��+���r��W�LW_:p��|�,Օ���k�3���u��8��xW�&�)�Ͼ4�<���O`� V��aN���w���b�_�H�q�l���4\Q"{;	O[`��9��(;���#A�qXx�n�y*B�/*�{�կ^���ɋ�I�;ʚ�Y'}xv\�7?�O߸D_���I�(d����(��Vmu혮�.۩��	��,���|����i��X$Q�(�FS��0IL�HƷ~}�u$�8���l ���M����er��� ܔ�@�g��/�U�x�~%&�q�0�vT�ߦ���q��5�0&n�}�E{��\��8y5]K��G�M@g���&�8����+D���<5��9�O%*[*4*)���
1�<�S��rR<#�)��5��+T��3ɗ���N�ԭ4�@8q>+(�4p΋��mx�mWz0���0bO _մ�,�����l������?1����Ώq�����u�p(H"�T
i������͛��jt��� 6u�T�m qY�c��V���ݾ}����Y�D��t���Ǭ��gb|	����w��
5��L�[a��8A;���=b�WY�ش�5+4�_`z�F]��|s+�lG('[lɱ��0�JCx�XV^�xAfX^�aAS�p/�����R�~]n������m?.��}��e�}�^:��<��w��D^8����E���Z�T\����u<�Ws�ӓ�������'��b*�*U[*��Q���֭#^{��YA�KX��Y��c6�e��m:T�,����aA�Czq
-�C;Z��g�=��5N� l/
�s�<>j��K�P�PLQ~�,xƣ�� ��mqKO

�e9��P�:�B��W8>���&*`�YU{�2�{��-����>)`ơ��E��JE,ï�7�B��9��C��Mg
�uI�w��·PK��j'�4��+|�I����:=�O/>�r�s� aS��q:�󙯧�z�S�o�^�)�������v�3�Zv.�jr��[��T��$�5��`�S�q'���v��*�CT��򐐌�Q�H�/��������e�;ބw�I��/���²�������;`ó������R�(J��4�<I��-32:���%
Xi�
	��.�IA�r,>g�1c?Fh���C�.C��x�I~�p^Ŵ���S�o�v �4�q؃6>�%l����,��Ӱ�����A�
�&���w����JQTnNOј}���R{����!���sB��l�t�0s��w���k��n+O��`GZ	/�1q�l�/�����*L-��2b)����X+kF�Ɣm�7�h�lx�:a�܊��F��Y�T��Wq����:��[��X���g/�c���xV�y��/�(mC5{K^�NB~���5r�3_g�	�6����)��=�T%�b]������tT	SIs+�K�!�ݾs+
ح�h�Y���k%A&ʣh�T�!�lJ��ELS?qe${�Qvm,fr8R��;�굖/¸U�u���`�p���X���H�(��b���"��]e�x}+�EA����[������.��iv��+��r���$�*)��#pK��c�D1�lyARu3}i�A��Q^J��O��yS~�b�QiFH�tk=��(��(+[[�bA�F9�~@�(\m���},k�6�s�#,�O�<�
�H�ѡP���~w��>�"�uU��i9��8����Q�$��oP�?[\��uX�iN�H�1+X-�empw{�`������o�t=b��SP�c��}�9c��劒kW�q�Ӕ��J�Ve��T�-cVͪ��pY���;����M~$3�6O����52p9��;[��-�������)�3�{:5-M�_7��x������rbYQ��]W�Wa;	k�F�d�G�8���}Fˬ YHTr�F@��RV���'���C��x�Q��&KD�0(]nʭ��ս�&4?y&Y`4� �ʜ�c!��(�p;Fn
d����v����Q;�L�BB�g�)�����RF�d+�LF�3���Rʉ�!����nT��%���A&*78|VP:x^\�k���
���� S�Hd3f�n^�|�þ�AVV�CU�h!�M@~�N@�p�x��#�q*8�
3���r�s��I?8k8Gv���������B(��+��ۏ��;�{]R�NAu�����d��+��q���Y6֤�J/^�[J�X�02$A��ir"
g1���`qy0E���$9���^t�4F�Y�)�qU �E9p�J!7O�:
��6:�{u��	�	���{��b�f5nw�e�N�RX���Dn8h=���WlA����Aq������:��,C�T>RW,s���C�zp�MX�^��o��M��ʃf���~�+*����D���
b�� z���-3^TU�Tb]�G�=r(�^����+��[$pv%n$1�(
��Pţ`pxW�n�&�k(6��J_wpTXT��*[�h���1^!��÷�/��-DQ��9 %��ґcCxo�b��O���\�)?�Pän���Ǖ����ft8F뛊�Cݖkϴ|��.�Y(yI��]zl�v� ��%*��w`�tsl�t?������7�gU%�
��=���NH��1RG��[J8�z�����p����[��m]��`��`!���I���[�	�P�Kv�y�'NB�G�����,��W�����m�R>B�[�ͮF]��q.��@�X;��S��h%�r�+~�Dל�6���D��,���΃��ϲ�Yg�-�"�BW`)��?�	����'ˣ�Xu��r�Z�4���������[�N�/�W/���_�L���q˳�l\�6�?�-��Ҹ��lWf�2*�4\Y���яL5A��Y�X��?QyE���iv�Y�Y�@�������	*%b�J8����.�~�6�V�����	�� ��� ��66�t�;*��G��[�0�u�Ӵ�ݷ^�ǭ�fB���_p�
3�UN8��~�qR�j�IZ���P�"�������#�3����^6����M�}CC��`�u9H���z�Ͱ)��% �W ���*|а�ҴK���T�lh�<u�h���*S�q�l)������L���dx�@�<YU枃��}&lcE8��>�26��WN�/+3
���M���@bB�X�W�?2����ne�峧�R���{�2Bem�yX*e!�wQ��z�%∹
w��N�;ԩ����T��^ZQ0<�5��**��U��<���(`�\����ل����1����'ʓ���	ƌ�0BX�F�:f�'�G8�Q�3ᡑ<�ğ=��^��\�N{�7o�g�L���:�!�P��C%'�1�Gě�J�
i���f�Bɣ�+��Nx�՚�9V�O?�w�P�S�����SV9jIt1��䧧���+C�yxAyj �_N�ת����p���.�0CCV�!�s:��37���,q�{�y^�G,0��n�~�o��냫w�Gv���*VY���#"��)�r���_r��4{�V�s�a���3@�����&� �/^��e~r�1�˥�p�u��z���|�̰3/��������G?�A���{�X-��Q'b���i��G���l�"� /떥����K sҎ����ɶ͑�*y���+�t��rI��N�z�7�ÿ��~q��Y)(�Y�y�LC_y�g���z(��2G\�������Q�I�iF�C򑿸�!��0F�+7>#\���M�Z܊i�AR��hBu�WU�%L%">�r�E��pZB�c=����_���A���
nҮtg|6���)�*�0O�Gn��E��o�A��(L��68x���I�%R_p۸�U`(�Sa����Ib9���]���n:ϺW�;��<�i����ӵ�y
<u�{b�.�;C�b��n�6 s�ژ����ݺ��cbx:D�¢�JcL�y|��N�fp���� i��2?�F�\�+���ccE�[�ǲ(�Ղ�9��u ���pM�i�6Z�,�i�L���R��S��?`PKH�S�m�U��~��������Ty�GW�3���8���Oq��M~�EI�XZ�^
+.��.�(��|���e]�-���{���6��3ɷ��?y�R N��#VJ�Ϳ(�
�
�0� �<��D��l��(��%'FZ
v�d��kq�!��^E�FA�2�0��[*a/	�ҥ�"�B��|��E��r����:��=�:XT�%3�H���X�
��h�6U�����9b1�yoQ�Qz3��ƒt8���&��r�y���uQo�'�	|K�A��=X�Q�k�\KCҥ��cZ�i�~�4�Ls��?� �<�?(�Gw�u�:�W���=�;A�)V�=��;�k�IK������M��]��z:y3^�#L&x�0� ��Z�A��q:yZf-;���d5��&�x�2%[n-y-��M=�L�J����M� �PE^^|/���\ƣw�%���O�pCC5��:Zc�d+K7�ӹs*
i�FTQ���O�
U+V�dű��4w	2�)�ॖ��C��B��>>M��:�=2�g��MG�jz*#!^���(���@���ƻ28X�weX��(��t�o�X&�`h2��S"�@~q��������p'Y���pJC�����2a}w�����n����$|+�@���K���?����mO�7_rmC�淍���O-{�øX�FƆ'��*,�R�d2t��.���Ғ�V�UC�*b������ʥtHr5��-�G+E4��L�~�e�
��!�����[7�/�b��p�C����8��&��L�!(L����4����zU
A�~���1|ʐ�����{�.�g����R,����n#�B�aS����c�q��l����T����9Fu�9^�
��:͹Ml��Ε�ᑤ�]��j�I�qFi*E��n��i��`p�L�5��lw[
a2DKx��9��YR�m-��so���+ݖ�'ls����mn��5z��k,S��c`�s����$T���ا���b�����{}]�<q'�a��ǽ���>k�N�P����Th��e>�u�����,C��#��o���*���?�,%_j�6ρ-�Y�R�a�\�2��N��1��nf�Rj�<��N��ς�}:XG�s-����)�Q��78w�(��2�U��3)/����r?󣰞����2AR��z��*O�Ӽ�[�;��:r��[r���e^:�c�[*5��1����EU$uXݻ��qD��a<+.��I��z��$-	cp�sb�xB��1�O<ˍtQ
�:���p�f�vh�WǬ@�d/��h�:�*��iyh�S/0���#=S=',�D&Ct $�̐2���[��� S�7�>���o?˯`Sq���q�R�@+B����g<�&Nv{��+�����/��8��o^��|~������ſA���6̸��K\����\�ZuoZf��쵒H�~1�~| Φ�AO7v}�g�V�T8� (:	���������4|&���S�!x+J�奸^� ��(X�U�rWy�5ҥ�e~V��QB��%_���Hk����78bq���	>�x�/6�j��,ĺ��IP��jEc�f�*a�!�<��
^V+PXwUv��/��?*eVR���C�<J	�y��e¨0�0�s���s��l�����kV���E�vڴ�Ty�gþ>V�*~j]r�ù���.������>�#y��y�7�?�� ˦���R1Z;��Ω�|;�	�R���T����X�WYV�bi�N�_�׭.���|�a�[c�P䱊�c�EQp�QdQ@���A���E�RT�Ǳj��`�˗/d�{li���Z.�Q���y�C��!Z�7*n��e_}�y6a��F�ң���h/�b�r!�,��*�Օg��<@J�4��G�Z0������ye~!Q�Op����,E�W�SGC�NQ�$����ȋ`'weܸ�k�yu��;����B	�0�m���哕�+��Ո޺*��I��ԜJ4�"��?����Yi�e�F՝�?�e�v�P<�ps�@�:8����J�f����̳>�#�2f���&��Cʎ�n��2�<u5�t"{� Ih�Eh��o�3�u��V�������沼���`^FL�hy���%$�R��L�C��_��x�=A��uB=r{�-���y�sSY
��f��L�hf*�d%Pb��w������ 5�IX�L�����Q�D�/>�4����L��D��7�[07��K�7|�B�7P4���\˳
��4U�v��!˗a�4'Y<��l�W6=��[�h�+cj���⣣ �����	�g_:� �����lؿ
`���1Q�t���|�@_�	8w����֠y�k�4��ɓd
�g�J��w
�V����~���Qi}P �4�����@�o�[gl�kxK��K�	G��q~X���� -Z�Jy��7��@yl�	��X�����8G	��7}N���U�0.���-�6;�p�;s��x�y�G(8�W�wI�
T-Wq��/҃=Y<f�}V��f�r����K�N�ʀ��g������T�� �˗��X�(-�!Q|Tf��*!�ou���;bC������@���5�2B���W�&���fE��
�J��R߹�-i@i1Z�\��9X/��n�����L*J�	���<��u�![o0����\M��T��L��a�t�`��o��Ƶ(N�F4?����)C������a��p����w�P��~�������7(a����\���|��%��ǋ���(���0e���\{(��ܟMK�u#G1��X�RJ��"��t:�ϲ��h��!:)��d��:.��#��zeD��:g#bp�|�
���:I��Gd|�mb���3iI��@�����w� [Bvrj�v�0K�����h&��N����A�P�������Y��+(���s��h�:��p�Ӂ��|\�*��sf��/� �
�����jܒ7f���21\�s��0�v.��Y��%���Խ�C{B��-���������eX�-�S����*Dd�u��[��ܮ�zÊa��;��{�����Y�6OE�ڥ0 i�t+���0Kr$��k�vK�e$���FabȻd*�������W<橽O|x�8:s7a��"�M�7^z�^	Pկ!|��u՗�SO�ew������K��4�0�:�
~NM:4}o!֥��4M�[��B=HX2��g��-jq�@�������0�X�C^
RM|�k�;w��y�梬�3�G	z�C�`�Ȯ��ͱ���z�2y��[E�ZT�ܰ���Tl���0�thG+��7@A���7�I^[Nަ4iS�r�9?��c�#�6ܮC8z�P6\ƥ��0p�稘�����hwzT
b�A�rb��|R�z���I�孲�s��lnzT�u�U��a�����/�s��R�@��<��*=�Q�/����eGN��+������)<Л�`�����9WJE�����
�;�1�K6<Uػ�t��U��tD����\+��r�'�A�T�o���Me�<QΩ�2���Y��+�%��3U&7�7��'l��f��#?L��f4�p���-�
D��0���y��*���g(_�jw�g��r �����O�F��b��0Q��q�	��>=}�h��J�#貌_`��<[�h�۠�E�=����V8-u�$�:	W�ƂFy�!^�QF��km�3DU� 4��6`��5WLn�'�讏|��G�o���򥲛����9i"-������U�#�<g^K�
!�D���ρ�����̙�9��x�
q�M�}ɛzO�l��sI��������XgގvO�&<���g8elջ�te�:�Re��6��4b;� ����/� >������Y�x�l��w����\�Q�Z>��b�K��!����'E�r�;0���h��SPƎ7�2�2�@7d���{B��8�2p�?�`ۡ�Sx#MM��H`H���HT�7�~Oܿ��f�
�ińX��2m)PC�1��3�ebK9)������G�T�>���^^�c��c����L(�0|g��� @��_��'^�g��-��9>�X`@�Q4 MC����W��>��t���rx�MIC��=��UZ~��*�K�u~bi��.�3x�i�:{����.��"�3Oc��8_�Fʽ�^3dv~�)��}l@�bA��<�P) �������D�ȡ[�����g��&b����2N�&�(\
�:)txɊ�cZ�w�����0�W+�b��"N�]�vy���ŧ�Q�d��G_���7�DYy�6�c���������7����/?���.�Z�T<~�c�\R�� U�4��׊v��5�/�/���gEr�4�����U�6�*�Z�đzMj�Q��i����O����9;�I�W�|i�vZ��OZ-�TD��\��Y}�������Q��#Z����g=����Ϲp*��>�yV�!ʖ֧�2�f�G*`�^_�|�f�N(f���S�A�%���ǯ(G�_��+���JG�*R�T����� �3�i����Qs�T�y��ʭ�T��1�+[HP�?���:��<�A����G�����_v=ʗJ}��'�j���R�A��z�P|7��?�WX��#�n���[S�D���`	"��#q{��{5K�͇�Ao, ������v$�Xp���(��(ܦ�:d&v\��U�݈�+��7��
$x���D�����_sXͿ?��r��Y��Q�˪��TЫ��T�[�pZи[��gv�j�NU�=OXT�0�R�OY�|�M�K?�S��L.P�������[��/_��%�s��ᚮ�S� F�����/z���6���(��u,{a���{ϐK��F���`kLЗ��O��d�E-�$
4˅Kʏܳ�qznzjG����`�~c�քۋ��%�􊵁3CB���%|M���tEP�xMt����+ � ��2�2S!y�w��H�,�T�i�B���>�мMP���OT�����R���w���Zi�;�����*@A@�Aɏo�ud����*8��[�+��>�)� �w���ұ�ah��T�W�p�3�D�θ�$uY��zV$R�0�P�(7�ŵ}���3Y=漣sL�&�D&-g2=���yAW)`*/�u5��v������^uq�������UA����L|&n���Q��Ė,㫌fV<2�F����*.�8�"���r�Y�W�\D��j9��n�lx ��{�.�m���|ʈ@�W�������_~�a�CJ�.;�on�aﱇQ8Td҈*@�럖.���ə�7np^��0w���;O���	�>>a�ED� $�j�V��9����՗�!�.��*��˳�/2����l�p��#���5TRTZ�}á�>�'����G�e{�J$/I�tdU�J�J&n���9���^_��z��#�5��(�C**ΐ��j3�Bf��]���V�l�''ol����gˈâQT�w�g�KŚ�Qeݡ]礩T�WR�h����ST$�r�%NE�U�7P���7_/>���(�6r�,Gl�1)Vs�ך�u,J��	��9;�sﺝO���a��i�#��e�i /#��h� ʎ���'�N��(_4&�c�AY�E����
��|�*[>�۸|o��8v��������8�� g��ȟ��x3m�:����~W��zLxV=��n� �Sxo^+ZT��E2igg8l�-�i�)ON�W/�qEFy�0��	W
����r�t7�tK���쪧�W�I����S߇G�,�� �΍G�~��2�ď ��H��2�Aݍ�f�Qyy�ԍ�;�.0r�B9���vډ)�61�k���C��G�Wap��!+V^�9�=��#�`r���*��d�z�������i� i @��W��������� ����,�7�4�͞c��'
7��0�H����
Ҁ�1ݙWD,~<q�Q��M��R(��o��^N�|�ು��Υ��T��y_��I�OC���N�M!:�/|���iR7���⮂M���d)�L�s~���.Y�]��\�J�j^I#�K�[&{W��WE�F�F�9S9����Ν�2T�!�?BDe���ci�<g7� ����v�믿Z|r�<
yO�6ܦ����KH��.i��L	�&�8���� d�1[��2)���q̼�������(_W/�H��_d���A����ʜ:�9t��2F����P�d���D}L��⅋�/�9_6��8�zA��*�h�������(%]��!�78��~��{�8�R�kq�:�<��أ���5�SSQs�x7(u��g�}����c~h9J>�,����x��(�Qc�b�������k��$e�J���	��o~�+�V���.�	��P$ge�.~��j�$,w6
��h+ҠJh���dk��(�Z�g湏�,R)t�I������6b����1[O���>�\mj|�_�V��ɪ�_3w��/���Zl���2|��<a�W��Ôn�jG����A�Md(rK��EA-�7�N Sa7Ԙ<�:�ut�ג���>�9�j^�
���o�D�@�o��Z�=�1)��%2�S����Â+��1�����:����*��W��~��J4�8��SW��r�����s%"p.�Z!�S�P�(W]|bh����zGy&@�_��q���"㎇9yf�㎬���R�	'.G�c�����ݔ2^ZV���#m�2�)%	S�X�7���E�Τ��j��A^n����P�����g�M�*g�Ȃ%p��"	Y'��<�Bc�;A��fi�!���c��z��-�U.�Ċ�3B���T�0]�)H���oc�D�LV@�ޕ&�J16���mc]++�͞-Be�D�~��<�8���E}�, ac�@����n�NKb����w2 �I���dbeM��N!���&���\���
B�'^߽ƣ>��x���l��P���v#�+�j��Sq/[.BZ�7���=�O��e��K�e������`El����ϼu�����*��g��i�g��
�gZ����λ�V�QB��N����ء�9_�]��WiԾb��o���:�-]ک�Km<��!JY�n�
L�+�3Ј��}�D,�(�(\ۛ�!·\�*��F�'��\��!sXgCL]Ъ�7R��>���
�2�����E�<~4��oOl)�	�L�5}�zƠ���|�8Ck���n���"U..`�e̹u��x��x���M��a�(�ĳ����Қ祕FA�u�J�>�42��ɐd����C��Ĥ|�F�q�rp;c"�,�Rx�u���C��u��.0�L%A��!F���d�Su:r�Q��I�-~�	Zy�qLl;�1P��n�Q��4G�ܷ�y��'.��)���������9�>FI�! ���/2��4H�J�sU��΢[�Ж=�|��}w�U�W ������m��
O�*� �w(���O�g��E#�$Dxb�����9��V�Iy.���H�g�ȇ���"h|���os25<�iGtl^*����W�ο��Oᝃ6��N���;�O{�n����C�>�8R
��}x0b��zefy�>�m8�z�Q�-`.�Lӝ���-�}��e
7�b����R4����"�e�@��I���[����r�s�ʤ���Q(���b�i�>iɢ�;�XE�	#b��z�+e%����ۆ��G���(G鉸c�	P�r5�n��aʚ�P0�]��a�k����R`�����r/y�e�g�j��� #�I�\�f
���2�DÔa
+8���wb��#;�KQDd�W��F��{W�o�1�V���k��$T7H����[���|�QJ�䐍�i���C'�J�1C��
�(���8p�|��%�^��������P� ����q
І/l5�}��W�T���`a�,OW	ǿ1�O�`��c�K?W#!t�`^�w�JyU!���'��Ub�����x��V̲j	B����b�����^V8�P��-����e/�13�(�yc����46N��KEYs��\��<�]�=��O���}��.�6�Z'<^&�m2�ᤍW�9/�!��۞����PM
�fr-)6�ul��u?vö�(�Z�WH�>w�9a� k���6
��&��ZG]�X�X������C�M�@�@KG[l�#��*�*p�ӂ����m�Ӻ��V)�ާ���a-��/o^bE{�~Y��֩,�DE$�q[�@[�1���L��1Ƒ�g�b�Gx�'�j�´��X�%8p~q�Ȩ8:��}��m�[��|e����70�<}�b�~��K���o]%���w�ֿ������]�/a-W�3�����CQ��ǔ�^8�K�a^��Z��\Ս��e�e�F��3�M�V�Ë����0T�q+�ħ[]� �&y��^<uˌ5��Z a����\��ny�v��=M�򽂋E��p������Y��2�5���L�5|?��sN�H�)�ʿ}����W���!R�c�!��
b!��Z����?n�Ͷ;�#v��
�4��;p��T�ðҔ������SJN�c���ie���z�Π:�2������M�5́�YI1)ӁLx�h����h���IhE��!�e�1c��0+ ��%8���.�+;�{����t���3Ƙ��I�6=`&�mp�uՎ��l &��XִX{��p��b�G�81"��I�*�+y�E��"*s,�_���\���U3&Q7��I��5�˺B�JC�$\��@��	�	gì 0�)�V[cr<��I�Ao#N�
��M	cdNz�ſX�2�3�� n�O�����2K�
R]��+�q�ޥN^��ti7�2x���⟆o�c�� ��n��U4J��D�w~:H�O}4�O��%�3���a����|�Ƿl�K:�[�n���  ���M/�􍥞�;��s��.¨A�*ÓBnWڌj�w�x�GGɡ�6c��AWoeO'�6Q&���9;6����^rȲ;Z�3�1$ �,�0�bHR6y&坻wP��0h��dm͢�R��jf�  @ IDAT�Щ�p<g���[��X��>}�����k�ߤ�R2��w뤻�?�o��w߆���3�%L�>f�
�SR7�SG��I&�3<i�U���y�nL:�ܹ�G��{���Hԥ2Q�<���[zH�^%mE���q�1��Py㷗����G\f��/�&���O��[?݂G��h��T�
�W�I�x��M���s�
U��{��A��8dX��1:RW;>��C��8����b���t`ﱠ�!'-�i��~��<	?)�ۭ�~���ӫYͩ,m�}����=-`��U�TX��{������~��3RrJ�V��w�Cҁ|� Ϯ|#��+-c�{GGh/R����-��,�rS�����a�X}���Kˡ��d��9�2<xG,�K�7�n�=�!�Eyd�(̐\2���+���6N����8�h�����\�RG�}t�������h�'�~�]2uǠ�/��B`-L[lu�7yQ
A%o:S*O:��rū�ĻJ�|��P�4�lb��{ے��W�����n�O�?-����0B��I���j/��S��@:|'/��|U�)��DIrQ(�|S��2Pu0��r7��4񝺃�&Ȳ���9T�PKG�Σ����QÓu�*x�t)�Y�.4M԰�%�
��:�L���P��	x�k���b���$)i(	�Ĳr�����&���L#�(3���	k�'��(����I�-+		o�e�JMR"lh4k�KN�{�%�l����s�)z��8�@�skÙL�m�r�l��6}��"�����	�*,p4 Q����.y�U�b�Y��\��L-w��5��3�ɓ��{�T��wX���AA-����s �s	����s��(�P���
]��KPhqQ!��yǢ(�Fm�3Su��O���4��#��WaTx������Eٷ���]�CU�%�R�TZ���1,��hx�^1R÷i�z�� �Bּ&�N���~�x�Ʋ����#��+x�O{���aϗ(O��8o'u��A�E�R| ;6�a��\�
�2���h)1�nt$�O��J��]�ٟ���3����e'�?c%d6L�p2���e7�5�l�_��_?���{o!|��hh����=�b��E��r�'��,H�J��'ԫ���z��]L�t�����t�	��BY��՝!5ʐ~*�������KWþ!�x���1O����c���]R܌EO�q/G@��/_�!7+?�ߡ_(�"~���/8O�6���pa��ټU��i �DFT��]��%���ߓ��Q��E�J��ü�(iҐH	���?��F���S�Wx���l
����%�;\�����?.n~�y5�v4����&�*O�������;I���'D+�c1�|W'ú`>О���z�P�ygʈ�[c��'K�C�Ұ�Ӽ�S�%���p�C�sAs
�a)Y6�"��X2�T �r.�Rp5^}����rk0`u���y\��,���Y���:@a�`��$�5y�n9�1ܖ�bE�˲#�a���<�[�>t�	<�/i�]%_�ۺͼ�Ȥ��bA�x�h+����#�UVE����e��)E�#*_Zj��j�F'���V�䌲bG��֑뗖c�e`���W�ј�C��4���I�Wh�NT]��vu&�;)��e��Ƿ��6�X�r
E��rn����=���+�Ҙ簎��9�Pn����mcG�1��J�$T53�,S>�g��c��@�O� ,��|2AB�*a�G�eƚ"*/���Z�L�&K��Li�'
]���M#��	�o����� B	O�*e��f��R����f��7�/wa`z��J�*���A`��^L�xo7��Әꍯ	���w��p/��]u-�e�~��,4Ĭg �o C���<WҜw`̐��_3�:<�Y��O% nK� ��
��(��M%���Y��(��)�"m�XN���vyZ�D{��S�ʢj�Ax��QA�UieI�Q�*-:�Ð�L�ܶA�»���6�r���t�5�O4ȷ��j�m� ,T�PK���Oӝ]�Q"�G�,-(���Lx��s6)��U�s���' ��_7�6��@aCf�܏Pr�@�d8짟��NB�y�U�Y�_:KQ��Q���sU|��1	~S$�G�J>�`Ԫ<�x*'���v��iAq�=ғ31�� ����v�Q\�:%�K�������n�t$|�a�g���{��V:�>n�x4�m^�x$��2Y�U|�B�V�W�YA����<�;GVA�|�������)R�o9�B\)h�Ug��g?�A�<6�Oy"�vY�P��J����ɻO�b#gx�����'_��>h[;��Cʱ\�ti����
uq[F����K�N]�쎢���!PL7�uu:,I�1'm,=��[E�d�����m���:�.*����W�m�1!)zW�L��g���|�4+�BF~��:�
zS��;~�p%�Y���gd�Z������ ��̐���U�L�rD���\Lf�ݰ�������O'���@��=Gd�:.�\&�k
C����U� �Co�G����Ȟ��P*��z#�2�{)�P"N���>�!f'ARGS��O~{�)-I�Գޝ�1�0�x�r<���,B��@��SI���Lv�n�u�gj� �θ�G�}+�ǲ����&=�LFe�;p�c	5Lᣩ;K�=6�
��ƿ��7�u��K w9 �&J���_e�~����2A�ZӦ�
��X�l2,�\6���se���F&8�d�ϱ�L��>N��3�T�tT�R8���iC)��2��s	��V���$@p>s_
����:����`M�[�g\	��at�k	3s4�LN~r������6�z�9�/�ج4
<8�`70��Wo�cCg�U���J��1\�s:�3� ��b�R��JEo�8������m�^Q��'m��U���Z?�os��6c��<����&���c��a��=�L�����-C/�Z`xV���Q
��k��Qw�n�چ�+��<:�ʂ�bf8�p=`�'���F$6�
\�lؽ*L5�6�*P����Qx�e�,/B������k��!sĩ�u.�8�e:Xa�&�'�zk��Y��+�!��L�'�R8LJJ���[��|�	qJg�Zm�,��v�p�-�R
�i*eݸMG�E&v��D�BHx��W�z��>�E�gV`_�<�:~������G�}��*��K��*���D�mZ|�=�ي��n���H�<���~�1i�~��EN/X۸@�e�%�!C�nw�^gY��rF����E��v-�(��Y�K���%�6r���úC�͊���R�a��$E&*)�i������*��*+Ĉq�F�u��.���w�7@��H������f�팞x��v��<���/8T����6r)Q��[�k�X� D��we	��>@Y%l|t׋o-Gn�lv�����I���O}���Q��'��Gk�&�������X�/����n���Y� u�:��PO�i]�d^+OeTV�4��IN�4m�wp����V-���!u�@A��}i_h﷘z�s�
�L�8\<g��:���U�m����F	���C�9���a1��h�Tt2q7m�Ϩ1jR����H�(h�u5��3��7�b����3�fx	�l �G��o	�&�7n���u�FHJ<j��:!�����W�f(ԥk���3�1���;T��j���}��[����Q��*fq!J#� ��
����.
6p�Ln��l����.�7��[@�b����o������#����L@R��
n���)�3�O~��Sy����,z���Wb�!��ma"2��ʂ=�!B�ur'q�{;�WE��k�UL��p���(]<���J�2T�0��fT�lЎ]�G�:���5Y�$X��a�3����(�G��@��*Ji���R�����
�+�;�p<ġ 2=^%T��*�U���O�[p���͂��@P�'����',$\��=��O�?�v�
��P����Y|�7��g�'3��|�������������W��O�a]�:zӴ�&O�D5��gP�i�C^j�l>�<��U���4��õ�U�Ze��`�U�V*
Fx����^�ԯ��átX���� 9�h�v}��_��rSˤ��x#O��|��mC���w6���/$�2�ܳ��&����.���#��pS���r��!8���V�H#�U���Ip���ߍ�T��я��_��Y�L���@�$���&�B�H�;7}���kNJ��_�"߭�>�_��]���[��q�[ڦ۲�l���w䦝L3�K���(�y\�\\a��<m/Z�9�\n<v�79c�E>��u�цmV%)wk�e���H�Oq����j���7�Iws����@\�=�]�r�Έ���'��\\O���n�r��G��*`8�խt�Pڴ�g�����L�*b(���δ��*�)K��=�cV�ػ�r��	�Z&��	�0�DS��D���!�\2E!$\�-�x� ��081!�aQ�hq�+�hΌ����fV�E	�C���+���{j'(e%t����ZH4;���z���´��BN�4�\��	�=J�JoE��3�0��D�˫~�+�c� ��"�3�w�π���k�&�S:~�Gv������r�T�Ls���T�����nEr�����0�!�q�<�B����<��.��FF
ˤ�!�`�Q#(��[��;<g�w��^{�*�}��!<��Cs՞Cx������n����B����ť��j�8Rj���ue�!����W�#��O]���&<8U|��Jw}w��a]�+�ĵ�"�q6��u٫�6M�φײ�ݗq5Ά��0�R�]4Ls
���E�^�Kz_����Z4)vJ��Kv���[uV���*ZO�i^�&|�a|���Ti�t�=�ә���j��Y��k�l���;W�
�&G\1:���6�lZ�א��F���7l�ˑ���ۢ�2���̡!����KnQ��f}��˚uH�D�8�wSe�r�_�_I���ΆK)@\���[�1�7^n|��.���k��8�cп�5��-�?aY͛.���Y>�k�w�9e6��G[.r��`�%�ct����,N_�	<y�*a�*���j�6?�'�f.��+�o��/>����sŘo��W�7�ÑZ[mx�	�ʉ����~K/�uF�f�j�x׭���]�d�J��#E}�b�#W�)��wa]�*�Z�,s�f@�BC����(��[�t�[w�y�+
����х�{�2�®,ܢ����,;��&1���J#���LBY��TB+�76d�H�[���b��C#{!{9T�� �����u(v)<	��L%���8�W�
@Z����eR��/( ��cp��#Ih�k�i`�x��lD����AS�����,/y�,I*sB~�l���PM��4��4�П󧘖�
�*��f1΃���3����R94��p�!�)8a����%K�t+^xba%-�	|�ߝ��҃�Ca�P�\���9�)��@�Q���T�����wf��a�V��/r�y�xh��������5�V��}�Mv#�+��wW��W�����C��udY���=EZ�k˙��-s� ��mr��)��2 �|E��2X<�͒Wg�����xV�k��񶂡��+b��a?E��;����:\ו9L�~տ���9ny�"eݫ���=���_|���K|6H�_��C>�{�w��ո}z��w�c��p�~�]��x^��J�TG��\)��w���޴�*�K�J�V);��?ʈ
�OWM%M~�P�+�W�/�a��.��Sc��<^��͓(j��/IZ��j S?�=x=BP�h��JM�"�m�i���|�����l��ů��_�X����F�5�X��_�/������� Nen�D���)	�����Ӂ+n3�M����R�H�n%���%+G��nx(5�?�z�Ŧ��W|����?|�ŗ��q��hw�b���W�UFh��
n�	n;�>�:m��j�
�;t�z�_�I2�C9+�W��������GÓ�(�uZ��p�$֘���._���J�V�Q��X�0����p�˱��㛋/��OL��ɱZ��X�R���0n����T7��,A��Kų�ݤA3s_��!�*FZ�j��ēB ø�w���������c��۬κu���	��<2�8:"Q�6�� #���n�0H?tP�^��u4q�ݢi�қbz,!u�Ca ��.OybCZ[�X�B� }�c�G��)��!x�_*��.>��X	�O�����pg���\�/晗a�g{�'c�8ˡ�A\�ժ*������*��}F�xt�R�7+�4����`|�GI|��O�l����uޕ}4㘿����=�`���3TÄk�u��lP�2��+�Qi�a�e�rQ��sc}1��&�NM����<�Lg��x;�O/��dX�gh�]��sp���w����xc��]Kֻp��*m�Э�o:u�xۭ�U\�o��0�򼮂�5��E��i<͋N�S��ǆ����2��p����{��i��a�/wd5"�a�S�w
����M�����(_����V��[y�ߵb�9��0�F��(��i7P�\���eD
���g/��h|�J���dm-��)H��#����J�#n�}ȇ�]�!��"��ora]%l&O*
��M�ėH����j���W���x�[�#2b�!-��t�J�#%�S��I>�a�.�"�3%G��n�uY 8}֛ς�{Гxt���_�'h1z��.�f��ѥ�o����W_}����u�MD9��e�Օ���x�M��WNQ��W:��)���f�������΢�d�`��,`��7�+�̡}�%=.�o�Q:�(_�@�ra�2m)��7n˼z�@бWq��)k��ʇ&��c��~�Z�c_�aqC-*_�b��<#�d�X��[+N������21��t����Y)�ƁVX��-�ff��!���4�q�T���WXVϹl���=�P�=�]<~�yrh�J���h������4㻈��2�8��Ź3���7鏖�Sˇs��3W��%��X닏�i�|� 	����i��$KV��<+�ri�:���{~͓V� ���̐�қF�|�G��2�V!}�0�^�G��S�����:��,iY�iŭ2�0b�(���L�d.�+Z���ӳ��x���S�/�l^���tNT�����(!�?����{W��VĬ+Z�7�ܭ�����7�#u!	�_���F�X��	!6�iX�|�n��g���ϧx}FQ����w���L������W�p���<(��N��2q�^��g�.ejT���H�p�tU��qTxqV��츌�����ns8a��g���_�gV�����f�CgJ���X�u�t��9��w/��bƨ�ah�ߠ�)*K֎&��CuU��в�����)k������p�E�юA���rGZBny�V��{yiTH�4�I�$���$߯�u��O�	����S�\�pw����G��w���>�5�-����Pǯ���i�A�u�wx�/<�"�t�x/&�Fʼ�6JX�Y0����$�o#N\ƾ,��"�x�Q;{9g�~�����,_���z<�1S�ا�x�'�'M�[L쬪/jAꎓ�����b��� ��M��w�-�Ϳt�֤���l���u���E�zʒ�,G�R��|�t�~��u�+��{�Q�tlJ���I����ɀ6d�
��HVkOܒnK[N��#DBؘ��po
�B �s_��rk5p.��E At�I*͝Xc�!�E��	�ٔ �ڼ��os������?��%�l���⇟n/����#*r�C�u>���=���7� ��9E�]}5YP9�{%;r$=��L�ɝ����[#�L�{m��a�F�h����o���'N�{�4cBf�@ �� <D�e[�#Sjɟ(}}�2��8��V�Fn������VVu��pBc.<k��4fZЭ�c��{���jO`�n�� �O��a��ߧÒ-�U��6),b_�����nJz���t

���s���cr�}�-���қ��_�S9�x������D.��5h��G�H���4�l���z)�[�H��Q���^p�M�5��%Avc��B|��(��6=�[tR��c�}�jۛm\�͡�3�����`{�0�)g����}�߸8'��>q��8�6�ٸ��x��{^.�M���{��9�Gq��(���~��+�1^��WUe��a��l��g��"l
���72z��a��g��#~�'9�L�.�M\Gr�5bl��f�hTt�j��s\�M�,���gƸ�a���?r�٦m_��Ƶ:>ᘷ�,�ŷ~눱�
�ʦ�X��*z�;3�^�����U�U_v
���X����k������{�-��/�鏍G���Xa�I�7?��a���.S�ë��x��N3�q��q�#��{�=���m��!��p���"��TE�����}`Ia���������|8�������;�u�ZZV�c?�({�.t���R��\���.�����]�ԾG�k���*[P�~�~���i�4ý9U�fg�mXlKs�Ic�M��;�؅C��y���;oH�(�{��5�3�{����۽�\��0���¸Bgf��mw��=���ב��/��f�N�t>±���M������hE�ǡF�*��'8�8����6r�/Fp��[L�
ħ3��m}��S��@+�My��5�{w��L/������ș�;7�Ə��;Ɂ�#��GM^�B��_��v��E�-�׊�Ѯ�B\ߦs�3iw�u����7v=���s�4�=���P�'��>�?~�`���O���J��=KB/f���X�y��pNG�ue4?W`t��Ic��3>���q���w�-U���`�|���u`����::�x���8.����R(�O}��McȰw6|�bC�|��Vg��Q�q��� ��F�e�v�bQ0a҉�(�*� 6��;��=����b��T=��z���N�-'k��)F=���#�EZ�?i������������0x��#�S�I?��V�O��2KI{�4ˤg����׸�ane��ߧM��fΧ��`sbЋe����v���x�}��51o�<����Η�pg���ٚ��h(X�C8�8�Ӧ�@V�o����o����ƣ&q�g��?O8��0	�h�R�Hc�����`�1ÁL9V��>֛7��eI���-Z���b��h�0�<n�I�7��Ѽ�9Y���N�)������:���6q~]�����dH��җ�7jZ���4�X-\GW�$Q�6%}
?��ϴy���ط_}���-�h�&�1g��/I8)��������r`����~|��t˫ïv����v��m���~�KI�7���)��t���'�-͒�e������T�����]�G��y[�����k�u��ͧ;���7y.k#p:�}���/���9�_\���ril�`e�v��ϭ��EV���3�(�V�1�;)խ�3%m���Ç���J
-�;�̀@^��(�7�P���?�#�7�??���`���������<��0�Rz=�n:��#�>���C� �pkAB��2H�,����6D�Q9qb1$���TX�cb����2ן��)��>i��;���V�A�8�U+L��t�hl��ѻ3��Ĺͦ��F�ɬ�&����z�6�cd�S��c�
�.�?�A��;����<����±�n�g�,��(��Aĳ�9y���.��;w\�{7�Y\�#�K#6�+����Ғ?����c��k��f�CO�;�� �Y�C�8��4y���M�[��|�5}h��٧���"^q��j\���N
�3��z�����/���Q,{^�G\{�{�Sޒ�sƍS�5M��\����8�`���[7�y=�1����ǲ�L�#�1��a1y�!p��:�P�(m�kZz� �#e�L�~��/f+��v�+3�:o������K+�q�$wv�g
�n�E��y�r�|)B�̪��Q��g�R�*;��o�4p �GC�IG��¢����M�鹶��?�Jh�����	�[���DI���g������h�tC��"~��m"b��������W`���S6�Ã�K$6���~~�o���}ȣ����>|�z��������`�3<�lO�:T���N��c��D?g�-_��w��?vm���ڇ�v�.)����u�� ���5�9��5�7���s�w�݄]uUa�'�㘵�WwISbL�.���57~���g<�+&��O�elF�t�RÛu�;�s�36F�+��"��5x��u�xS����y6�̀�.k*����2�3фBY5�K�W�^��\���̎ ^8�
-�z�
7oE�`��[�|�Bz�>qp�Ba��#�@��ׯ����6�hc>��:
r�{���狚�u�3{�[�<G6��[y�{����2���mzw��R�DuT�\�+�a�Ux՗9�o�ȼ�f@��Z!s29_ķ!��{l�aN( r� �t�3ԥ1���I$���ۈ.`w{����?g�F������PN�e�����tzhg턪���Դ�}D��kx�qai�״7�l�/�P�s8��i{���ڗ�8a�ױ�;����:����L�4×��#���,:��ZL;UF~tjn�[z�<e�|.�	�mꮃ�9)H����Ǡ^>�A�΃i^�!�Ph�Nwa� {�Ӈ֜~_f��H�����F���G^��q�W5����ڄmݾc?6��d(<��l���Py�g�u�������fOiU��C�2Kd�3 ��,<�������9��36���0���*�mXy߁��W�����&ޛuaN>�|[;�_x�AMfǎ����cO0�s=g�F9�CZ�h�ݛ������i��ɟU>�.�6pr�4sS�u��O�H��(s9?cSs��ϋ��%����S��s��M/� ֟7�������u�X遼�3�>[.�P_��~������tW|1]��6��&:K\��K�����_��T���o�Ue����m�o�n�����)�<c�U�;g��[�oǹi��S�gۯ�;6x����؜2+����5���u��SY�-�r:*��k���|1���}���ҁu�p��><����R�kgϾ��x���\o�����]~�AEFe�A*�3s����a��&�
\$��jU�BV:ū�J^'K�Ё�����6�o�������v�T�V�Q��<�Πx�&{�p���s_�:����8?��;����=��|������������i��7~G�Y���T�q�TN
��-�\�&�IX��Ұ���&�֨��c��8�?%-J�.���lb~ %����BR*C��@��R�љz�u{�������O��/^��љ'�����VeZ�nNą�;並j7u�q��[�y�*��w�nG�Z:`΂�r�}L�"�[P8����t"�q��n��.�>���K��]Iz�2w?6ő�|S'T#�H��ZI�AS�=/�pΝ>i�.D#�0I�̍�ّY�A��Ya��̓��Q	�Yf?�ɓn��EO������?gӽ�<|/�2�e���Q<u�Na��M��M���L�.��w�}��]�.�a�ZK��r��'$��#7����<��N� �:`����R=�F�-,�X'��Rof;c�6ވ��	��[�@C������2��ԛog�F��Yg�җ�F-Ҷ��:_)��4����!��wtM[��zɹt���mUD\�E��r�-c@�k�h��9��Ie�0�k�<��4�9��N��~Zb�9E�%�r�B���W��+��U��U�9������$��~v�5�]z��~Vu���_�Q�hۋ�"�O��fu���Ȋv���>�������������~��Oa霹?��W�9׊{����~9�Y�7o�RN���Kj�Y���`�L��ø��v���or����}N���X�7�4~�}0,\hsd��͏�gM��s|g��ܜO���m�ۼ�u}-�	8��C1�欝��=�}�s9�L��D4��5�����4�N�I�E�*6��� ��*��:�a1��uz��������.�4z�]K�u�0Oӆ����O"_RxÌ�G>��Q\BR�P��}�؉x�v�&^�5_e�ձr3��O��R��4�b�#������2��ߨ�Z��ʍ�r�H0�9�e3�����\��O9/�v= s��s��sx����v�V�'��VM��u�ҳzNI�6\��?�6��Kg0m@6>�jB�[H���s�����km����{ =6,�Q:|`�����,:0���Z�a�V�S��p�6�f�l/�x�y�޽� 8������s� �mҒ���4�5+i�[��=�͜6l���Am2�?r{o��'�y�b?�-La�t38�����+=�_�ᘶ�(���2^7}�m��u�n@�g{&[�j=k�����N��S�8\ا|����ۿ�h���^?�%@;�~�I��^�}
���L���9h)��˟���E{��n�M�]����㬻��:5y��\�S�Y�y��Ù
_X�yd�`�&��
��%���WX
o�	�XD�����]��U/vB��ů��n���O�9�۶��\p�"m��!���OT8�˓�x.��O�@��_=��T�)�W���pb�S���7��x���鐸%S�m���C�f��e�m?R��[���J;�B˘��Q�m��&C��{g����7<o������ ���.�<���e�Zݼu�7�Y�~�'W�D�����3m�|���L|�G�di	7�>J�$K@h��U��+%�)CFH��y�����'] @��˘�sx����{�9�U}��<e�7����}���È.�.�)�W/�����U<�=�m�թh�$�D9������>��4|�rϑ�5�vX�r#KP��4�LG��ǝ�=�A�" ����ƣ�i�m��8�x�J{�g��܌a�{ϣD{p�;�`�1�醿�X��o��y�B����u�T�5!�R:�W�B�@���CS;���كzt�q��g);�]��&,Մ'�j�\M��iF�ςug�L��a���@9}#�P�!�<��� :
;�2��GƷF|䌙0,9��~b�r1�y#T.gL;��c���u�`�>�����'�ЯP��gf��o���M?K��_�~}|�*���l�n�j#�����_�6f{��S���r��h�>��t	Rxg��l�,�轈��l�Uv���L�q�'�>i�W:��O��	;�<O����r�ܰooSF؁��e<������,'�Mͻ��	�"���Ÿ �Q �8KCc�ɏvc��N�h���G�"�����9|,�	3t&����u��j5�
�M}/;.��5g��چ���/�n��i�_���Kֶ���k��Ug����/�#��_���v8��ۙoB�9��[n�P�����Rț�	W�.�\�su������������C��cB�6\s�>p����3�Qh",�ѐ)r������s�'�^���d���~�[����C��?���}uP� 'T\��S��>دה�g��1�Ȣ]Z_�a'[ګv��>O�\g����8t�|$�S�8���љ�'g����w�3Y�w��?���`f��P����`�^X�B��4��/��:e񟿹qx�X�����G�Y2���_�V{�Չ�чm��O|��ɡW,��q㗼\p�ͷ�}S�����wb�aNu���LO�
N��luVt����n�L�Ҁ|��p槈T���SΔ�9ˤ�������h�Ml�7�a*�ǎV���lp��5(��Zn��Y�!��w�f�WM���x�(p��|ƕkOWx��g�(�WWU�Ӆy�C�*0����{wٮ��z�wྜ-��CR	��E�t+�-y��UPgѭ<�p^���� �t,��ˠjK~.�6�%7��������4�=k�>�-�Q�y�W�ez5e�78�D{I�O2A@�y�Gyq~u����g�i�P٥1�8�\C]*}��}�ƫΗ��wf�](씰S��"�T@j�uņοN�e�6�Ƞ򑎋D�b�C��w��k+�>}��eg[��8L$���m�I����1��EEL�L8�Ϥ�9�Å�сy�<K�z�PP_{;*��&q�r�ևV�jC��1�'L����a��G�������gR
7��|�
�|�K�9�r���q����[�Y\:'sC���\j^u%Qm�C�z�����pFlWʑ����4˷�Û�U��b���ݾ]'�A����kՄ]�A_�>t�|�ț�̞8&�~���:_�u�X��M���:m�"���͋|X�ɈJ6s�iW�la�2�.|��7J�:�#��r���E�ʥ��+4z�\}�Kq7o��@�(�z�<'����'�B���&p��М�Q��=�6�؆��ɺ/���'3�:^LR���N�:��Z���w����-�;��ԇ��9n|�K��k��9c�����?�O�#�5l�[~ģMJ�-�n�x��%,�l����b{�����ݨ�yM+.?>��F��|����&���~�0��84�ƪë��t�|�����?��	�;�nY+p��3�ʪ�������x=�N��4`��4�\�������M��R�>��Jc�r�l�f��C̢R���$`����3\+_�;��'Oy���ElWy��~��\���j4*=�Lߥ���� �K|2�{�b�$ڦ�߹�.%w���)��yQx��À7����.;�_�o��f1D;)�E�tfK2�(EN�f~�"��8���k���f��/�ʺ3�%���ςF*�4;�(I��̤#���ׄ�
aJ؈Wy��ν���̂���~pe���4�"�ڋr��2ϰ�$� L�~�سE�Z�<��Ɯ�r�7���O`�v��(9�P�������4t�֓|��b>���tL���u.]Ϲ��2�Y���L�p��I���.VVN�y�TwnX�	ѡ����%��[�#�uG���|k�������f�V�{yMk��)3j��i��䍓��2��|4����O|�,��-)�����rª��@~�~����rC�7���z�K嶼�8��\��Y�����,G���N�f�/���^ԣ������_ʷC�0���M��fvV�:fu��Y|�h�G�����X����eĲ�����a��kr��r8�޴*�os�,�Q1X�����j�:_���A�*��
7���vB��[kي�~A�qPAw���S�u�l7���.3)��Vkʠ�?ꁿi�d�4J�dP>%�v�}������#R9v�{��><o�Q>�"Ox��Е������1U>�|�����s5g�8�S~w����?Y&ɻ����1�L� �u��ٟ�<�zϘk�ۯ�]�M�)'���{�N;�x֦�����o��妝�  �D~�'�F�fO�j_���u7�f[�3�~��\g�%�8_�c�GhX�[�ŉ�	� t2�I���I��x������3n��O��-��/Q��@��K�?�p��f[c��]&t�n0It	���;�iK�'�������m-1�[�)cs������U�TO�gʾB�80<@J��\ t�������[�0y�/G���-�^~?����޺� ���@��|Ya�����A!��>���PW�+��{��v鸠��G�O۩���!3/����B��O
U��!JS�U"�B%QA~����E�N��(���8�W|�&}΂� �<���`�ߥNT�ڇ�a���/�|��f�MH�Lt�ަ�˛:ױ1(F�(�tf������3>Sq�E�:`s��@�SXz}A���'�CO=xH.Bs��Ӡ.c�����,�˲��Bh-<��Æ޿��G, `����eP��7��������t�>L3~�^�|�����u�6�����@{N=��u���{�g��γ�<)�A�<�Ԥ��(C��a��.���X�=����2�1��o�������Ƈ���&�t��J�  @ IDAT�q��I.�߁;��_|�HR�Tf_ rV5y���3�������R�Tn�SC�tqy�	//�L��c6gu�'�X��f�B��,��?�u�]�˿i=q�K~2[�2 玾��v�;3Ut�W���z7�3�F�^�t�>��23����;��Q%��ǈv�O å2������^͑�H!���g�uq6�l�.��MeG%���j���{%�I�2e�8a�CN���`��8�L7��O��b;Is^�[����ї�^��Kmlϐ�x�JmK?@�u~�\���8�)�ZZa�v�E.���<v�"�	K�Wܲ��}��Ն4�Vt��a������댧`�\��Q�F�d���0;
�;�Vm�2bo�����v��-�v{�ef�KpS.~����e��s��]emZ&x��� �M�S'�m�C�p#�|�pI�6#v0��_��r/�A�QP���qZ�i�8�g�`ț�2��R<g	p���㧬AC�k<B���GO����,��s��2���`��
��&�v�p~5:��.������e*6S�2E!=bw>��y>��]�:�A����~�����a��j�Eo9g\ԛw}>2�]�2iX��2�p��h���G��c �ȏ����^�w��h0�(άwXuh�X����4���1�J��:�gԿ�Tt���_�Y�x�;�Kց�=Xw�.�Q�����&}%�dZ:���C�8�����`gDSd���蠥�� ��L�a�����-Xa���e�A솼P���Pf;(#|;���RI'���9S� ���ɟ��\���9�"���c֙������&���^I/�heH�<z+��3�ߟs�K��_:GJN�������sf�A���x��4x�e�ec}8 �>lˮ�rO���$X�:2��q˛n������4OmӅ����z�j~��������!\leo9f.��ϖϝ>�,: ҞS[��|\���d�e"[�7#��~EĮ����u�A��E��p��n5���R��f�է��W;�t�ȳ��֞��z,�0�6�����R�Z�6��ЯdLs�2����^�R`���ǎ�8�����iɋe.b�4�V*��z6�KA�gg���B�QSw���'<m��
�:<yى	�+�[�{��mꀱ�6�^�4OK��`1�5�W����-�֍PqZL\�� �l��~f!��4��1��BP�ڄv���)��)�WK]��G�����eO6#ǟ+��R��QY�yv���e�O����˔�Y��r��� ���NzA��΂2��9�^f*X"�R���~��
��^�[N�e�4�� 5�Kx���`�i�6bz���»��3�[wY��oTF�Շ�:"��;��@�oa��d�C��y�WށXC�2_��xޭiQN�v���G�>2� D=��v|P���
^g~����'Fh��o
��Q:#wY�(,6&�$�D)P�*���m�n�{�����>�$��z�Z?bK����A}i
]?b�z7i��y/�zD.��=��=[t�=b�Θo�ܹ��p�:�n"v �����補SHV��g�҃I�XƎo:�>��ŧQ�u�|�ӑ,�vp�isө�(�;(95���o�Kao<\g�5�=���4M���~1M����2xSb�GO���S�KsAF�����ʌ�6(�8[3h�e�� ��	����&���]�[�?4��-'��Ws��E���zh��69rW��߾��><�nً�堿�����2^�i;:X:O�;�UG|p�&�=����8�5�͋�q�vh����	����NI�dM��[��k�זI�F���#N�}P���]��K+7ݰ�A�����,�D�E�.�ύ8|Z�>e�/������>�CJy��#�rH��G=��[D�E�e_�n��,��N��+�k֖�������5�Ŷ���͸��MW-��ۓ2��={ݰE&!��sG�cz��[r{��w�9|$�E�:�%�R&�;��(���5o�����־m~�q�%H��O��v����.�{� ��P��O��_���5����96����t��������'��O�$L�̾��^N4sr���/�JM�;�Q���*}�|��:0m.��K�����x���'����h1�CIj�8��L^0��M�e��v��	8��r�f}+�g�8:�h�]�7��vj\3�t�k�[���2�w�O\?������3T��wbH�<��%h+�+�)����]���X����9��y7�^'�3o��	��(���{,���Qlk��c	Үve�A�P4�T$|x�w���������7�t��g�u� ��W�T�z%����2i����y�{�l�~)l��K �tꅺ��>��֣�Xl7��%o:Z����月[���1�9�#�����X>��[9��;��}�rF����,�a���+y|0����oA����˼}~t���7����k�b��,g���N'���Z�1�j�画n��ȍ�ܫC�r�}Ӊ׋�`���Do�<J����"�n��y&��z�]�s݉���E+���e&��-�q����G,\G~����2�_�Ţ�Z�mXn�ޱ���i�(Ny�������씟Y��8��G'b
_��r�n�% =K�u53��0��Cs�gNz�e�2�����9��w�3���S�i�\� nCO�n��׳�[�-�]MQ+�n<в�E��V+w�����Sf�_�S��7ȿ�/��L��M�BS��:/׌NtJ��ei�<4ex��}��orP7�Ora���%��Ǔ'O�+�]������(�\�8�K)�� m]�E�?�t�-a���<M���L����.�J �b+��5vt� q]%���[��z���s����3�ЮϘ�q���;����8y�O����1M=T�/!�	Ǽ5�e<`n�ϣVyl�85�c�eH�3bC���^����92��b�R�	|���Y?g����	�<qr�NNI�xiq�~2Ê}�+�B�GB�pmE�+��l�1ABE�6Xa����0FIJn4X:'w�����Q &wP���iGSɥ�w��
v��u:�q��1���L�e�O�O��˗��JW�s��'o4�Lǡ*��)X੡^�Qj^����?��#�y�iqLSA%��.���� +R	\�s�G̻1?���?e�vۅ���G�6��~�8h�,>��$I�I�����*��vxǰ�S���)��"zը����\(N������:�[�l�����!3`/�;����nb��u:y;�=�6�U��T��r<GY^ʛ�� [�>�H��*:b6;-�l=׹\��GZ���B��1F�:bm?���g���&? �`�+hO$/\+�?����P��/ }��J��g4䙮Rw��o�ڕ�v^U��O��>��&��Ƨ�<����#����]t%��>f+��:�\㠹<bxY�S��/��9��ѵ���,<:�.:_��F��C��%N���ӗt^t�]�
���*o���^?�>:��}���T^=���6c�Ö:��>��p��.�ԏ�A�sڲ{?�n;��tK{�yt�e�oUf˼a\�n�:�`���׺���g�LH�����-^�y����w���IH�5�.e���@7h>��\�x0Y�:��N�va�����4�!ev0Ҟ������7��ܡgy�y$ɍ�{�v|;n�pD��܇:�V"�µ�7n�o!뭜}2����� �!����>s �b�x�-�4��/���g��u�6��2����ͥ�A��iBYU6\��/�']8e(|����C?Ot#�xq#�֡ͺ�^�4��
�q�߼ ��.�آEF�x>�J����J�ɫ�Ks�	��i<l�e�|d�7��}G���؎#�Es�]�,�;�s_��9pp��#�C*/��	�W+���Q�L���Tbų)_��DV��Y��5oq�·������\X���QJ�p��E�l>�DF�ӓ�kvk�ip�u{ɚ�sh��)���H2�ͣ7��0�����gW�FOC���<2�-$��������D��]����<jC1|��g/2����P����_}u��[�̀�J������dK�f�`;���cʮRw��cZ:b�����8��YPn>�ϔ���aU�3�\0zT~��[#�v��A%uT���@�2#7q��I�<�7���oADbm Go���c,��}����ć��}�V\mo���K��Hse��:�-~�[��G��n�u&_L���f_N�O����0��e|p���Z>��1�a�x���{��U9��X̚-��<�1g��x?n}����k��w
�!�O�6���ڠ��x�|&3q̣����SL��@��I�5l>�4�i�ä,�a_���{l4y�=��І�����:Uὁ�^I�B�C�������7����b�![��R��C�y--�r���xҿp�}�K	XN�s��/�0��e�g|iC[�}�o���qL�`u��!O��
�,��C��5
?�ô$�x��K��/&����K���ɂ݃$��O�t ��|����>��/�<��vWWXä3t��:�<\a��e�b�á<�^r��Hg��d���9�ߜM֞�/6a�K퀓�XP'_�O�[|��.D������/�}��g��Т����k���1cx����-�!�����ӷ���:rKt%�]����q֯��6�ri�G|[�H9� �\��F|����օtJ��W��sڐF���������׌pUCJ&ia�|�qjnA7G�ұ��PLQ��۹���m/��]�V��λ�*0�j\}q�������i���ʶ�s�ۗ�����:�L�[l�LC��U�Npy�q#-�BH�u!m#N�������&a�=�R`J��l��ӣҖ����_�W:4�)~1�3�w�?�����᣼�~����}��Wt,��@f��DL��D���t({[�e�_��mPN'�-al y���ǕW��T�W���tή��[�,������K���wx|��-�>Ju���:�g��6�|U��K������AF���d�f�JZ�緃��b�4�&e�I�t�V?s]z�~�q�̠^�ű/3x�,��c|�>8��Y�It���=T~�k_�X�l+t�pC��g���ym���F{=�w��~'�ِ�P�Aa-o�p�=��^6��g V��_���� ��ψ|sa�]0Y��9�h}���.����c[���U�y�6�5Y�fsdn�m�o����*7�<�1o�+[n��m���,��r�+m��{t!�A���Z�+�=��n:�:�_��s��[8/�1����|y�
�ԡg�3sD,M���*)�6#L��
���d�yp�zW�$}��<p=G��sm�VV;T'�E�����K]�����:~_ױ�9k�^�e�����y���&���q�rë;�����P�K��@��aa�XmF�s��l���gܲB���';({�np�BGY�������~1,>&�3�u��E�|����6��-�T�j��q=��S����7�CdH-)9����Z|G�候�J����j��=�m\o��ZIu��i�k���x�w�\��:/�=��b8��g��X}�
�٠OC�r/ٷ�$C���m�kpRE+N�Z�&߬r{<�gw/q�� zɻL0��7$I�c�/ʔg�1i�5*6��|�@t>j^>��ꫯO�tx̣�wܙ��s�3���T��G}�E��ӑ�^���~����O@N.(�B�ӍsD'���b�:�ՙ��}��G��w�$���ß��=[~<�S��c�/�}����缁ʝR�z���6��Q^�Lj&�s![�]�p�s�ԍv�f�4��$x'�zF�ډ�`��8D�� w��l<�]�ݼ����=�Y�����A��V�ؕ�`p���#�x��o�9$�J-��d�C0�s�H_�)�Y@o-q�3���s)��_t��r�Y�����L���y�4����i99	;�1�~��e��6�BL�����EZ����Ô/���x.�:K:*�W�љi��S~�ӡ����S�q�);��V�^��5_#>�5���_|c��B��U���Z|:�Փ����O ���_}��������-So:��lXf��l�q�2���?����?�)���ί�o��V&�ʺ۽7y+~��733���ml���&m*o�)�v��f��!�1#u�b8��m�{����g,k`h:��/�=��E+�Ooq"{n�1�=(�LF�o�::���Z�NY,��ʞ!g8���~p�zqLZ��y�I7�}�u����ӂ�S>�~͍�OZ|��yT_��ߢ��������@�7�6�_�U��X�<m��.�脽.���ͭ�^ڐ���6�.]Xwډ�\���-�Am6�s���Xn�>�V���3*�p�%T�mG��xd��:�\�1:�׫���3-�v�o���n!嶫�4����2����y^�<�N�b./���J�I�4�)�%�3���=c���b�ҚC��W��n��ޤ�9�S�x)��(Ϲ;s�����
r�+���<+��Zl)�Ԋ�q:���*���v�����	��_n�3�,Lm'�����4X�� ���]�4W@�*����1_����'�@����0���j���#-�� ���cԨ��Ց��3=�k�k�ܬ�ż_|�M֔���GitW�W�؏l��;L�S�[�E-�l�F0��H�jt�#w�`��S�%�8l�\���{w7وO]�p9k��7_~������M�|���z��L������_���c�?m�5H�k-�|�@�)�&�.by��ߟ'^����[ƺ��ci�o����2ρް�C�2��'�*��7��E����ܾ�i�1�91���iy�]�Ŗ'��f�5]�:����s�?������q�tfԹ�e��2ny�=[�C::^nn��œ�b7Ό�/܄�&	��i_:��,���>��o�}�+h���@Y�O
=�1֟p�=zx���x�37Q/yĕ��I�#�,��.����6��V��D^�Ag�2C�����~�wCd�0\	�rN�8{�.h��5f����.gLr���Q$}}�l��#lxu��/͠�@W��|H�d�;f�ذ�s�oNp0x
6�C�xZJ���p.�kI�v|n��&�~}��5ov���r����sm���to��|��&�`W�0�-%���i���W.��ʎA\¬��eێ���m�������:'���H�HM�yb�z���F=9��,[���D>'w��A���+u�x1�����@I|w��*czt=�gG~�O�l�7[�z�hAK��97�sb�ą!��^Q�+�x=���=SҾ�:��ҡ�� Tx;�zɹ�S�͙a������b]̕��J��R�Ѩ������@�)_�:�ߩ����C�G���d�g¢��%@�9R��t�Jr�O� �w�ٗ���N͙��?��z7"�ų�-���;4�o0�HŔS��4�����"��Q->�V�)O��kH�����.� �А�ۥ�ٝ�u�������':nf�XS�#�o���������*jt�e��\��W�* =*����/��d����-����6^re$7����[�f��������;��y��8��W����/����7�=��3欦��?���`���Y��W���Z�r@Mۛ��7�4�QDL��,s1lm)�]J\���)��Ói�M�A��(����?|�e�b���~��N�iCR<˺���ʾXnOc�c����e"�u��7����?��t#�=�N�p+�q����n�3���}����ǡs�ćOU!�x�[y����o�ʇ��^>O_���O����?���O��c�pt���S���������	rs�-��c�4̍�#���<߮t�X����2)+M:��f����'������xlj���<�T������_�/w�]���6�btIC+r��C�%l�"�O�'��/�"5o��ΓfƦ�[��'9:�OY��ca��|�<���_��ߺ�����������M��2��	,���~��$��#s��)�)jq���3>vZ]Z�>8:(.g�x]{F�G
CGv�{rdn<rQ���I��ˇpp�ζ�����ڐ>�&�b?�Q{�$�2sQ���Yw�b��M�*T�+�X+�B���$�"��� 4\?-�E�
͂��?^�N#8�����M쯸�OR�4���>l0d��¡(v�"�(3��E�L�r���Њ���#2H�h�E��V�Թ.��8�'\ͧ�.z��a>$~�&oKy�˴}:�����Mc��J���|�_Q���]��#�S���,�!��ȚK��\�<��GVg��њ����!d��q��`��H�����jf�X����_�葩p:a��f��Z����%_�ɡ�mrə�����E쌃e��:�.��6�7�6,s��u�������e�y�o��_��,OR��z�d�V�A����l����H܁�v@]�,���hbs�]���c��b���u��l�8����Ҧ�b�Û2���ҙ~���"����k�`�>o�oϻ���Oᘴ9�6�~R����e=��O�0��㤃3�.�9N��<����s$ΔWfΰ+�A:��ěE����)�$f��ch���SZ�?>���H�=��{�%q�x\��������������Ol���ͥ#��\�v�.�v��3�h����Bd�$O |�[{�Y6�j�ª�M�^������W,�OvR����M�H:<}��Y����U7N�Ο�4h�+7Fbl��� #�|Cɗ��g|�E�V���<��M���EBA
[h[,?��䍽8^�+n~�[�:_���{��_oX��i�&�死�s�e��7�2L�`PWo�_D�ώw-�4��9G�j]��<i������Y2&�4�~�f�wc� v�Zp����J���Bc�B�L=B��N�u%�i��<1^*���"���U��G���d�Y��;/<�С��]�v3e�#N86�����C��F��D<K*���\��ď���ij��رۂfJ ���LT��G�v2MP�UQy���c��r�Wi��b���`�6��9,���X�t��8�z�j�H��k�FCg�L�ӱ�I�ȯ_�7���Ŗ���B:hy+���R��إH���::_��X�5�������=���	��K����NZ�q�rvλog�|��bft�\���G����7:y�����_3�u�]��|W�K'���;4�����O0����F�sP�k�ox��`}���ʇ��8`z����;���|�˂8kG�8+�>l��AC������;>�
�'�y�}�q���?�TꇇH�ӚT�����3��Q����w����E`�M��	�`'b�y70�sq�Q���|���I��{m�2ܜ��'.������u1}�M�E:s�9|.}L9g$c�+������ҟ�ֳ����ۊ�[v�s�����Y�:^�zL|蚦���#f9�p����>.9��I��n-�$��r)`j3k1ŕ*ڰk��G]�N���nsCᛋ�z����n�'f�]Ю�׸�̓��%��o��v�O��MdxK?�,�a�5�3��Q��ζ�����״��#M�\h]+��V��P���>�go�����Sf��xxq��\�e;��g&���G����ߖ�A��RY;n�'�]lCÑ��Ro���*!��Up�q�SF�9�O`׵�E⾵שׂ�����S�7l�����?��S�4�&�]w��˽/�9�~��[���KU$�_��B��&X�_І)��)�D��O�P_�9�Ү�%���1^�Z�W��X_D�^��a���|�ߧ_�N��h�ιM��,m}�Q��>�4��Mx,�[Z"�����r6�]������`�q�x���⋛L����S�aގa1/��nC�[)�����oO"

&R�̱�b'���D�X��P+���'�d�L�#ox��,��OC�\�7�tr ��n#�:��t-��s�`+��<��;>���8��v��)|a�vSE�K(�('א_���J+�%.�{]LG�� ͓�ʟ�M�t�����fC� ���2|��ɣ�,�����	�F������o�a������"��v�A��{�F�#����D\��7g�<�+��e?�K_��ih?��MU͋:��������\�u��z�C�3kc���6�c~��!/Y�|=�n����\�:3�ؿ���/�Bc�߻H; �k��AV�ZW�ӱC
���1w� M����ym�����Aۗ��-WX�E.�&߳i{��'q�L�����3������H��ӝ��=G~q�v��E���~�:�A���1�A����d/�i��8q�� ����f4?z3 �4�g���{y���.�G�u>�^]�x��/��w�!_����d�_��-��F گ9��cE��ə��\!�ip��F������{ϫ4m�)����A �SU@���M��@���8,Ϟ�f��샶~���n3`��$iӬ�N�L�Xg��\�H�h��.w�ٱ�^o�FL�I�?uZ�u�q�]�7>�cڮ�rv�ud�d��z�Ƹo_������x��/�|�#�������������FPF����$����ʰ���~ɿ��:~�r��𥞣0����K���>�xlRR�������#�k���1nl�u���(ȯ�$]ļPoE�?�����Of�N�X�CWa{p)}����_<�F3��L�;�c-I���m.~M<oǸ~��k�3'6\+tU3Jj#� 1��<$iP!� t�\���Y,ȣӠV�E��WT	ӣ�"��B�5���	rIɎ2�fi�O���:7ʑ~���/������/�#���wםo;�v&��@D
G��� :N~�����?g��0g/�+l���r�����y�a��B:-��Q�#�鬿��s��/���c�����_}���W�������޳�c���~�]�y�x0br���rK"���8���+�����-�QD��u�!^=��\:��,7�y�*�vx�Qn��}���h�����{����^��|:C���J��Ƭ&q����k#�X��tS�&pa��qԔdF�^��X�mq�6�� �i\s�Ӵ퀿�� �p���6e��SF[1�SW���zmhd�~��N�OmN��o/O9e�Q��p��e�N��Ҙr��F����T�wM�uh�F@'ݙ��?tG&�=,ӛ���o�N�7��C���%�o֡�N�^���O�~��ۨ[Cy�~��Eɮ�-Lu�,}֟Ao�-o����'��^}���ŵt�FA��=Ə,���U�`�C� ��Q���q��}ڎ�`����|����U=��mޤ��yx�@�}���^&p7�?{��b��V/!�o���)'~�%�Tޖ��.>4g�t5ra,�0Yθ���^��ϱ�)6a|�n�菜!��o/x�����:_|������d{�ܷ��3�����*�Q^��#:�+�R+��=�0�n�p���+�g����K~���/vhJ�#�^�����ȅxS���d�5�8������ O�kz��	;���Es=?�P<�C�xd�k޺FM�vzN2?q�H���p�L&���-υ�c^;N�h¨�	v���*)������r[n/)4ϪҮ �y�o��џ���x���c �5��-1�(W���ԉP�ͨ�N^4^·w$Ί<�����^���_bA��1�O�P�V�/��h��k�ċK�֕�eg1δ GV�H�t vP�ƭQ����kw[~΋O�<ς�G�|9|�da�l���x��u�G�!b�Й�W�ZW�c�^R$�p!�i9:'M'�)���q��w��<3R@�l��<uL��茋�~�~�0;s��y�B=e11�H���@����$Dmc��	*�@�ӈVJ���-�d�7�ݟ�!6z���/������ڂ��r��f��㙸��K�-�� �`����x�G�m�^+S�x�7|Jlp��4��ڲ���E:�ۗ-�7\��i��,P�G��i|�˫A>'�V������,���ɲ��E�ʬ��8.�W'�Q�����C��Y|d�lP��G����Z羱��u[���#W_Z���������DdË��Y�2�)�"����z�~fti_�4����{,+;%�X0�'�lj�O>:��ty�N��2��J�3���=�]S'���(�~�v��>u�~�7������BHi�"��s�}�i�M�L��/y����6G}�����u�����z/osSɣ]0�A�x�yc��.x��_��=�2�[�Y�ʋ_��^��9~e^����������VD:�"�F�-�ܪ���Y�T��>H��r$�t�����$���<�'Z�-r����LX�o��@&�{��X`��|�yKم�TS�a.-Jj���Gl���hޕ^Hկ}�I=�X-i��Y��ôHMe��r7�r�D4Hi�"����^PC@8oEW��XUS@�������l�e�N�!7��;�B6����9��"�<*�q�\��C`�L�i�ȟ:�m�߬<�	�滏<��ŧ�~8<�n�;��4�,���@>z�MR�X��R5
��c$Vl�J3�_�3�2�F�V��MI���O�tB�ʵu����<�Sv�v��ÇOx�3y���_�`��W��;��#X����S��\�_.čUw+�e��ަY6#��e��4x{�+أw��|��(l�ӭ'��YT����G������5�"A�����wv��wP�q��FJ\:�T� ������:�Y���*�	������Lj񅲸ũ�� @�bZo^	�3u�`��u��S>���ȃG;� `Ay�H'5smy���)\��l3�r!�����5+Y�L�i�x�Bm�ΚGJ>s��ύ<B�����:�ѳ��V6����ef���ҫ�8�9�':�MA�2�"��G}ȇ3F�z�[�y��8O�Y��
c\�����.�$��]�G���Ǹ�ʦ�kg�Y�t��:޳Tm��o�7va|l�]�1���i��3��q��3�ul#'��#��"t��$�~��-\����+�aO"mu�^��8��Ug�lG��H PBm�h�hJF��9`���X�ئh����K,F����;�b�q����?��S���@��cY�f��+`(m�#�8�x���N''�ܴA�/A�m�1��J7�N;l˶|���x�i�郩fP�`5��bڤ6���L�~��ƣ�x|��Ẁ�7��|� ����!�1D_�4۪r�� (|R��'���~!u��&�1��C�;�1�a�����h�N�Pi��%��Ħם�+1)��9T1i�fc��q6�'"�s�&zH�=�fC��>I������NI{������z9�Y��ęԡ���&̓*!�0��9�F.��\�D�Y�\���!�r�@^+���1f���Mـ�S�UL�;��K<+,��:2�"'7*�F�Թ�dY��5`4RɅo�˯�F� ��i��P.30�T|�����a0�V6��k��9���|�������g��ө��z;��GLr�iYy�#m�����ʣ�ѐ?3_ʛ�}ȶ՝4���s�=�����g�)k�q��y���ן���m���b��/��5���܉!mZ�zS/2f��n87�a�$��#��U`���t^ޱ�,�hʠf:T�a�3�w��[����S��~��X�ʟ��N��w�l�Z���!)�� ��Η�%e�����,b���@'�䜶!����e��ú�clͨ��H���:�L`���B)���ha7�9&=�,C��������@��q
qҀ����<��9��u��UQ(�
�әg��# .Ӵ�����d �8@�K� .'g�<k7�\98�=�u3f�NV��VY웪��v���#CU/-�νk�޳����t��az왴��Յ������5O�:��h�Q��{yR_��3��QƤ��G���׫�t�l��m��30ࠥP���d�0X�, ��˒�h�����s^��i���MN�B�x���^p��c6Ⱦs�m8X���8��oI�MwlBG�~x$j�*�\���'ɹ��f{@��N ؂�*�u��姢��̼�l��%�=�֫Ns�|���̐�W�}��>;ܾǓ��������؃v�Z���tV��pL\,mi�iŋ<U���>\�.�x�s���7g}�6���V�KWؐ����ˡ;�!!~�1TDݰ������/����VG�~��R����N��e7�	�{�v�Z�.���Y�'��@ؘ����b��~����J^��	�=�iڊ��Hõ������1��ZvX6���	�~�Ȅa`Τ���:T#�l�z�6�:_��\A�B�5�r�)�TZ�	�@.q���/����˨C��,g�,�W�6X#@�!��/�Wg�:�xr����b�+wO�����[6Ht�w�C��� >:��?ϰԽ�J�Ngk>��[W��CS./��V#�@�X���ܙs�3p6�}���Gޒr��o�s���w����oY��'N��r�}`'f~���H�+������1N���7^w���T&���%\k��6(��j����S~u� �D�ջ~�h��w��.��,u��wr�f !u-��'�M�U��V��`�i;��-
qx��ܴհP[t��E3	B���k��ە����0��{��6�X�N͕?��X�");?��$��73guxjS�sy��uz�^��s�۫�uvv�C��㚿L�èb-��i䷎ZO旦����7�მUo�6%�9,�V	qΛ�#�-�E�&�C{��[vf��4XwH[|�BkiEk�޸Ξx6��QB^t�>ӆJ\�������0����u%α'pE��Y<t�}�l��_gQ=��$Pߵ	�َ6�ЖG�UN���<�����&5��I�j�IQ�XUқ��9��!��m��c �7�^:|�@�4��ow�=�_�x���v���<|)j�f��~Pg(vо��I���>�MO�H!HtC^����
O� $�#3D�p�|��Y/7�΍#z"�q��or�ӿ���/�d�/�4x,�zg�ԅJ�TP����k�zt���de<��+{�d�������n��9��ܤtf�-a���z�NBMn�5{�\-^%i��԰/�iXɂd0w�a�#��}�z��Wǎ�����&c�e��t�3}�%�	Bv6c���["���kr������P]r�R�R��0Ha0E���U�0���l���:Ep�
���=�3#��krbz@��f�*iV�`�9��p����Bh)��-���Rf�쨗!k��Qk���M�W��r���d�T�7w����|�ٔ�x~�=�[{g9�G�tXP�Y�[ q�K�b��#&,u��l�j���8_և�Y79�)w�;����S̯��z�^_�E��­{�>���&Xl��7�Ϋ��t�|�quҫ!�0vaƾV��Ja�)8К��ԜH0+�$�6r)�:�E=Xs�v�IDn�w��!=��og�m	�ࠑ2��rV� ��7W^722W�@&�x�:0Q^�8ez�^�3D�@�@�`ʥ=���m����?j��������$52�T��-�$f�ǩz7��/0<�T�ē����;N���K�N��ԑR&Q�$N������x=��Q�1�<�L������E�mc!��c���|�mhy�Y�qN,;���p:�CO��t����^��e���hY_(ɌO����a?#����7�z֦�ڞ%kЭ=�[[ɆIyQ_G}�O�hm��L�4p� �Bj�Xc����\��Rz���i0]G3>� �[�k�/�e��{����q_e�X��"~3o��1q6���N�xՉ}JdF���֫
������.�f�c�u�Y�Io��M7�}��`?\��>r��Ue>	��Rߪ���~Y�.[n��뜙�|^I^��Wy�l��tX�dP'u=	mֱ��U�� i�T�u��O�[M  @ IDAT~����7���!?����|YO�Mu�'��3���Zބ��h��s��&�ϓ�ů����gB�Ʉw��i�O$��������+<١��͙�O-a1�R�����	gz��`���~'�p)v����uy�\T]�/CB,NZ&�5��������G*���ش���>���#��i�ӹ�8��i�V�A�J$64��l|�U��6��z�tt� ����y�a M#PW픳&�4�G}�շ�p�S:��̂}Ϛ���rgv�u&�8�4E������1'�:�^��,ro理�r-1���G�<����x�Ѹ^�yx���x��#o �F�����;/�����͎�7n�c]�9��{�ȸ�V��AH�}1�iC�T��P���e���PWζzt �ެG��Y��H�l�`G��8
֑H��K�}�Խ[q�|�iί��|$`'���w�����:a�6��8�˥��VyS'ᷢnyx�o�#�G��)e�N����XP����h����O���%����$?�Tvy�#�N6�\�-"����;~�;d��5�HN'¼�o��э����>�St�YJ�v����ި5�(�!r�����7�h|��8����P��F��|��a�ʈ��v�=�|�B�}3���7mh:��@d{)��o�M���Gtg��*;���`����:�>����r��\��\=v��~Ŷ:4���:��$��������X�t�Z��#��xGފ1+���,T��>���C���[����-�B�a��]�����r��H��aP��(x��ߺ0����b�(w���3���t�f�:K��.����Rr�ph�������].g�|��&�W��R�7_�r�
7а����7?խ�n�|�@��U�v�ur��(�K��0��VGŗ~�����v8O��1v,�>�}K����O�wo�U���1-oycuhȄ�e8�@�c�;�]Jc��j�����	��6�RӀ�ϙF����_3��6�wu��z�D ^�B�8g9[�Ԟ�o����e2\p�*�x0I�G��-^�^�dvA�I��w�֝�6q^4�2&�<�B�����,�ͽ��v�����o��G�L܈l%M�f[]����3)^g��|/y-kЊ�/^�9Gny�٨|[��i�eFL���[$,gk�W�>>g&���>������Ā�#��*\�?��1�1*�K��K���Hg@'� g���ź�X;񂽃���1^y>���l���7߱�!o;���
;0���eF�QB�U�2\�+��Ea�M���r�^���s�HdPv�8\�e�I�q�����
���H{��6*b�"t);w�q�a��ԁ>75T}�S�],>��+�2�!>`��EO{��4�)�(�r�2ɘ� ��`�������I�"0�<��$�r�-�C��6q��Υ���S�Z����j�ߧ�BV8~�i��}�:p;Tx��ɫ�9�olbvA����*����U-�=Y<��#]����2..���C����e�2>�,o��~�W�*7�C_xym��e�$���@������n��ٲ��a�\H��\�&�(;}����U�?y椏�ϥ�f5N��v�Y�F�P��Qpj�����0����,C��f�uƵs�k���nw��WJX8�������w+׆]w�Hm�괳�G��$~�oH�h��anh���8���᳾��o�>�	:}LR��%��3Ɖ8\�F�u_7x�3/8e�=�x�ޑ_��.w*�6Ԓ�xn:e.�DUJf
�@����7�}S�J�ӑ�>coD����������.q+k��"�]_zJ���P��֬:m�b$��7���+���f�"��7�Y��x	l�P�Fy�O:.]b�3�ެ^�wa,���C��yjy�c�x�H��z1l��D'=��٘�)KN�
���,���:x(X[p�8j��ù �	�qO0���^G�
!�sl1D�����u��<a�i^ٷ��aK+���/q�D�Av����uUG�X�ԭ�@>F_\��8�����H��pV����e��ec��sq�V�̞�F�/O����eQ#o^1E�B�t�1َ_�H��9"�BySn%x�f��띃�up(�ޙ���{\�୛�8\Yh���l-A�b_�s��?;��?~��,}ㆅ�l7q�]���%:*{]�D�]+���%����z��Du���&or�����w��Σ3`�֣2��3����4�:�������q����5be�^� ;u��������7��5 g��g��I3Ծ���]'�%��_�7��[yD�_�B��{��p:�w�6��uXr%�Ⲅ�-$.S4*a�ܕ��&z,���M�B�5O�Cu��8!`ne�V��p��iG��e[��[���K{O���P:*��PN��Jc�͘gW����~�X<�c�����p�eP��a���8,���Aǳ4\��:V�̗a��Hkp�V�4_ܮo�~�>��7�$�i�k�s� <��z+���mG�/:����ᚦs�͈1��S�����a��8�I��hg�L����k0�xe| �����NfD ]�h��/s�˽�]�1>���5���ǒ?���G,�����yK'��"W"�x8�[�������̞�B��G��·D���YV�ȗo4�.��8�s>+tg�N��v~��q.��I��S^o��_zT��7�W;��s.�3vsL
~��.1+�+f�޲%�z�|�z�������?�6���oQ�k�k����M���w=2������д���e&Pe�8�Fcw�-�����G��طng����S�g�A��^y9��vs`i_n��$���|��q[ہ�f�!��#Y�Bjҟ�z�Q����Yq�K;�����*�jB�8a$R9�U����i��E9H^�m�5�)�Y���p�"�K�4B����G�u������ |�[�,�ف ��#&�wс�rd�s)+�b����o�W�%�x����HM�axg|�#���W�m`N�fm�k�@h��A���(����U�:}+ҫ>$��ݛq��	��:w&]P���z������w�:__~���׿���x��8dqٻ1x�V"O6���֌�d�ѕW����g��"���v26P�'������7ƨ�޹�X�#e�DTX����G��ֶ�u��9z7�'�ĭ]��Y�6D;fg*����p���Gq�Lխ"����cʆ�cyo$ʔ��0a�9���\D�����1^������:��0�a���#C@W_����Al�����4Wg|��x�?��ߑWq��5��KY��t�t&�e�8\���%��q�&ϊ���޴ˮ�H�=�A�I�V�����`���Z��D�$�U@(��yߌs@���Ϊ}��)2"222rع�,ﺁ34�\��G��7L��*=�q��Su�i�[�/�őB�3��<��b&�8v�?�ۂ� �e�'3n����F�� ����-����c֤���CcpO]���I<H�HI�@M-�B�}�3���2�]���^�M��c���=���v��������Xgn�|���������:oV�����U�Hi�[t���n��xcӤ�9�!�/֙oc�;��NwYr�"�#��u�L����w�#�}�ȯ�I`�\����M���G�+_�����Q~u@��H���y{͋YW����8K��X�u��n�b� ��S���J�t�?/���)��	("Ɇ�;m;s�W�7^5�D��l3�"�VΕ����mɥJNH�I�=�/��B���)�h *����Ȫ���p�Px��)��E��>��
��l�!�s����g��ҡ-x"O�Yc����8a��������Aص뜌��!�<+���t�EO�L	�/�eeh��7¯�`-��ܔ��<S��u#|� �r�	y�r�EՆ��g�/�㬠(��6R�o�}[s ���]xtx׍�_l�x+��[/^�W�_o��໒�Q�pU�*�|�ƫ��g뷍[Lݟ��vV��B�,Ɯ��y�RLg�Է�J|����s�2������H��2M?yR�0Ԣ�僒���}#����l�z�z�����c�Q�mdv��?���%_̣�KGH��h&�r�m���.d#&�sƇ�?��Q(K�yy�t6N)S�jy��p�4�Z�r�uN�9#�?o��C#�*����	B\�5��\�aIf��)��.��UF���������F���c��ep�/\��<$��z��:e�K7iRO
�gU
�:V	w����6p&���)����neEg��û~�^��X�w�˳�]�G��8���t�Ng�I'�wqʌ�z�ۃDu�JC�|;~�'�A����3a���3dV��=^��|�W�,�g�i�9���O������󲞽�C�7����g���i�ã�H���
�Q"��j��F%2~tN�vY����+R^��V�K�'о���[uQ�ʵ���O���/�ԋ�sζ`�0���s��=x���_���g��o�sΠ��T`1#8.��x�A��_����UjݙNl�+�@"�� 3,~c�=jw1���u�*C���}S5���Tr��J����9�-�t�;R?����{}�+̉�}���a��>ξ��\�Gyyy���w?�ǟ2X����]��7!��SF�5{w��?eD}{x�@�~�|�]Zx��|�o&�EF��T�X.�M;瘑�|�������.M�Q��)�Jւ���߿���d��"�7�_���'���8�>�%"Fj�'n�[�h�NM|�,@'�L����,�A�Ɨ3_���f6�]3��	�\"��Lѹ����ܼ�A�L�t�"_\�X�U~RN�9�]����.�4���%o��	N�DS�>�-����4⫅>gj�l�t�c�%g���|��*gk2��4Jݠxי0�=�G_��t�%�c�$Yܼ?zy{�^�F��\��;�\��C���0i��+.U�tT(e&X$����`����f�'�~���W~H�K�
�3���H���^��"�T\�B�_ʷq���Â����m:��8���(֛C�$8d�I��Ȁʤ����Rj@��K��D��3h.�~B��ůXr� �c���!��1u��?>�7�<6��XU�R/������"w�Xl�*6��{�~`A���NQ
w&�u���t��Mc�ܷ0ġiVJS����oe�#<��й�!�}��Y�q5\df�8��^�8F��?6d�Oz����D�,����?��Y܇�ⵛ�Z�D�45?��_�4d�k��,���Y-~������Sy�i2G]a�7���j�i|�����|��7�i0΂kx���'�y����o~��	�y�k����%ߝ��T�b�į+OJc�n�U��t)3V�/���`Z�u���9À_�U��~µ�ȃ�Lq��o񞰍��A�}����2��{��|�c�=������>�;�+�8���v���ن�7�ڲxB9�S9�x���/�~,�-(.�z�q�*�� #�����޶%�^�J�_e�-[�V%���1��L�S#�MH���耳�m����B?�vM��(:={��*��	2ǡ��*Zf�җRХ�~�D��!���}0�	��E~�H|S��
����%��	pp��=��IJ��O�±���aip�� ����o����$&-�ɺ�L�X��R?�����-�+�E,.��h|�l�5vh( ��xͨ�:�H��7�
�Є!!Zw��(��img\���H��d^IU�d���N+L������%^�7S�S�(@�#������l"�����8�bxn`���T�4#	ՎBS���4�T*�F�	12����s@)�G�~�m>�!�a=�@Мb�Aa�7)�3Yy6�is��W�}�Ye�������pr���o�9��]����͝�*�ӳOHﴷ#+�(=ܕ`�A���I9M���J��֓�����o�ZΤз �C@�w�}�����K�V���Q9̡��r񞷺F���1�� ����KN�~�	o����F��.�5_~��ͣO����~���tV?r���ͫk>��m�شq��E�A{���<�1IM��k��(���=@�G��2p���Rb����e�
��O�=�(@&�1����xW��l���yȒ?Ϳji�tMՎ���<�6�����A�ez͖2e?�K���V���sCg�r�Cj��S�i9�/ӈ���줧��_�pl�83\>:���v6n`�#/a����~�^�_3�����������1�zDO��o��6�L�m�?�寛?�៹��Y��s��P��}�=G%���ci�bH�cB�N�C�9�}�q�s�nM|��r9I��˯\A#|e�S�>�86�KKwٮrt� �7�o0�n��X���{�|�գ"4Z/��o9bֻ��{���u�I�P[z=�R��D�
9�3��n��T�l�	<ed�*��s�=e��|k:Y1�Ê�M�ޏ��b,�	��8�Y�)J_nL8Xx�f��������^���=��v�%�v����K�<_�g=̞ghqv�-.����Q#����f=x���,a��3���A�9�#墘=��/�lS�ҤAX��?I�o��=���3ϐ�#pJ}��mH��2ox���ȯX��0�~(��PP��5l�8{iir(�K�\�J;ˑc|�2	H�T��I��
B�=��i�u� ӎ�q�!��lk��pf�3���;Ò�$?���h��''�"�P�d�W�C��r�]AUX�E�ĶӰTI��7��ܝ"�2~s�$���|r�f��f�)�]4	�t�ࢸ��K{��u��tfD�ŏ�y�$��M�(��Y���|��R�Yξ�93_��)`R��;4@Oh*QbH�8K����y�& �Tʋ�}����~��&5��8������f�L�nO��j(����lP�{g��ыw՛�҉��Q��s���=����bf	��G�>�|��7�˷��� ����穼v��~�q�[Y��q�G�e/��A���0��m��\Mey�}Џ=��Cx�h�Nʌ"R���?�g�c���mg���e�(;�O�)^�ڪLp��M_�l�VM/.S�,�ʮ��K7��^�h��M�x��S��5��N������5���ih������Or�2��w���LAi��d(<���]��9f��,_�������~Ɂ����-3��+X`��R�uj{��*q+�9�3�����x��mn+�	o��ޑ:p���['>76�5S�����/1���
ZO���{����I�e:d�9}�y�}^���Y���5�탤�x�2�N�k/�c��agЫ��E8��c��y�?	�U�?��89�!�HB�Г4C��i\��-�	N�	������H��L(m�:ֺ�z� ��Ebl��?�P���H�9�?;vVJ�[�����?s�D�H'��jT�c���`�}�]\�֪}{� ��O��-#��M����]
�\J��D�_nK��(Om�O��<ߨ�4��5�����h?��t����O�x�y���Ap��+4LP�٩XB\��-�`wg��{�:���q>.�)�27T ڊ���)<׹%[\�y���>��F�O�ɐ��/ح�p�4|�.-Q�� ��1��ڴ
�N8g��������
W�Lc���z
��Td��3ari�Z�����Y*��~�Jb���Ĥ7W;�����b�+��(^���f�����c�!����ʽF4����^<������ZNG`�C�h����xi|Q�Z���=1`"^܇�%a��<�e<�~d��ԕ�z�
��׺�P�pO9*��Wy�~W��5��7�<nå ���C��5�����ͯ~�EF[�;��tX.���*�u�xɾ}�:D&Z�%�����M�w���+�c0L��t�UIi�Q��"����g�UeȦ!�W���-70�_�q��`��}
�8��i[��e��kX�Ƅ9��E��o�Jޅ���g�_��?i'|�f�Qz���?i��+�H�=�]��)���o^�h@z9 �/�I7i�C�r��8�X^��	����^�AH��X8��qʻ����i���s�!_=�����}4��\�i��W�6f2:T�ճ���>��;{`�S�IAgf��2�:������T��ȸ]Ч��]d�As�Aa��a�C��̀�)�}�7'�i�g7���7�{�5�Z�7�-�֍y-�0��ȟ���0K��V�ֲ�HؤI��&��@	N��)G���<� )�i4a$�/�	��q%����1��o���̺ʢ�X�^~��:wō�O9?�����q���o7��{f]?{ >�e�q�����6�#K��3���e�e��ϒ��9����/������WԎ��G?���n�� �p�ؚ̬*���k|���A��� a_c�h��b����6z�GǼ�!G}r��^淡TB(���t�
Ӟ�=_4��deZ ��{O!_Z����"����ְD�4Y��%P�~a�����M�]�tv�hۑ9p�rID�$W�0�.�ʁ���b7+�Y?��1�Y%\����g�ӈ��-�(Ǜ­ņG�T>�'0	�k��QA�׬rEaX�3J���NA��yL~��,�0C�gRS{F�eiֶ;h|�1�i���	�-Ii��p0���6����[�f�n\�'PW�}�4��/��N	��	�M��
�����S���]~=��[�W*9d���b�[d]��#7���Rrh� i?��~0_B����,ռʆ�W���S6�rn�S���"��)��b"�1��S���ߦ�s�ŷ8��<�/%��0nܶ�кʝH�Ӡ-,�d&M�g��t(p!ńq�>I+��8�|��Jy�(1i'�ܻ������ײR�(|��̂�r��"\�-��^�ׯ��	{��7�<���U6x��t�吁�Y���78��
�����1��o�{ĀK�.��v�:�=��1�t���q��z��%����,��̂y,K\l/���x�w__�g�����<�K}c�2)F}d9ʍ8e�+��<�5ħ-�A\��鵛qm��nG[|	�(Y����I��h�?yl3+W����VW�g!,���	n���s�=�Dޡ�"@2��>�Lq:@)�GBr���W:o�O|���/���J��u��O
��!Ӷ�ݡ탬��!�Gg�4�Տ�h] , �# ^�|����.rs���7��<��2!�:	�)�c�����J}�]�K� �e�o�*V�v�~�F;�x�pm�Q�,�[��c=�DRD�Ӟ�g����Q����<����X�����1&�)��z>z���D�8F�L���B���1@��b�J��:�>y��\a
\���	�d	[�T^�b|kƊ?�{fJX��H��ٓ�]��8���fM;a,Ż�sVNFc�[�-'KN�:����XvB�*(&�uM�ДD��<��hd�����������4$�I�_\xV8"0�/���*��J�O8��x 	�0Қ�k�`RL���>A����F���-�����2
#)i^o�8��e�������~��R6ܸ��B�P�D�Q�s��6�\ax�
���*�N�ǂ��C�������'�4n��Q�N���{g�Q�A�s���Ğ={J��2��N��|�G�� @8CK�#읛�yB�����S:��x�ϳt{�3��y/_L�ո}����y�C�|5|�cJ˔���϶G;���x'շ��h� r.q�YCżg�v�5���i�i�3aG:�c��1��%��ye~�2e�ߙ �^�1�\�y�)�T]��'��-'�H��7NMx���i�L�^S��3�z˺j�{C�^^e˂o?>|��R�ٷ.I:��
������A�o8�"o2�U�_�x4��O�M�s�a�syfע{ҖG��,��ܹݳQ�����"�n�����P����m�@��#3&+�5����������̸UV��&h��"2��:g�<�
��J/<�<i��^��~�t����z@Y�i�x���m�ʸ���@�uE�#r���@�(W�s�y�g��9�D����#%{�N�]'n�>?'��,	^�����>]��Z��eC��i�_x.���gB�!�ܑ$�3�@�n���4V��6���U2!v��#��lf�ɫ�-��0����&ixc]z,�G�d/1�3�a����gi2S�[�~6����+,K��-R� 
�*�( �L���I#-.l=
Q̃EI��P��;����
SA [dG<k�zEaс%;t���=l.a2B�ܝu���wt��:�<HJʘsEb0X8�.�<�C��T��g%�J?Q�EFpGw�G�|V��!N�Yy	H>��5i�0:��&��}N>����+-b%
&&<��"C�r�$��y�'����gs5��)#��2h�`g`c�O׬y��ۈ����ƭo[ҭ�>�|�Y�q�S��u-��b���ȫt*X7����G��;�o��gD��6���ExNf��<��������:�0��pF�?|���/��u�dCc_)]�<�@ȸ�>r"� %�MX9�mx�йM#=�k~ӶS7_�WE����[XF�<ɇ�ߡ"<J�v���A�(9d~h3KK%�4\�=�>a5$��a��{��a\�.�	�4:����|���ʴ�j��/9;%�xGa�3��S~��[�&|��˻�:q�6�����kݰ���D%����������52�p�gk���`b6>�pC0��7N}[:zlO�: �_�-}���dk8���L7k�(3?�].8
�V�߉+߷���5|�"/y&8�(��I��oxi�fN�p�=W���- �/:�	�4�)q���f�2	�C�J;e�*@Vi��q�LR_����TPa�]���e����O��9��[��j�3;��_`�]�/I=c9r�f�K�]��7O�s���&P�w��ס�'��+O��T��<�m#���?)B��6m����>Y_ 0���'64}����g�-2}�A�3����c�������7/7`�F��%'�s���_r�8�Pj$�`-3���8�K�����pߕ��,n�#�����p%X6R�|��
Bm�f�(ꈽ6,?�i�ڤ�|3ʥIq�buZ���09e	:'�ju3k�ѹ:��fq q*˼:+��&i(�������_�T�9I�$(�pf�W�$�j!A�8�#0��%�
Xệ�d* h^_�3��pR�q��#�o�@[�~���<`1��yAh���:mjb�i뭴�2�`�����>x��gS�?��n�N�E\�~��e@�[W1�hW�����rNXLQR����j$`��f�|��5K��~zҏ�2�����B�k �[o��Zh˞i�eh�)��##�U^H�s�la(�*����?n#���Y���"�堗� W�2�\y����P'�+o�_�JϾҲ\����L;~��X��w:,��*C_p0�0���0���4�y�Y��w��}g�|���|T������
߻�ǐ�<q���Ѵ7�>��tC�aCM��8�NtFJp���=�'�1�f��0j�W��C�e�q��z�fw������8��LzB{�=��0f�ԩG'��]vr��E��A��g�b|�{~��[ȬH���T�.�ST+�	V㔛�NhI;�I�SF�
fbc���Hp({��AH�k����K�E��`W�ܶ>�l&σ�ǩ&��b�3M�ӯ���B��7E��W�ʌ��}xV<		?�0�r&4|��b@����#/^�6I�ӜÏ}aC���a}4��L� ʶ{ި��W����6��r�S�_�����ͷ���W|O��oz$�e���	�[��5�ӕ�2��&����b�����91v�Bg[aI0t�@��=Z�N�ы��w��^�6r�$���c�L�������6�F���=��7����幛E�9\�U0�,=M�>Sd��dܥ[F;�g33o8��l��%�A&؋1���� �vl�vN�'��E�S�(�=���f�-
Ԏ��5kԑ�<R]�u^�?�AD���Z��|:$ʻ�S���O9��gX�á�5��ŷF��@D6���ӂs�GT>��l��EQw�G.u��2:b�����T��;#WW �)Y�-.P����vQ�31?O��6��v5�pS�C�nBJ/��"��m��0�)��9@�>D�;�|�o-�Rt��t
������e�\3Q^se�z�������p�S!+����P^2f��+ζ_V��#O�A��(��<��P�	qa��HZh0
'������O�W�ͼ -�F��IL�r��Y2�p�����l;��a���]�i�����C����UqӺ��+������14acH��X�4��,/	�D���I��8�M^�'��c�X��u�u�6����)�pݔ'��?�E߬L��|*v���|-C|i�'m�Ƒ�	O�MoYſu2a`8p
���-(O��?���e(E_�]K�r�M����+e
��q�0y�q&K�8h�Gg-N������3N��qc�M�+���w_�b�&��>�[���Цc�m�� ���b���&A�@~I��l��ge�� ��DJ�JТ/��ʼ0ŷ
[|��3	�7<Z�CM�:�u��_����Ls��ҷ�Տȫ��o���U�̄��W\���+�j����߫���K��x�cR<T\�qD�|G�9����ESՖg����r��^�7��i���|�+A\$1
d-m��<�� Z,����-~lܒ=`��3���0����\w��;�M;����P�g���:��; @�K0��F����V�~�ե�k6�k4��h0�A��uZ�v֧؃`�Q	��{�^�f�[ޔ���ҽ8ـ���M�Lo�0-��@�:B�L���/�)��G��d�S:�#_7�a����>�{^��y��
?��o6��ӎV�y���kig�aQ��Hl���Z���6��th��C�&N��PJd�oq�h|=[�����5 p�h������(0��('�e����D�@B�pMR~�k��W�3�,����Ԧ�[�w�>N9	����������̿�r>��͵��4&��F�|��㾁C�Gi�Z0��̿ƀzŲ�F�O5�i��q_@��q� ��p���#@Ҡ�o�,I�`��U����~����X%%�qS��S[�[g��E����6����W>>��n�-�y�𲳗*��0�"Ò���nZR�[�u�
<���������0�t�f��Nt3C�8�ƹ�i�f�#�uch	��-^�>Z�p�f�ʻ~g�t�ohZ�X[x^�u��+|��2eN:���,��Ѩ�&s�i�'�Z�8� u���S�r_�8���3��	��,M;�e�Qo����V_f=e82}�w6Mک3x�ۓ�{�L_�z̀����v�GX��,N˰͟�|n�?�c��_�"��x�Ih���KU�M¤�y�S��gx'ov����0��w)?~2����;X;(���G�����_V� �y��V��8"���ꍁ�3.:�W^�J>���/�Bs�����GA��ѶB�L��֏[���K{y���+���$�T���?�ɢ�O^l��O�����C���C�~��/0#v�L�ݧFY���n�'ʓ��훫��EV�V��:5��A�<�����<�|	!P�o���}����{��W��;`����[d���xY��>������~��S6O���O+�,�zN��MÏ6׼^�>��P-VRL&�.�
�LӤ�X])q���ۻ��sȹIL@� ���Ɛ�����v�z�jv������«�̃�&�m,Û7�[`s���S�_`�^�1�k:O7�R�p8ܖ��[��j���Cu�����|;�6me����3E���s�/����u?�lc��J'��`B��7�ezQ����7��q>7��O6�~9I3���\��p}�Y���;�ﲑ~r�r'd������`Q/�|���X9A���H��*�5H4J:{���/8悍�6e���c����y�z|��K��b�,�V�T�#�H �*��w�{*�7��(����H�I�����ȄY��ʀ�¨3,JP���"O��I��P���`��CM�2-��|�g���Sa�S�k�I1&��� H<C�$4�eq�a-�6���-��v�eLg��`ڙ��q^�+�0�ʒx���(����3����s���}zL#�u��rvFQ��,d���a�Lo��q�����K|]B��Y!H>u��8�)��cXD10�����;�0�N��#��7_��[��H@��'��9U�s���#a�1(v c�r0z���y�8QZ��r����o��ۘ��^�Є�9HN�{���*�<o �A����r@���i[����t�czq+����W��vp���F: 5`�-���{!�l��oԺ���j�C��*������ �^���4���#�����5���7	9=;����O?}�����C� ҈G���1�1�L�`�ҁ�2�~�'^��cm�Ѵq�P*l+��3��������{�����j�:`��9�
����E��4l��"U�=�S����..^�<�r��&]�Q���v-C�F����/�%S�z�<u��c�ğ�H��S1�$��&�x��:&��C@Y�:I'��Q�J3<�rB�s�[�б~���|F�%ƗUp���G_����9�ţ\͌��ƓƗ^+Qh0���%�̆�Aw�V���*���J���5$�_&���R${K����A�٤��%i	lY?k�%=){O��&�L�
����*��m��^��5{�.������"ѿ��b���6.�� ������rV�5��/����sF`~k�p���?eFԣ#<8RP�]6�" ~��%F�%#χGԩr��p�Y����v���%�x;�P|r�Ͱh5_R��>����U��/�%���̙����!#E�I��%?  '�ԁ�qD���E�mWc,�|��[�0����k���mI]�W�e�C�+��5\c�=Yn��.g���2�:�2^g~��8�ޱ��c^aIC�M�1_���,?T��#i-NQ��(����7�#.>[�����:����9^�%d��5F�i�����i�6��O�'~�X�~��q=�\	�9��s�l��u6��1�+_�)զ?`�SxF�'}e�G����Ge*�"�����3�~A{�����/"�a�z�K�r9���t�6���z.-���v.!�F'��7>��XKN�˲���&�DI����)u�+�/�Z�~��ه��{n�==V��K�5�����ǅ[h����l�\{��q���Q�׭Q��˗�	su��s��{=R�s�l^w�,�Q�V����4Z�wMԋ�.G���?Ğ8F�U��3l���'������2���分�>ũ��a�@p���[�ez�Zlʎ-c!\��S�$�k���Ĉ"�m�H#��L�a�!�1��1e�S��x�+_�g�����T2y��oY��:�Kd1H����r��YU�����9���+��6����Op�@K�,G>�z�+��_���g|@����x��6:Ox?Ā|�+\e�B>�s��5�ҩ�Y;�:C��+(V�|���-cZ�<k���-����҅����Q�N�k�q�z`Ɩy�fj4�n��r<n�/�LT�2I������(l��$�٦��ᗠH���.�����l!�ɥ�TRa��em�a<�V���7ԽˌO�����2������1h=h� w@s`��b�Q�tj>��Q��� ��PG���������{�������O�8�i����Tv�⣛4�B�p��G�
�J�S�٨�B0�6l��@J�l6���9kPV�	ǭ4 ���G�LG��%P���m+q�	@�ᚴ.[�Ԕ+�d'˝p��1-�� \y'^�5��1�̫�t֍u��'�1���mz/�BE:���k�οnܾ�?�T�?�D�/��W�Ieo}-�st  @ IDAT����L���1�p�5����ǰrU���Qy�=q�6��Z&\�}D�hK�uU?��׎Op��������/�7��`���>�f�����N
�a� )�N>'�	��Ji�oJ�ֻ� U͵���]h���$f�:�A�0g��+a�1�� ��3�/�'�#_��M�y���8[�<������L�02�B5oK��c�I�ʡ�8t�F��~\^��:�l�����LW��h�3f�;~�gg�����Y������+f�<w�3<G�V>J���b+��_D�v)�_�O{Wv�.��o�P�C�t$g�s�dUf�4��i�ȺMD�@���5Dt/��	�<�-��@�lh&:as�-@<����������F����5���4�z�L�PZ�u�Z*#JЪ<��$��(1N���P��i�aT�� �X�иz�>����b�yP�{��4��'���wz��b=�K:@�{�N��^B�&�O#,]F��ª�2S�:�I}h�����JR��SE%_T`^��l˵�$�G��%˥Ё�B|��yB�w#'�����S�N��^^Y�"솏��k��jǄ\��
V���������Th�wO�|Tx�wa�;��YJ;T�����S�ǅ����1��bH�J�2��@;�c�K!�C�,֙�?�� ���:���x�c�1;���fU�>wÓ�� E7N:�G���Gˋ��xӑ�0�yH�s�ӀR�ЖT�il���M�օ3~0<o��n���y���� ܰά0hX[ĻuX����*聒��l��P�姸��V��|֙~��F^��z��K�n�-ď����3|^:;6F��7�K�3��mY�}�˰(�_�1�sʕ�S���_�q��f���̕r~$x��1��տ��	ø�Q����iۋK��)5ͤ���s��R��q��PL��J�;\$���Sv�.�,?�c����6�s�����r����Wꕳ�M�4��ƚ�k�>�+;�����Y�0�2�1Tms�G��m���������q�8�܄նyV�� %��2z���\��#�q��ƥh��7�����MyT�z(�}�%Wu,�t�1W�0G^�%��*r᠐Ze���O���l�(��줌/y�C�!<Np��]���l3�y
_H�6$aʏ2�,��;��Qѣ�W��RG�<@ǃ �*ޗ��SJ�/���EF�a����`�1��H93xB�
M�	��-�~q����F��v��K0'mb���-3N�dp	�P�4�6f��a*/�Ӏt��dv�!�:���b��#t2�N��%Sf2�l�&Nq�T�
�
�
{�����؈M!�;02R�SW	P����K�6˷�x�H�i��;w�x���Cʸ��AOI���
�H���
�0���;a	%��&��S.�����א�M��¬=�齖�f�(]�`qo�m꽘��RL+���&�+t�[�I��#šp��#u�௿�Ӹ�2&�O���f���DR#���7�|7D�&�����$�t�Q��(j���B�̚Ldnq�23T���^���z��|k��ѓ��޶}8�Rg�?[7�ǩ��8�-�$U�5�|3ӳ�$��
?a��d��ж�~�Y|�"�>gŤër�mg��<�9���#r�a��@yO��S�����*����n�.v,���'z�Io6�z��Y���q5�l��=�ŉ�k[��y�K�,�P'��6��c��0Mc����n���^���R�I?q�c�g�1&�<ioҪ~�޵)3�2g���7�Ҭ�Uv�����i�����4Ts�_m;7�՗�~�����t{FX^���Y��$~v����Ù�:� ���7�VD����^�� i�yZI�8��i��Rv"�«��V�$0q�|\�@c�$�,���_���Eְ�9	�w?�Y�XFL��W�Ջ����
_��?���36�0Q������ �E_�E�Z��-��-�v���4)�s�$�|!�Yt��	�����!��`�"ƈ���֙#2�B$�wY�C�Z.`a��j���^�O�	L�G�=�+ļ���
V�F�apQ6��=Ub���G�1�2���OhY慢 \�^m�w����~���={��L p�O��#g�:��b���ѵ�[��#��ظ��yè�I!�
�B�Zn�	U;e�IWL�Ya��,A�4:�(�y&�3`6>�X����-hqz�8�ё�t����2k��7��\��#ъܝ��쉆�:ʡ��|PyZ���蕆�*����	�xP8Q�Ж��#S �{5��.=G�N�4���%L�n��#y1F�r5j�8nE|/���
�`2�>����<Ɨ�o�pr���I�3���_�4��ȡ��|f�:�k4I�vLy��:�B��t4���ұ!!⹜?䜚;$�6".�xf���G��hP���b~$3��� �F�P)*�Sf��a����k��Y�gG6�	��5V�Tm+�H崝}�[\P��߀Q����^ӻ�*>��㌛#>g��z"5xL��T�\j\\!�17�ov�$�O��?Gӻ3h>+�12�@��?�d}w�8�RW�R�АN:#p��i�����6�,��<����WN�����f+2����m:˷��4Z�N!Ӿ��|�vҖH�}�
kA�/㽦\�x@@.�u��8�߇��\#�e@Bҕ�@�gW��:@���\�8�;�����<�-3�i�	/aY����Q���S.�x�_+mۺ�~d]Q�������sɎO�!e���ˍ�ѱ�� oG�aeP�I0���7^�C�9dAC�j�8c5�f��bt����o�~�`B�b�%��r�-�-�S/)<)���/���Hn��.A�X�n��6����<Q���
�|���w`G�|+8�-�k�� qѧ��h�R���m[H�\����Ǜ���n'Bп��R׷��@6��Ծ�y��`5��_�����z]�I	��r<%��dW�,��M}�wq��`���٬|�ǒ���K�4I���EF�(\��j�ۇ�G=XL��B���7_��7�|m�U|� M��c�U��f�nnT���$g�(��qtre�FZ��{>j��l����B(�iP<ddKD�%-D�lQ��|�W ̀�s,�	��.�T�
(����Y�2Z�S�ԩ`��Yg�~�I��,K^�A���9Q~-Y��a.
E�+e���&u�Y���	
��|�Ε.��q)UVdd� �7K�Yz��Y� s�eɞ��J*(�d����`�̶ �#x�!�a(L����������_��h��K�b��.B��5�^�|�۞�ّ��\y�������� a��l8��-?uoan�Lc�g�X7��5��rΐ��и��Q�@��X8�\��Ɋ܄���ǲ�W�L��{o��,ـ�;K{�X}s��}f�X�ޤ3�>�rФ�8��K2�ªIZ����Oy��^p/��[q��#g�p�3��-L0�i;�=�q�Ǝ��b��G��<�o�1 y���C?9��gÍ��QxG��9d���7�x�af7Js�w���|��g�R�S�a��f��g<�Ã���48}2��j�n��#��~��z�3�1�V�5�w8	cg4���Ӟ-M7�����k�̣�D�y�y/�m��0���e񠰄S�����`ˏ��q��}��8���/�����2�-_J���O�<������Ů�ny#Ȗu�2�w��:�/��L��z�/��.���8� n˖_�\�L�.U8�.8Xs%Ԏ�Γ;Q��+�$]��` ����k��'~��n�$n֕���J���4!���ؕk!Ҥ�֧�'��\�˛x�P��v�&P8��O�\3@���~]��l�I����.iI)����-M\ԣԙ�hQ���[m��s��37�n(�
yu�I6þ��=ߠ������KuP6��Rs�����@v`���$�e��W�y�Dq�;�>jl�/�Dw�Ft�a�q�Y�O��qO��z�ǖ�je������[0�MwM,��[#�e���['��Q���0��1�ҴȮrH�1�;l\�p4�t�a�:���ʡj����k-�0��]�>�Ip��'�3��{��#QB62޼��%8�.��CA:�;i��:,�a�/��8�>L�X�2s��u�y�ۑ������x�)�<��^?k`Gs��hGL�HM� p�-h����
ؠ�a�6(��ȭBT�<���0�8+]C��%I�����4�:�i�^{W)�����D��y����L#�h�5}����'x�Z­E���������R-/�<���B����T8�.sx��ߚK����i-pR����-;(��Te��f��Է'l���O��k;�D��P�,G����t	�"�#gI�����J�����=>���g�p��'��R�?�3s�@���G^�����ΔZXn�:޹�����M�ֳ�� ���i|˿�!x�7�3^�#Whݫ�"��^��S�Z�m�%�⊜��4L� 3\,����0�PC���r�1�愶��_"ۙ���l�
������5�O�i;ޖ!��a�ď�S/�S��Wq����@0r�Ѳo����e��3�,�x�������ǁc�ɫqd��������g���~y]~�@%I�cY`L'�2^�ʿg}�E|���'��K���4\�1������w����������_Sv��=�0�'�୶?��/�����o�]�o?猣|��Rl1�v��3�98\EęU�v� ��44�Pzd���vKq~�zs@�A�Ȍ�[�Y��O�o�4ʇ�g$�0���8#��z�ᅤ*��T�b��������H��*`'i�ZI���w/|����[w��y�ʻ��K�^#=8��w���o8���-�����Ke���U��@f
�K��_��z�x�(�N\yz�C�2�񞉍w9s�����Vl�,�_5|����<d���r�I��fReX�~4��?�hFj�e.��5�r��K~��(yE; C~&?i��a���f �uav��i^�+n��l�0�' �;��k�FU����y`������Q:};S�L�]kՒ�V��+�@]b�h�9�sse�R������l輗);A� a�(�*�a�"�r�/�ۨ�a�!��_*�p�?��<��0!d�C��R�Fؿ��ϱ���ͧ��A�U][��/��0:�w�{P!���)��[��ۉ�N��N�.t�2���|ү0�F�)�����.��M�*2��
�
�Y�ܩt�n�2�����"dy�|rw���1���J��*I�W𖡛t�o8�����+G�t��1x�|q�(�_U����P çDXL.hd:5�Z�*_�t
�}�y6�~��(<��'\�?d���~����:��`����;�l,��T���S��|�����5�6��	G�ؑy`�#tF�����ӟ����?��v�9N;�z7�p�&E�G�]�+��u��?*Qg����f�l�w�q�"u��8+��m�&>>��� �vb��1�]�Ҷ�\���9Q�{��-Nm�c�E�#�ޓn���[�	�k�ӝX�#�M��g�����ĭ��Nb���5�ܥM:5�&��'�|����|:�u�����&<��ƙ�3���3 ��'x��S��r-gp�4�T\4�./}�Zݴ��/ܑ/e��Lp�)�8h���6���}|��sfP,[�>����1��z��߂|��Y	�/�١���t�2���/�^0����s�����3�q0��w��>��+d�r2 w�P�9[�1�,��:u���W�U7�� ��kG�����啳����~d��	P�^�n.�[7e'�	u&�x�����y\H� �G��� ��Ҫl$�֑��f;?�1�+�������)��FX��3ڨ��=.ľ�R���K����c�̚�l_�p���[1��\s�"��3�2�ň֖W䑖w�|NИ|�A�R���6HN9pR�2���7�����l�� ����Wu��T�h^a���O* طR�a�ѓ�)-�b}����$����7���岼K���5�0#|����{�&p*Rb\[5�C;�4:):G�׷�Φ�7l��kN�� ��\d�:��-C"<4Ĝ6N9�ᣒV�M����1\&�`
[k:밾�H���<`25���;�u hNgzd��Nx�k_pF����k������?�f�__p�}2̄3R��	�=KJB��9 ��O�VFZ�F�ޙ�J�/��hT<�0:�|��e�$DAW� |hYQb�S����
�#(�sP��޽t
�(`�h#HZb�Q���l���(�;"�6�����![��H�Gy��@4}������/B�c���92D�$W. �`c�s��n���Iy�w�	�8�1!W���`R:#����w�}�y��)�}��+��rz����C��+u�Q�ԫ�B;�-�Q��ڱh�m6_<z��O��������O0Ȏ6���l������i��2Ҵ�>����1?�3;��[�2�<l�ʳ~ɰNxH�ү��O�:!^���_���N;��NHO���/3_�7bԛ��<7�Ɨ'��ي��(.i�"�#�ڷ޳��l|K;�.p��"���5�K�����ӑ��.�$Tf�&Ot�`ؤθ�rD����4����2�\�����|n�i�I�h�r�?���!��^�~��ҍ������<�7�s�g�ɧ�8��<�*cV��V����ن�o�]�2�e�C�[����{����z �kF�6��,��8�����d���s>s�`����i��5�Ϋ}�оU�a�=.��<�9sO&�}i����3(���>�RxD���JD��!��*�Md�L=�*����G���Su��W�ؾ��>*\"�~�B���1��Odi�|��\d��Bi�-�C91�[�zp���	PU��J�8R
�#�P�>j�Z�Cv�۱�*\i�������|��>Yٿ��Q�ٻ��F�a��Ҁ>:$T^��8m.}*���B�s����qT�L�m1�|����mI//0���dF;��|!Z��A�BO�D�|�7x�/	���qB.���L����=Oe�ϫM5�}��+'��F�)�1��xv�$y���F�å%a�'ܣ_q�Kc���eti[i����*@�.:2�K!�z�frXv��/�ݷ8�C�}����Hh��ک�s���`H�3B
�HW0INʟ©��X
q��ȿUD8�8��u��mF��&7�ޙ�F����i��';�K?���/ן}�����r�[����7X��r$��Pj;(;�Lg��E�A��[$%,w�3�^H+��oc��3�*�v��$L�_1�F��g��0�&w��ǥߨ��X�g= X^��qϬ�8��8��hgj���f;z�(b�)0��T���3��2�Rw�Q����%�tǔ������*���\J����N:�0F0ʎu� �}�;�%]X�6,a���������\6y���[�6�9��ԓ�ƀԅo�o�*��5��ю��7�UV�������-f��<S�h�3_~�%{g>���UTm��=F��ܵ�&#)7�D��>YL��x��g_.G�����G�S\��-^�p�b����k\���0���X)~pٱ-�y�>P�p�g��Rr�g ��J�Y(h�7��$�؏7�&^�� ��3��`�a\�h�F�ǈ0�񦟻a��U��e}�+�LP���a����s?�M^\q|3������4�l�c��G8���9�4]�<uuɇ�MGО~�7��y�/|�0?�q��?�s��g�tIv��~ÞJ����r�FE��z!�8��x����%HZn�	���}q � Ɓ��Y�W���7Zt�o/2x�S4��Y>c�F��H��D},-������[F8(�ʼ8+�y�$y���N����� ��8>�O;�'EE7�����/Y�<�zW?���k��oX��O�ÉYw	�z�i�CS�/�����r"�chrw�g;zG��$��{��7�^9�EF+N��6q��1���6�����a�L���q�=2���E���G���9���94�-�DD��+��Q� �چ�=ˑ��k��E��Փ��j�ҹ��xX�#�\ew��뽼mH��Dˍ�YAF5��7�Wf`s��^P�Od4g�� �΄mD�N���w1��;/
Z�0h/Ca�uF�«�u�~>½y� STP>����1�سu�A��->E*H�<�Ԣ��sx��%/'TΐA20{�8��#����}�zgH�����H��)c+'iҁ�lc����c�byzv����������?��cv��-�)ʱt��)ShȀ�茑�P;����#�ħa�}�}�4�x�x�6�o��48ff�}.6����nd|w�lR�i�*27��<O'�{)����Ox���*	�s��ө�5a�$)���uw���պ��7p:������3G�Ov�����y�t�y�.���л��v�(�7��d�b�t��-��z��y�R����x���9:��8d��#IN=��{���)�9�;�lʃo_e �߻w���t =������0����ٳ̾��@������h]{�ڍ�X%�,�RpI��^Gb+r@�wx�ՙ�:�dh[>��v�]x�+˰����NÙXgyb�kx�� p�4��*>�gh W;��-,GW�}HrA�Zk���Ӹ���N.�v�	/�����Y�#������8����]��+�Ԋ3���C�8����r�~y!�l[��oZ�錷����s�=0װ��
����o�L:��
O��N>�
;^��û�C��&�4�H��ozq���La��wJ�����%�YJW��<������,5=g�c�s�2+m�io0Ag9���_�/�z��`��=�ΐ�F)�a��B�׿�������'��>���}�o�_Ő�A�A�1��.�A�T�5Z�I���g.gy\��qmƶ��C�Wu��9��Ph��:f�t@h��"�P��W�����a�V�-w�hoZ7r*0��:����iSn\�:g@����v�,��óS�8����yxtM�����'2�w���m:�S���|�m�i#�w*~P����O��E|�����݇�w�ˑlG�u�r)���ş���Cgì��f�y|�	q�`��GVm�4+�|��a�k��S����Zd�l�4���}� ��%h�?a��#��ˏ�Ґ����wEn���LҺ�%{�G���vx� {� ��e���� ��C�9�N�9����ێ����DM�[x�����,¬򶑪d�$B���)���H�!kW�D�U�0�p
����d��ă���3�;=�����շ����u�)���F2�C![4�Wy	ߎ�ƪ��v@�x N�m�ĦR�<7��C7r�t�B�Ғ���2�lҚ��Q����A�a�zъV9Q���U���?�{G��u*����zF�"E�(߭���|�s`	Oځ����x2s%�K�M��o��0Gi^*y�9;�a�'��t`��-o��n�%-��L/�Qx~�+>�QD=|��a��/
�oi���eq�����8r=>�İ�ᰊ��c��@.m��!tz��)��y}� �ۢ�����4�������S��b������a=��63vʧ�[�X-x�W��)Ox(׀�R���_��s9*ƪ�3��3Di�#w��V`;��=��uF��Q�Lf��(������Y
�Bˊ�H��C���i�(W��IyQF�O���/��[��#�cb"��`��Qa|-�p�4�n��8˘�v��O��)�W�xn���I��ؿ�'<��I�Wa�@4��p��ׯa��qѓ� �y�������?�~ʔQ0�4�˪�Nl�I��y:v�gT��4:���o��ټ|y�y��S��ki���"�Q�k���Z�"��%��hп�46���C�3~��"F�	��3�QvL���ċ�/6�h_�0�������bI�'m�r�7u�}��'ԥTg���Ȓ�'g�Q:R;Ju�Ƹ��1����=;�P���[�,��9�Z����7�?e��:�3����g~��5���2��s6�ιG>$~;��e��K�����MG����� %ϕ3eU?|g��@�K8�^�M����[�6���y�N�EHN}?����]Q[tWȢrg!�[��<X�X^�y��p]��Y_����\;���� ��7���#��]M�8k��[�R%� ��8�!�| �Ě����럹�W@�-p?�D"���5�.�P-��u��-6���X�("�k� Cm�G;4����"*$�n�T �L:�\��{*?	�8GV�B�]���1��l��'M6>��@����C�!Brz�*yc�s�n5��yXzw`�N)�X��4�����F�HBN���c��l|��jX�o��ܿppl#ng唹o��x�7�o٠�e@H���*��^W��=<��1�2�+O56\;wD�l#bKðq�zx�=���kDA+�Dd���Q��:ة�i��\�W=�E^M�R���v(e;Rt�5��Q�̌YV�H��O�`��r`�p������=s*L��}%��,7��e��%�U��%�J�`
��+>?�+�G���,a�᭯�{�h�W��;�a���/�剗���9����<c��o��[�݌//i(E7��f)�g;`�(���P[VI�"�H1\g�i0Pԉ�F���Ef�!pug
�_5��ޞF�o�T����ٍ��wFg��e�&B�Lqb��6eǩt�QQ�.�w)�ـN�_i޵ogx�&l�U@�נ���gg(\=�vf�6-l�5�H-�*TO��u���^e�x�R��bh�)���7lw�Q\��s���!��.�tyJE��a\ۉx�x��F�gX9�����|�-j x�v�E�LS%ݎSx�=N�:y�Rϸy����z�_��MX��*��wp#^ܤG���3��lxp�o�9�9�]Y�'�?��!uo�0�V>*�ֽ"�~�nlߝEG���Pգ`�U��:XDV��_4t<�ӽY����:z�^��<t��$KV�r���<�Q~)��m��s_/��Y#C�\P�o1\��J�{���*ɑ��z��;��cy�U�	�=����+u�����3+��[eJg^�@��ʣ��|�N�q=�d��:�!T�0�|�~=�wIA�bջY$1o�����߾1�<�<t�W*1>R�J �ge�S.�4����-��Y�l�.��KW�H�D���)����5�a��.�"-R �p��i�䷍Yu�O0��	��^�N�*T�[H` W�������K9�w�i\ ��g@��4�oB�u&>�	<B	�K̘6*&���� �CS�-D^�E�Ë�ٛ*?���1&��*G��T��	�
I�b�)�*L�f����xiV���I'�<�H��Ί�8+�r�K�����/iMO�TS*�
ѲFP};���s6f��<��Fs�ޠ�^(�4fᙗ��6�T��aO��PS�<;r��8y`@���QB"O^QV92�(�*)R*Y���X5�F�T�!V&�|;+��2�@[G��"���bN��]!��)��I<D1аT�1�ds4-qȀ��s�s�	�+�S4�o(1�0015I�<a߀�[�pT:�i|ppui�cOJ3_t�X1�Xj����B����6y���/$a�Dv��<��o%B��FÉq��0`D���umr
�;K2^��Ӿdi���U��e7��؉��8�fK=�C��K�����0��K8�i�:��ҐK�`Q�& ff0Q�~�E#P���;��s_���5Q�N�q@[
K�ʮ�%�5N��6Ki��t0�tt�9�.:��N8�+���[����v��,��|>ﻌ����!%Q��	�� �����	O{NZW궕<�:{8��|��(C\w`�c��+c�4��+��<�*#���j�jͥM�4�e({�=Ï�;�� >Mt�m��>��"��Y'���e&���0�5t���<.Uwc5KL������@Z�ۑ�Q��s���'��W�	�hQ~�� 3��A䠙=X���K��o�/�"q���7ܥ9�B�.s�[$���̜d�3s |b?��Vg�a��;a�ڣ�4��Š�_Tx�ЁAp5���	�R�Jf��笘%+�i/�6e�.5ƼZ7ց8��3$�@`���}P���S�WW�LҎ��/0��5�r���@U�<���mg�����#�\�MK'u�x��ҭB�&˦�#�����}�M�ʀ���c����ҟ�o��~eb��L�:ɯaJZ	�y�� qw�L AP�\�Gn|��Pg~�}�7%�Sl��+ρg� ��т�ʛ�,'�%��_:)���tX����`'b�t���s �Md��Θ�W���0Tpn] P�dC�P�[�@�t	�@��T�~�����I a��ݳ����5<Nf+��s�'F`�9�e�6�?��B�����;�R�|�U��:#�����b�b,�hC�	%ܺAÀ �N�9���V:��5o!> ���G�W!�`Bg�P6Y�#��s�����"��SH��!�k�̼1�r�C�D��ƈ����de�A&OT�c�ո���3y�'�2���o:+��u����5<��G0��(,�G�-�廜t@'(�c�pp��NDe�[w};��@yr���%�tT@���rˑ
��4|d�Qݽ��!y�]Q�B%r�U�E�t�����P����4NF�4�Q�(�S�?����,E�z}����!
^�@P�H�-I�0P�<�B�rM�".�x���� @�	']�#�4��sv�h0qp&F��6j�c�v��3�˴���w�N�{�
a��,��R�޺���0���1a](o*��x�������;� ��rk�	�|�>���>a��/��'e�fk|�������ɫ��򕳈�-�<lÛ��N��Ik��0�#��/�ݺ��x۫��^ۑ�<�[�C�L�����o�1�B�_u�&
.�_3I⚍��5�p�������4�r�NI��p��j{�>� )��(�3��j����v�4ִ5i���ap��wpu����{�Q�>�ޫ̤��o=� �d����I�aٿ��=[�15b��[�5��9�]'������G_$<F�,��\a@0Z��ZW���X�����cg�䙙���~ ��%��Hg�#+�vF�ȆsTw���<�HR�8�-�[̾�v=�l���t�����K��P�·mN�8����@
j�}��;o�sA����%�h��� �����Gt��8y-��xt�Ç�%N/�� �U��D��:����ma�g�/��Ɖϔ���7 I�w+8���7�4�O��@<W���	�w`ʅ�ZW��e�EQBn&����s� �Y�K�>ԂW�!����XA+�:!.���;�
�k�h�D���sx[2�<\��o�;���	FvG@c�f���?>A�8��A��6��n��y�/>����P�O!v��50$lH��ˌ$}M6�
�x���<I7� !3W���UZ )Y���H�m��״�E�?�PZ�����G#��5��e��� !��WA�'ql��όR_��k���]�I/͞2o3����/�gxKzZ&��7:ʃ �C!����F<����Y8�*O����o�I��+)�l����m.E�9�G�\z�ꙣ�c��n:MFe*#��/p��|*y;5h����|�A��;%	8:��l=8���y{��ǀO��N�@�K�����E��v��w�u;�}��CI:���V�کa����>e�|�n��u�/����_ͧ"���^�&&RUw��NCX���G��x���㌜H���Ȅ�~;��2$��_�����5����������&�����0�|� Q�LǷ�g:ydϳI�[��j�����[�b�<\|����+nI�Ϥ�\���C��N�C�<�#�D���� w�n�)^���\�-�����(�LC��j�F}�S���|FX��Ի��l�A4X(�g��w�=\g)�0�33斏L�(�S�5����=�Xk�;e��Ç��gݪ�k��E{GO9u�>�O���>�?տ7^w�����%=f$�s���ͧ����_a��R�y�)xY/��V��ꫡ��,�����쬞��u���)�W�bH�C��,�`�1��1�"S�.=�a��֠oH�Z�Ϸ��r�x�҃F�����ejx���K�왳���4��DXD{'����Ϻ�^���1{6O��i֏fE��	����K\S��/UNx[RӪ?K�m�
���{�ĳ�$�1�=��$��T�� RM�����HR+9�S��1]"V�ᠥ�]"�Ʒ��s�|�nf�&2�����t�"��(�@��*y�œa]~�c�1<R�@q�+��4���}�3,!�Ҋ�R��o��W���!�XM������°+�������l%�+��#������?�ǿ�|��G��qF��lM'����:9g��pf��su�w(ˆ��jy�����XV� �D���q�f5^�uv(K��gC�	�ӎ��r3��M�Qp��j�]~VԠ���o7�s#'x���UvPv�4�=�j�����@;�+���XLVD��)3��"��Kן�]r$	~�A����Q��L�G\�������R93�]ݬ@������ěY%*2�=�涹����Gt�b^�~};7;��_��s0����O����^���h��fj]䘪'c�����;9_���p�;�ۚy�����}y�!7t��̋�Ąfz̸鄻��X�@��u?[Q3����O*��k�ʬ���8H�xрm1�3��=�md�]�0��܋r�1���_���ơ�7��G�#剦5��(�H�i�Y�vv
ȁ�uLg�O�!�.���J�V�Gǎn��pT����'�3@/�:����S��9:��+��8s�Pe��A�/����ٳ�m��O[��^p��|�{�����Y�N:]+w���=���pp�>k,+�<��֮t�Ҝ����G�C��x��8��r�z��g`jw��p��f�����\^���g�I_����f����7m���'JL�����d���e�j��G��D����8*7z��No	�i��VN5�7�GN±u���m����i�g�]iͧ}�f=-�B����S�����=k�A��E�p���F��o
��~��ɘ���}�S6���%��q��{9����q9��"����-�`g~9��y+/m'�J~��z#��G�t��qr�p��+'�snK=���x^R��9x�{��ڵ��k������������us�+���5{�(�ƨ��+�*�K$�WYf�a�������Uh_/��=N�V���%�2~�	�}�cz�Q���d�7hR���uO�9�t��g<�~�������O 	h���`ͺ��I�x^��4Y���UýBO���>9�	�,����L���-.���)&�c��x��2D�Po�Ǩ$�:]
1��)3�(XؒΗS��Q�Et�s,�Cx�̹�Xp�_�\�~�z�{��o�W��B㔬����X��z竿�cz�����~��&r��{5�:Q�W��s�=i�f�z�;�<�: �U�}��4��zIhq����°'�A{-�0S�۷7{�2k���|�(	�'5k���䭝��̐�Fگ���sHyu��ؤ��I�_�R
U9�Tg������:O��K��b艠�$/cX#5�������sDQӈ8ZBn��YE�N����h�?�dMT31��W���m��駟������{��oQ~�hgP��Hl��:�}�����C��)�+Q��=�y�5��+u��1�ŠƷ��ּq�Ffь&<��;�pJsvY��k�����4r��>��td)G9���d:0��R�y�� #  @ IDAT	'z�I��砄�����J���\���>9ӇՉuH9�$�S��&@��5�4�H�X8ԡ�q�k�<�Ì�uT��zv�ެ�Y8:'Q�u�N8:��o�4��.���`�PX�J��<Ҏ�Ó�`�}8`Y�V��|�/\|�:�.{�w��g���n���p��.y��e�F����W��̷O���\��}�ZK�^�ܓ�Om5��O���%�P�gM�H����]�xh���}������"2���U�9\�)�%�&��a�/gdk9�^1�;��x���w�74x�z�^kͳ� ���2CƱa��,�c�0��<��vr.~zh�[���^����6o�^��7�E��g����d�V�*=��^�^���Eo�7��G��^ۮ�vɉA_���@O�[��O/�ة�R/��t�ʙ�mJ״�%E��J�Q��^g�Ǡ��]?5X_z���ޅ�y8��\�����Q�7�\�fk������٦@� ����to����_���|~��G�S}ݖ�`N?5y�]O�:��I<jv7��ΦP��yv��hp�;�샻���s�;�;���gz���cѬh\�YOδ�50�PR0����N�����`-��I����{�ŋI`@C$Ϣ{�Q������+�O���n繎_�	�7�=M��tU�?aDs���O�s��ѿ>}��jL7Owq߸s/ƶGO;�����rhz� S��&��|�(m�1]�i�C6ȳMC��X��wx1#ʘ��]0��ٯeBo�v��N�sdr�tb�S��6�T~:����ߒ@I:��W���";��ȁJ�ð��3gޯ�zP�����5�rL�%:�rd��mR>�n��@��>ݣ��2���٨N����)�5�����\K�9�댈'"�:�ւ�����%�Q|�!C�C��� ���`3h���cD�W�5Nq��<h��zu�h���%�]�nݛ�0-]�D�8�u[=�:�P[y��������>���c�~N�������_W���ȯ�8�ވ�A���:"\o;`�G��2e�~x֩lf#^:'Fw�"Yr���X�QgxY��	��ˠb���!�T��CS��z�+��i�-�t��Ћw�}:p8�0�'�q|��m܏�.�=?���q�o�����f�g�����Y%�����3hﹼC���c��p����ﵫ���$/���hv@d�F��q����.����`u�q��[��kk�x!j�djj"�!2��+����� �I�N@��C�[�BM�8��8:�'-,�mK;��e��������,�xp�V9��W��b�Z&���8?+��^=�g]�}x��x���M�����Qk�o4��n~س��K��7sَx�_�h�[�hi;k����h��8[���m�Z�20R�����%�R��]��� ��C&x��h�S�{�i?�Y�r���ɟ#�sن㵶����q����Oy+���e��<ܞw�'��\9s7o����[�Ӷ;�������5�v�5�����"p�ݝ6Ay��K�ηs�iR�c���EBBݵ�q��G����"wh��n����0g?�W'��8m��vF�>8�c���9e�_ ��q���p&���T��9Ø�iF����{6�P,�@
/p�ո.�m�&ғ�U#q2�o�a��^��2x�1��Y��pJ�i����br���0Ω�����g��	�S��[P�\%�<K�6Z��_~zz���������d['SCx�V?=y��' S����ߔ���>�:X���&��Y�ݛ�;]����@E[c�:7����m!P_�;�el헲LN�>ǚ�q68=�+J�?���zB�{lv�{C2r:kS�1]��|���t�W��r�*�<]�^���|�L����6�Y�-�$o6�7ы~�áF�:�th�0�<�e7�G�鍨K�6��}���f�L�	�����񺷷��w�u+-@x�F��::1i!S)�|���3|Y}F�����B������[9�C�z���x�x���5�ț�a2Y�=�R���n+X�c���໏�p%_�8��E3����1M���}D���)��d�Y�i�~�����"������%��}#��2�U�=g6��!m�B|\�KE����ш���D$�ع�o�����T���;�����1�oih<�ɇ��N�v32X��k��gx��۴���iXOy�����m�=��u�+p���(+���W�h����r-�m�Wnm�gce����.u���%����;u��i�w��-��t�;��q�0��b�K�r�g9Em�~<���-A6�n<j)��^������^�k��Z2q��0v�V0t���൛/g�糖/<o��E���y�,(�>��^1GM�o6����_���ӟ�����P���7�������-:gWf�6v�mZ����D��ٌ���� �c����r����T�A�U���6pFxx���#z��eN��ͮ=�lQ)��V���Aqm��A����z��������|�{��8Qn��RM/
�we�_ρ��4rӱ�1����s�Q��}������2zؖ4�^����hM���<�������M�r~��L[���SV��iN=��k���H��mm)@�����NJ�uW�R���y�j�����^r�‛?��ӡ��8�u}�L%!'cDqh�	OXc��k���~'�S���=0W��0[D6�
\�93���$���sfj	҆���]G�r`�2�@���?�=�3I�[�+�:��A�sz��Q��!n|Y���o�}|��"}�z��I���I��w%�
,z���mS�3^�����F�w���V��ܹ}sxv�����x#���I1v���/��E�P��ְ޿�Ti�в�6��MJ���>��\�D0�ã'�_�/���z.V�Ck�6��-�~?_D�A�rp����ZSq����D�ZU#����ȡh�Fp?���h�� Xt��O�,��HҮط�[���h��duWo�Z�Y���;��+
�^�8��� �aG��U�:?#oN�Q��F��O�F�C?����8C�t͵�x�4ǻ}�g�|p������a4��w�뻐��A���na�/J���0�qVM�k�dDI�ֻ�5����q�
�X�{����c�ǘ'��6�F����2��_���C���֚�T8^>Os�߀͈|���DZ<�]�cx��я��"��E�����9@�L��N�
�n������E�x;�e�m�s�qp��L�8�)/<w�8�����haz�q��:Vl��2Ҏ�`k[�z`��<���'�ql/��`��{e\�(�Q~}W���Յ�Kt��pr�ə��w�K*���G���l��k����b�t:���L��p�E�M�Ygt.����;u�:���x�+��	��o��C�К�V�~���{��������e�� �C��P޽{�z��۾m�ܠ�ru���fkmW�1�{�U��~x��o&^�~��O������k1�����=뛭,�x>��Mī>0��xr'}��"a>"~�\�����j60�cKk����w��O�]��o|�;���͌Fm�#e�X2%c}Ë��x3~;�R���p.}t�Z8j+��&�+���8��Ëc*��ܻw��� 8��gv��y����Z�����kڧ��mC��ק�}jH�$A��ágE�t�����1Q�IGY���%~�{�p%/(tÿmW�=~'�n!:��G^u͑2T�[����-�N�{T�k%x�({�~%(U4��^n~EL���l�f�����Op}&m�����YD����uHu�:�1�1`���e��ǁ��A�`�2���IG����Ne�ï�C\�N��w8^rM=tx��z%���D��Y��N��M��L�֝��S�����M;޿�k���5d����!�)/v�@������7��Fo
i�y��H���,���;��ۗ�[D���sR�M6�2��3 9E�3fuz9[��0�`r���x��Wƪ��H^8X)*��Ƽ���ȷ��;�,`͎vd�u�3E��s�j���e`&U��1�l�Ҍ�x!a�����"�#��ѴA��Ԁ�<�'���l�������>}��Ftތ�F��;����W�Y������#��/�g����Ah�D�1�j�G�p�4�6Yv�(c���3��!�]w�(�]��ſ�����{F4�|��>��G�M���RA����KDBc����	S�ciZ�L���V��&׋E�=��ⷎ���k:��8��nb���������z�Kb\���F�Ө�'y��%0ޱ���S�h�k4��(��@vN</����f�3j_�$�	W��"�X�j�e����Y��9�S7XSO���q���>җ��|�!�8�=ל �ڀ)�c�ڑ������������s��[t�m��ș~S<+�AO��zq_Q�%�S6�8��|������-aԭ��}{���;6����ճ��5iK�]�o�d�؅'��e����b�Ѫ�À&��ahpڴ�g��s�����h�/9\��ZO%j�D�5��bs̼�(��h7����'-��1�w�BN�n*��U�rp^�I
��J�/��D*��8�K�ڭ�bW��E��g>�u��/��ڱ�rm�=�l��([�S�/v�F�-��ިL���{��E��N3#	&�v#Pb �!���0������-G���@�g�ӕf}nN��|��������OO����?�,��CS�߶�u�u��ϭ��T�1�
m�B7�<�����,����@P��v����u��#A���cq�����V� JC:ڎ���BG��x�����:��{���cJ��d�g����kmk��D�����I�~dj��+G��)1y��RJ�w��|�Ry#%yT���E/�:�W�����3/�ܥQ�)7(�<��Aُ���;)�tػ�M�)&m@"x���"���3��zL%r�P�\(�qΎHط?<�y�Y����Ӽ�R�k��V�jM���4�z�Y�l�Ҕf��<�%��������
Q?���FK��[�a��I/�b��Om���;O2�:���!�ۋ�QV�FX������c�˧�QW�e4t�I2����q��[��Y��y	/�U�i����j��8�FK�'�&ʴ�@ƈa>7:&*h���Q���~f�[��\�����x�c;<OH��kS,p��h�޵�7�[x}���p�&�pr9��X�����3���i #�x�ߨBt'G��02����_���G�>��^�u�SxuܿoD�h�����?�Y�{�b��(7�̈����A��s;��^��W=C�D}�����L��L9R:b��hxU^��q��X��s�4��B�QvG�{�|G�u�~��y�8�I�vt��|u-���+;��t��s0t�p�gh���D�Щ�8�{���=���}�>���G�~x�5<8A�o��k�`�vy ���l���q�z~\�w�k󿑵�|����-����HYp���,W�~Y�/K�<��-x��j���_�r"D"���V�A�_����ٜZ���x�Y�n�]6i���>6��3�M5�&:
����!��M�7��u��/�1/{��������q�H����x��n'�k\�D�9/N�6�f�v�5M~�I������YCz�H؋l��[�,��J��%��A��u�}���=$��dt���U�M[�ߝ{����<�>��{w8�7�B(���Ev�7��"��9��Y��U`�'1u�<;��Bgo_1��?�I�ɲo7���h_����w���<|�������i��D߉w�Π������v9\�~��;w�ލ���>]imܫ�"bW�"8^�g_Gg�k|�X���>�q�ȥ�M�k%Ѕ�yP�u��c ��O�`Vs��ca.�`��  ���x�]�#Û�S�"�?��:z68ԧ�`�q��9��GN��G�[0|�u0e�΋�䮚�aH�N�7�0��1g��+H�W)�|�)�W0Q��9�[(`:���^$Q�5xG��cpL�#��o����V�C8��y�}�Z���8��M4�x��^8�ZϫyP��RG�������wN��Fe�����O��D7n<�h�v���|t�xտ*����s"ne��ܽ6���������ӳQ^�x���ӻ}T�(� z�9Y��mB8�s7[�45i���+9R��(�\��۲:����|m�'b��zD9^p�� �xfd{��ae�f�ܻE��w����{-��M�vl�ի�r�^��I�F�9�����jp�e�w�Q��Fx��,U��9'9Q1!3H�C�pށ�j��巑�pֱ��9x�a�f����F����<&ݰ���3��Ǿ	���Qn�Nyݛ�x��ոFD����t�06���u83�(�&�j��v����M�E���C���H�~�%�DK+o��8�խ���r×x��jq���!�G�;��c�Tv��t��;��/{*�i]��I�<R���Fp�vh�r�0�ԩ�S����S��#�_x��upV�\9��t���P�qώ�o~'��=z�4�CX섴*���s�XT�/�����~��lK�}Ԡ���ߟ~��ÇF�Ϸ�������>6o�Ϳ�u�M}��ݣ�<�;w9S��)���3>E��Ýh�cd����&I��o�9tE��O�X;�;���Wٔ4�u\��x��������nQ�96j��'�n�j�#��u��4&��N�D3���Tr�"l7v-[P�ed0:�Sv��kE��gfI��6О����y48�xR���g�����V۽��h��8��!���t����ϗ�Q6D*ߧT�I�~8/4Xo��&g�Z��r@3�ɵ�[/
X2��ڞ�`W�n��An�w�[�co9�"�f�8`��#�7p�����O8����Y���C�?��=/��BH]N�%\��E��M��
� �eK�g}j�9��|�S@6��w�}��c�;g�2K.����EM�+����uX1�\9$�7c4�	F!����R�@4�7�*��p��ԅ��=!N�}������Ӌrn妆�W�<� e��{0��z�SN�Λ'��40��7FF�A�;9�8����DZ�\n(L��V��X�nm��:�+i�� X�/�>�i��A��:�{�Z��^.Ϟ>�{�����6<�����g�'?������a!��J���<}��5O��)��Q#ON��B�܈�y8��I!��ơ�'�(v��jF�2����3�I8Zg��5��! ��O�Xe����n�x����zS�.�}���7������Ek���������5T�t#C��G�����վ\�z+�n{~1�Z�x��� 8�K2Y��3l�A>�m�������}7���K���~m����?�K��ӿ�ͯN?��'�2�h���:��_=�F���o6�-��o�]cő�9�^{!#ʈ�d���x���N�Z�y�}�d��S�N��0J�r>~Qqt�ov�/��F��t�uD�ۧ���h/�96�@b:��pZ8�o��ę��g�fӏ��hO[�:g�?�?��-؁'��WݦNGǻF�4y������+��~���K�G9p<�<��w���O>ц�au,wʷ7�����|�v���Ӆ���K�8����u��e���Nx���;�|�Iѯ_�~��_�>��:ZQ��7��Sf�O9\)��Ͽ<���������?����ʃ�/��ر)��"[��ܨXHu�@vD��y��[j@�ŢC^�)���e���!���ׯ��gk�C����4\ip)J�ێ'o�/��;9�m�Q4�u��/�ch��Y�b�γY����Ho�81wr�n�i}do$�hZѨ���7ߞ~���/σ���F��"K��C��]C���iR�(��ė����wf�fPO�{�goL���J`9WE&��ޚd;������K���O6D��������m�a�缨P���E/�c;i��񊜏(��*a��� y)��gBv���}+/�@c�4v��>v�'	Φ�w��@���,�e��{*�YOϰ�ݫ�1�$�[�$:ҡ��y��\��w�^�m�/��.�~:<*S�9�����C��w���\(T�*�,^��&��gNA v���9�϶�l4 >��ￅ���;� y<���.��]N�#��}��!�?C� ���s`Ĝ�w�MK3Gm6��k�q��Dg@Дb����W�D��ye:���ڽN���a[�����G�<��&*�l�Wi?��}��楾����~v���<}��_������O�mV�RC|^���szҜ'�?���F�"i��͂�(����h���f<N�T���U膳<�L=_��z2�2<^g�(-���L�D�!�Ҩ0��k1'�"��~��Ӌ^����������sLS{1<�ݟ��M�l��{���������G����J�MM�/�-d��\��r�� Q�s#����v˾�|�tI�K�c�����9b��X��>�#`�2�[�j�B��cGy�/�u4�Q���g��1�i�'�B��+3����Y��|�x3��&W����������/E@Eqk<�p������D�X�e�#kDnT��D��^��D�B��T����*7�	�kx��#v8e�8������u�H:x����G=e�X�L�\WV��q<p_�Ҳ�I���S��s��x��1��;_��W^>�p�%iS)׹������-Q�S�Q�-ѝs$-���>Lo����1j�\��t1��,�*� r�{vV;e��ta���:�ɒKw�s~��ʊ#�ʺ�2��p�5r������C�>�����:���! Y�sUÜV�M�GY����E�܋���},VT��y!થ&��ԾiTӱ�0Ѭpy�MF{�o}�ǋ�|r��H�0�j��`��]��/�����0���8$��o��ȕ�?9���Aof��`/�+Q��g�]Qj��~q�����Ot�WOvp�$+�8�k#�� ���Dp<,����uO��<=�W98��z���� ���Q*Pt�8��,X|�����o%����9�0���Z�O��q�)�Ӣ��˜��lz�r���a^|�'d�u8���ޢ��j^��ţa����J�$�������_WS��N5�s^ÄE�r�� ��[��-ܮ�֨�aZm�r�N�F��3�M�PfJ�##��,۔�����C�pxz�|.(<�E����M�52��n���k��3b���7N~x����T_��j#�[��|�R�� �*�`ِw|��|F`�+�a �� �����#�b���8y;o�X32(a�����{Fad<a�]��p��x�!�2D[#��ԕF�>� ޸������?6��h�S��>e��l�0��Ŏl S�PÏp�̎�2F�ɗlb�����I,E�{�c�|Ft�'�����|�t��5%�Ua�?��铏>8}��G� ���EΈ;:�aC�W���m��\/=��0lsF�Q,\�c�.�]L'0�&��u6�¨�a�N:'i���Η��]�MW�xNǁ�_����Ct����!/X'�E-�/�a7b�|�޶t�.�^W.�t���8�-B�<�8�(����#��t�������U^��\��^�M:��U��������s0'l�r���CY������s�x)8�����j89��e��%k��)Rá���?�e��Z��~SQM�U�(�:��:�ױ'���u���i�@(%��P|��Ac��-�{.De�0Q=���q>�[e�k���hSaE�p���i�`�6.�uo��7�Y��z�k|b����9{k=�n��椇���
k�øt��e�B���X�8m�R��T[U���㬭[��AӺ7s\mS��_��}�7��CW}ǧ~,�nV���Qn��<;x�pя��t�Ν;����^�N��|]�ت�w����M��>�@�'jf�F�=�q�������.�P���� G�8=�Z��������*�l̍���۱������x���g�i'�w{�t��q�F#�Vg��爓�wٚ��湿rk�G.�k��5�.�G򖶛��ޣ~��D?��a@�D
{a�{
�~'�g��3�,C���7(����9�$!8H�	d8e���~J�O�ʫ+�Y���(XP��2έ: Un���P�b���Յ��X�P48L�7
9w����@�:��	}��o�')����\��Z�3���m:i;Q�l킊̷ߺa�;u�Z'�[��<��]X�"b@ա�^����K�a��o�L�(T�2�|V-�F��vD*q��lZKq�t�7�l|����䠗��v�s�D���3J���R�Rc�ڭ��O>������cE��ѷ�%k����8y�N���z��8���E��ix'���tְ+�:1���I�4i(�o��ځ)Zہ��So}�}N�_���6�=�-�~����o�i�陌�:*��>�ރ��X!����Ӓa��=�Y�N�A�L썒�Ҟ��.�Κ��B��1��(�܅��G�o���E߬[\��Mg��a���Vݔc���K����#�q�n�0�2k� NgZƣ�Αz>y~��ׁ�������\���YT�sԥ,�ݥ^�,����q��G���j	�=�9�;�<��.�A�j�=i���w[g�<_�{[�`�5����V���=9������k��Eئ����������7�Mtw�����񑽃��%��j/װ	td��;�=��e[�K���%��6i�7����E�\Z%$����3�6z���4���yt;����2q�
�D��?v3�����ïlS�
�|�5�i fo�q�g�A�q��wӧ"���KsN�3��l��mS&�%C�`�gn:�9�g���R�p���t�m�'�>�cR&�H�9患�� w/T<ID��}�*�l`�o�:0/n������\���|�Z�i��w���å.Q�LJ��	���+���O��E�Ǧ�B��Q@r�}+dw�U�����o�5�k��78�kH	������	��3�}�������6�sSg�=���a섚�e���1����Ax�u�[�h-�}f���Q=߼K�=̆5��~�����oB�ԩ�L�q�6�/�_���Σs�	c�PhY�+�l����A/3�o�(��X��?u��	�Q�|2��Muǣ���xqLC��<�����?��Q� t|W.߉��N��\.f�덐.�ӱ�;5�w�N���8h���&��ِ,<vp_M����08:���},M��+�\�8Fc�5"�;�J#���0�]��3z�o���*�ń9E�2����MK�𽍤S����c\2F�]��h�!��F�/�P�nGj;���Ȳ�ŭ��땉��<�j��P�L���'�Տ�c��sj=����t^�5�uz�����[c߶���������u&�T�ut.��>:��&|~���1:�G��9Q��:�(�0}R�pr�,�_��� ��]y��.ã�y.<��8od�=�	�cI�F����}���i��%ʥK��,����*3Z��3��n�*�������9�s���y`��_��h9���{�M��t�۩��A�_�G>��9�����>�-��'����0��"W���:ԋ��w׎�����<vn�:���Y�uhx�4u��s9my^*��p62*"jO���;-�@��A����M=�����iޘ7�޹TH~���0���A�w���Y5.���9Rl�V&��*[0�X|�;8S1����]�OJ_@YK��Ǉc�?i���
٠���fV��y#z�����쫦�*�Y z���K+m����{�w��C�c��m^ή���=MK�W������d��M�-��#��N�p׻�Fd�.�fF��|NGjm��-{��@� l���{��#����Jo��t���i[m��}��3,�n�����䲲�o'���$|�ζ:�<!��N ����K��n9[%ǧ��5|�>�%)\��%��S��ʱ�"0z��e��X�-^W��(ѷY7e`�|�{�1�V�`��| ���Ըw4��BT�-(���	�2�WFI}�(�i��TD�0���h�~a�Z�~��X���W�n:)��GX" A���i>KS=2��>||\��0؁i�O{Kd���qpo����a0��< /,F D��U��rZ��>K4����|����O�0P�4Xj�N�#�:�e���0�+#���&�o:(A�؅�����6�<�sX����E�C�v%�	�O���_���~�f��� Vf�,Pmx��i�2'�uDi�r�݅5X���1Maǘ�t��zk�^f$��"��V�yֆS�?���fn9���'c!M/�s��W�&���4;6�Gk`H��o�oㄕ0��dɤ�&ʊ�����/O_���E29]_~���{f�4m�Q��8W]���ѥ�f���C���o8d�ۣ�i�2��D��xk�ƀ,�GǏ�_G�vg.�m��~�j��6D�W'���c��a
�N��n����o�M}��s��g;򊦩c"t�m�>����'>�)�n�@z{��;p>��s�w<?�����mSo%��������C��h�c�����K>'X�����s��9�oߴҩf�61x���H}oNx�����:�ySq-7y9'[�!�ܗ\�U�m� �a;��kk�����|��-D$rʮ�H�W�z=�8�Pں�ѿQ-�N����S��y��pljy�/^�X��7�D��V�P��5;�~S���L�+��aс\w���Y�A��<��]�i%�L��Л���f."��û�^��$��!=j�&�9:)d��q%|�qp�o�=%U{sFd�W��ľ"Q��7i��M�6�Y���DX��d$�}��E�>�XEy=W���r�wNZ @�\.�/�C��q4u����搧'��=�K:G!�(��9����T}��ck�$v�Qفu�p��8����a�68�.���M���ڛ�� ]��&��� �Ǖlݥ^k5�����.r(�3ߗ�Q�����׹
J��TP��>h?�'u4���73����i !2a�Y�����3�G� ���
��S��M�9�O���1_TdF5�	Wz 䨓��W�R�hFW�!f0�t�TF���%�q�ʳ��2��Czz��=�p��#�s� �:�����sW�B!=7-���ƙS1S*��� fѨ�M%���NI�/k&_��FILA����q���c�:8?��a$��I>����z����o���5���X���S��V/ظ6�WF0��Gu\5b�h�i�x	��E|뵷��\r�K��f�i:�`��� @]����gu�Ρ�YC���Ag�/^�v�ETs�;�\z���j��*IsM�17�N^��"���F�3{��b>l�Y��7ꚎU��6?���������UN�f!�,	��q���ap�a���V.=w��J�&�zv6��Ql
����'e��O�dؒ߱@|�z���޷��*�w�v�ڽ�જ�|�����8����{��;����������14�8�����;��׉/p<��|:��p�t�L���h�A��	�{�N0Ҏ�5�o���m^-��Nux�^m_���Gx���/������H�ܥ��þ�փ�Cw�^[,�8���Zyv3;s�����MAM����[�]���3���J�g�@��ۖ��Mo�$UE�xm�u�cYь]<�O�����'�{3�بu`�c���^ijt����"g#�u�3P+}���Qvh#C"`h���ǵ7�:`و"c�bK�̇�+m=��uD����>v�;��>����r��7j��/��	W8\ɑ\l�G����ѭ��t�|��Δ��ѡ��3:h�d
�t�SFp��=� ؋Cm���}���K"Ϲ��]��nFw�������T���Hᠤ�@���X���e�׷z���,�x���l������~s�JNث	|����/����̦���[2�����.��L_?�������� ��>�V=�Szl-8������;�Vjr*�;4�#�Hp
ݭ�J�5��i�գ�焵)g�򚇮U%7]�Վcso�17*w=�;���:FPex]c�p	��}�&��L�Ӣ�0	�z������I_7�f�����Q�2'�-�w�lz�C�<��b��l�:hMœ��`�� �>��������������Z~|A����k�l�w�oG��N��z+sV$��bS05(k
Bw����a���S3�$�i��C���)���oy�:+��b����>�u���?�|�	Ѭ΅�fnHpч'5�í�<�Y���
F��֚��zL�����j0j�3�#�s��i�()�q��#����iH��|D=�/�L�Z:�d�	����kG��7k/Jp�gS��)�ީ*��,�$C�[�]��s�尕6�P��wQ����p�Dg�'�:��@��u*'r�e���� ��:`tm����H�7tw��6y�W�Xc�88���	o�:���H��h�����Ҝ���q�]ε�~�k��g�s���z<[X��^/\�<4:���|���gp-c��3}��	���=� ��Z�/y����ߖ[}B�t�u`o�e��^ݵN�%�l�i
��6k��-^�\;HP�'lA��}��6��>������
����M�D�)W�F$�p�7�\����N��ÑR.��^[�}���gP�C�ӯ���Ի�T��e:�NN^L�3ч�-ҏ�ã돯�T�A�Ցs���ϋ r�f�٦z�I]0�qG��r��A�s�f`��צ�w���F=�M�����f���Z��hX���=8�n��� m �W��� ��<�\����m����`h���_i��8��|x��W�� ;���^��`tB�Q�m����/OO�$| %�}�����E���{�o�'�:���W����1XI|�Voɖ���ᩍ˛}�2[��?�!�L��yk����O4���Z�7%W�5m�)daq:ϱMH����Z|�g#�h�5(�n~�6�0gIBBY�9�F��3%�0W��z	�k�z"`�J�A��SBF35�='����;J�� c���˨�?̨3f3g��FE���� mp|�(�V��v�`�s��AcTh�R��B`x�ty�����rVH���Jt��@���N�w���s���N���4 M�n ��>�����p6�#t���7<5:�Է|��留�k��q�d���r;�m�C^�fկg���:sS�� ���40�*C�,ae���U ��������$�h��k<�!eSׄ�{�'���)\�bH���-Y��J����d(��sE6�afmG���Δ�%<�̛���8.E�шՏΉ��
�t��x��0@ә ��o��	���#��S5���0�{S���V�5�ъd��i�.�LA]�g�22��%Bى� $�螷��Dw����֡�+���?�x[fe �.v���ۇ�c�s�m��:���iҏ?�sʷ�N����~��/��ci���q��4��uh�(�i��a��m���?���(Ǝ�'�/�&Q�I[�&��HǤg����i�Ξ�
��-xhk��ت�~,{;6f0ˊ�`g�+����c���B�|��Z�hvI�Օ\��6�3e>O�8m��k��녃��9�-Uj�
�p��s��pt�������q�!�>�z6/<��Fo�f'�y/y�RoE�9P� }��Q~�E,>=��=9U���(*8�h
[<|��n�*��36|���(e��F�rӾ^�*b��x��~��f���r��<#s�]o��/ǖ����e��6��=�;v��8�fou9/�#���
9s9�6�Ӓ)�S[XH�&k��Ӌ68��y���W?��w�����?=��o��>����rz�ӓ�9P_V֚�l��z�p��� �i3�X�=��G��<��6t�*8f	vy��W
h���A�-G���Wsت�ٓ���2Kn"_ź:�}���[o�Ns�-��	{к���`����k�  @ IDAT
��ϊ���9h����[v�5�����;+]7�G;bA�6���D��28v�G���l�s�߽79S1{p]��b�qxN�_�(
��\`R�*W��~)jW��>�a��¦�g�@�1��Zpj�5`����A/	�3#��C�S�]���ְ�f^?vZ�6�atTX��8����H��Ո�P"a�c웃rI�߾>S��7�������rK�-A�$����%\��)�8��dv0噏k��HM��h�3r+#�t�ѝ�͹#a��Q�}a|��&����n�wS��CVg�!z�<�^��̌6'�"�tr~7��4�/���?t�M���I��˿-7�{F_z*g��oLg������tl+��=����d�2$����p��,Lv�`�#�u8`�*#r����v�P���3r	�|&�S'�>�^狞nG��(�@�"��)30J?�9"�:���}�@Ӂ�g?�:�g~u�����حS��|9p�:�����sx:�z��#�=;����q_�mզܣQ�`�w��tx����ۙ������u����w^��4y�p<u����O6M{����UN�CyyG�/=�ۥ��L9���I��UؿP��-�g9_�q���K^D��){���,?]oQ�0cG����t/��a�]�Q��>��2c?D�v��h���T���1���r�*|��S:rF�g=|��wxr��Y�[���x0���:mO�;6}�O�Ms��e�v�oM�ȃl��
L���n�x�!���>��E�2=���x4��E�|J�e6e���j�`3������8A@J�is�8'VT�!�@'$h������9`�N�w�����r��^�I����oo�[0��m-��˥��_�����0��U�q�k��%��ܲ_9��ӿ�t&��֞���_��OD�l;��8���3��wM��F�)Ho\.Rt9g���>��Le�x�G�3s#$ZHx��^�6��ˤ��32���)}O���e�5�Fi	�TM}L�IY��ǋ�0�@d'&\�ٕ8�S����8N\�	�XN�����}j�٭��YJ���(. C�4��A�[U�z	+�ퟦ!O�F�F�`�	�Ӆ"0}�����G?}�i(e�귋1�{���k����/G���Ֆ`_�3#���Ys�2�u:��`�m綆)�(��=x�:cS���#W���z8:;OܟA��b�8x�_/>̜�k!�6,4z�?F,�����p��r�C5�2B[��/
��O�(mv_./��>8�a&z{���1\E�з2���F�<rp/�%��:6?��Tjz1GŽ��8��a���O�W�a���3Ǳ��Ę��}�Y�rLU�:��������i�:�F����q:�4`sJƉ�؇s2�.	��ҏ�������9E�8������>}�8��4�0�J���my�F����3��3B����'KY�:0L���
t��^>'����3�A7z��<l^�ހp(��sL��1����)}xsD��zL]�<�#��Du,�k)2�Ц'��?����s��3���p������Թ�cj��=J_�����dZI���6d��a��Td.'%�O��66�B��t��i�f�Sx�耭Q�������2S�W�}���(�wg��^�yK:�9��/s�;���5�70�\����,��l���O�����y�����̋T�U�o,zAM������j��f�W�p%��_��9�^������+ߕ�[�O,���S�k1�����7_��Gҿ���~�]F.`gM�����Z���>uN�i�%f�Ȗ�`��Km�6G�կq�L(L�]!�[nt��V���8�Iy�#�i���̓��B \����`��B�s�D(E���z/i�j���������ὖ�u=x�"H�X��?�V~"�K&��	��|Vg�	>��!+��O]����礮���۷ �*��{��Z��H����^�>E$�C{���ɞ]k�����"ENy����Q�g6���7׼���|����c\GLW�0��7į_�-V���}��e��e=�I�>�0�C-�K��Åd@�/�&@N�FZc�,�&l^Q�0���ה��!K�"#����n��:�4�[��ncTi[�C��t=#�c�͵�i�?�(�	��Ż)�z�� ��Q��`ME�*�t��1-�������8;�s��g��7�z�U��g�x�?�3����x�����f �����rlm�a6���c�C�<��DB�g����?���}�,�iHr5v�.?R���:fsW��G;̗b�l���|x�`�G8,eHB�Ps��xr�W#� ���g8�Iipvߟi�,�.ȋz�@;���JTv�w>����4U�;�r�!����\�H�~R�����S��e��N`��弭#��ʐ�h_����&��G��ј��/j �hrs�;~�)��l��O�aS⠢�ы�1؋�{u��=��Bs=�2��p<=;�'��D�{������ڟ:��;�J�u*ǐ����D�n��8u����Tv�r��wF����8嚪����v���	О����\�S<M.K��H��!k�+�3�.oUzL���>��b�O輮���M:+��c.=?t6[+gp��wQ��ٮ��\���{� ꋯ�9�����Pِ,@H�k�\HU8v|(���R�B�|�%��E�����ӟ���O+=-Bs_�q.����yց�#P���B�-��;�ZGB]��U�>�w!9��E_�>�s$�_f�ɅsK� �=Qn��I�ҟYj��y��o������;������l�!ĩ�8�`s::j�s�d����w�O|�x֘�9���5^0�/o��K"��?ҁx:�����W�$�G��`�7|���+��zM�v/7���j�~���V�;\VN[
q/p����?��OKq�V�շ���_�������X<϶�pģ(8�����
����p�vit�m���{a�KW^�;#����\��P0���c�B�O[x��n��I s�(���l�1/�2g�#eO����s0�·��.%)�y������������i���iILH5u�\r�af4�ԞX�������������'*�N�1a�"ҩ;ؕg](Nw#�i�n&Euc��ᜇq��54�6Q�����1��R���U�x0#���`<B����l�+�Z�������3d�/�3�������nο~P����y0�3�m�ɿ(�\#ه{�����eXc�.�1a�/�(�T�S����DS��%k0`��M#��#a�7��+:�ù ��ʰx��+d����_{����8��q�mp��W��TG�hh�0�mg��L�e���z� �������o�*RjQ��Ђ�!c�џ9���쁏a}R�Ͽn�!�,<05zǴ��zI�8!pq����Q\Z:NF��	?���+�ժ���|�w�26�.����ښpma5�16�o�T�t�=\�隈]:�?��3���E���Y�~�>����D�73]�{,�Ao��F�;d�\{��:S��[|K�I^/�۲tz����N�NӚ%�z�;]�������v.�<j�:�<~��i���xq��v�;��f��3�����أ�94�ɺ�g��+�Էxh�ڡ�tŏvQ�8׫>�v��z��zn���3�U�}"1k��gMU0kJ�c%�O��a���������<K��^o�Ă^B�ۼ��2`���X����Q�$YW�_������v�O�����_�yl��+v����ޠ�R�0Q�.�܁Ev��r��̝��NN��_#�k�G?2�����ع���8�Lgp�I���I��Y�P9��.�_63���7?��s���o�>��~�b밊�h�֩����g+{:�ķd6�[��c=�q}[�0�o`*G��(�2xuPs���?������� �/r�)k~ɋ�'��"a질��=n5������7��M����,�����?8�������Y_'yh��uXޥ�l�`��8n4Cxx��N���'�3�9-T۩��h3^ ��9t3��n�1���@��֎��/0�dI�h29B�!���%fԡ5Bx�B|R~��v���?ox?�[�5IJ.��U�"6�02"���/VW8�C��)S}��?3���x�m?��9� y������AW}w�EG_�.-�Z$,e}�B�:���M�xvz�$R�r6�y`Fʾ�Y�Q!�Df��������t�ЏY ����鋞�9o��ʃ��.�!M��G��>G������q�0��0�^�����HJw{�D��28�?��]�:�>9 ���j�k�Գ�hyi�O?|צ��?{?G&xS��U��b���c���ʤS�j���� �iw��I��jp1�^7�Q�D�yi��7|B�H��[e׌��yg��̆�5*+�s��<���N	s0=�c���;J�^5ʻʻɞo�$�9�>�>�K��D�e�4:��}ϏN�������q��N?*+g���co/�h�R%�6�H��Zmv�tc�ϰ����pf�Q���:N	�.�8GN�r�O�^x�8�=?p:i΃~��s��sx���m��s2��W��.�G�4�_u�����2!�u�ӯ]U+�܁7\��Q��]|��S�����p>F���q�Ǜ�ނc�n7�����ki0���v%�2�Ygi/9M� �ڻ�]R�p�hl����ϼEۧnr�*�
�?�o���w���Ӈ}T�˧O�~�ׂ�o��:� ���$��Z3�h�ӾPQ���?~~�ݿ����?}��h����5010h@N�<�`z�"n���������꙽%�3Q,�{����'m�����<�!�1x'�'��(�]yi�3Pw�]e�7��Mѯ����o��~���"C���Ӗθl��hr;ς�x��-�||���w?><=$w�NN�b+�n������Rݾ�DS�T��љI��6�n�Ѧ��Z3u%o��۷o���ӷ�ɞ���G�n��f���A���sp~�٧�{m�ml_�����F�(exm��6�#�ck�M��Δ��o�$6�zT��ѣ����z��#�{�����~�i������^����l�M�K���C�����ztz2�)Eٷe4
�	�B0�f}R4J{2W�̻w��VG�����m��M�PQ�u�t&�Ncfzpx�C��Ή���1�:94��l��K��D�LER��՗��8E�|(�r�g����z�6���j���T}�h;���sF�p����r�o%E�<j�h\���`��SGO�+E��뿞���_N�� l����k�).mtl�H���,�ș�R���1*�.��uy)�O�����.��|`����\�g �"cdXT#Ռ����_�n������{w�6�mT32�>F��U��Huft�P�[��h�u��L�g(���_N��~w����)C�\�mx�qt��`�ò<h�9��K��6���Ot)0�6*�V�q�ۮ���i�����H�K#_C�.6Ч�5�6*SX�qV��<�2tx�-�;EOt`�Ч����=8:�u���.������:m�pD�	R�X���B���%d�n��F
y=iSOߔ�f���F?ѭ@�������s2m";��x���ҫx�=x>�x��E��|8��,��p����Ɂ������W�+��Z=g,�)s����W|��p�N�r��c�&�d��9Nep��s�U���#T}��|��*��@x��e�d�ި�M��.�X����Z_��vK�)���8Üuz�m���UM8�guQ}��@	?�dmm�����2~�4���hjo��o�{p�����qz��������t�����F�m1f�E�����`K��z��ǜ��f~��-R�}KD�sb�9��_�m��Y�u�"�%�}��?�Z��,�Ù�)c?�P���v��D{0�L$t�
����+U(]��ZcD���ԟL�i���Q��g�����^_y���E��/cK�
.)�����ux�N?����˯O������:}�(�%=h��i��){&��)��{��;���8���a�ҫ�~Q�����E���J�{���;}���"z�>ʑ|��w$ܾU��<komVN����b'��O���X�B{r�K�w7m@9מ��QF����Q�~^�#�zi���9��{w��l_e�����,��O6bF�!4Ҡ0��J|�������������R��m��u2�,!���`:$�q�f�͔��"}ktx�4=�鲎�Y��s-ZL7��l��?�TxoG�Ôg��p(Jj��H&�l�9~�mF��1G�_��Z��ej`ι��w:�\{v��o:j#�=���ĝ�u�W�`���V�1�/7*Sc�K�M��zg��S�Y\����g�q�h�{"�i�(�?2����Zܟg�F$�_;��u�𘖅�����25 ��	�@Tg�:�a����:aX�I?��d��X'��d��� ��K/8�]�Wr��������fd�����?���]��cЭ���������g��L]��`�'S��_�x�/���|H�N�^��r礓��I�.��9b�O��JE!f���M3�܁���ov�>ݿ���Ӿ�w��ݦ�n̫����N�)�a`u����������4t1�q���y�󳙆,q��i[|�u`u�xTi�V��u�{��`L�]�50�e�����;�(������������Q�����=q媶�����D�z��gx%�(0j%s�x)�MN0�:�>u�+��=w�2N�Ҝ[��Á]xCG�%�ͣte��ߑ���|Nuu�]�(�3���![��1%:���������];��-�e��<�RߤX#[9�M^����޼��Ѽ����O�0���{�^Ѩ�NT�:hS|���Ш�i?ᨾ�O]���5��ȟ�4tx��'X�,�^�wK�A�ŋϿ�Y+����{����/�A�gGۨ��i�h���_����"_���[�������E8��`�%��K!�+��'�v?G$�c2dL�ي^䣃=�n�U���!eo�����Lv3���e��i��ԩ����>��F�D��=k����8U�����o��q��f�7�������н�����{�������A�y��v}���k�����m�[=�m�[]C�( !��9:Q�$�w{�s6w�^���xf������n����m*��g��$��~�Ͼ��Ř`��6:
1���1��6½t�z���t���!	�ړ�x+������v�m���[�N���K+ِx�tVw��|�k[Oڈ�������X�*�us�>�Lh1m�f� ��"޻�������Ӌ�u� Nؠ�5��o�@4D��C�������n��]�刕��Yh^靈Yx<hJ��_�p|�����C7�vF����Mv#�)�=K�� ��1t�����b��u�9�9_�T��#[�;*)#�����#��da�t��"�B��=}p���5��_[�P��o~֫���C��S0B3��o�5IN�&���m�/�G����?�,t޷���%��{e��+��J��oO{@yu��:Khn��ԯ26@n�h�~�Htγ�����zd̹ģ����Ɔ��_Y{YT���9c����(RX�t~�G��h��yT�����E�����?���wu?��\�dTnAcɌ+��e=�.���ꙺ๸r��$���@�Y4�غ�x�;y���G�_�������ٽ)�����_ݟ�q�ݷ9�?���/�6��5��:���p�J�8K!Y�7���Y���`�1^��[Z����`N��Ik�tL����Q����Y�<�o;,�(�#�o;`S�?t<8ܣ:�Ku`��㙚��l�E�4Ù�%��/�a:������qp,8/�k�L����)������'��u%;y��7��鼗���y�3��ӈ*��ˈ/xfpk*p� 7r)��ᯌu�~�Y�8�n"����*��:<��yK3x�<��'z���OO����R��n��_��T
��_���������?'2��~�.�c+ʳ/��쉲ѓڊ���B����k���?�f�ګ�9�.ϋ4�j]�0F�u�_}���?<�_O���?��m�E[$�t��<��ɡ��ʯ[|oI��	N�lf[�x�ۥ"_��_4��g32���<���Y/_cQN;��|�s�j�['����f���a�WN�ӛ�M�=���=��_�G��}?�H
T�K�.@*��=���צZ���W�=�����o�տ?}�����Ѯ��ݷ׹{<�6_~����囖�<)������Ģ B��캞�I"�ރ�@�L�2���W�hCk׾w��闟~t������/�I뽚Yx�U���ѕ��v���Կ}%p7]{c�u\jjP�	0����~�
̯됙����t5�p��#�����i�t���3;7�(}�7#k˽��~�<o֏��D:$�p��h��i��*�����5��(�}�^�L�
نY� G
Ԋ���1�!:�kS�d����_)o��nq�l6��3�X��
�}�Ï)��)��w?e Z�\i�QH��F��zp�d��b �H�s��{�B(֋Q�4�>8~/k���{�7�<c������5u��Y�G���H^�̏N��×�2
�������+�2/*�p���\�
��y�ُ}���M;�����h���Ӝ�y�a���� �{q\'�u��rN�+'���\��o��!(8���>\�RH����/9���!�16�h�{��FSo�ڔ�2�Q��'<�����ܞ7ϟ!.���88tpF�9	E���)3c��������~�CVj�1-P5�,B�|ɉ��� ���W���}�Y�U���Lѣ��ӭ>C��[��}�a�A~���y�ͯu��t�{�f��x����M���o��s@�|ux�	��5u�Ou�]�+���/��l�?XzάS'�m��H;~�408~���]ǎ���v(��N�M�e�(:�i�mN�F�ٓxUy��w�)w�����޴��)���8��.ϧ�ā: ���˓�G}SF��Ӝ��^H�w4������CGʧG��4{?��������:��O}�)�C�tN�����u,�3/�s��\�]v��BM���;��R�.tʌ���gs����Gup��mj�3(�p��u����߭|v���^����U�"�Y߉��ќ����z�������*�f/ʉ�[��E����
</zuQ&�_>x2m����?sTl�iP=4|�|��Ū�m&�S���c�̢��wZ�5g�#��X���3X�h��?��4ʳ
��HN����z7-+�1��ؓ��:�����ݸu��\��Cَg9(@�,R�O2�4�@P�f�E�`_����>~�`������.���������ѝ��d�����v���ZO���Wp�Dt�v������c)Q��Y�]������~lx��z����ik�.��߽y�7��Y6�g����}r�)�6���u��3u?�����R|g�虈<ۥ��n�O�V�����M��CH	��7p��brM� S�F��v5Zyv� ����v�}еu~<ݺㅠt��e�{J&�� Ps緋z����!߂�������YP%�����F#:�_SS�0��F�Z'x��ʵN��$�a��Gc�C��Q���dJ"��*�e�<�Μ�XE9��x�J9)���	ׇ��yCiP�g."g�Wkrz����*/k�/jԳGI�,Do����/�E�A��8F�Å�=f�g!�?}�Mk�͚�_��[H8#�pZ'nxx��n�|�H���_zm���w�x5yٴ����paxL&�g�3ru�#��/�S��0���v�n��Ykd�A�Q����сD���ˣx�a��A~�UR�P�7��}�'��������?���'��~�g�9��1a�k^?O��~(��(g��/����2�<�����0u����:��7W%�;���Lg�<~O4�g���H�҇��Uŷ�s����N��7�,��,r}���7�\FT�p�ţ7J��1���ҶޠB$F��q�Rz2R��W��y������q�ݏ<�7\������!��ن����/i��e[�#v�\�3oz_�eZ��4��a��W�Zz�Im����ͼ޻���È��V���}�#AAI��B�
v�F	F�̽n�_�$
2x��w�O�p�o��)��vW8��WG�Ce�!�2v��ʏ���/u~)�L�?<�}_a��i��g߁���v���&��|�g�v��i.XxN=8�AX�:�����u�A�'�6i
�|�N:xૉ_��=Q���A�(gKNWV����	oH�~�|Ye�p��w�ҧl�^��^%�|Eg��(g�]�ܖ5Wo&/+�s?�l}���S�X�FI��j�y,g�_x[�b�[zp�;C/o����I�|u�Ƴ���+������U���_jю�6J[y�gBK]�Z���g|}��֯�F����+.����k�4:����ʀ�5��!���h���|�w颽�=KV>Y��]�<N��k��-�%>9�M�w/�������$+��}p������_�m����JQ��ߖp��+=3�_���W�d�����+en�'l�'�E�&��N>�-��u9�͹,TY2֨	�H�F�u���X��1�Ç��rԮ;/�߳���}����������w����l_$̌��s�C�_�V�\��j)ʕS|͏q6H�]֩@3n����Y2rE�*�������N��)�:���4��`,Z�>�v�wf̎�\e\���m�|����E���Z�Y^�ʄ�@b��y�
���SfbV�+���gv���sE���	�X�aS{g�
RXuS�D
��T��� �`z[~����W_�Pw3؄!1����C�1���[x�(ͽ	/R0F�����mB��E��{�8�\�K�vk����D�3m/��6��Zf�6CZ=y��������G����ѻ$�e���K�{����/Of���NcY�p��	_"�ɢ�K���9�W=�gY�f����
?�tL��������zQ{�C�ݽJ�dޟ�ʤ V�$����9{/n���_���aa�$�u?Ӹzp�G�����x@�_�}��©h�~��rс_��!	��@Q|�#�)�����S�?��2P'��u1�'9R�����ngh�o#��>K��&�
�W=5���sv\��o�h��ǟ>��Q�8ޯ^֪����5tq��h�7vzp��c~�aW�U���:�|�AX�:K��4Cy��Gބ?Z8�{�`����u�S�#he[�u��p��ȡ^on�4�B�a�~>E�@�d�R)*�c�����M�)c�Tx���l]�/�rb�����[��x��g��m��u���E�].g�J�luL�e;���WH-݈1���G����޻��b���ؠ�S�0#��&y��R��r5�s�ɐ �
���~���=�;�Y��J��{����{��\��F���4������� �<��,|�,`y���\k�i|�Y]z3�t�����������9���L�:���
N��4yK	��5��[&��o����t!C ���BȒEk��p�:��,-�cc�qdJ�����Z4���O 4�,Z/zS��ᴆ��M�����;ɑ[����Y�UV�G��~����_Gv��QՏ[3K5d��&YR_�zEA�����d!��mu�b�L����d9JE���}$�9�f�����af�%�F�{7ﻪ+���#Z�˜⒤��I�NK5e��I?>\nR�{��w_~|�۶��W�>����^Kp<39':Q��8<ii'k�q{R�M��@�����˸��Y~ѶE�ZߔL��Y�d��_���7���� ���כ�W��S)�����>F'�Y�ہ�^h�~
�e�aá7�4�8��j���G�?�(f�,HV~=���+ε��ə-HN�X��� ����`����٠�,�3���]�~�{=Ű
9���5��I�bh�5!�aSM͖���+7�����bg-�7A�P����G)_�~�M��?��'J�C�t!������T^��Jw�A�U�̉����bx.�h;ǆ�|�mX�� �7��>מsT�,�L �J�R�j5�G�/�������;�?}w���o�G�Ԉ�)�,g��L�X�1�����*f`��ps��[�0JV�z�k��Xh�ڴ��O�At>��]��*��	��h�$��M(�У�;��W�g����'N��L�d�{�o�o�<l��O�.}�c�^�ۂ��4V��G��_��������zC���Ţ���s!Aïc֬	��ҝ��f
j�S|�T�FuWZ�8k��<�sx�E
��5\)�˲Q٤t�Oa���ow~�y����:O�n)���-ț��A9:��wz�S;��x���7C5�N�2:����ڇ&wr8����7�P>�c�V祷.(��|)��v=)�`�\΢��1�e�~y�k �ԢU�*��I��M�L�E*�WZ��(m=S��]Z�X\��F�M�l/��:ໄ���K-'Y���O+��;��w��u�ZN���^κ.Z,�(��d�$ͭ�I������� ���G-7S���R��v��]��U���M8�?;KJ���~�_9Ȟ��->M��믫,���T����x��k&��V�b�nx�~��42V�T�٫79ι�B����n�|.d� [k�O�2|YH+s�"wCz��Q��|��d0�0�Mk3�R���?.y�lz��|�]�O�����)%���)�L2Z�ѱ��tl�Q���d�4�Ay�.��!�͗G�ep�6}W0E0x`�)��X�|`)�V�����Ѹҋ @��������3����6��O�x��C"`�#C�[c͈�4�P�3���S}'��^ʹ�X�rLa��I��X�[Y��$���Wʮ�Ӣ�:R�gu R��)9�R��X��oQ�x�1nh�/(�V%x��a�k�(�!���?8���������h�����%e���R���Ȫ2��	�Qjn�zg�I�C�ƗY�W��ĉ׆O�%7����+F�Q	Agu��=���t*&H�*�U����BqZ��0�)���|P�5㖂x)E��u��&�6����b��yV�w�͔Y�k쭥�T*��3�nf��)��kEV�P��h�𓏐Qx��x	Ǚ����~*JYb*?�L��i1��-^OY� g��!YB8G~���a��������\nh�Z�f>����'h�|<��:Q)r�]�F����V �)*���vF���Q��cMI#tXPb�h��k�>Lc��3'<�/��8Y�}08c9��I(c VK̌��E�֑�Z���#��1 >���K�GSl�{a�U	9�S�^=o��&��b?�3�� �iV:K��
��u��Px!�n��zn�R��
9�𞼦��m���}�8�~��T�kU�"u?Pނ%mʴ^[�-�+A��d�p�t��W(�zx��6��R����0F�+�pE?k�=|����?$L^~�	�Ze�J71�E��]
����Ya�4e��!;��><�� Ȅ^��s��	������Y0�CHvJg���y�O��}Ხ�Cޕ>�Ari��X#z���ş*�&c�"�Y$J;�ŷҸ00�R"���Wx�	��Wa��5�Ki(m��xxu���úG�Eӭ����0�>�;�[�K=������[q(�+�Jo�q��]���Pmx��p�Gǎ?�ga��Q�������B#P���0̄�}�݋��?p��܏s�U�p�P���̭9���xZ��ތ/�돒�w��[lZ�'�u� ��K�����H=Ҧ�o��)5�R5≮#7W]�o�K���v�6�-�0!��i�:��52hJ�0�/�QV]ݐ�h��Y��\��7]�����F�4��D���v8m�)7��1��+�	0<!��ܱC�9z5�7��e�N|]�����pΐv����aE4Dg�ʎ5������Y��x`dvI��S�! ��Yo_G��z.�����1�)<w��/l�F�Wb)���Wy���L��W"�:������ڒ�s�y����,_��_e�ʑoa�^6:_�Q&�OYuI%y��wɮ�&�jٔ�2=�����ܫ�˥���(�H�\��`\l�(�!��`o�!�됝ɳ�s:��i�������*��J�+�S���y� ��7�Y��0�h�!S[5x�����RT~b7Z��9Y�Ci�����	���)M��	����tx5��q������7�t��4����>������ׇ��|\W9�,?�.���<KA�lz���K������䔙��nL�u�J6ؿ�����SK\<��#�Rӭ�4%L�MhP��0��)+#�6�Te�`�e�	��C���|�Tv��5֡Y4� GQ�QN.1G�T��*�K9O)���\�X<����Fm�����P�"��P�q�7�k�m��lKU�=BB��P�w��2}���QA�x�G�� �W��J~�yx���>=��4���j���2y��T|x��]o���*hH�\���8ol��Z�Y 7:\L ]��-�7��؋*%?���e|P]�%�bA���V#��S�{�*l*p�%�=>�)?ΣV�6cMϊ"���l�'��������K!�kiv���c7�"QL<�[���� �vF�	��GkX~ŠL���hY�j^��A�op^GG���px���}i���°~4�̐�� Qx#����\�Y�;��ua<����5N��ຆ��v�@4T�=�ȑ7�n�=w������ яg�F��γz	_�����n�Պ��;O��4�ۊ�8;�P^����Уp��}�Y�6<q<��Q�{��� ��ɔ�2��p�����dm`:R��R��p6������ͺ����Ѳ�P�o�d�0���2Bh^�|�4��W�!����c�b�)^H��k-�x����²0�*z	ςe�Ays�g���7�aK�鼗��4�␃u�z��F�q�Nv������s�Q:BF��g����b�k�ڣ1��q��fP5ޡ�1ä�M�V}S��js�	�� s��?�z�E��+\��4u�U
X�Lz��'+Y$��_����YR.�l4�-��9�W`Jפ����Qc��o�|�i'�4�r5����H�M��]���8VV��;y��V�������|������N�cF �����xY����{��\k'��<?^���SG�1�2SOR^7�I4����24�֪��r��h{V;(~a�1<�c�N:����ž:-�mh���w��0\kR�.�,�>�F+����j����iL��fMj!W]� z�?3[�<�4*\C$��[耥P�>���v�^�}�D+;�~k8���[d��o3��k���F���[�]���Ŝ�d���X��k����Q�0�(`����.�H*�񇟦����p��g	��A����RL�8/�XAa�N�S.%'�4ZR|SE�Fd�`:%[�upgz{�MȄ3�}�U���	�YX�<���S��-�Ğ��1������*k�B�����y�o���㭫�P�xmL0��X�Rz��^�#�G�5�x]G��2�"�9�_��7�Q��,�	ﮢ!r1�*}�|���z�1v�T����J�\��?���_o������*�T���|	��U3�o�F� !:��գ���.
t���^[fV�����ʏ�.��w��V�Q��PC��~~�������ƪ�JX��;ue^}�o�[�=z�����|��+Z��4�2��$nt�\(Ք+�t	0���w��\���o��`�7�h�v����J�����4R�f%�F��b5d5�#D��������O���1�x������q�+pr����@�����bʅ�s��J��>�Q��\�'��V��*`M.OJam|Ye��w���,��MӍ��?I�I�F�l]�u�E�
�X����kX^���If-Y�۷�������J1�I����xI�:�  @ IDATp ��й��4���-��M|Y���lQ֭�T��T٨�Ȫd�<��s�F��-��G����V�޽j��Ң� ��Y�6��;6C|��5�Y~+��FɌ����G�R��],N�$+�h8�����Q>6�]���H�V��_�=�-�4��J��=}h�إF�L`i����mo�ܷ�3<��ɠho�﷣�.��6Ỗ�'T���	Kr>^)t����~�L�%Xsj�/a0� ]��i�ϵS���|����k�����j܋�0:��+���t����2���^�6{P�z�R����GiI��+��֘�Ž�q��E�a~������^X�z�*޺�`�\��ת'x�r�p���X�}��1��zr�ɺ�c���{H�ۮo0-k$�4�����i��]oO�,`�qh�Y�JaS@�$�������HC#.d�a���OL��V��:�<yp�����y�G�Bd���c��՘���3I~x�����9��zǬ�c�
���J���/,b��s�/Ċ�1����nK���;����s�������|�p��u��Ѭ�l���%aBQ-gz��/4��Y��]/o��r��O�� ��1�ZB��L����*ؽ�O�AB��sQϤ��+.%�"��/]��U)�!]���sܼz<�{mO�1/����¾I ¥����Y�%(+�۲z�ֵ�Hʪ�t�4G�g%��J�C�b��p א���y�3��&?����,�=e�4��&;�A�B�%C�8~ȓ@��?�4���ɣ����]C0<�,��Ś{�+���H���e�UZ���\�m�+�=��l.���̧��9��*$��V��uufz� F7|H�m~]���:���ΐ�x�
=tD��w�X�(,��-�A�N�V����;�����5.pY
�x��y�U���?����tn(��
��ݨ�jgJ�<j��?�®�R�4�c�P'*c��n��7)pr.X��=�u����ʋw�]W9�[ԁ�oߜ�BV����O�GiZ��t}���~�ӧ|�	g��,���s���ϓ�#\��:Xӥ�rN9N��Ą�ߔE|KT���r�ǖ�B3nx��:0� |W^���Eg?<�\�D*Kk{]Ih�gq�dG��aO1*��\I�7&v�Ru�|��"��^�s�<ϵ��N��r1z��Y�w�����h�[y�����?r�F�1\{!y��ס#��T㱦�A����8
-�DG�D#�eލ��^���rʗ$+��,��Áf�Z���E��?Ds�7|������\h�4��B���skp�n1қN����/Fl4�SЮ�/�M_�/
0yQ��\e3��S��'�(�(��T�T��W݋FGޜӕOD����C�g��uY���,��ǵ����������o�q{{��Y���Mt m��^C���ʉ=E���C��E_�Zj'i�&��Zq�A��ɣ����c��4�O�;V��,���.��'� �����<�l4���LL�l�i�`�W�1z���e4���!)Х��$i5�2b��� @!_fт �Z���}zTN,��ڳ��.&��~�Ne9w���̟������03���>�������u+�~2[��B{�!�g�!��\"R��N�'E�F�ŕ+1'f!���z����i�)��<}t�_�?r��.	����g4��ǂg��w��¢0v|�>�Dz+x�=��M@�guz����y����ۆ �rn`~o��/'wP
(Y��W�-<��z!�X���w�};����lâ#�J����)NU��56
�Ț4�tb��D�B��o��x?�3߾�y�g�߄*eOP����S�p����70ä���v��࿄�
%�N$�(xevx)�{��4G��֬��1$J�����$�G���ɨ���@�z�$�f4�� ��܋��v�ŉJ:���(�xa�X��-�K�.�Q�&��E�x��2�Ka;��	�#�]�	��)� ��ۢ�YH��G�E[��@uW�	>!S������VD�k��`ǨwYF~J9�\9��"��6��z�4�=�j~p~(�����+���^�8��:*��nu� �/Xh��Fg��G0]<��z̨�=4:���vv�{�ߊ�;p9��o��L�.�y����X��JU�����SZৄ9�X����-�h,e�[�Ճd�\���XvãCw�"WX�8ᦤ�v�������L11<IN!�2U�!M��hhmup*��WoɕT񑝣6��{���b(���O6��
J���o=��"[t�����Y�W��5yR�����T@����ߴ�ACc�Δ���ʫ�VY����7�a_aCY$ˣ�Ny�}����&@\Ȃu��K�h���ڪ[�o��gW�����n�{9�,�_T>���G��5�F.�M@�mFm���Ɨ�Y����׆��yx��,��s��ɧ�7yxY��_���sqI�I�����Z�����W_�_�][�����z��A��hۡ,e0ʪ�{�`p]'�������OF��+o��%L=��<*���P䝇	����Y.���x���Y<��E��knƣ�Y���U�S�@�9ĜH��A����L��R�Ű�7,	^��u�Ƃfva��_��x����i�|�h��;?�p���o��x�M+?�������|��˯f�~JCD��AD12o�p�
���F7��zG*���4,5.�L��͘�ݶ��ǯ��Y�n ��2���a��/�m���d
����?��������û�k��{����'��ܬB����cb&T�5��Z1b�/OKH���,�F��71�a��v>A|���'�?<|�Ż-�`�h�����
�7+�e#fI����)�>(^�����o�_�/�Aֶ��b�ZV�_FV���Hؗ�5C����;��Ɣ_W
���xx��JR¥�n��T�3~�)C�,O��(�jHǮh��ྰ}U��kz����w�%��G����v��FT�:Y�ш��P�K�a�(��������7�����?�d0���^�-ó�g��8s?<�y�:Oу���rthlWCUz�ZPC�k͉��4��)�¬���
�a��s==}֎u��܁!w盍<�-���l�����X�S4M���ʤpc���>�E=��݄�U��mZ��xM�#��N~���Z�a����o,cC��P��=�⸔�n�3����<�s���\EX�>�~���9��n'�`��%��_�`yZ�����;�k�r���{)S��^0H�$N��e����ͺ�Ko�L��;�J��c��^�P�(�Sx��E�\=^6K6��gX,��v�:�ر�Rc����,T�V^�L���ʯ����"�¯ӽz��)+�;b��eh�<�M��x�(��(#�}���\�K����X<�@���Ƚ�f�����ޏ�q�R�d�۬;����+�bX��f7+؍ç��v��w
Ut������&CX�2��,8�|��/N��-�)Y��*H��hx�1�܈`0Ôt�^�Lt�����Uf��XG����g2� ���/]�r����s�����V��$���5m3��U��j����э�˒;�U@�}�<��巄/W�W���t�_�.~���(�B��P~�_��s�5>���k�eWge�^m����У��L��n�B��&�qN�M=�}m�F9� ���]Ĉp��~�Z�f�����4Zd��f��)�t_�Y�9��_�G�3V�2�띟F��U�7_���x��~?k,�enFO��q�ED�G��)�q,�_�@�1d'!�*�jY�K^�aJӭ��o�_��Ь1��(h���q��)ORy�����-]΍
���o���>�H�z��Q��;�'[t���jţ�5�����)O�F(���$��d�=��7�f�JB�i�k�ɰKY�.N��%%�����]8|����Ƿ�>����;�-�4�2�՘�9�brϻa~Q~^]d�v~���8ܾ���QK�5���-�x�H��C9���/#
�ߔ�R4'~S�g�S��Lz۬F&h�ʌ;
_R��MP�$�Y�"��%)�A	ש@�9+%����FK4M�V��P���rY�Q�`�υ��U��ëꥨC�~փ'�D�2�����O���;Ǣ(�uo}����xқD]:�9�wLw`���QV jF���m���?��
;�v/�R�i��R�ltO)0l-����az��/.�=�&�Ļ|�$�KaJu���vx�2\f�k�8���N�\���1q˗+<�p[���*4Z�ʓ|�N��,en+J;.�N�pxm�ܳ��wu��֮��0��W�N����������;�X�+d(x)�'�s��m��Q����N��s�S��y������;9�GW��(��k��}-@��u�-���ث���3:DY�/e�9���ۂ�|������"o�ꀣ9
M�~����~�ZNo�]�Z�Ec袳_�+_�����NL{W���B�\24���0�5.��<C3���{y���op+<T�.�K,�Yћ����e�j�b�O��}��<�24����2͕h(R������\,L�x[�C9�&�R$�<t���3c*����	�E�x.�o��7�q�M`o�,�*����Q�p�%�z�z�hZe�N��;�k��/�L�q]��\��-]r�Z�K4B7����_27�-z��J�C��]��x��n�^�a�gaU�ޣ��$k���"aAO�6y����{�F�׬���(�~�_�´ax��� ��z��c�h'�*81�G�w=s!A������J�
w��V�z����eKC<l	��Y�ndA��Ï�������ߵ�^��Ye��m�.3�G�b�Ic[�0�@8�ϓ�8)z��`v	�U��}������Q�^����5�NLV :K׫�{�t�������徿�_�������������?}���ΏߏRU�x6������U����f�@����S���zQwM<h������Z)3�aR��M3��NK�T��	+�ہ;����,V�t��ƲR	��,�*�a���>�;����
���=j4zߤ�l޼�����m�z����򔐰<�[��`C�ZID�c�wݽ���� ����>e����u�Q���W� �j
^V�f.�l2Ƽ�-N�ȇ㹙��Й"_�n�c=4�i���h�ҍ����wd�<��#~�.�*�^��U�u�g?����U��1���Y�\�����Y���Y�5��΁g׵�
O5]�� �Qr�f����vA����A��7�3�1���t�R$�����Z��a�hRR�`P�,��">1^�W�մ�-Í%�ʫ�[�5|@����2�]����y^#{��K��;�`���>�c�N�Es���a��n[ռw�#:-�c���躏���ȫ��m�����	�8	�ؖ4q��qv=�8jB�@gJ��������b��w�X���|����]W����釶�P?F4M��/ř�X��HO�p,�:uc!��W��_2��깎Sۈ@!�8T���J2K�b�qf��ԥ`���Y��,Z�k�(HC~;��Ka�Vf�����G�(�y��⒢����ڏ���x��C������D�$��i�a�}��&�@��y��g`�.�;�7�$��0��/u�G^�/�O�%���[j�^���V�c��>�@��^ɶ�ReN��~�$䈦���K3��k�Ss˶@���)�� �7C���V��LnN�iH��c,��]Nf�m� >������j8��5vK9��B�UuDuqt�W�#����ɄY���I5ί_���Y���M;(^�-���� 3�Pff�Y��Ě��a���r���׸�(�#�C�>��$Y�r^��2֛q
����Õo��ո(P�)�O�n���cކō]����&��`AXc|���z����X�r"B�	�iP����1�{�L�`��q�'�)�[BO��o���i3׾��!�ϟ��d�U��A�Qb�k�[/�9��y�fK��ޯ?~��χǭ\L��|3٭
'KN��@��u�Q+�~��K�{�=�n^j��L�MBPQC.3��[-��0����Z󝒔����2��=�\���BL��-;TN�����\	�׽{���K -(|�T9V��n#��oT�!LE��2�"h��EP��K�@/���U�UO��Ϛ���}ݞY�8�����V�b1��>Oixf6��@��?�ܼm��9����.����ryf�Z���,�x�`Ň?>�m�ߌ��5x�ʛk�����Q F�����������
��%.��G�ޯo}�yKht?��Ѝs�U��Q{��C����b��(��w��!+��5����c��%gp�~Sg��}6�n��i�=SQ�0a�-��)����B�S�
����c�XB	O)�]��s��g�����"&�e�\<�t�SJ���������Z�(��X��g�(���!�u{�!��EW�!�pV�*���)��#�ʼrЈ�_�\
�ă/��!���X�w2��I|�?��i���z���b7Dh$yr�p;�OQ�Ή��`�kڈ^W�d%|���g���o�rZ�J~�)�gib�uN�F���+K���uʢ�*����� [���^�5y;{��{lj�[�P�}�$�X����x�vp/s1yQ>)a&�P���;I���2#G�/zw�3�<�Dk;��?�4��Uc�+>:�f���e�խ�V��Ћ����O4Rߖ܇��r�s��а'kM�ЍB��N�-� ��a�^��I;z92��w�);�;(~��k��`���#��ڪK�VY��)5�Pgߔ�������*���d(*���C���ď�M����ڬ���B����rFV�L��׻�q���P�(�SG�&4�H*��Y�®8��-�1-�i^p��aw�3���+�')	0+�=9i��i��7��G����V�O�5y����>�pzr�߄��5�L3:� ���0T'�1�U�F�R8�A!hX���h
��N3!?N��	 �~j���~���R�����o��`�́�|���Ɣ/U�?j��w�}�=��J-^�4��⮯�����3	��z���\O�>lT:��G��mgۇ*X��r�u�Z��ULQ1�׸�x5
����r̮���w�M#ŧb,��4+�O�hN(V!�Ǥ�
�2]�x"�UoXc9���]3}мt��d�o�xk5&�`Ze�@�Hք7Y��������o?�i(�E�ԗ���Vx����-O��P0i���T��I��y��LM�YJ�4Kh��QӸ����:�D��teQGb���W�~��S�1]�͌�� ���,�xaY2�E�ȵhr�[��O�p����P��1qL���4��]���A�t",��6+�U��7Y���ߐ�
8���V �i�|�l<m�M3}>�Z��Yzh�Ooh�����!,i't�Q4�Ƃ���K���l(�[١ ɧ�2�k֊K(�=d�����p�k�|[8�w�z��9(M'ep�++�g�B�)�>w�"�N�u�߂�z��%��Y ;z\�V,HEr��;�].�������p_u_u�µ��42h:q����mL:d���,�&dY��|��"��a���fĤ�r��/%�^$�l���Po�J�{S�K����>��~� �zv/�$��He1K3G����[]��\�zӚT�~�-��7�]X��֬Y�\V��T���\4,-φ��LO�
9?R��&9���(HB�0Rg��B�<�h�X���������,50��2��,��$zn*���Ⱥђ7uZ��^�]DS��d���cE@�/����X�u�Ս��8�^��\M����X��r&�o�.޾}+>Y������z`V��s��-�W�+�]�C��z��\��ڟ0�n�9�FU�cud�G��8~8��J�/^��)����֑_/������A���Ba�gp�垯�z��MȢ��3��m��Al��1!�L��-V�]�+L�B��:\TܫYUn7�����T�R�,�?=�!%x� �����^l1W�Vp(�p���y�"�"��˒`3ԫ-uqk�o���7?��i!��b�Hf��֓zUc{��fY�Q�0C�ر^��-�a�K`��Gf��9��Խ��_=of��u���<ߩ�S��D�a��f�/�¢�����^�ߥ�_WLC���T�p7;��X
�����^@i�I�NM1�P<�A�d� |�����pz�]z�)��/S&���_`�`(3�'l��Gq�y\��P+
�����o�6���n��^�7z��2:Z����E+�/�b�	JgJ!C;��ߘ�U�0����
߬��
r*�Jm(FIC�kxZ�v�^��J�u��SQ�="٪K��A
��+ܷ�p���	 P� p���#�`hY�c�(%[��1D�2E!j4���c���®�|Xܭԍ#z
�,��O5��~+#�C�`�E7|�E7+aoh�50�1'���Q�ܱ�<�s?�=N>JW�����V��;�z�����V�4*�wx߄��M�����0[1��L8���ݽC���w�o��x�_�;a�бn��://�{���2�E�Z�Vz�|�s{��foݏ%-^� ��O���9�S�W��z+ٕ2N�?��c��R)'Q�	�r<��^(M���&��^nV��N�/�;��f��6di����(�eS�?d�[.k+%9�g)��y,�)��űM�~q��>��l�wn\l�KV��pዏ��ً�����!��Ǘ�����_]5ɧ�K�r�� �O��oa:�*/�?~0��In/"G�!Vy3Ԋt$���<w�x��@}�\&��u�_�\)>�>��]m��u��Y��y#��7��~Q)j���`D�C�ua�"�dӆ�$��$����ob��5
�6�P;u���pcp�ed��#Ȓ8���T.�\�B1�Ni)����S�1�:�OCh��9��s�m�t)�㿩��$?�	-Bg��ގW��;v]�+<\�W�'x-h+�^w\�+�lY��d��G�]�Q��1�I�7��­Q��#ھ|�hA;Fޙ�O�/!X���z�'졊����S�&���@6�%���|@�ՀEĞ}'S��	P�6��i�㗓ՆB2�'m7�}���xwt��������;9F��%��	�P&n7m�����R�Xj��)i�R�l�a�v��b[�����T�[ͪ Mg]�a(e�
s)�۵f�ب��k�,�G��
145<��@a�*��r���Lb�)�U���9�2�;6����!�2��R�GK�	!�b�m�:a���z�T��ӳ�#x�e*���Y�����۷/������om���h�8���y�.�)}����"�W�%���7tCC	�-��@�R�I�N9�w���z�b����E]z�0P������eΣ����#7*�b��)����w���,��>ܻww�$��]7���f��;֭�EB!����9,��G�u�t���Ց8�Q�f�Q����ʷi��f	�:R�#��l�mw��_���z,W������@�5���.�z������:C�)p�Á�䏕 ������Fa��xƮ�ܹ��u+S`�#Kޜ��7��X����/�]�UF�7�l�2&��S%U8��4�l+v����,K��ͷ����Y��^>ܓ9���H�����ZF_�Y���V������Ф2�\�pd��z���w���a��cY����󃇏�'��}:��YF/_n���%��Z�͇���Qr�"|�UV�癍^ש��2!�1���t5>��(������*�<��:9�U;��G���G��%_(%��uT���k�+����E4+%2Z��ד��\ˏ9���K�,���}��[6�FC�����o�V�H�݆�6�*ou�U����5��衞�����/��~����Ky��G�Hy��bX�F�Vg���:��|�l�~5ڶR��o)*��J�V���!�}/3o^6����i��{��Wmɹ�P�'�P>!����JqgT��#ȇ`�'���> �r�3|�mX�9zV����ZD1R@V��3X���ҝ]
#�/�4��Z�\D=���:·oRw�~���G���7m�8�݅���YSN�p�t߳מd@���ҩx�A�Sm政��!�S6���1x�O��?s���/������x��* +���L��f*ؤ�sZ�4�y�]� ���L��K
RZi�C?�m������:��x�Њ0N�����1��z�C�P�0�
���q<�����?V�����ʽ���./�FS��ur>}��^�E
A�'&�x���k�3y�CmJ�,49���~�
s�e�/�V�z]�j���Мn6O��zO9����,�#{F>`M�̚3	@�G`�C'��#��*��ʖ#�?T��N(ǝ,�&����Ð0Z�*HaL<X����	�K-\�(,	��?�]h�埀S��XN�P�����q�ݙ�P/Vc�lU��|�r���?I �5&ڑ�^烶��d�{��;�>�)uJ��۷�;�{��S�um(_�$�M"1�⽔0��� ���k	�')M�)�vF�����bhzSw�jꃠ[)�q��FNxu{	C�Q��NC�����gED�,� �ƛ҅'V���(]�J�JXA>��yT��uuhuv6�R�4���(}�LYHOu�Ӿ_����,�MQ��	���m�C���m��m�t��Li��}��V�,:�hp�Y���ʛo�:��u��6 ����?�|�l��q]k�������^<�$�~�����{���hBҭx�B���?���>�g �:��������dy�zC�!P}d�T�n�h��Ω�O)�Z
�3\�M�tM ��si��7
rtKy�K��O��:�t,���C"�߉*d6���偅��O�NȤ�A��AiT��_[��j�`�=e����<L�˧�Q2����4k.~���ѥ%Yu!y[c.�!�X��	��}]�)G
�N�7�_�`�~\��R5L����&�w���,〞:?#���]ꉖ�����x� �'CS�-�B��k�%�r�7��tN^��Ս /}�uL{�1���%'�@�D�q)�řL�rb�- ʖA��t�ф�i�^(5c����)�`�g W�Zẟ�h �>�ߊ�NY���>�4��An�l�]!~�������AI+������1�bl�z<���B�$և��1�"ܿ�5_E]yG���t��L�m�,��q�����8=�2 S��юb�� yM�%-�0BY�8�����X�z��s��xMXמ;(!����
5&����y��|�;�2|4~2UN�2���y����7���`8��I%y�;���Y��V������K`ގu�VC�NÍZ�iqP]�S*�!��Z௪��j�|$ޘ
]~��y����C�[�y�C�)NV��p�O��%:�)�U��SP�i?Z(��-��|6f����L](ok�G�R֟z[|������<z�4z��g�5_�}[��7}p3Z>?��@^$)��u�X�X�����'��4����]�%��W���\�෷���9�nW|��b�5dcV׃f�~��O�?��������f��s9�E X��O��O��w�efz�͊o>���Q�(b��zy�����`���wm�ug�BStp	�nvn��QhJG��슪ή�����S�^6�
�1��hX�%,L��m>�z��;�W�v���7H���<Y�&}��x-ݱ86���"�p��P�,�a��U�t�NW��\4�m�k�]�n��U��u+:�a�w�#��>��|�����������q\7Ly��놻�U�6
;|�s.%m��T��U�+.:P&V]H���xuLr������	X�Y������)aדO& �ey���U�r�~J%u~�Ӳ;-:mY
��{>���o���NH#ё�`-"�ϧ�B�Ϝ�+���P=� [������~������RJ��}��>	��@��^M1������o�z������f�2)L{�2F�sgF?���t��q��_��O���9|S}y�Qؒ��s�S��8���?X3�Y uZ;G	����3<���1�c9�u��g�a��~�<���m�Bg��f5�����������O?��-��,u0��i�U:Ao�g��&7�`��Φ��s��o�}������I���
CI
�pT8���1�&%c^S�*8e��Lvߓ�QQ�*��9�^yW�¡�#��{|�h4��Â-}i��:֛ �G�ߎo�}��ر�S��A9c)�t0�S�(B�����1p|a�>�v� ��<���Vh�'�|Φ��P�.s�M�c�#�uY�~&��� ��"Q)C�\�GgWV>T�]����x9"?ְ�?�y� w�����+�0�<���Í���i��'�%rv�����|f���s���s
���ځc���7�q^�m��
>~��S��͔/CQWk�_�]T	^E���r�54&lUg�4����;A�|K� ��/ݣ�ƿ��Kb7�FA��*�p���G�Q
+u���<�NE"G���$_����I�hcIB�q���L<������	��<���T�&0FK��{OB�MАp+d�e�ʇ�z�WK|��f��Z��?���E����Q�o�c�(��ߵ���_���f������Yp��z�ر4�Fx��h?TW��!{��aE6�����]��c�(�s��_���A3y~��ߤt}��d�����z߷�*�d(��XlZ�,y�K{�࿫w���w�ޯ�:A�|��(�xOJj�ы�����A�r�ձK۩'�g�ǄP�ESW}_�v���oFPv��|�Y>�0��.e��g�V�C7xኮ�Q��l>'o���	|�czΥ� &@ٿ���Hy�s��������NW2�~_��=6���Ci���CyL���9��:�ܝ �����������m��t����,�U��X�&�C�(<y�����=%���)^�ƞ�9U�Rʬ�d����S�,#4r2K�唉��e|��G��>��M>i��{�<,7��rp��c���B�0qp�!��ᒲ�=e�=!]���HJH�\�{���������ǹ�ċ�>k,���(����IQ'�ܪ���8�'�|)9q����r�p�a��OR��Qz:��v?����ɚ��R�X�]�Q��~�?�绘�U���:��37t\���c�'{�P�*����_�����@y�{:y*�H۔x�3(��B���q��ۄ����ï�~~�4ך��k��o<A�ƨ��VYh�����P/�΅����: K[r�J�fu��l_�!<:�;=@S�כ��F���x��1�_^&�Iw�]GO�}�� ٣�Uw�=к��wV֕�i�+�����_��Y�1(��w�����O��`�OT0Cr�#,��n�����5P)<S"8�Gi�`6!h�8�:Fh�dd�ۿu?�*�(�|��W���{T������2��Cw��$��͔�[�<hHq]����نea�nf�IJś���ԙ�x+GÎ}����?H���Z��,}���a�p��ح�!��B�`1�����]H��wh_�G+Y!+��_�����S�E!�A��@S��\���p?�9&-��X�s���(g�ԗ�!��.X��|�)`皽9��wf椖�]�F:e�Y^�x#]8���^ή��y�w�S�R��	v�滇�>�<����3�	OH:,���Ͳ�U.kh5aP�7
4>�6����4k���͆�����|��|}&��l�ː�S��e�~�/^؄{�H�H0S�A�� ��;ӓW>��Es
��cʮ��ϱz�G��	(ܱ4��\|���T�ޠg��Gc�{�3,[��`yY�z�JQ���	_���O�$��s�ՀD�wY��~��c�,�9V��� PL6�`�m����#`��!����h������I��E�vx��Mg�@߄��N�,\�'���9��"^�p��R���ʣ����$�Ҩ���g�%�N�`�����v~J�2_Cj,���[t��3IKo)?���� Nѹ�
g�#V0�~�����O�0��ۃ�Ω�*�p�+�a�N�����8o��|	u�~�Oi��±Pb���ҠZ�>32s�(����������>����Ϛ�n֯�z�1
$��,�A^�B���J`����&�����O��X�+^&�=:Ξ/��W��El�8�JΨ+dڬH/��w飻td|\fbs�:�H�!y���d���^�����]oʫW��dc�,�C<��݇��3�[ۥ��R�Cn�<~�뇇���&�}���n�Ϸ|�|�x����y�|���=|3�+ܖ'�.���!����	E�XO�۴���rE�ű��E�:V)�����+�HĐL��t����wC��+xo{��(�/� �|h�}�VV�s.�n�l��C\�γ<��W�8��/��+��.�w?�֛������V/mՐsH�@�歸���,t�������8RMv'�E�?�;֯�#N�ֵl�v����~�ax�@����|�i 2�&��hH�uLak�4J��7��x���̌F3o$<���"�ShXJ�T4�=F� U�)h��U��"N���"t�V�O�*��Ih�g�^�d��>q]�|�-��NB�z7���b�%4�����4]��j&
GK |Y��͚]���@��%�/ue��N��vx���5"��(�W�C�؛�/�(ٵ����x����o>��!�������L���ĳz�����i������� ��p0LG�қ�\|�!�+	���+g�3��6̢~���~����Wxe�zw����tش��:�����{/��ӏ��o���f���H�!������/ʸ�������2>�����0N��A�m����Kw���w);�Zƕ�$��ߖ�S�
��5��3�1�q�bJ�=攆�c�x��9^��_����$��p$,W�����b�&�����i���w��ǹ�����|y�^p�l���CZ�h�V��0��V�w��JF?嵆Дkx�����y5ޔ����J�4}�Ѡ߾yZ��j|�ДY����g��������B��;����خ����YÃd��'���t�5;�e:YKNZ����tl������T�Q^��Sk:+�}l�KIgu�J=v�����ͧ-�a���*7�'��L�g����$*�kd@C�O�{�)��~8�,?��ԡ~Z}�����!�XqX�u�xXZb0���&ϑ�Ƃh�f�w�����c�Jv<K=h3kKi)�'n)`��X�E��w����ګ��[[2�w!e2����yu����Φ�J"^[���sh_���X�~xp.��s���ە��i\�[�ȑڦ�3=�pxS,u�$��]�8^Vrǀ��}��NO�O��c���\?(�?��n�~��:;fQ�B�}�^��4�|�k���9�ٍ���y�3�1x�@x�I�q�֊ݵ�^�}��_�5�'?+���I�,����q��ڀڰȝ;?��*֋�T���N�T.=0=Ĭ�ö�F������_���W/����f{�I9�[���U��U#j�ڰ;�쒕w���4	��U̥�A��FD̾i�)�	W��5CoY����o�A�`M�ߓ4����k��n
+�u���L^��|��r�f��e��ҍ�R8���7MᦔQ��ऀ]�.�.�٪�/��3�Vk���H�c6+.k�3�_��OJ�_7���'_���pC�z�˷���������]3����z������q�64��d9���h|��֧�~6�_>N��>d�yu���[`�a��#������a
N�7�1?H���c��������?�����?ܻ{?���GA�h�i��E�9�^���D�)�^h���O�=A�LΆf�X�Zt�j�	d
��K�Y5�3�@8~1�b��`����V̈k[x��c+%��FI����#�w�>�8;��t&Y�����,�����7su��\)2�	�  @ IDATx~+��ga�� gp:��������(����'�>=�46NA;�Aa�^\�,_N�೦�'����~:P�5$:!g�[i��Yڟ呕�����Q�K�V��F$̴����?&�3��r���N�D��q��^�4�
��Y{.���SY�^	���1OO�j�2y�z��݇՝�s՛���f'V�c�ExP<���0����j�Ү �f|Q=��c���M�f����a����,.��2�6���߼Y݈/Ə��6���������$���12PVm�cc����R/�l7����.VmJŞ<z��Ǉ�~����?�?f�©w�5�T�叔��D�������x+���46�hr�B~^��,s��It��J���/��w}�ū�x߾����һg=�����+�f�����;��p˧4�}�HKm˼�H�����N�݉�|�&���A4�L����-Z��4�"�����w�}$${۹@����*�qɕ�d���H�������~_�[a�6��/PZ���߳�Nn�g���q�Iʜ���c#�q�ӱ~�Zw�r�����|���g�ۻ���jr��۩���m�Ú�E�/㮄�8~��½ԫ�N��8�|=kW{��)�EVjwr:�ζ�)Aq���e�X�&�-8�/HU�#8�Q�Љ�u`�R���M�0�	G����e���/
���*�.sx��u��sY���Le�i��D9a	�|q��\��()X�&��bC��˗�'4��	{V�&Ew� �f��Or��,'T�F	O�y���]?����O���_��n����𭰄BTJ���欱�����Q����?K�t�_L�FV��kY�D���v>�7|�8��̴�(8�F�d��y?ڳ�x��p���ǽ��M��wa�����ǂ8)�^��{������:Y�X�j���:e ��x|2�
7Xq�S�Td���������������x^B���`����\W<wy�}?���y��~�Э%V�țoN�l%p��3�s�6�g+����!mpۖ�����{0]Ͼ��~/��,7��p|>�hɚ��ݠd��R��%�ao2�Pk��N��u~�d��@w�T���8�m G٢@<�"�U�^��)DfS�f�ǔ�+��J���=liiP�;Y������~[ϑ��_�,E�r8C��0�C��Q���㔗�Yd~��~��D�᷍$��Hfi�8ߤ�U�zՂ�o����%~^>>����h�q���dI���+�Cwe2K`��\���$��ri�^�@F��	��ӧM:(��Æ�fM[���j��EX�`Ѱ%;�����6�k:�a`���d��7���\�Lr9E����ʋ¢͡�~��Oc5�:~���NmC�)��$C��ް��@F��.�����?8�̺ym֩l��;������W���y�p��jY؜ʤ�����t.�G'y���1|��W���|���b�7�&|�"��2C��}q-���;i�<o�[e���
��e.��R�꿀p���pǰ]��:��p'NnV�w�����ެ�$u����L��À,@�
4�[��zo3&��0=}qzw�/j�t����n��yܒ_}�E��a�x~������A�RAP�*�Y6�gu��U6�`��
G�L��Xu���nt�؏齵cR.�5^_-8,5j�b1ԉfKC��y�b�U���1�o���;<7Pb��w�ߏ�@��	�7�Wa:7�hT�� ��Sq�L��H�g�F�T�{�5���Q+(A�!��J<��B�i�b��!��[�ҕ6s/�j��v�i4[
�5{,�fR65�L�~������M�}�r�)E�B�/�-����b������?;w��Ǉ%�<|�͝�/��w��_k�,`����dk����gŽx�BÝ/?|��*/�Zk���B����'94��пm�¥�8C߭���:������ޔ���V|ȳX�G9�-76��yV��=��Q��k 9��R �R3��0�'�3��_D_H��((;��y^�oKp-�;fgRϱ��y�0s;�(���eѪ��8j�v~����	β&����F��C��;7.󡔅��5y�Wҧ��R���5�q0�GX��wpΞ�-+ҳ�(��j�t&�Ͳ|]&W&����Zy����j���HgY�����N
��;?߭��|���NP��²�'��$���Ck�u��T�,:�ӝ_��0��-�z)���c,W� z�n`��b_�b��0������[�b����ƅ�u<k�SB�&n�<2)�l�NvǷ!�c�0N��
�^}���8��c�G��u�,i�^����_����]��iuh������?����yC�WS�X��Q&l+�l�	^Z��AR"Y�w>��������Z�	�);2vjzy ��5E��ݻ)�f,6�l ��� $�X�HE��w�Ͽ��m��:��o�>�*���f�lR�6�,}��%�h����ﰩ�3#^�C	���ԏ���쐶�lc�#"��vZ@=�S�G��\�k��"�u@�v<������$�E�#����$�_<OH�W�ɧ��<���HK�Q&C�B���P܄_���/��xl�������N�|
d2ч��j$�P�`z��h[@�LIp�ۓ�'Cǜl�x��+|%�_�,(s�܄�� ߞ��&��m��b�8���|t����*���M�}�%K�c�����|�9�U���W�����hih$X���#t9Q�RM�X*Zy!���Na���}�hs��<{��0_�E���Ꭹ��K O�Z �A���礴�^�y���Ύ��k��b�9T����_�0ed*Q�cm��ht���g54f:����P�_��|)��zB�e��������囆I����
?3����4�b&������-?�9ߔ��ǿ9��$�*aʴ�n����:���%�Ƈ ��[�m)a	���i� �%�EVjx�y�Ʊ����}�����������e���Ɖ'\�y��M1Q��(,e��ې�~e|*�c+�7RN�	�8A�f5�G���y�h��0]�s/W�c�Yy\�T�N�ࠎ:�r���#��}_��X�g��I!�n�G+��u과��J��
�S��C���l蕷[���
	��:g��:3��8���g��qR������93k~��,:Ū����p�k���G�¸�A�N>���c�SX��,F�V]�:�5&K�t@���z� ?I���7
�((xt�&l�%xO�e�+��(C�R���-�W>(&=@����9\
�桡M��j�yb���&�_~�Y֡����H��_Gy0��6Ys'϶���n&��L�w�MrV����s�Bn���]�X{�)�08꥘ڝgmv���{,������Y�>au@��Ɩ��ܠ/Z)������7�y��k�Ģ�-�{�0M�U0���B��;�ߞ�_�\��i�n�8����T�aY5�馍������N^hy��;�?�Ky�,x�1��~?!��p��7��?���wP���8�� �|Bk�l�����j���n[ {������)�sW��8*`E�������x��~�,M�s4�P�[䋱J�|��p�.���f�섽Bu��K|��v��5HG!9	���c�~Z|�~��c(��Z�vDO�Ƭ1+��z_�ĭ��6�M�cs�|�J��u���w��Ai_Ih�+`�>
wM�f�W)0�*�Q�k/9w��>�B�"�]��
���#Ay>����+0朆>�#��*�No^�{���}���)�ҙ�S|��T��wl���~	�.��|�b[]���6�p�i�	v�N\���
��'���I���?����Z��׆;2�?m�A�2�`��ψ$g]�P��ֈ�̔�Ӽ-�F�I��r�%��z*��+��	6� 1�,!B�����k������w�L�Gi�|�hh8jFY@�!�������og0e��_N�y�y����/�+��B�ȼ�ǣ`u	z|v6]�Rk�� �~����g���l����w����r������!�]
zV��V'������b�ő��������p��t����E�B��m�^9��3��
����Z��6�gӖ�M#��o��o�&�T[��1ez[��+))��s|yP����g�ps��#��_9){��da��=�v�?Hެ�a�fmfy�۰�?eQ�5kMÊ`��V����l]��uJ-�����rh���8���eig	��W�/��s��G���ׅsF��Ŝ)'͚�o�\���_~f��+�_Z�����٧7Y��Ѣ����:[83��a��y�0���l�lS|(Ĭ��A�e�J���4ܒU�� ]{�J���W���Q�<�uX_��`�r��!h|�R5�}�~ei���!lx�hx�b
��������ډNm3��i_Nޮ����M�L����2�d�{xz��=��m*�,��i˹����������c�N-C�}.@K����X7Qr�Y�<~��I���_=Kkt�d�,�֒<ڷ�ǆSYU�^hg��s'P9M�}�2^��c�.��}y���������\��уĴ�B�#Y0��uz%��y��(lMzR��YP
0����de�g
q�D��-���/}�a3��ұ��R�4��)`�����H�/Ĩ�b�E�>C4	�q�,�X����YCmǄ�ĸQ���pl�RC�^��p����a��'�\^��o���V��g�Ne!x����0�{_�*�"�Q�Nz�Iñ��n���Fѭ�%�}Ch�v]���As���D�r%5��Ʒ�B�ӫ��%%�����TB�a�ҷ�};����0���ǘ%{�I�`���=��2C�7)vа'����E�����Zok��*��]�H�}zކ��TY�K�x�d��	���(��ʭ�
1<,��4�B���2�ǲ�#�O�>+��/��N��8�V�`v�u@N����=`���2�?,lƂ^��t�n�O�'�ga-�4v����'�ql.�p�_�)?f�f���z���N�����1t��9���|x�<i�φ�"ܷ%]���{4=�r!����wx�.|��݁:�t�.pذw�<����pGYk���Q}�B]����X�B+�_���k-+����ʷa"Y�œ{Zn����bO'������f}��1�0�-\��k�x�j���fcÐF�޻)k��bu��`�&W))���:0�E�t�/�x�_=S���w�{��W�M��X��6V������Eio�lQ��BΔK�1Lg�1��u��8���#y�-�JZ`�hK;��E��#��[Z.�9���x@-Yg�<~;?�k��X8J��F�7�c�]�}�)�����hl��\��������5q��;Z,�b��х̊充sq͒�������U�VvCpߢ�B�U�[M���: �fDC�߽��O�/�&`EcW��!����J`�R�v�;�z;���`ւ��X�*���ԙ��[u��>�Z��n~� 4ҁ?�V�̲\����໏ӻ]��~����������O��rP\L#�����n�~ˌ�C�߼���Kux
�d���<�*�)�{^��+#���0ֵ����g1�*�Ys7��5��Y3�B(+�7�َ�n�-���e��E�X��S���zp���('�KA�k���[�J��)TJ��M�U�%�(�zN
g��d�7��c���}V-ȴ���90��l�0��$ ��rh&��W���J��.��z~܄ �W��gذ[I�q9V�^@t��򳾏/`��3d��x|`��A%iG�A5C�f��g���!�k+t>���rv&�qG�n�	އDQ�D�=^����������%Q�O @�Ǿ��M��}f���<"######����؊پ��e��հ�[c�H���0!�iD66S
��΋�*���PĜ'�m�R�QX�LO*�y/z���r����^�c�RA%ϸ����
���`$�	�|�& �C�Udy!��\����l��
� ����˂0����y����w���/���K'�m8�P����o+tQ��ǔFac�Q.nZG����U���W罕re�y�w/a���.�	�AA���ǔ�n��aMS�Ʊڙ"h�.�~7������qm|��r��Kt���Y�OÈ�O��7�o�.���J��s���noj�^�́w�l��n�m-��<ZʭZ<������~�%����݂º�r��?<b�}�Kt�y�"q�Q~���ɓ'OY1���z�0%��� ׬�,�̤x�'�_��N���ir�$����k�.e��b�3V�B���9?1}�E9�d�u����TT$7&�L�_C1>��o�Q(��}ϢLP--�������{�m@#8嗼aLcq��Λ�WeV�y$O�=��t�����=�s���ef��F����Z)N��O�<��ϰL��,"�o����oA�=����4�b�&gs~�Kۆ��,�����˜ϫ%/� �7�g��.�����ʦX�����
��~�T�݌(�ϐ�DL\�;c��f�
+%[�z�Mӫ ����(D��)߼��4}WO���K�����%�� \�D0`X�r>��/P+#?A�ߤF<�+Z��իj�^��W�}ű�(�H}�LZajҒ=�+"�aLw�E��9��3��ɤ��j2Ҩ����5��Üo|�!��䷸��_%�=�����5�_�n�y̐�+��8�{�6�j���^DWXm���*+�N�j-K�� 2�ơ+VB��K%9@ �@0�[��Vb�K�)∺����i�xI��e��*���o��Ϟ�h��6 ��d��[�k��g�����g"��l�R��)��<t�]��;�r�Χ!�C5�H\�'&�E%�!����^����N���8N,��"�s*�1��⨥̊X��*@�;Ŏ�|6���Ort�穙n5��
�e��%(a�a��9q-:H�MǰUV/����P���)˂��	�{]��_�k��L��b�_�!&QYx���dJ��;��o\�F>�ϓ�S�:�W��]��Kru�"M��u�--/��	�=���k߽�����_��Nɫ���~��j+F���4�"Wʙn��|>T�z�RԄ+;0_�a��OG����3�ˤ�΃���$���Ά5^+`����e#��t.�+��#lu}7�]����|΍����l���=��[�{@I^>1Y�x	R��%����d�mQ��
�҅zf��������N���%&�_����@y�F�*�*i�w%V6 '@���
��`�|�C�2�^���*eʡ����W�i�C�kn��.�7��$�;&��.���D������ji;y�X��^Z��2�ft��1�4�B2���஛�B��׃��K�i�s�q�E��]�����I�w���9s��'��vr����y���n��!Ɔ�}F	�Yǫ����=�?� vՁ�7�Lt�-��Яb%�ݍV�Y�����Pu�G��,lA	Z@W��9�$�T����}��O�U�š0�%�ʷ�*q�ڸ����Q�u��m�i��XO(<�ow���&:)�1$@����h�;�����P��+�I�:@ې��̢&�X�{|�@e;�Ή;��
S���('��~T��;����]>�d&a	<ʔh�h���މ{�ܸy�N*�.˨O��d��`���𴨬b9Q�s^,�2Ǣp��� c�b�w�ǻ0�K�u�O%2�oi�}����V�D�	�%N�\/��d�7L�0�����0�9v�3�Qp�h|�eέ�����Ь�V�zN�[	��T�(_%G���L����B[�k�l(a��U��..V`��J�[�x�=Fw�.*�w��YW���q���ޫ�Xi �	gզ
�K�]��p���j�J&�7Nɜ��V0�/��w/,3��2s�N	Y�
6�ƣH4��M��wo˘�^ҡ�~�9�N�q���-���?�ۧ���Oᖢ.�sD����Gi��4����`�����J�>�KNa��0l�.Vg���`�#�xY�s��?��[7���V�,��e^��v*U�i���V^��ҹC���i$���歴�o<oyM��|ɭ��P�Щ|���J���g�)��GL�Έ{���Ƚ�T:<6�Xv��?��<���kQ���a�*�-',�]
�iQ�P,ߥS����~����U� �g���쓧���+6+���M���&8�UZ7�W��`1Z�"��킣��<Y�&�<�^;m �|IS�ܯ�c͔��*x�e��t̐�
�4�<̣�uz��H�=�G��H�X�HOٓ�Iك�P��=;�Ν�B�toH���y�tU����$t�v7�{�=$u�a�T�驜��s�<��&�����I�đN��C��b�?b;��=F	�Z��KL�Yg��G�O�[��?��n��.�;g�1FlL���������1e�²��j��Gg�N,O�Snhk��S��*�P��c5�yA;���Ǧ��u�{�zy���yg��煦�y�xBf���3�X��k����++:��ԩl�8���E����D\�Φo���X
	��}}6`%U��eJ�>�%���}�Y]�z���3������_��x�p���O
���3
�����|�� g?!I>�1~�]i�8�������{,q2��N�_��H*T
 +��]�R��9'��G�h��`����������¹'*|jil���H��;�BϢc�ʄ���R2+Ct!s�rf���� ��;O雹k�@����B{R�r�6�i�|��3��U�Lx�l�Q��_�yZ %��%�fOIuRrP�	,-4��|�P����>�_,a*b�!2���p��=C��� �Ga�
�d���0�(R��_�Nhp,?79t�Q��"z �xJ<w�>��!�]%� �U�5�~s�f��J�'����W�PJ��O�!��:��?0��0��o��nx��y�l��|ŭ�G��g �w��m9��Q�����[�JE���'�΁�gxP����4�țy��f�>��mt��H�r�����_�˧���W�+� �7�a���~O������t��{�A$�aw��k>�7���g܎R�~wW�Y��0���p�1����5ia6�BH}�q�8^�R��'|i�<`��'k���ιו�ccȳQl���]��������*0n&j���r�*�ȾS�(˷~��.�t��zb��On����i��wglb���]�rCl�p6^%?5Y�F\�����u:�S>�w�� �+���:��c�j�+,Z�U���c���_؉t!�y8`(��4�#o���2���YM�Ӆ+�,.��ǣP�ΦηQ:�4zSEH#�Rȸc�B�5�<,�锇(��d�%m�x�(O��U��������"�I��U,K�Q9hZ*k��?�j�J�CĞb��c�U�G0�[�|N'�{�"�P�m��l�nd����hP�6� \m!��;<B| � ��C`��3l`�f|�\�Gc,��-�0�e)yP_VO�5�hy򓧮^]��������0"Su�V�:ʩA�kCH�
�x H�d����6�p�H,;	���o�7�8����Mџ��O�;�|�BnL&j�'���[f2O�%�Q���
��0��*A����#ٯ�^���8�w�J�+����ó��t�o+����b�� 8����#a�i��^����~��/��r�h�q�]��H�������E�F��T*�N�]�O�I_�ap�r�8���s���/��B����?��ϡ���$oZƇ���j%��p���� S=yOck8ER�$"�è�T�x������(�&'9HՇ?*�4;��9�	���*t���tmJ��_˿/�D�R����w'���f��-,�j�o�eLE(G!ll8v>��<}�t��{��E:�"����=�=�����#����6u�#�o���F@y����^;*dG�2����gy��r`vN��ѕ&%�����B5����'oZ┫,2��B<A/W���=��hX+�L�`�4�B��3��u�FY��69p��+G�t��Pg�#&��*|��I���'n ��Λ��U!3�5���/&���ˢh8~%m�W�BT�~>]��{6v^��ͷaJ�]7�n�xF'ԫq갆��C���2p�p>$q-��R"~^²���t�-�·�U�p�w=��"6P��A]Y�p��:��hy����]�OQ�ܻ���,�_id'�n�	��s䨓����ON>�Nv߿�|d.�yY��B]�{�}�W������4�nea�m���]eu4)h�q���_�H+{�ԑ�X�\���󮬛f]ˣ�Xy�Ʀ�����3\E�!��l
��{DjM����(� BDx���rfxtV�q6,�w�nT�σ�7�!���ByRђ���Nk�" ����89��0����\fQ��3�du��n9K����o�в�ێ)|h~s��*|N̷�*��	9����6;���c�B���&���\W�l�)���D)�6�hV�R��b{�	h�� �<*�=|�h�ʸ�v�{�nr��
k�8��N�J�r\V�Ŗ�N�{nyl�<[�m�_�L�˦&O=x�����'�G�����8T2��!�
���D����-��%ec���o�\���C�|'��}�2<��Bb�@6#a
XF�d�4�0;e9�dޓ�2�B
�h�`�Jk���$�}'��|`�4wE �=𵠻 �� �T&}�" �04�ۧ��ׯ_�>��nE���C�r.�L��h`͐&٘�ɳ{���a"� ����$~�7	b�`p��
+�ᢙTt/�� ���,��>��R��]�'do��2�C�K�f,�z�O$�Ƃ�J�Q��8׍R Ut�Ţ���S �M��s�Yp���4��6��c��ζ읋E����GWL���x����Ә�����^�bӀ�"t�{�H�1L� ��t��|;�OK�k�@Z>���` �}� �a���:�)n�f��onO�� �����[����{�F�l��l�w�PEh�P�!CTs����4C	��+t5x�)���p���5�V��K �?Jv��g��4�FVA�yx��3�
3٪t�k����P����ǗO�J�T�T8Pʅ�������
P�J&9���5.>����633����p���޾�?>[�R�w�+u�p6��k8��4T�Z	�4R/�DS'[��y�ȶ����I@�r�W������t\~��'V�ߦ�î�lŢ�
���6��J�1Է�m��0RX��!�sW)��Px���?��]��١�
��v�';tt�>�D9r���k�K�9��I���F\J�f�U}�l�`u�c��q��v,�[X�����ؠ���*O�(UF<
�wzK]��egi���ޱy�	v�_>�z��)�2�:���2yJ�������q�!G-r6�*%˔����W�S\��D�@?Ş�K1�K�"���8��gZ��K泂������y������\e����2�����z
_&��9w�w˝�D�N��,��ic�Ë�=8�	8%���:_
�bOI�H�K�P����י�a�v�m'r�|a�0,%勍	P$�C �&�p,�؀R����$�}&�;��!�(`�eS1�vNe2y�(��h� h�$��P�%��/eU�#)'/��s����!�/��lt��ixS�p@<������s�*c�E���f�$Ñft�jj�426�����"�$3�g M����W��VS��T�(�!s`XO�/�}*�'�?�ܿ���%�-rt�)�q���]��&P�rkU��n�+0��6/��/%�\J8+a5)+44�'���i��1O��+0��� J�$nl�x�1x��ɹL`>yZ����V�SY�/I|v5�`V���T�,Ky�+��t�z�M���*]���y�9��)}t���'��I�$�<��*Dy�?���]��
�_�g#(�-�<�'�|��/�d��s3��=d-����	�Lf�I�_����L4�S`*`i\�WH��W�\g�����'
���j=C�ѣ�ˤb`*�ȹ��g��%��T��U-y�I?ʛ�Po:�X��{��AڔO���ԩ+���o��5��w�?�c&����VX��/�Bk��0�W�3�v�H6�2�^~#=#����g�3�	��L0ˍ�M�L|�<{�}�"�����W�6ĥ ����jZ��|Z˿���+S�-�]�So�(�U���o����u\����̯,fZ�׆����C�)f*r��F�\l֩�b�ۗ�����F7���<�;(_?�����#�w
wpp�a����-�����R?���66�¡�B+�%|��2������_0~}�|��m�O�y�!>�s!Խ{��[�Y��
Ie�5�-U,VQ��L^�"�>M󔣉�}�I�w�c�3�S�y�',ߟ>�a�����`!�Q���	C{�����=���o2��������s󖍷JL�r�=�*ݶ��[Γ����>���`h���oװ�����5L���K�r�$�zeCI�\x_�fG4xP��;�QЪ�^�J���:�29���a{�\yx�)2M��Z
F���Kq$�o��܆������He �f�������H��S~�+�f����VC�,dz��5
ބE��	��o8�����׮?N;By��/��D%��П���<���Ė�1�C�,�� _�ީ������4���
ڼ���$��7E[,�g%kJaC�!]u�$n��EZ�*��[)`�ʇq��f@�ZӍ�?[� s9�-��Ũj�C�Ԥ	i��0Ӕ
����?#�N$]��=�f�{)��*Q���Гt�xV&�W��7�+�Uk��*�J���٫�=<��yG�{�f{�e�'���N�g�����M�����j��m�,l�R)Y^k�=�G�+�wށ�?��U*$+�����^�T��� fE^� 0y���w���/+�� S�;�4�1�(��gv%�0�N��7��{��� @��J��!�O��V��o������� ����twѡ9'冁�B�|V7��f�#'���s7e炸����8�a�[�mr�/�R(�({b����i�w��>�no_��b�
�����J�p�i�L+��en2�y�t�ܻ��{�[ehұ�e�=���ΙA�C��K:Il�n�"���x�g9̮*}䯟U7g������oާ\3��N�i:v�K(��������G��A�����}�%�d����n~���T� r�%�BΨ��Q�a#���_��������n��dC��h uk��^�?��E��2�8{��O����5k�`8iSq+�ٻ߳�$��[x���h��37��6��`�:�#��g��@������	��ʜQ��n�Zz�����M&��+��g_�),eh��ЕͭX�D��숡1:ӳn:�㜉��L�wҺs�<��yAZ�0o�:�^��t��yh�]�鈹X��7$̿���	�P9�����l��p�f���@Y�F�E��
/���5�8e�sͮЙ��'���P�B���s.keh)�%_G��I'�0u��=��/yD����� �V(i��(�JU�Ǻ�lޤ+�8TA(�.�B�M�LE� ���y඲�x�9t���ǭ�2��2w�~ɜ��҈���㠠�e��m=��x���m��y�Lb��P�[�%Z���+�����,x�b���?D��v��zNݰ�D�P^y�(�|"�U,W��'ϫ�$M	#nMK`��&*�*_'�y�m�|���
m
��T�����]U/�	����R^�VPv��QO�;��I�_��MH�z��2�����WY�ی�$��X���;�[G�H�R9W�����"�q��%{�8��
x�:+3��f"�Y:�0��P(�ʧ�!���^��*2ɚgV2��;�ڠ{2�3wTg%��3�9e�2-`?.�^�����ke�9�9���v�?~� "��\�V�X�b�H��j|�J�u!�D�
A9)͚��+�_�:
���ˤV2�s0�V0����x��4:³r	���[�Hi�b����뻌l`�I��t�|�'|+�_Z��2�t:>Oa�
f�$L��p���k�
i����.�&[\۟l�C��a�4J�g(ǻ�ֵ�}�������Ϊ��P9ܬ��/��A�>��Ƅ�� ��P�<���M��t��@�=�bM�X���pɺ{I�s�ÊQ�76�'�ԏ���(d�7�� V1�A�2��VRR�^���JE�<����f�_e�24�>����S6zX��?�Jڤk�ʗ�0HM!n�&�Ʊ܀G��kZ#�O.S�i���0=_�˴�g��R���;P��i���k#�啺2�*,�U��c/��\,ݍc�Vr:L�i�I��u���^d�,E���iY+]���{%c�O��,X�<*��#`��eL%�p�W�W����� +k��|'�6.��\Y�l,�HЏ2a\�h>Tl����KW����j6'����v>�� [\Xw������{��ɪ
�h?���\�bC�P��ə���z�=:>�鈕��1Re'�;�g9��Q� >>�p^��`�k�.V�#d`ؑ��k���`�g���]8S+�:�
u֡�(�`'�ao��r�0�Q�hKj[D�ʘ�"��"��
����ߠ�ék�#������!�)[&K'�@�IQ�`9���6��
��D� �
��1�yb��)v /����8����R�}|�c�b��@�1T�z.�%/�r)�*�n�M{	%p�U��4��:�t:E~/��������~j�?��w�����nd~��Y�{�� ��
���� �*״��[?��pn�s�Bv�U�(`��2u�`�q �تc�le�L�O}��$p�\�E�3�DO��i'���a��a���]��5VX�o'�X�
�  p�L��]������h߄7ƍ�)�B��0B��b�?���,� �$��A����A� �C��'��X�~V�j~ q�X�O:� e�M���;p���c���@��c�S�p���4������^@0�(��V&PҠ.c�>� �}�Jf��dn�&
�>�kES1��JV��<���"�Ai,x�a>>Z�93�����2�W��O��q�Tz{q+�3aV���$܀m�m1�e&3V�	�q[敔��yB���=뷞�{`��`�ږ�R��M�"�(�cfOr�UVN�ux`���n�7�H�����!��!+�8k�t��o)WC	۳�vP��2���Uz���t��An��"��
�b/O�0�����p���%a��4��z�c��	��?dU���|o���MC������(y��O��<}��������UPfdv�.�^]��%�*o��^F?W|69�@�ɻx�\�����q=�o���t�Oi�v&����`J��#^���8N��\Z3�zk+��m�m>�YܦU)����ز��[��p��L�j�JX��������`ަ�Rz�G]�f��Ȃx���s�~3�xU�TŦ��W[[7���*���`a�3���A�*-�0Tj�������q�:��$� ]ȩSw>�/TE��[�G澋J:-Q�.�f�
D�Wo���fg���H<+3gy������MV�;�6@,Th�u�lq��w�w�{���<���T�A{�>Q���Gޡ�>y�$���a�2Ľ=�h9v�:{q�Y��g����8�X�Tu��4�"�f�D\���XF*��R�(w\��P��Wr��>��
��uѐJGtH�`�.�|;b8P�k�w���(�o�ud��?�2����A�ǲ�z!-�w6���|!2
��3�GɃ�����-������R�Ik�����S���EV��t�(/g���Yfw�R��q�K������z�M���� +�l�+���<��Z6�@t#|:��q�V��3�Ȍ������
핆��UWn� f��x��v
E��.&�6��l︶����ڣS�qҧ���q�7���`$[`�F]�`U�L¨�8Zo�F�<�b:b�^3���9-bN�\E����1��I�Nk°�YP��yƎ��f�Z�xf8��1u�܊|�I�ݻ��ߞ<c��p(  @ IDAT^�[�Ƅ��a�+�w�\�*�y>�熻sP<]^�˒�/*��H� R�
�n�K�D�)�1��}�jo[���'�L��.��Ĳ&�;�h���Mz��F��'j��� @.܀)#�3�z��ec ��K�w�������_
��{_�3�K�ڛg+����p�v�ؕ�H��*s��|�Ս?>b���ە�aa��
���q-�(aTD����;^3���ǿM^�e?"z���6�&W��Ln�=�����*��Zv5,�P@`�"��Tq��C����E�{�nޏ?FadcJh뜴VQ:_ ��
��Y��^�&��/q�'��S Ўr�2�'n����R/���v��܏eڗ8�#��w��iZ���s~
��:^租�F�w�����;��2�����s珧�xVYÓ�v�(�eUh�Ip/��}��[�U�Ώ�p�e�h6����F�Ռm��Ҥ�K��W��i4,��Kw�~H�;nhI�+k�s��/��Y�-By�&h�Ǳ����<��kC�������["sh�A���{&��o1��s��qy���:%^*:��;wJ�ҁ16R�(�]C��=6���r!�m��4�:O-��В,��E%�s�p0sɻx����(�DrA�e��?���?�Fg�C䶖�k[��ġ��){�g{�2dw/�OZ�~x6���Y����r����۷��~�9ُ�!W�͑J�G��1>�6Z�,Sٖ�o� r��� �u�Ӽ|$�J���>2��|�k}���槱eٸץG�c�i6s�a�c��0:\�R(��/^L~{���
�Y)c�M�$�E~�pd�2�5m�
��n�������F�h�R��By:�8�a���9��)�<e!�F��M �d���{�_�K;$ϻǻ���+�G.2�&��af�G^��dV뗼�tG]"K)��YZs�l�e岰����u��&��,�����������9z��y����qJ��!���#DV9�1yAӱrF�JL�ΙBaS��|hY��F
V�������^ y��<5��,J�®� �D��Q���V>͈��$fDS��`N�s��ֹ�gv����RVGR���S�J[�p���7�w9K����ѻX,.�v]��:���P��֨P�X�V�-���gV�P1�`��Sѣ�<_�-E��6�ش;ܹ��[]Ā���aI:ٵX���H2���aA��)� ��|҈S���!N�����2�bP�`eN��O�m�e�A�|+���jF�k��7 �^u�-�����d������ �:�m
n Vڼ����phR˧
�x��Ff������� m��heL������iun����0��>G`EA �'4
��=ZE����6��_���bFA%�E���'�|��+��LW}e@*JC���N}��L�V�Y�
_�ipH�6I���(J8]f���t柺{u�����\��t(C�R�A�N:�8��J�	���W��qh���x�^W�y��)m�F�����V�����ʗi(wT(:�~������*^���c4&�����.�XBҨ��Y<<���*Q
��
���&
�&S@���Z��#��ƕ����E�Պ�p�v}���C�40X�D�S'����=�(���0{��PpN��w#&�����*����;>e����ƗR���:�yf.�Q1���!�R�'3��p*G~�����M~��	���$�I7��v5<�I�/� ���'펖�X�1��K�������#������-Gi�<�]�O��lǰ���U�-Wk����2]���	�y��o-/��W�X���"�3�_��W,��p��w�U*J�(���c�4l8�*������=0�JSҘ[��wR�dS
�O�"Yn�%��l�|�� �2sd�Q�_p<����}��:ܨٓ;��O�m��s�j�#1����Sٗu������n�.;���p��"���
c�ɹ!��ω�H���c� /��� Yb)pѠ�a���m���2zs�E]�{�<��$;�`�1#�'*� ���uij&�[IRQD���/�L�K� �-1$����(a}����($^Wa�c�35�:���3���� �*f�!���� �
�̞M�̗�׆]�Z�X����P������o��/�M>!ղ�!a8�jݞ��z�X�����h�B7A*�V	���e��Y����7�w_*��x1}���K�,�r���⻔ 5�-9���m����D�Ø��
i%�� !��N�bd��^��b!��)����*�������M�)*6 ��P��z}�ǩ�<���0��L��� �
�dY�OcL�W���a�gj���aP�S�:B-��(i��9�yʖ~��/�)�v��W���p��V�s)Z
o{����Fr˷^�Y�<s�4��򐬌K841��oiHn� �)|K�*���������([>�����פl]���>��W��4�{�THp����-o�<�M��+��7LgXm��q�F	A.��W+>~��y�~�����^��<,�̈́�e�S�M�������V;㉏~�d�R�����g�n�ѧ��
�����ehޫ����_�i���z���]u�IG�r?�p.�i���U�w���G"�d�m������Ml�
�)��r�<��`Ag�$_ԧS�&�tK���d�]��9_7�8��I�����i;�ί�	����L=����	�z�ܷndB7B{����xx�1�~]�W�[>q�@��)�	����6U��T����;eW�X�����g�5��W�˘|p
�߼I�ʳC��]����^��ڍ*(J��C���(n��0n��o���,�x��c(,/�N��>��v��Qڎ���5��U��}����l�a��U�3)U�ͷm��Ϥ���޵s)ye4�<�W��0�i���X�.hcl�	�����P�KF"�P��0geSE�p�N��38�lys9��^�.D�R"��1�	�����q̶]QʬN�Q�2��V&�F~�7�&eۤ����؄�҆جg���:��1��liD��)��&��YB��`�T&+�h��.J$b/RB�G�,bj[RЃ��he��bFf���Ț?�-���W���	�F*N�!�k2���G��f|N��.�2�	S��ǧ�5߽Ĵ�#�3%A&�����關���ɳ�㧯��Ȝ/�/�ã�#<9~a�I~�"�E)(���,����2�)
J�|y�*���d�h)���3�D��w�=|�k%�r0����4?��h�/�8����x��峅zz0J�8�`I�
5��4d��o��h�<�$x�:/Č�O��=�|�ŗ�S�<k�:O� ,L�h�<����۠p_BߢUѬ��8�7I��ĥ���-����[N�w�UW���C�o�r�-�K���eނg�=}�|�ɿ�tbN��·+�]��F5M��� ZA%��TY�t���{��0�7�B%���y�i��.�r+8��t���I�4c�����?Ҵ�e_:��`�{�ӽ�~���8�7M���<n���÷<���RVh�3�P�K�sM&�����.�|z�`4���i���5>��_~��袿���*�V�ڽ㚮����3�v���a',/�{5���J��a��
礋���;��k��\����o�x$�J��"��xR�C�@L��� �3�����T)�f���-,J7���Y%N_e�0[�c:9;Է�__�fn��g%�3,�;XeT�,��P�5�ΒC�',��{�)6������ϞM޼}E�)"�W�)-:Z�=��y��(te%e��!���u�4�;3U뗊�a������;�X2��ѭ/l�U�̃i(w,��7��é�(�Խ�TU�c�V�)cK	��^c~��0�5O�MB�0p��C�* �W�S2���J��P�gn3���1{�iQ;G�/9�L����Ox@��r�[�m�m�����6�*Iy�G���j	%���J*���j/�/<�B7�%��v^��s��na���ܞ.��h��y��ŧ|�Hک��L؎���|����߅��{�D�P>ó?RF�@��'9T0T�4\(����Gxe7#+�����.+痝'�H%^`i�
��@� �����T�炐�d�P�Î�Q 5-_A��&�)�zӁ�䎲��l:*ZV�̉�4Y��8\T󫍭�Z�'#�Z٦U�����7����R��S�)#ib�G������_�:y�{&\Ҩ��;����4KĊG/���4����	C���%Ҭ�I4�P��Qq�.2�����N2C�A�Hb�K�K�z�ɞ#�a����6+�W �x_�9���O��ƅ�>�T�J[�C����-��R�(�f^G8�7.�TÔc�-���:O�QAC�Y1�}��U���@���'�׿��g'Tm�A���rۛ�ؿB|���s?�;�8O�z㐶�"��Q^.��W+�����$�4|F`�c�3si�
��U����7`�2(�y���U��k��E�aSX��aX�'=�@���uQ���T�/��9f����ٴ��%��4��w��/^�}7?T�R�<?3|f8N��5N�Æ��n�*V�Re�2��v**}u]�ؕy��S���~{��m8>�|�����-�V����J�0[���k��G@��86�i�����m��1��꫞���m��v�T���M�za�pJ_��
[���嬊�s��6"���<�4���M�-w׷ZO]y����[Z�_�|��Kq��U�X�~_e���V('�ߤ#t�yj�RdUp��WNWPArh,ǅ%�<?3�ǎ��V/yJ���������9�L?��Z��n`��H���p ���2�;�� ���9D*����b[V��le��2�I����<7J�`ME��R�L�Z%�:0���/���4V(�*眓�N���AN�gԹ��ͩL�{�6y{4��������4���.�+�h`8'i�js���o9(�0Q�����<8��0P�N���9�s,����*v��O�J=�&��8'���K������?�?�������{�Fx^CH,�Z���"Ǧ�NF���rLJ�qֲ*=͒�b�dZ�yV��V.B�=�2��R7����θ�_��<9ԫ�-��w�h�~���;K�ߣ;,��{�p����bD�a<�����ahM�*"K$lAY�u�_�$��i��5�E����CbS���J���6K�a*ͅVJY�%�nLWK]��U1+�{&��((���������-�]�>{9����A�R)`&�o���aò~�F���6�T.�Sa�B�����S�
6�zYYLW���$Y>�-A���&����u ��Z`�3N����4��#����s�	-�Dˏ�eJ>�X%���j��cQ�a��L:��x��%���nJ�>�*��\J�|Hy�|T���ۯ�{ ���Q)s�K��*V6H��Ge�孛eb�+�� a�2m�/{�5���^��ثV	;b����'(�;�%U��g���?��A�<�̬��V%�z��y��I��6B�W�j]���r^4�?)�|��U�.}ķ��9݄M�Jl��\� ^��n�ICO��,�����ɏ|m�.���n��Z���+:�����г��|�l�M�����\	U]*Ư��PD����5|c�j��?|6>�r�wZ��z���߭X�#��F�a>�7l�4.�\ʸ�Ư:z�tP��&�MIU^,R�q�'y���O�SF�O,�«�_��"�����y4�a�r �W8)��o�����l=S>�;νT�n�������U��7�nt��N�W���c�������T0ٛ����#�3�����#(=<+M����.�-��/�Y}��l��-�}7���L�wT��Q��Eǽ{4��]k��d`�ԁ�k�ISփ��̡`���`Z�TX����y	k�2���_�;Fny;m�*'\c��M�e%�a<�۬(ߴ�{�s�.QR�ky�C��aA�6����M������Mn�	�	�:�>a`p1��n渒Wq�I���,u�R_�-��i�����)�!��H�se1m�y��_ܘwm{D��j�c��O�G�:��p�M
�,nnع�mX�̫e��٤ ��f޴I�h���^,򑧏Ѫ�<�V��/y�V3��ߊ��@ k�~e�O���϶E�e���F��8��Wr���ׯ���� �!�!��;C�֭{�t/��Uz��7T�A��3jahf�2�K
�ރ�&�;.j��k$kࢰ�/��^@t?,:*��o!f>��H;�*.�.������m��_�|;y����9CKoP�>|t�-�Ι��j+���Qk�	���n4�*���<�)4�t�S`��౽�-^
�g\y���צRi�
נ�7�?_���{}��Jb�T6�w�*(E�����r'��8�$ 0m0�
X���_3o���c�J [����op�C��c����5pN+��"�4���S�(�(V������O� ��{3Փ&��`�? �f��\"ބ]xN�K���7o�s��d�f
|��`t�0��~��#��1�_��L�|ˋ������#�SpWSXF�aEտ�l/��"r��﹄#M�5O���}vh'�*�I2�޴�k�
�)̤� �'����W�5	�K��U��2������0L���Э�J��o7����t>�U��@7��#ʊVv����_�WڕH�ğKy��Yx�i	��J�4�0?�^C�_�T��ڿ�Ge�a��Bb�糧�y5��+/��߱�G��/���i�����6�
�S��C����q���H�4�g�RN���1p�s�=�*Y?�8�Q��G;5������*�2ꡬquS�q��Y�X9��Ў/�ЎH(�<��Uh���[��^[�����(n�a���� �@���<�
'=L�!�Cb�ʦ�	'#3�-W��|��{�S����O>��V��k�AkTћr!ҷFN�W�e�-�Ӟ<{J<&f#�<�1rya�;��}�E�-� o2�y�=�\D �3,O��ͩ�R�2���`�n�y�ese�j�o�?���K:���S�(Mb��|DNC���\�NQ��4���@���1u<��/*�.иd��6cò��K :�x,!k�d�=;۞	�ϩ����ٓW����{��c�ݛ7�b�t3l��.` �?@eǺX@� �OVX�!w���}�u˝'}�^Y?���dc�]]T�̡��GF�J�`�|��#�ې8?��1�(e��[��g���k��^����� �+L���JC ²��Qo�N�
?�7���T0�6��W�ʕՀxh�~geyy�/ʊ�K
�cY��$<��W+>�XX%�X��h�X����F�Pd���o�c�r���.����E�0X�,K�E,~.��x�Ƙc�IQ�+��W&u���g�ٚ���0��oV�feiS8Q�bۥ˻��׏/\8U���-s	�s��	z����8F�U�*S
��߂_�K$#J_�I�~q�R>_,��\��n�������������Ȧ P��VHe�~�+o�c�'\�o$�k%-����pr��ޞ�#+�LS'��O�:X��@��=ϰ_0t}�nߔ��l����o��X���i��a�8-{i`D��&��ĭ��KoNy7O)k����栍o\���j��]�7@E�	<Ǵwp��!�}Ϳ��y�]5n)�ԥ�|�����`�yP0^)�����[�[F��E������}/x�i�ÙF|	�����_��g��a�m��k�W�'@m���(e��W��*�y#�A���4�~��<���N�uY�+��!H��L�i�=[�Ȱ�tB��~ZO�>���������	h�Ȇ_� o�U �]����8g�a����4▍=Q�̃{-ma!������Q ��E���e���PT��:;%ALk�
��:/J�ICi��M�س�̟��]�-��X�\q]�hw�̍��Mn����5d���ӧ(�X�����[Љ�*wI4�|"�N�����I*iQ�p�>V��V!��Nr$ Z8Lɔ�UV�k1\pu$tvj�{F�<}�Ԝ�(�(���4��K�b��e������6Że�_xCz���K�Pjc��U7��ft!
�Dſ�S�tg�/(�.�p����t-��M6Ig���0��"��'�΂�^B4���~�+�+��.Xv���5:9���3f��u�;8�rq��Ա3^&���|�hP��'���DGA}�iMNm��,&�4|qbO p�
��&(���T�MYbnS��@`�?D58�S��:��Rs[w�]��;��p�YP�6���xbe�'o�矉����a��",(2j�5Q;���ܩY�ƫ��Y��!�X��I��C�*^3�|Qq�f]��+�g��X�X�G+�^���F{~��'�������w6'xxsre�Z�N
P��BSFm��:,!<i=ƕ<�} t+�ٻ����O�� �M*Zx�v|��HN&�r����"IU��?+��dx�;�`�Ц���05�;�(T�[?�;X9LWӱl�b�5�x68���ݯ1�/\��q�L��.n��h@|%$4I�RO���Z��0�;�ZFZR��2�o͇s�6�(eN�M�G%0C�/���a7C<��%���!��B�IY5��
^p 6�
o_���A�E��]����F8�*6~D��1���O��F_�:����܌g�^�^�|7��S�	4Ż��_
��o�g��s�7�v�~v���e�"���a}��%�v�A��;�C�3��G�e��򚺄�������cƫ���Ѹ��eܾگ��[҃
陏��Ȥ��=&�~��$���`��x-�xH7��6����3�i�h�3ٚ�+Okr��![ dc�kU��ZFI��������eK��Ǵ�#|눲�����V��-�h�o�yO¦�3Uf)+�<�ᵟ=��`�O����=7��D�ve�Uꔸ���\,�m��А�$��߭��GJ��TRh�T
��W��m���^h-ӗo=oVe�FZK��!�m��U��b�o�.�s�++��oq���w:��v��2c��@�4Sv���bO����ߒ}8��<U�Qi��P܄��o�'/0P����*#^�(YZ�����=u�|8��X������j	;c�t��k,n@A���:�r����:��E:�o�]�X�y� �X&Xd	�d����W�����Ï�#�;�D9T�!�/��mX�/�pY{�*��E.
��=�n�S��GYe4Hb���wyeu� �l�'�����y��g[� �&4Wn3ُպ,���0�@bj�rb���S`�d�N6�ي7�"2C�v�����aA9a����D�2(a�g�p%,�4��;Q����8�~�>���|�i��D#��IS�[N,16���iv�9o2�1�;����|��RdVV҇Y<���i�1�.�^�<�͞Q�[e�x��X��Z���P9�W�-�W�we��& P�a��5�]i	�⎆玡���_� 3z&d�^���2<�p�@/�A��s?�4�D>S���w$�>-}n?M?�!��>����D*�$o���3�i�c����S�U@Xړ��}sgcO@�9Y��19��|<���Ҫ�X������H��iH���y���O����1.��,6�۷R�����2=^�C��w�����e�]e�PE�����~�G�0>�ֿ�}7^�z�-�Bs�(к���hX��1F�����׫a�����t�eg�����@�8U��W��*�\�7�W���p�*yJ z���U৳d�`}L)�T#�ʙH��¯�W
�2�sR�\P�h�1�F��f�o�<����!wb|�����K�<e�-�Zgx(�2��H�Ќ�rҶ�5��7���PF�@�����-�r<q��2=!-�� �ݬ[��UFk�PJ^Sz;TKO���O뎍W�>�l�R�zT�UY|H�l�Eu˹7n4�	]6�$��L�
�,T��K��;i+b�m'�r9g� V<Z�}�<��yl�k��B�A�⾎�̹f{�.ݝ�Q�d���͊s�o��%��⴯��J�h�4J��}|��A�ٷl�=�(w7I�D�:OX�EvBC<�6I�h4���8|�{�)�$�}��Ӆ���u	�E�P�U/��ʿ*����Z�ՊȤ�6�}°Н�c��y��oĩ�M���#&��jQGN@�i��ֵ�F�\�&�S�&����.��
Y�*E��J�����
W�x�Q6n�a�����BZT�-8ӓZ�����O�[��ZqĈ��%�=�[xTݖ�ͪ�q�+C�bn�B$pz:�a������fZ��`d�t��\�Z%j�������	��oD�e�=_��R�M�j��
���Q0�rJ��r&W*�=4����T�/Q`h�V�
K��%Ll%����=(�o�rWhͮ���MP�����2�B`�����b:^���FF��']�{��2����B����e�ēYɛe  n�rS[V��=�d-�$g���^��}�	;~�Vf��?��ި�hG�4�� ���T�A>aW=]�U����r��U��sr�q�/]��0c7OD����N�^���G?<�ˤP�2���jLWf�)czt�i�)�/��^�x+�@��J�z�r���ZE/I�e�e`�*Ǌk}J>���o��&�I'_F����ea$L��K]�F7���F և�0�W�����&^����[�!�	G�/0�u8�~7,a��nZ���o�{ux�ۯ��[9�-����G'����V��d�n�����-��޸��9*�����Ze+����r��+�m��3J�B��9^|�mD<.����F�LH��/�8OI��V;I��e���Z�O�Ç�ɣG�T�Fg��'�X*��1��vv��rW�!o�ogڡ1i���'Up�+s�����_V��̰�T`\���:bՅQ��?p�|2�'�J7��7s����S+�A�	���?�̜a�T�M����>e79|��;�Ca��v�����PF9_��2��m����*���7�s����9���(����=oVY%y��F����{e���
eR�5}V(Y'_�fd˥��]:a����1;��q@��ݚ,���&����GQ�;��vB9�T
.1�\:�r[�;)Io�I�����m@�I�O�r��U�Q�� B��$m.lc	O`MN�3,� h����"��PI�!n)��%+��i�c�X���;ʎ��N�;b%^�iE�8�o���P�I1�� k,ZFv޵��SZ�����Z��ڹ����	��"��2"PQ4�jˇL2>�r���;�0S� � �9]������O)��nΩ)�e�!�BnZL� �b�#�2�M(�h A������Y��C��QKC�9:��g]��\B�rr��r�!��a�T`�����CM��G>4�Zq͛w$Ѣ�x��Z�'�k\ޱ�ʫ��X*Rx>�4�R¦��
2A ���L�a�M�R+��0�t0�Ἄ_0J�����I�ʆ�,�(p̏~��t��/LÄ�|�{�	ůhPU<���|��U̪�� U|݅U�bѠ�(�D��*�j)�u>����HYZ�,�%�ޗ�a(��
����ۻ7)R�R���͐�;�7;���3*iTܜ\�Er�Ϡ� ߍ!`)+xh&�ӛJ��cY�ws���(�.(�[�J�xE���H�h^t����7l_Ӳj��s��@d޽���������O��{Z�)�9_����^<l�~χխ/�;N?�kw�uo?q��`�Y��i��8�խ,�ǳ�6��w�u\{��uq�y��ƣ抡����:@�1�q��怂e��3�$�R�B������u%�I��{0�n3_ȕ�쟅���ݍ��]|�.ei)����D�M��XEZgD;Xn������f;���8����W,��x ��X/<���XZخ��r�y@��l-���o�M�g�!=&n��"r��7�Ñ�i���?�:��+�̦��7,x���\���������E(gW�V��~)�LV:؞e��I�N��(��%��JOw��Ӷ�6HeU��:Dy/��_B0��r����9���t����1��w�_���[#�ƕ�(��{�]�m��w�,J��(��Q�C~x��*���6��Q�r�_���%b�|��hX��@���C �Ӗ"Kq�=���S~$�m�`��|U�>�g�B����´n��c�D�+�m����:�C��-�"����ᫎ�`��<H�o~�+\�?Ƴ[��xR�rʓwr�|w�SA������F
=�@�
��P�$��c��
~�����n�> �Vb)��ef��L��n�	�
�"�c��|�w
��i�l	��R��0��U��%�Qq�#=٥B/����ͭ�%8�|/w�_��,�Â�ͬt<��O2��a%�ְ�0�� ��U�<x����$����)P�և�U�V�3��W2�w�������;fI<�-Z�^�V* ��fx/�e�����k����{3eдl�q7 V��|4��g�Z�����H�3�U��E���ޤt�QB����|�BRy���%��<��)����;��F� !��pw�sV�,#�Uj<���L�Xc%�����9��v
�
#x�~i�=�����Q��L�1�NzJ)���W�vӱh�b��<�0�<x�kf�!���tWq�:���~�+<a{��0�޳���p�p}G>/���{�_���0��;�gx��|�_��S��U��k8�޸X�"��>\�m>�v�Ooi�e����NG�����{[_;|��qS�r��4�/�V�M_�e.f���*4v\U`R�M2�(OKŸ���T��#�*_��W�ׯ_��f��� @��dbO�p�]�{�X�i#P�h ҩK=��>��rt��C��3�)��RssU�Uk�
�\�bi�YTA�MPQ���]�>��m$@?��Kl1��:C��9�3Cso���y�O��,d'��wnL~��a��V	9x�b��91�������g":q^�[�]H��y���-����*jT�dY7��m���͞m���X1x�<����8��X~�!�����uFm<ڈ���"�?���x���d?K;uZ����m<����s5!�2}����u���㐰\R���|�#���w+��z��96*c� s(��]�R����T����Fƣ�J�t@�H�gD���w�=�qM-��o����V��״�K�T%�p���a[,K���,:� �t���qS_U����k�nHe�X�Ι��ǃ��m�.��!�?��vF�S��=V?�U5p{�wtޗ���2�0���-R��jc(A�2$LgO������X���+HY� T�(_0_���p���~��Hl/�f\�4¸

��=�F0<��\Ǎu���׆�4�0�?��m㍕ޅ�5L�N���.�B�3\�wb_8-^<�_ �~�< L���M���`e��w�o��H����;�u��(���0��m����CG3��*�x�w�7�+,i�m+8�q��a�z�/�X�eO�����n��0��+~�I��_P*��H��)Pt�L��N�J��%������a��ƥ�P8�H7�=q0y��Q����i�.�v�F�p����wƉ�;1d��f�[X��)(z���qI�(`���R�i��E�r��
/qB���I�m=��X۸Y��׆�xQ4Nؔ��s	��5=�Ǥ����5�oZ�g����U���K�}���4��p����B��Ȏ،[(��O˶�7�^`�ѝ
c|yux��.���i?y�� !��[��-|�[����p��2n%��Q�Ϝ���T�J	�����pM�-N<�,�Fs~�Ő�]6!U�z�����٘�m�C�טc�5�	Ӯ"�=iPg��J������� �����L�^�~�m��`w��F�9g�P�Zo�P�T.m���ez�,��i���X<f���3�6ω�H�Ϙ�,�iR?��\ö*��/:,<~�C���٩+QbU(C-J��i4��ў�K&Ż�{lE�A�_%��%�BH��Z���N���5U��X0r��,����S�q��8>���%啓˕�Z����E�ds�>�I6�ժ��|(�N2�U,�lT{�i���1����	�OΘ���&|F@2ej��
�v�w�:�zSz����u�
��jd<�:�OlcɼC�*�Z�l��T��,��"���FhJ�������� �Vx�+��O�<��5����r�R���{�~��pj\K�㛲0�`���A �6�w�K���@/�n��g-;�~�Y̭!N)0����>I�@��1C�c�T�V0U
�BT�6S����63u���\�D������|�A!���hl"&n����d�Vb�0dփ�U�djͯQ2(�4�V�K���%C܂�f{��4��.I�g�1�W!���{��H�5}l{� 9p
��f��$L�.�rx��!]�s���?��,4�+ص�I��>C�>eDa7�H8��x�a`�]�s1�x�@���+t��]a}�>
�����/:�Q�md�xǿ`������yu��C<)�@�J#ƻad�����[=6
����~B��=�gI#i���K�7'�=�a���c���H��o��NJ����\�8���P��/���&`y�˯��L/��_���0�@P��<�����4+�S�E�(�����M��k���k�e�eztK+qE��a>�L����Ċ����2!���������A|y���`gh��ͫ��%h�G���fPp祟�/8�-�O^�q# �r���p�o���
F�uS�0�)�^U~W�O㏴:M�^�f��:�����?b]HGx�1�e �F�i�����z�.9T�����!G'߻U�:礮o��R�������r�}Ҡ���P,r8�3N�2��K���I�i'X��VcUGގ�ʒV&-P����ʑ-LZ�b��o-�n�|L�\ m�</�����p�p�Lngn3C~{X}��U���w4*�U�<�BH����3┡a;�$U���x<��n����6�ho�_ [�:(:̻�3]�rx�Y��2�s���F^(g<�֓^6(�Zˑ4Q��B�Tҗ��gpQ�/�lA�kX`�� �cd��|��CF�L_�W�2�r��9�ȗ�d{(��'T�#��(/��9���`*M����8��r	H��d[	,]�SC�f5�ε���B��_�7��E��(���� ���u���3��K��#���[F�ˇ4quh���U�Tͦ�˷2Ȑ	�p�]�ҹ�.���e�/�r���8R����,�_`��?��:f�"vJ���=9<+��k��
e�-�3��I����-L�"�*�f&����\A���K�CW� D�"#fӌ�MR2�\&�H
rU�VƜU��bc�ݷ�V3�!��B��Uh�Q�b
P�[Šz����7�40A0����c�j��A�Ѵ��������4��0��Т�6����RM������z��Q�s�²��2=)���ʖD�x�<4Zj	�M�)"����4?����<Ki�4�g����]&�>x�pr�9W��K96�\�i~�{����h������/qi0yC�:!�,kPw(�eӷ���������p��l5�4ۓGE�v���u����}iz6tN�e�k*���_Qx�~j�X/�]+�MG�N�0�q�Ǐt�g�m�篂��5k�K�c8���A���a�iX�囧q���U��;w������{�ǉߜ�|�Ns�.��m4��,����58���r��;L����]X�/2��z�<��������抬E��;nw�@a�K���/<Μ�������O�W�7��_�#�G+�G��(��h�p�b�o����W�(ױ��W�8���t.� �v��%�Ǯ6W	�B}  @ IDAT�4�f1+��H^��*><��3Zۘ����֭K�+ߡ@�Ѿ���}�m�V0;��G*@�}i�ȇ���m�ӝ�����>��<�υ�5�xi��VMIh'�p�:�;��d	�$h}y��C(HU�|�2c ��¨,X��2,�:y*a�)����.b.�:Z���SX�/-힪aU�ᐴḘ�������~I��f|������s'������b�n����M����(x��e�|������(ܪE�Đ��c���o��6���gm�h!KY�D���L�t��Y��$n}��xW�s�@���ԓ0��/�(V�O�x#�8U$����I+Z!n�=��x|@w(��z�`�ىw�#�s�bt����b�L ����p��H��^�&[L�g�J`+}�L�f6j O3�7���(�W�A��Q
���H�5U��[�����@�R�(\�{�o�e�ꉀ�Y �<G�J��*X�0ə��|�ਹ/3���(,2|+cѐ��|�}�9�+�A�N���"f�
K���Y�d"+���TX�驲�s�+�U>)��'<q\]�{U�@ڜУ��^��<=^��3n��哜�6�f�����JZ�F���W�Y)M+���45������O�&��e��-{u�_�݊7h�-��fæ�z�y/�����vҖW�y�	��?| �+Ƀ�>���~N&6O���<����<w=.z1w����;�a{���?{���"�`{ʕ����0B�SXL~$��P%�!Oz���~���� 3��Dc���x�T��?�@�zVY%�W~��,/�3��O����|��a�����\@�Գ|���kp#�����g>���O���a��;����}~���"]/���*�} �a��g��]��8UO_q�[?�ޞ���&��,l�Oi�������w�A���a�u(��/����=gH͎�[x���>x���w����G��s�>������M'�F�F��N�2q(_�lӐ'bJg0)JH衸�'J��������W��s:��|����{.)�X�P��oL��|ݹy|�{�F���.v~��|��R��j��:gF������(i�e�E���f���״F�,]��d��ƍ��߅5ϟ� _OB�;g૕E�S��v�T��rSZ�͟~5H�@E�7D�s5��R��]A���7��&J�{"���f�
e�UN9��r��V�qh�Q,�h�Kz{Ǵы��a�P��	����]XX�c�"YUvI�:���]8[r����kt3G��L{K٩e�L`�r:J6�a�%<��l=�B)��=�w¦]��R�wȤ�	z�o���o=ڽ��ّ���쑼̻��i2~�?���$}yݲ�ϫ���v���O���^�O;Y)�0�/�� M�P T�r� ��s]@ ��B���u�ô@�`*S
y�7T�*`SA�Y�I*��ďh(k�+i�f4���g\|'3Z�l�J	#��U �~y͕J]և"�xqO���W,q����@�|�ԭQ����E�>*^����_��k��$I�ݐ	$�Dʪʬ�]�3���"/x��	ι9�3�TB����{Wus�Ď�f����Z���WK����&��<mū �[�6�eC!�5��z#}�h��+X�&a+��'T��Vn�����{1�m�W��8	�+�3����A��=O��S���8�4�~�ȧ��<z���Q�I8����an� ����5Lxw��e�n�;(����q�����v�\j�Q����&�+���D�TDq����:T���~����a��������y����aN^>b���]�~���I�r�!4���7����ʔ=�]�+3͗�]��QE�.�(I$��H�L��-C����S�����	d<g�[���n��[���2���o�o��7���?����q�m ���U��6��mz���ģiδ-G�C�Ӏ�"Q�ԀR���[ ���F��}�������yL��	B8ʅ�E;�a�|�in�648�-�;��"�����@�'���5�پG󐎫/�A����s�Jc����re#�\�d�ҹE��h���r���F��G΀��/f��5u��-36œ��o�Z����9��`iys�%�˯�J����(p�C���ֆ��l�%){ �n�^L�{�~�)����6^����ܣ���7_=��cp�>b��=Un�jD{ׯ��+�MoNu��̨I#�#�����y�1QÃ�d5�����g_<�~�s��ㆎ2lvʷg>
���5\#m8�^^�McE&Ȥw)F ��NYN���ҙ/�*�x��G��W\�S�`y5�QB�ֽ�`�q�f\eM/Ì��y����t��&?��P�J]�[Ă��d��}o�Lo�~��h����H y�⅏IM��Oe&�dF����\����tڐ��sx����5�8`|�U�Z�t[���ݕ&�FE�U�9n"h�	Xt Q�&ؔ�X����7���
»�k��F��-��]�`�@:�D6�#|�$�M�B��4F��z�OQ6К�G ��a"8H�H�$L#ݎĕ9$��I�Jv���b��j�]������W͌��ӊ��pk�%[EI^\�F��L��C��tWQ�\�lL�%-�y��xyG�.?�����4�>�)�*tG�.�e(����o2l��ɷN2�No��2���k���mMj<���-��W�D�*�V��u��/xa-�Y�Z��;B�d���L\=�*�w}�0��P�=[�ae��a%���Ҋ{�	�T(ۏX���9^��th�={��`�]0����{����T\GL&Va���§b��ɲ��ѫOiI�&�#���5�g�o�-#e~�d��#�=u����F�,i�'~�����GWd����&���TFӥ��p�oCHN��5�*��x���{
&�¯B�L��7�1ބ��L������t�^��tťʴ�v�i�Sf��s�O�Ό3�ϧ�-�}j��_|�{�y62�]:�%�,g�7�f����r5�<��B�+:�-Ñ��z�����^T���;�9e����A�FL�P�cnv�Yg�X���O�D�*]���4*쁶a�Vu��7#�T8�!9���ix���/��l�Oy�A]����`�y��{��)2�ޡ{�m���rk��s����!�ڐQI*�B�Cm��'�|�T�����?���?<"�zV.v��O��!��yn~h�Z������K��鈅:�S>�X#o�h�/�������U�|Bg�e߯co�#U��bգ�o<��nmT>|���,�aя;�W6��0��5�$�����U��2D^��H>Y�X��Q�[O'�!�?�"#�7�#��a�������y6�0���U���N��o4�2���"Q�12m���'-�k!����ƋX�=��?q�Oo�L����5�� LC��Wb���o|�0�.�ى�ni��n���6��J������L��`�G���8k_�UZչ&ej�I�������0�l�J�� ɗ��pPX�3���+�RA�Y��!��C�۸}�P�7�������B�2s�ӌ0��kl2?n��/<�I���E�5���D �'����/{}�t�LqD5���d㋧"5֤#J�|S ���^ƛJ�ol�[���HX��4���{z���AH��5`ZH�7�I�!�-8�D���C
���J�6�챚F�ĹI���Wo��߲��!HØ���B�SL�l�i1D!�����t
�������^�爐暹�Q�V�~�ਫWw17ƽ����3+�ޓ&�l(�#�q�ҡ[�]!ۊXT��	�ȹ��
sL*7�yZi���ӹ.�3c��R��h~��U|�G�\�U=����u4��2L�\�b<��
n�����}4Lӽu/�;�N���|�r��[��'*�1Q�{Ӛ~����*��������5NC��<����5`�o4�u3��]MOٶFy����ʘ�Uވ�����eJ]`��lhi�/�i�^�	��$���t"
�rO��n�H��C��@o��ڭQެ��s������v򺧉Xd�x
�� p�|W�_�+��4�!tq��w�*��ϩ�f�HBu��B���>e�F�FX�T~b>+5i�<��0e�.���f���cO1��[/6(wY�qN�81�:���Or��K��y�r4��2�����ޥW�r���C��j��mq������)������QkN9�+�"���yNAH&�R�<<��n�1�{�����#K�H	?`�U�� s1�&��ܼ;�w�S�eG�H�Ud.�&�Ե����ǥ,�����KZg�i��3?��\�g���X	�I� ���r��_/{��U6�P a7n�����g�pr�'64� k�G5\��q�|/��UϠȗT�;ˏX�P��k����%F�9�?����%C�5O�	ބ��|I���t�c!c� �^/M�FL�� �?��J�JS�
Y0��)�(a�A&�Ό�6���ި�dZI4��<y�!�I����dB��=ё�c��8�\��Vs�f�5��o��oӎ#m�8?��|��<�M>�o�P�iz��n�(g� �m�%�I���2��<+���O�h���Oy�Y����2�嚕��0�P
�Ɖ�]�&"~��&��KGi��|57���h� W��A�s+���U��W��7mt��:�ѽ(��z��}Z�.i��g4����_],�E��I���`�>k���0D��m!@�p�Iŀ�&?���0v��,��,����+Z�:qٍ_<���H�@�T�Jq�(�%Z�"�d����RT!nI��4�K�]r�a�9�U���7_m	��.b�w�M�����4#��<F6����xL���	Ty�LJӼVÚ���f5l�����3������{XEU�g�>'~�ƙ��U�՘ţqf����/2���a&i��y���*?W��.�%���V�ܸR�����a�<F^�����C�3_�|���!O�Y�����L8��|����O9��p<�����z���Q�艶�`_�t�Ӗ��l���o���;�:�-{��b�|��L�*���&e��.�;��c&�x�!��g������8ϐa6�=w� {�>YWa|`�q���3Gr#�[{l���{�gO�İ;=����􂱝�%������=�؎Ek`�� z�>��>w���)���	_[g:�j�Yg�/����^�l`��n�0VQ���)�\p��	 i|a���N"�6�L�p.��Wؠ�v��xo6�E�Z�G��}2��ow�R��P���Y/uP�@�=} <Z~h���1 4��`,J�����ʹ��D��9t���c�<���z`J��pt1D�5G��_^�a�&��2������Y>r�q��gCD�ȫW�	�U�F�n~�c���I?d�
z��(��Bf��*�1�"M��MV�W3����Ó`�LZ>y�������K�N!~DAH�����-5qK:'?$6�o$�`c���I8�z���Hz�;����O ��+�I8����XNxVhSQ�r���(�m��C���/J�N��]�&�/�
��承��w����س���a|�k���ۻ���\�2�Y/��?��Ƶ8�(�Y�GLw��]�����wK#���;"��k�s�h�m	�bI�d��=6l��JCȉ���z���\�d�/UX�n% U����0��J'^���#7����/Wm�c#H�	��t�
�Ù�8�e��'VJ^��M=<*o������5������������3��g�4�����#���ౄ2���]��PV�*�A�
j�k��ʷ�����l ��m��j��6���3e��f���H�G��㸄��3��[�̃	[�f��/q�q�S�g��e��{�W.�1���u�~����Ca���ʏ�B>����O�1uk���oRƲ�"�s��]�7�i�7������t'�~�\p���-_��t1#ď홦�e�V&�3��3A�a�������,�9�>:�>f���`�W�W��7)c���K/��?�ǋ^3V	�Q�F���[.�Q�3s�^s�Vd߯S?z�b�c�E�vu�glB{x��8��D�h��+��ιr���p�.�P2<{����in���t~%��!���$�e |+|M���W��嵍;{�l�ً�|�S�L�?n��x�yk)0t���B�!*�W����oR!�������O��^��l�iy�k]ᖙ���^@� �2«h�/b(<��N�!ˑi1�"�bhj�ޖ�>b�|0��dLQZ�߰^��(=�w��қk�_+��Y��mK��W��)7n�r�H�`Ty �a%b�M+ƄCw�=�Ғ#d(�&��m*t{vle[�8�7G�%�&3�����_) ��d��/G��Y�	~���� u@���B�g�q��"Ӓ9|6Ôx�!ޒ��P蠿/x���gķJEC�`�6M��d�7e�����D�gұ�"�^^�4�A��q*v�g�8dYx���{�|Up<r���#��/y���B+ύ*�U�9U`���5Y:����/�۽�p���ځ�ud�~��x:`��&��{w�aG{�֝�A�C:�ջ1|���=��I����x�0�@e����˕yu(K��fŗ�EY%�wa���C�ޮ,r�y��&���}A+������,|p��8>����]>.��'�n�> ,�:+��v}M�f�Gy���aJ�
L%�;y>��<A0��/q�V>oe��U��_��#?j�oB���m#��u�eh�O�a1q�߆���	'�*��*��^��	�p��Lg�������8�r黽��q}_��zͰ>'/������m��W��3l� �M7i�.��˲���e���[������}��(�����jjY	�~�J~#��b��m��G�]sue�{�ql��)�-gE��e�v8�hB�q������i�X���C��t$���!=a�0��hp�o�K�Ḥsv}ϫlBzJy�`>Z<i!'�Y�v�k��s٨�v1wH�M�>�|��7��5t��+�(�w�0ꆰ�N)�6��@\�=�>go��i���Wʵ�]�:�x�&H{DN�{��S�'g���N0��OѺ2uo��G��a�VW�{uj>�!��$���l6���]ʍw����u<�� �&�7|�C�pʀ�ȇ��O��6���������W0�8�wװIӹ�-7�'�κ��H����tM�2_|�2��g�%��'�!"0ŋ��-��^�v�F�y��v ���8M��W�)�i��(RA���2�fe����.׵�f>�B��nq�=�@ZF�����鍸�z���13� 2��ZU8+��o��$���_��+L�U ^�'j�D��6�X~���#fF��NB(��! U�d~A�Ci�8a��|*{� <%��a� o��BRX�#����3oS�hϼ4��,��X����a�K�� ���1�+�]�o>)Z��@�q\>t)��&a'���=��D]Y���e�̤{*	W�nm1�w�_?z��=����Y�}b��N��0�p��`�K���9q^^[�Sq��0ɮ���ixu��{6�W�>����-�b��`l�?xp���}ʑ�|灹��ϔ'�R-ؼ7�ˣ>�O��o�e��u1���2�4�OD�Z���gU"
$Ň��X?q0��L#,#�OC��qX��ܭ8���t��L��A�Fz>�G��.�wӜ������U��=�Ű�n˧0�i-��f���Ø~�>'�ާ�j��������2l�e9[�c�?E?�Y����OyC�w����m'v�3�G���'VC��a(ϡ�44�Z�ָ�eAٳ'V��5I�Bdk��`�8����_�#��b#Vה[�Y�b��e�iv�Q�����\O�C-�v |�0�H����ao<7�vYW�ih�cX�9_ǧmO�=�a��k��#�%z2{cѐ���E8��n�53�\$7��0>n��D�Opq��!�&�{�@����^6˪z�$_H)|ǑK���5�bl1���v��B���oN?�@��eY���|��-+�eީ;�7/�'-��zs��N)S9�}��֯����fX�Ы�u�+p����I׈��ȼW=�_�N�q�Z�j�)փ��-3���I�0��R��x���-x�$L�?��L�[��t��*K��<8Ʒo���-���x��HU�R��#�2Py���Gf�E�1�a|�V�\U�I���^��D���|�-!/N�I���D]���ʿ�/��&���t
u�+�x�ݦ���8�M����s<��+%����G����KX~oiq\~��l*G��/"Y8ZY,i�{�_�\��
^�V��ij�����BG�	ch�Px3�@�vv�ǭ�]1� K��O8)�n�*J�hja��͖	�
qc � %�?�1V��
_W��r����,=�@�r����x{dS1P!�����}&�j�y@�-�S�3W������;f�/cX�|��+<[������qD������a�e�_��kZ����;�EY�0��a����g������Y�(p����|���o�`VE�;?���+
�\�*�t�[%��1����e���Ȼ�����׌/�P=�W߇ӌA܆U��{q���]���^�4&.��n}W~U��G���>iҚ_���Wq����z#S�x��3^i�-L�����~�k��v>�$��ބa�yMx�i\�yMw��GƟ�|V.��nؙ_�*i���p�Y��K������ӧ��O>_<|��愞���/�^G��k�1]�"�yU���F�5��]7���A�b�N�'}��7�8��`����Y���z���E�<^ݥܱ���1�;�yj��۾��Xl�L���fH��/�s�1jaqʾ�鱶�G�d����P]����yRg�'�	���
#~�Kh]�A7¦�Z� 3�`��[�o��aZ=�捽�nMa���)���gC:EA��C�V��o�VC���|C��1��^�7�o��/,N��#������"0'SL3�=��@�%�4P�n� �l�i(Ӌ�oH	��;y�LJ\��q�JGF��UCiD�K��f�L^�{�L�:ι�k�d�G}���<C����<X~�'ߒ�0��Uf�c�7��3T�n����{H������vp7&��|�4+#q��pH?A�ho|B�AЬ��)t�9��
���"���5�|r��ϼ�`w˖�g^���0܅P@CD��X�C��P���K���7s���߿�H���@G2�"�U�L���r.V�)@U��'��P0��O#~�p7%�5tz'��ý���&�0��ě�,Z����3��<�s�&>�K�)��=�2�K/�Sc[��g̰�Sf���=�?��W�+NĐ����݇`�J+J[���r/"w��0�]�v��^�(V*V��!��������r��C�۱��J��-"+�Yʁ����U����s����2�����y���?�å�������W��t>G{*+�_Z�����_EV)�V��H�sލ��&@,�w�h\S)�o��#�5meo��Db�he}��?�V�����[�ȤiLx���֤^�}>������m�H��]3����x3��jٓd����.ˌS��3���l j��m��.�m|,�F�N)�e^6}}��0��B�'�=e[C̡{w�w��/�}�\�����k�@C��0U��Y�W�n-�2��A��e"�&����75x��3ı��-{��ۡL?����/O?g�-L����g!�K�9=Bn�`/�G�wi�=�`|��[8�*�M==��:�r��AT�9�By64����)nv��B�oǄ��P/D�_f��a�� ;=a����dx3�4�Ҙ�kT��i�p'A W��9�]���@��#a�SÛ�/������9~J����.됔i�u���a|�����,C���.����[7��<_��B�x.�����_ox�x��p�4ѹIK�oM�B^����w��@�H3�'�I�r%��M6iJ��}d#�w����3�����g�<n�
#�zP�ge��~��(A:˝y�|�&�k�I�f*v�m��1����� Vf�V��h�����aV9T$0�Kx�����V�*��ӄ�;�G,^{���f�D<�xkZ�BOt��4��N��	p'��O42��eN0��b�LI��-�%��#�g ����"*��%G�tK�'�����RQ&|�%?�73���";5���>{���J6-�j��g��S����x�/]�B��c�ҙ�C��0C��� »�Օ��?20i��R���W1й�qx�䙭cy:�S�D�قf5"C{�����W+9鱅��m��3��
+DitX@c�#G���!g��ƚ�^}�>X8�3r�aI��X�_�V?xC6��U7
�t[��{x�!�{�y)�Q�����˙�O9$��+)�u�/м&��,�O�z�+�|�o�p�����;�}�S��F������/�vU���8�W��ϧ��9��m'�¬�ֿyl�?a*�f��Y>���[��s^���tk�eXy�e*5�[9jX��P���0ꟴ���8��%8�^�K}�tf�����T��o�:IjX�@]g�5�a�[�����2fϊ�H�C좖�M��o����CCYޅ=$�X����x9uDz��ObI��T{d��樘=e�
�<#���Q^���ş��>���ހvn#��[d�а��~�L�j�#C�/^�Z�퇟���ū��ؐ�
����+u�@P��nP�:�U���;I��o�Z|��3�<���T©[�4���t�2��p���;oӃ�D�K/x������f���Ј����w��[[<ek�����K/!a܊"G��4���C����ݡ���?���kI]�>m9ZI��mO��L�@5�-����G��/B���F�N�W=c�^����r�*p�[ҕ�|V���Z2�7dq�j�@��R�9E��=bֺȹb �\�x��U����>�w:�j^�;�5�-g���e� C���=ˠi�|ק�Ip櫅vk\�ߗr÷E ��!��h��6*"g�������J{6N�)i'�ĻX%��
q����;�|��	� �9���IC�p��iŐ�m���Z��̦%�^�#�	�����:�q�$H:Aٟ�ϑ��M<�S��K�(�Qb(ڵZ�9	�a�o���M�!�f*x�;Y�HCzEi���A^T���ISP��'|"M�:����������~�����Ƥ/o�|ȟ �a�8�.�j��G>EnL�7���^��!���r���^0#�yVT�D�(��S9���U���јtn؅�����_<}��ϞB��`E����K�t��.����s��$�]��<V�{���"�`R�C�7���ሯΎ�h�T�"��
��+�}���u<&o�_�p�0���0Fس�F'����p�E��	�#F8�>��e%���2�3�9���,N�FY�"3�	c��sOH,�\+[������jz�i����'}���O�u��~�G�IwIUc^�ch������ϙ��f�<�7�;���}3�?�+#si�d���N/��֟!�D��^H�w��lx�aB�[A?��p�x �H~5o�.���Dh U��cSk��=6F~��A�!) ��bˑFD�/{D�Xn���n��z�x�\�~�q�����Wv�g���J�����琹�ҡ@W9�������8�5^.Y��}��p�u�(�: ��^3Ϧt����g$��S_B��9��'M�~�����OO�6��Ɠ���O�1�5�ڢ�x���u::p�ƩN�g�xg��_�Ҫ��W�|x@������o�b�e�D���Iػ�ig����'�x���J�Ӽ5��4,##���/�d\���k�:1�d1�`�h� �2�F�+�5��X�4��{3c�'&�D�o������ܿ6���9P�H>�~ZU����ҏ^��`f��~k$@�aU����ɼ�-��o�NsFt�<e�-a�	տ��MhNB�6H���'��ZƓ�֭�1L����m��]\�@�3�����[��+��ΰ^s<[��`�
�-�v�ꯠ��6��/0���-oH=�|�!lV8U6�1�39��W���3U>��yR��7���]�Q^���y��3�p��>'n�_��e,�-�%!-/����~�h���+�&�ȷ� "V�*D[�(
��dHOC�}�SE_ȀVY���u�!�*&���������s6R<�'���Y��c������(U���6���ӳuD�����L;���,mढtC^^�i�I�(����&��p5�p����].���SN��T��?e�|�a-��I
�
@6�-������a�(τ7�6�	7��K�"��ʲ^~�{��s�'����O83=���
P���
lq�������L��-�p��-�q�m�'��K�Y���<�w�İ�sWa��W��2͙������P}0+45��)��8�~�+`�Ox����)������I~
��p*?*GW!����u�	F���k	.M叩r�r�Cnu��bEf���0pO��h�q^ ⾀.\�t�~&�?�[���
ٺ��_~��'α����`|�Q<=��J� �K/����=�{����;(��|���}����p����Y��[�zA7ez�o ��uʐ�#�O}b�\�!{�1v��8�C_ x��|t��"[n�B��jS�$[�(,�'{�7��-6�� :���>`�D{��'L�V��>�������9'$��v��O�+�� @�H:s�|	m�Zj�/�[4��/^�E/Go���}$$̷���$���i#<r-��y6 YZ���ʡ�e8]xƱ���P7#�D6d�������Q�V����u��,>�=�i@ !��[PbDHa�H��X��	�Ba"���/\B(K�w�HP��_�0���k�J fF"7[�&����z'-� QE	L���Yѹ��8"�[���^�QEk3=�b�.ϡ�,�Fj��� [��_\�ސ�{Ӯ��*��R)w�E�\��?�W�)�H�$P��7ᥑ��?�߷p�߸���$;|���i�U�#,7�򠊶�l>�ӓE�چʲ]�
�s'�_�-���wQ�SN�5nrdT*ft7{˴��ޯV@���w=�ު6&�rT���Gq��me������ �a�����^Tn漓��1�ز���J����bex�%��'�Fn�#�9����.�k`/�52�{���(�Y%��ͻ�ǲ*�^y
ۏ<�v*��)��͇6�H��q���7���	0}�����`��t��V��|�2᳴	g �s���׌�{+I�ʋކ��*��e��[�L�&Pnb�y[����'�)+n�7��0$p�r�zM�"�o�G.<�{5f߅oJC-oA�����l� X���M^��h�AYx���˘e0�J��}>u������o8#�v�MP�Dߘ7uy�X��g#�Jy���Ǻ����Y�| ǷPv1��{���ȯwl�����U�3��kzo�����;��H%鶧%:���:����
^ஞ_G�WX��~g��V��ۆZ7��K�䕟˸~�o	6�'q���!�~	L�*6,m�	��N�HFW�&a�|4������w{�1/��[x�
�}��r��Q�Us>���>��0����R�J��$�����������Mb1^�\�  ���n6��ɴa��Y�U�ԗ\�,|$�g� Vo��ԧ���S\tM��"�'~�q�e�!֧u�6ʫ�%��T�~(T�����Z�pR��/Q�v7�?��*�� �@sb0�o�L�bY���Gt1�O����2p�a&�y�"��c(��1�@�6S��4��
��9��4H��̄%܁�C��y
����`8�3=�I~e�5�U�u�O2I���IcK�$(�Ʃ��� Ş��,�U���a��m��o��,^������w�����&�@\~����w�/�N����r!24pkp���&�!7��G9���
d��s��aR`#5Z� �<��Ъ|Uvʂ-w��;�ӭ~��\���s��q�7j�gN�;c���v�?Z�gO�W�^Di{���>���^+qr[���`s�Il����J�9��^@�A�g���b�dA4?4�>i�b�>�D6�_��r>k$�q�H��<�-p��+�T����!2<�T0B.3��FK4�j%D8�"Ӭ,B�I�n��0w�V<�2/�,J\���7�yϟx�8�a���tMB�Sf��eJ���i����~L����:!�a�jZ���(�	lu��r	[~�`��^ ˼8I�jB����.�%�b��W���}�����^8�����x�_��r�ߍ��+��5ЅP]1!��J�h7�2"�"'D��vt�c�@0P\Ģl�0̡�ʐsne�������h,Ey�I(�򑷔ax�i�G�Qp�A�&��u�2L������"݂��z�����N[�%?�k�Q����X �.I)�9x�w�� ���px��>W9#0�#gvy+��\�gv5Ky��|���=�!g�φ��~	wp����9L�ﻫ��<Ò4/���0�ԇ�O~�\���ss��s�yT(��=���d�N��-��A�e��s�������\<s��w0�v�Sf͏�=V�2O���y�����[zGϲ��36c<��[�i +��&=��zx�aF*.��:�/G\�kd4�0yA��#��K��tR%I�� ��^�I��|J~��?�2���WF�	☆��;/a�Q�(�~�>�!>�I>��Z���1uT��i� 4sQ�kH�B�V�dc>aqY�6~E������!B�K�����
QF�!KhC���᫃q�i��7 5����/]up����Z�>�.�1��h�:�4���X�#4��h�.r��7���QX�W�j$�"�B�p��U)ʤi���}��+W݉U��i����,��V�=yc���P`��:Ro~]}��LCG+�i�2J�\��V���_�gX|���0�"W�*��Q�˜��8	��=_w]�u�0�~RQS��O��v��礱M@9�����ᇟ�E�bn�B����z������8�y *x�H%$>΁Ȑ�3$�CX��G��Pr���̠Ɋ9[������s`����[���/o��]��aw����Y���|F�>MY(�&��{��\��)���JJ�L�&��}O��^ʂ��N�J�&����iv������c<�1<�6��3�lM�s�A�MKG���M��C�%�CO`�[�R`Sn�.�I缍�%i���M���k���w���6D۸��o�&��D�[�RJ�i=⩿����zH�CW��v�;�1�ps��i���,?o�{zzp��D�	�P�!���!�2H�)����u�'\����SN����e�+�Ȅ�|u2p����lV�
r;�Qzd��h����A�ċ\8� �:Ԫ�F��?�0�.S��|�%�ܭ02L�Q!���>m�'M\���"{�	WQnwc#1p�%�N��tLp'���QF�M}�崇��dZMI}R�3��!��(Z1F��}��kO�� �sψC�CJ=%��)i1rp��Go�+$��>�m����쿨�#��S�M���8�wÚ����n
��zӴ���<�_��昞�4.���O%�|J��;�U@�fj~�q��03HB�b��An�^fNH3��Ij��Sf�mʆq����m|�1�2�߼��2Q�>e�i�Q����x�X~�l?)���kQ14[w��_X
�1�J�X�*���!MZ�.�\����)􎬔���  @ IDAT���5��f:"=�+�*�(
(���@�-M���ݞC74�!��s,,-�� G��:Pʢ���Be&�EE���|rrْB# �OP�_����-4�<|��h:�ۊ���R��Y�W����V��:FL����4�+�����B�(*��yl3���I ��m��T����;��U�m+�M.tW�o������{��x�9�.CW�����e>��6�����������n�z��}?z�x��3V!}�v�����f��ت��[���D����>w�V�k�k�s��Nnx�^:�B���4�5�B���m�V����UX䃽5��u�$d�{��r�y��6��fRn���ee������"C�	�
Q�(l��Ω����)�3a5��Ï��柲��y�gp1��Y�_�7\dLo��!etaEQ�!aaj,릜Z��|�����%_����,�Tq���k>�lp��k�D�K�|�#��j>xԎ���ebj�u��8Ϳ�I�,Q��r��qUe��'1~�=D��{��o�oY��r#A]b��aK�%�M?ޝs���̋��.�lK��=cҚ����_��c�.n��"Q��Xʞe�3�s���ׯhT���r˴�{6� lq������)�}�c�/vz�y�{�cU?�{P ]��M/{�\n����ǜ��>~����kd��6/{D����'̉:ff����X��.�4y^��o��r!��]�l�������,�\g���/Zֲ8	Xl����s&�1ƫƤB%��e�������+O!`����=^|����Ê�e^DM��$����<ᝲ�9����w��qy���i G>~"l��*8������W�&�}f�����e�2iĕk���ƐzI�]÷t(�#ܓ���0���W��qu�v�>�]}�O����E�7�bg��<E�XG(����?�S� ƹ�����!-
"��w�s�ng9��廑y� ��f��i$'?e^�y��e��Hl�7���K$&#⯒�f�Ad�f�$���&ў{���7��f��ç�����e��n��U�#�����M�Uy�K�.�O�J���$���EC&n
�>�:I��*U �7�)������W����ҿ���L��m���/�c�=�����~8).���ŋ�K�콲��K�Y�`O��f�]�vyk$�K(�� ��8Uy^��4���B䆐��,���zq�!�_oPB/9#�=G�:@חEҊ��ty���&�LF�o/>�����/��|�a�OX
��wjC���N0pN�$�\r���OR
t*(=�˼3�%g����#�iG J�Y6���U�P�z����R�4$U��Z�G��0�������Jag�*�S�&�k�c� Y���̸���O>��)�C�����^6�L���1�.�)��)� V`�F��vA�3�Ө*-���LOb~
c��9h�M���ß��'8[�(��_�r7=��YƩ�%� I�IK���\Z��d���?�Mü�r����d��S��c��Af�4��\��w�E=�)�P����(K�{�n�x>(�ʔ��(��-�%".��_�
�ߏ�K��7���e��4./��<b�ի�Lg���Y�,8q�/�c�:�{�����w��W�_�J\'����I���I�t�i최��WL�1���[t��%s>���k5�t)��-F�eꌞ���6�?C��� �W�Y���������{�~����,+s˳ñ�U�����濂��`���V��p��$�'�V~<��sr?g��'��r4@9@��p ���J�� `;�=�N������rR^��2���Op�5�f��I�J�>��7�<Pm�&�AKd;@_���b$֢ x��9o��pǨB��o�i/�y7d�&�p���>q⧂�.̢��oު#M#�0����2 ������4L�9+7��Ej�y+"d�$�.-R�r�$$0n�@(�y�%���]���d/��H��-�N�'��0y@D��?ҍ 8�e��
�Г��7�Q�ͷ�x�a`�&Vv��#���a�ўZ(N�vb�
3�\d���q�M�̤o2g[��Z�|	w�IM+R���/ O�Of#��X	+�b�o�WZB+����
g�\�VnP��H�FZL��_�0]���k#/�T"�� �L$�b��%Dsɑ<��B�I���a葕�[����e)`VR�]ޤ{Ƽ�3��p��R�[����?t�?������H/ث7�ٹ���ǟ~^�A����xV�ں�^��۾�㷋�������7������ �x��ܺw(��i"����rX"s�4Q����?at;	��ɪ;*&�uH���%��
۳
)G��%��)��|kl���i�828��O��e������] �O�`Ȁ=o�8�("ȎF����{�){�h�d� �:����:)�\e]�T��L��a��
�|����G�� ��J|���(��P~/0���r���xI%p����񦩜N��8!i�^`X��Wi�gB�.4��+='�}E�Z���a|/��w�N�-�L�~pP�	A�;���8��x��/pt�a��ei���&����S�-��	��c���2F92�8�2์ɕ�<�5���Y��ғl���V��yx,.�%NJ����H�Oy=�k\�e��\O`�C|�g��W�9��U�/R����)���:��C���O�z���G�i�`ϯw 9������i�8���:5�A�[(mιJ9s�Y�����_c ��٠��>yq�'=F�7������J�C�/1�~�]��v�tfGGl�Sg6D����H�e��a��T�Ѐ{��9�lm�f��,���L3աO�W�H|�\�cξ��߼��5u�zU��|
C��������O0�����0�7������C��eG7�wp'?1��H�yY!B^���nz�kC��W��.�� R^��9�X�?��p�?qR�Ut,D��>'�}R%$A����� �P!�Z5�[�����&�!r�iY3.��TV���H��Ȳ�Eއ"��D�b�ٻ�NUՊ-=`"
�Kn�)2��o�i��� �1Zo�� 1����i�*b$�K�33G���D㦕]:�!F�! �7�)��^�R��'�aR؟�$O<�̷j�"�\�� �:�+���d4�� �HvP��/
=#��\Qɫ �?�#�Oʹ-�s
Q'��@�����-�)`U
J!w��!8(���I�U0�C��2����TJm���^�G�-) ����RHǲ���*���|�^q0B칲�_�9�C����]x�ٍ�p۹ (��s����!�G�ޱ3�;����"���=V����B���{	����G,ci5k���'2A��������}�����/�`;
�]���R�X��+����j/^����dY�}geJ��,:�C����la���J~�+������[��W��?�!//=��c7��P�2�������UPDy
����Bg�6yȻ{$Ik�^2F9q��"b�PBM�0I|#qQ(�/����*�2l�M�6:`��p�R%��i����K�҂�5���|��/	�K!�_Nbp���������y��·��0��
�@�!	\�*��_�= L��Ѱ7i�S�K80�X����\��/yR�xb��nx��ޖ�R'���_z(��ʑC~�iZ����o/��/�����Nᇻ+��<K�H����H�-�G4��0��Z+:͊9� �`�������ۛ�0�4>�'K���|Բ7-��=��~��w���?0���	���i4�q��s4�4��4�^���#����oρ�(����ik��
?�8��n�A���9e���7��P�G��YZ�5�@�$n�Ue�]��!X��J�i����×��t&��U����ГՎ�������Y�e�
?���������M^9i=fO�tzE�̇C��:�pBV=�S,3��"� �y�Ӻ� ZA�w�2OB��L^[~�ox��X��`0>##��,>>�P`ʿ8;B��8����J4~S���u�v��
�ɵ!}��EL�/�RBȦW�$�!�[�k����]�GH�#���l~���H���ƫn�M+@Bl�Q�ЃlHTh <TrUt~������	�TAZ�-p�@e�����$��f(1�T�|�3`�0^�K���*n��U��zt���xw}qtw�ؿ�~Pf<�q��f����w�Bz�����D�`�§��$���K��D(��U��q	�UƟĒ�\�������N[�!�8p���ĳ��"d�L���$�?=|�s���Y�G� �0�z���/��s���N)q��N��;�j�O�'����h�EKw��g�[[������8Ű�e�{�}���[#1�ɐ��Q�{3>��w�f�ʣ
�y'(�W(�������?<_�~s��q&�
�F8����@��rn��x2o�p��l���`t�^`�d���N��<�Wy!mV��=Y�J���9��Q�fAz��0U���NV����ar.B3��-��{_� U`�'�ଌ[��|�pk���=�b\��B���\3�W���Ҳq⩜{ٰPV텷h�~2'��a���`�U����;/�*z�<�;4������mzN<_��H%�L<���,o��m:T�^��R�.y(\���K���y�N�f�4��NϚ ��ƍ�ʋ0��r~{��OS�=M~'�@Y˒΁�G������԰7��Y�]�����[�wp�Mvτe�t:�Ն��֐���&�K�8!F��o�0�T�O�!�%�(�i�:u���R'�7�:�������3܍-|������^慆�<���q?�3�;�B5z4���^!yG`eG>9x���^�utgh�����OH�e� �g1A�4�0�K����؃�^<9
�f�����Ve+��g�>}ʭ�)+w����F �W�c�0�\��,��B����	���_Ƞ щ<c�����{oя�G�k蠔&�x)s���'����\#�4o�'���i�VGZ�WfH�zԼKk]����y�<(K�fb�CK����t~6hR�BWt3��"��̈+��zɇ�0�dʛ��`��rzG ���oC[[g��:���	m)��ɪ %�;���c�#��T��r}΁Ǘ�t�q<���_�3oE�V8_�}Vq�&"6�"3
�*�*3J�`�J%�f�L^`ja�G癡�]ex������7��wS�x� ��w=�Gߢ(P
�1��?���	V����ps��KälX��K����),��+����4>��������?k��˿�����iȄ��pȷ)x�L�J��jV<3|�N�œ
N"��m�f��Ŀ�E�o��V�Gv������WH5&0T�7k�[��b�����z�M�^�g�U&�bx��[x�v�>^T�?���ޥ�eq}A������V���:�ʦ�F�����\P]��_z�Q�n2�g���_�ắ�`��굻�SIx�YW�Hs����;��0����S��%�\s��
�<QfѶ`߉��/U�V�r�
ݗ�������\�����]w��.o���0�r��f�CȒ,�&-�?3XE��3 ���S/����c�@�͐2"�JNz���WeH�ۥb�R��RAA��1Iؼ�����|+��ȯC;�n@����^��u���8��c�S�S�IY�Q�g7ohQ�5\\\��2=a�]�Gjϭt�o��$DҲǎ��N��@�F����Wd�z�#_�SJ/ ���V�ʸ�T����h2�Og�ieM�_��S���iw��mvg���ϻ~�M�=��O�N�3��Q��._����У��-�^[�Ũ����\O��'�w��hd��9�vͰ�+�c�Ǣ��W���@��{/���G����{�^�N}o����wc{��_Xͥ�c#���ꜜ����W�Sq#5�%���e�������O��:z;�o�ApL`��ĩ�d�$��<UN�_-����r��70�jԸ��8R.>}�ۑM�#�m ��Y��%�p�"�?l|u����!�c��"�Q�����{���o/`���'�|ʬ	q3���\r�8��\�����@�N�(\[?�t�F U ;�6�`C���C�S�c/Q1��ˆ�SWLZ9A��p����,�!�#e[FR6A_�N0�,�̀�w��a��w@��5�2��P�?x�=��Q��eޞQ/4&𬓴�+�WٳH�fX=Zt�eU]�D�3����ad����>� 6���aK�L����6���=(6�O�<(h��h�F-�|�BR�(�*$w��P2}$���i
����Af]�����Sa�̂��-��kUR�L�ʂ��mFY�p\#�-[��wG�OǴ�ޯ->��^=��f����&�v��,�E~ �
\��$(��q��/s+<�b@�WnV�C���*RçJ���g�c�# ��Pq�/Y o6�4���N*D4��`�8F��X
���k�Q�'(@���������
��m%����u&�2����n"�N��闗��/>,^�>�|7zڥ������{�ܫ&�c6d�f�аk����J:��C�R�J0��1x�Ѱ8Uy�|	����?����ū�/�XYt���u����|�T�T��U�jc��5
����}�u�A����t�d�G�R�ާB�g��� {R5t�	�`a���0�S���՝����5�v؟��G���	6�]{�\�/;�^�̥P�������u��TdHG`����/9�-C �o�����{�9�q�,^6 �'�/@)�{,fp.�}&��e�i�^B��s�����_�8�U�N��AIy_Èy�C�=�8�����,^rx�K��z��~W䋆��~��8�d\�V#������]�@���A@�oQ�ҳ!-Vj�b>v,�k��؈����Z��OJ�Gza��Wġ�O�?->�g���Q�4^4F�y�G�K�eS��,S��^S9h�R�� ����ߡ6d��<���,y{Ȟ�ω�a��5s���0����L���C���(����g��GW�p�q���>w08�qؽxJ�����#����h����JP�x	�;<�k�!��
_��gT�ȡƅ�n��O���҅Li�-���u�i��0�����m�yjo�gA���u�~�X�Vנ��0 ��Y }�i���蔈�����ػwi(��M߫=-掠��~�k/�e��&m�I[$�R.=�_��2��g}ku�_0lO��	�m�r�A9'�|��%�i}Bo(�f!ð��X78��.��5�H�Fŉ�5������9�\�hŐ�Q�k���"�knu�dD��+�]���z�
8�~�߸x�x��P��S���Adz��7��K��u>�����E~� �B�>����6�9�-2�j�w׋������(�W�R������_3gL��O��ȏ�(����X���E�ߔ7���М�	x��-�+5.4�п������F4������P8���	��|��QI���P���(��i�Y�!J��q��Z-�2��7m���Sf�fA�`VJN��g�/L>D�m�^-�&��Vԉ�+�	��4|���k��M`� Mjf
�o&i� �Cqc��2�^��/魹:��^P�	���Q�m�(����b8_@>��O ƍ�V�o+3щ��(�*'�g~� T��X� �,��/��i��4��f�2D��ɯ�޼5�a�k_
����4��z�*{4.�S���4n�MZ*�j���(�+z^��~s�x������p���Ұh�j��2���.���S��]��Y��I����GV$�n�g����1N�N�!���1=j�g��L��P����M���x^j�Dޣ��5e�<�[g�o���u[9��T�_~�%y��%�����&���y+;+h�S䣻x[\����[�����2�B�&�ȿ�x�!��g����! 0�y0�<����74�/ʖ��(��r���'w��p�}��z<X����1$�Cb��,7+G��42:�������ٳ/3��^�m*[�/0�^�~Go&�`��� 7R�.��X����9|Y����5�0y&�Ι�'G��
����!-�_g.�2��Ӟ9pð�(�fsd���T�q�J��J2s��c�:��<ý���������-4�%�/�D�a�21�(���!�w�J\>xL�'��+�kcl�4HN���@K&�LyB����Q�[d�=�g�r��b���ǭ�[):���:�{�|����=H��F�9�W��ߤh�� ҵ��_�z��	xR1P���1�+G���2$��[�$�L�_��QrVP�D@��W�\[�R��H��YCD�}�^|O������#ʚ��4���a}�6:�^ � -����L|�,������H��A�5��)O���=���{�g)�^����=`���MW;(�AJO�yԟ A���4p50�W�
N�A�|1}{�cT�N�0��/�5ڙg~i�S�\��ch�����9x�E�"� w�����.�{��ۡ��:�F_GW*���zO�;� �K��^v���@�r�)h�^o��}J.:��Y� �z�) �m� �Y s��#ȍ��'���]]/�l������O��؍,k8�����ͫ��k?�:����M-�Q[B�]�9����dT�#��%�D����m�ln0|LCt˭��3p�9��䛦44��{qF�¶��6�sh@"�2K������9�a%�c�VRX�ɰ�
� 	�^��I�>�~H���E���@2
 �hM&�<�NѦ`�%;|b6��CH����K5!���\���Ui��2ؑ�Z(�^���U��7pjK��9���-�0Pd��{0V����;n�%߮d�-2V��!T*��GH�`��;Wg��.�Ǖ7��7҃��b��K�es>��j@Yz)��&�*/�nR9�q*Q�unF^�0�Y�@ �`���X��y���P��"&���kz��R�Yu�
��LK�����c�����PIi�&�1dy��[6{T^c�e�,�}�P�Ǐ�1��῵x���w1|�X�r8�pg���)�\`��@�l�
h����9%�uM�fK���d�:GѹՈ�B�� �,l���̐�	�88�h�{l����8{�m.�h�k|��K��/��S���mZ��{�~�����/1B�>�P4�G3�>~�$��)G�h�Z�kx�Pag���H���+��C���6;dR�}�cW��y����j{b.����p��Z��4�X-�9�>d?�ﲝ�b�ܙg�o���]��S��`�ĥ=��
��g+���{,���᲏�s��|���c���(<�o��fQ�$
᪈A�)�VV�]���Az����Ċ�[cW���F95�ݱ�i4y(�=A���{�]�����(���Y)E���0�>�v������3<��F�����2d�|3��Tmf<��+x�������6+o_�/�s��7��R	�<|����S����-=�ۈ�q�p�Oa�Lp����G6w�~{�]�w��c��Y��!�ֶb���{"[�H�;���i�N�b��.`Z�B�z�	໛ ��?��⛯�LΆ��٤�A
�7��ϲ.ߎ~N�Ɇ���6N�c6~� <մ�|.�1�\��%����oH������l>v8Z�{��1
K9����%�<�3�d��_�Y���1AYB�8�f��{������L�)o��olm����2m9U�jʓ����ke����^n{�6il"+���9�h]&��/�7�+��W�X�Q��}��cu�˗���}�$�������*,h��8
S<U�v���<�e."�	iR>g�F����� �D/v��<{Do�7��=�E�p��m,~����x�(�� �EQ�W�=Z����h����UO�h�)�řwҠ�*����bu��U�!�pȘ���l#�gw�"�؞�uz��6��f�n<����- �Y4pHS�1n.�
��j&/*1��mE&Z����NKVcI��5��J(�{Z��w$ӧa����q�K��!��d��\�x�y2&8�#,�$.�Iq��$~!nN�#�kJ�0��ܭ>PAX��0�J�J�ʧ��X	ZA�W�ML�7���P���ӈ���u�o�DΥ-��0䛷�q�MH;��T�����il��!@Z���Sn������<�CLxw�x��0�(�m�^�\A܆W�k�2�(�-�IGG�(R�BV��3+�k
�7QD���s�c������կ�.ޱ�㇏0*82���Z�w(���*��Xe��p'�����'����x�p�Z�.�>����aAWa�[PJ^c��#�����AZ�#��-s��}<cx�nq{�Θ|�(
ޝ�?1td��
;ʙt�y�\+{�4�����1:��n�a��t��h|�q6��5�=���m9*�{wl��r�#L��R�<e�*G{�=^I�ǡ���}�����G5Z�U$��S����Q�#[����s2�<�|��ӧУaѼ?e��޵�}z�0����QN��J���^��h�a�ػ��z��Q���2�|���5O�
�p��a@{�Y�u�Oq��lR��N{cQ�5x���F��O����bR�e��r�Qd��z/���`ʖ)!�n�&����WϨ�0��]P�?f��m���--�-�#�	�R"E�~y*�3*c��{{̜U�����;y���o؃*��0���'�s:�!�|86���� �?F'I���kl���٨����向
6��P�yoX�UJ��Z�M��<��e�$���|�+��:ņgz����B�8]�\�a�>�p�OO�]=��Xtȟ�"��o��vc�^���_�{���zX��1D�Z*wd�r��B��F��hok^d��_ӱFu�4��K:O)�������q��\+{f�	o�p��6�$�S��@Ƹ��>=����"�':/=�`����F>(�u@^;%!��
��X��o��ߒ��0:>vC�l�O�=;�pN8�"y���Ij�d-Z}�\�~��޿n	b#E�:�d�{KOt��4��F�8"�G���/�]3\j��B�&l�N'����#�o�3������Q6?��C�٢����������k�y��i���"4���[S<�QyQ��Fc��p��q����_^��l$6q�?�ޱ	�����e����5.p*h��������䯮�46�����L��AX!��w�ۭyE�|���J-pG��%�5v��7�X�$�G��)`rm��B|,�oP����q$�$A���g`����|��c8����%^���Z6ܵ&Sq2=����1��iU���7���(�iX���cp���g��B^�P�!�!ʹ,�`L��f��$ݶ��ki�r�SAP�i��Ǹ�8,��|����/aF42R�P�|��_�\C&�^���$���f���C�(߄��ch$q�E� r��0��;��ďa!�Q!Z�g� :L�A�a�T�w�9z�f��J��������za0���?ݏ�p�AE}B���!}�w�ȹ`�t���wxw���,{���5+y�I�ʌ�dޗF�&wE�+7�3�v�y	��H�+g�M:�zG���m&�g>@�#Hdv�׶4]T�\�z{4"홰��ՀcN��Ç!�-�%+���H�c����g�1�1���H�9\��N��?��y��k�>m>[�\�gϞ-���������o�p�G�0$�E��3�B��1�p��Þ4��n^zM�t�R�ǋ�o/�;LDy�q[���(C�0�Ϧ1�-��"ֈ����/_�/A�8��J��*�F��~������F�����\]�����t{�=�D�z���F>OX���${F���C7�����E�o���I���=�nz���?���ſ��B���9��	�w�5Ce? ���59snF�����|@��=<V�����?��?1/�aAz'�(��{�� �y�ea��F��?w
;fH�|�Đ�;`NFخ����WE�En!����4&�`�9�g3���e�ѳ�/=�Vp�]6Vv�N]�������+��G�no�������k�tn�JNܜ'i�[A����h{%�m��BTȹ|���`7߭D���2c �����'�՚�c\8j�[�9��y��S$t�Je�S>��9	k�U�m �츍,�)pIQf��qa��G��T�8�"G>�R���p��q]``0;/���2Mu��	bB��ʣ�YK^g"��ޡ,R?���Y�8%�O��x�Ec;Yn/p�"psn"E,�[�U^�x�c$}��.��[W)Y�"��<�`o~���u��wV���t��s`�s�o�\axQ#�f�
����	)~_��Q��E�#gSK��� �z�E=�T�ȑ���J�rhXt,��:K��5�I���] ��&v�zTH��y�x'��NTGEO�r��S��7�j�-�af0�F��N�Wv��`T'܇2�2|�B�R��n���5�*(� (0��b1���
9��q�m.���a���+YpM��gE�YmL+M�J���r+L\m���������H��<-)\�H�������)�9�ъ���2h��C��:�b�-�uR��0�<����-�N��`����ɸ��W��<؛��̃T�D���5��L$J�5����=�pg�Q�6��POLK!���������9;g�Cz�T��ƒ�`^��F�Q���[��A��K�h0�-W+1�r�~2��zi>�Z�Gp��xhqs��b���J�>}�G�����^��xO�]�+�j���m @��`��� n����i�G����B�p��M��}�H�՚L��?���X�I�Ռ����� @�F���<2`�Gf�U���������G���rr9�/Ӫt�Z��m�x���YU���5� ��8*�W	�G�v?f�G��PXCY���T�"�L�y� �}h#�ֻ���$��m�<�؄�N�)�0�<�GG&�A/���)�Y��b9���p�ʄ	�~5�l�qs����o7t�NÁ�՗�.&���n>O�G|@��*�[��aJA �k���o�������W�p��l6< ����L�^K�s�����-�Sm�������G��p.��4�N��G�G}��#�n8��a���j_����P�fK�<	�e��+�a_�������@V9C|7õ!�3=�h~�h-�R^V�O�{��,�	um�7����(`��y�u*L����,�ޮ����&Սv��g���J?e����M�x�E�?��Q�����8F���F�g���-&_
��d4�}��%X���)��G��+����M����o{��^^���.���9X��xrT�C���vX?�[�_�*�WG�0����EmcEp��¤^Ym���	�`B��j�X=�^�rﳶ��|˦�Y��uL��'�:��[>Yɐ��AR*��<,]z=>"<\�����m������R�ɻ���:.s��j���)���eK��Qw���Q��}�O�
_�P��������;�.N}\�m-lM�x�����^�տn���(<K8'|;�͢�0N���QX����[@���0joF�.�۔��(N�X�sW��W3]�O_iׇu�n�9I�.)a�4��&#}���vL)���D&ތ��ؔ���^�=�?˽��,�+B�e�፥+�_��@O��0��ALDkb�[�.=<ydz�Z�L��i����W*���6d%��C�`\�k�3g5�W4�3�0�ҷ!�d�,�� /M��!�d״�.J8��Qw��<Hp;�4"�@i��P!Ȓ��}��z��y~Zc�5t�t������+̍�$��(\�бp��
3ļ*pt��OC�/"���@�b��������~���l([,Uk�-X
��e��4�ʎ��#�)ץ%)x<�}�YTө�F�<�#���pz�!x��A?�Y]5�)b?�8" 8A`k���;�"?��N���~��_�8��6J,gM�����,=�	�/D�-\�6D��R�z�-\#�i��q�;iaU3���~e�񎂜��q-Fq����ҟ�p����efՠ"�Ë�FA�>/^	@��Y�N�MqBC��q�N�ʖy�pp�g�*��R�mՂN��`�-r��0���U�`y�NJR�w%��R��ZJ�{�@��b��,�I��5~�׏������֖�h���5`��૲+A�r��b��f�cd&�z�EÁ�.1�g-���D�`L#����t��{C����z
̓���P,�����ЬN�ȍvk��
S�TǄ%�R2˃�;�G[Z���X�QJ)���Q�R�œ?�s�s�7e�-]�q[I}��e�����r�m虶v=�ޕ�W��?�sCw)aK�2�n	&x1�k8�u�:�6��Rf�.%�����[��lf�^+���r���o}Ck���W�{	J�!b�^�� �����ǇX!X2	�����|���)�w�b��O��u�������r0�Wt���C+��(-��hF�`Q�E��QT�b�m"}�mG�����D{vj���}��6j��5��[9���!���Y�,|f5.�n�g�n��,X����q5�����+�T�o�(��AoV;e7��eS��Vu0��}������U�¢ɡ��t�u��)�����<db	�±a����o�v��	�pp����ӟ��̂�Ë+���p����d(��or����oGq�Tɓ<����0:�:.K9UG�}Ј|Rf�k���W��ۇtt<��.W�:v�G͌�)�G�X����a�D^�1�]N �<C��s���ذ^�wT�,]&0Q��3��I��0�M��7eY��8|�p?�Q��}FH����of2��f���L�B���Po�
>�~�2<�l����5Iɻe�J���N�U�c�'��2�Zi[z:I��(��x��6�4cy��nbE�K9a��7��<r�*j�`�SI	[{�%d#�WgC���U�%X=S�j�%���|�`�󼟦 x5��un��TqiL4GM'x���!�(a�1C��3yQ\j`�\g/)�j���=5M�ж7fW\>�`+@ï
Z�=V���.�u���N`�g���VK��U���m��qೈ��|1�L7�oN��Jˆ2�4!0e�`�x�^<Tԉ;�ר8>�h؈C���b�v5�2���R��g1�Y@QQ#(=�^n���h�'L��QN
���9)��ܶ����5>����RxEC���u6Ci�[tP�0C/�ӱ3re����o�P�^��Q^U���1�.3��R��Qw��0^����3��XyR<k0W��_*=K�Lg���v��rbS�Ü���*G/OQ�7X��*ȫ��.,�!5�Xa�#���Ou���o�Chj{E1+��6~'�K��������=m���|�6ŋ������\~-�M�b!�H�JyV=5�/am�����r���x�k�J�j,��	[[9�p�bC�Ж��C��g�v������:�OJ,oL�6,��\Kㄒ)[�(��fDa�uJ�ӡ�+��͚l)�|��e�nʊ%T��m�,Q��m���sz
��hD�4�5!A'��KI��ә�#��^"s����6�s��XJ��ưyJII�������Z���^��o�y�����ŀ����GښSGC��-���<hh��o��W'|$��}�m�x�xuf��e����Q�`�����O���K8LQ�� ���}������í�5�U�R9�y�"yTa��G߇g�2����/�Ȅ�o����7Ѫ��Ix�U:����G;�x=ȍ�/�KB��A���?䡜��,T)`�*��}��WC
Cbd�o�������i���Y���}���u�)4_O�.��]	S�=Yz  @ IDAT`���xҷm}fy���Y{/��0L�ʮ68�?Y/����-���?��?T�ߗ�R��udl�_~u���r�}w־od�z�+�%��˾��,��m�G�Y���tЉ�?囶��[��GuXWY���Lg���Z�M�`/�����6S��5�W��:���:�M����+���i�O��Y�S��˝���~����5x�'
x��[fշ�,���P�O�Sr>/���d���f���vLG�W��aB����+m���R�/�S����j�u�I��Vr� )&�"��J�	c�M��Kװ�V��0G�����Ӵ���Y��!w5>(#B)j��vKp��1�I�k6�8�b`i���?��4��7��x��i�F���Ĕ�����a�F�[��$K�I�[%S�e��i�"�Zv>̱��ٯ��[�4�iH}��x_i�Є�;-�������/r��`�Bd��X��i���c�
�0�P�#L�j����j��_~Ջ������y��i�w�0c�*�B�b4�����e��2\�H�&��~a6�1j�����e�e��|P��z|�Nkv�+��>��W�V׿�����R:����T���ʄռ50�kVr�)P��@��!�������+�ѵ��b�N�	/m�
��~�̶+-��$Nc������c��������'�^3!�����F;+ó*�acȲ�������x���V��7L%��x���i��D����q3r����fv>i��*�y�޹y|��Æ�p�5|���ɢ�3X���bt��^��`xvQ��l,��0C�(��RXU����*fs������c��uJ��&Ȓ�2
�SJ̚��0Kأ�V�����f��T�����m�;.��l?�a�����naZ�t�"������NZK�rP`5���r%�Џzy�R'W���᫿|�E�Q(8�����T7|U����Fq{]|kB=J��������3;	��ӗ	�`x43OR��k
e��ޱ���oQ��Z����7�~3��R����G ����r0<nF���{�kk����ۄ�_����X����N1�a��Qcy�ǚq��[>iX���aF�7�ݫ������ʚ~�`q��6���
�(a]-�=��!��NG ��}��l;�%�r|��$)���7p�
3��A�t��ף'�I����(�ҋ��Yϩ\�� ���n����)a����0J�tF	�T��{���Gp�R��1�1��ju�	��N�FQ�y�:��=X���
���9eж�L;+����-=p�]m/ʁ-G�ZuY�io:��C$:���*�d�b1��Yˋ�Իr���7��W���U�"���
)_+�xr�i��8ٍƮ��E�W��L���t-��S퇻Ï�ϥL�k瓸��u��i��� ����=��9�����*wm�u��*�@_��W�-����έk%~x���w���a�� +�E�Y��N	?��?����Ȳ����I�-D��09��;v'��ь�ņq��^}��_Y��3�]�L�Y
���с�L�9�sk�,^~~�pC�]�ʞD%X"235�.��̐��7|�Y�B�zʔ*�l���;Ș���O �h�[�q�h��q��0;�c��S�i�M�\q�E+��Mi���L�5"�
��J�B��|`���8��$�d��k� �)b����Ҫ2�L�����C���AB��V�^�2}?͢v;d���������}���텫����w)E_����@2��MD�1a+P�xb�/��=[�i��,ƹ�u6��n>e�R�͔1�v������a�Ű��~y}�㟿s�5�lʋ��P��.�1A�%��n�f-1`���¿�Z�N3�>Ȑx�p�ɫ�ó����	���8���01��˔�sC������@8��oj���ŕ�R��B��0�ՠE�D8?���]/ܕ�37��;����٦֛y�Yu�k�/�1̳�z{�#��
��b��X����5/�k�,m����*Sl��_È�j^�^,Er���WL�]�%$	�_G ���ĩ�f���5x����X�ף�|���3��vg��4ef��1�')`R�!��~�H��)����Yy�a�oս�d}=�R;3L��Ű��;�4_~�p��q�X�Jx��aC1mQ��h��5���0�|�Ѿ4��m<�Zªa]�@�8��"Y^W|���:�ҋoX��}���͊�^�eM��+�j��Cb��{)���srk�MG����q��ݬ_ߥ\=��0X</|�u>��j��`6hΚӬM�!��S��w)_w��z��"�SҬ!�z`f��N�J���˿�)Z�WY�Qf�F~^�py+���|�2��Ѭ�6�ٔ5������U��{	'�(�1�úD������%��0�N��β��e��ɠ\;�ՃHQw?�1��>�}��?4�<}��p��4$��p�����%^�Y�Y[~c�Q�>���gȨ��6�σ$~�0�N�-����	��:��I�ţz%�(J[�KZ�V�~~�$�u�@׃m�(`ҙ!��`��R���Sؽ-RD�*�ᤞ�˩����e|����I��J��X�������ڧr9Jv�Un��"T;M��Z�:�E��r�+��~,����|O�)�W)`�ɇcC��-�Yj��$�o�����k�x��ן6��֨kˣ\X�8ͯu�Um�+}yN>�;y���S�������u輜����*���ĕ���N'ϕ�$��Q�*�:R?\N���T����'��-�Dnu.�c���A~^��J�4�	���o�����eJ�y�kL�A��v�i2qx��y�w9D��� �~���
�Qp0�1�n~�F6$/}���i������Ǳ�A3x!v�aη�̣'zb	�4��|=R�fx�Yw���[σ����b�k�����|�fx���ݺy�|�J޿>|�INǑ�Ŕ�mR����_����a��T�"VV(>.�6%�hͬ{qژn��gV+6n�꥘���a	�R��AXf�����?���y��Ə#|�Mi@f�YO�Ņ}Ť\ϑ��L$�aAz�x�����&LGP�a�VJ�F�`<��zK��-�;3���j[��W����㮗PY1s�Jo�J0��*<�R/��UӤ�e�H��p~��f��˕����G�=����aF,$7�UgX������@8?�z@�ڬ�ի��廓"w����4�(V�W��P�4ɩ�`�|���Cݖ�Mh);Ƅa�ԥ@_ɯ�f��α��J&-�
_�j&\�9�g�|���M=��_��u�8�`��UH�)*:-��',BeO���L�a\����d��L�����u-A��RKvD?e=�k���H+��:`y��!�Q��MZ����x�(�dV�/�;�Ͱl�d>�[��y֡�u����I�U3���u�^|�B��]�֯�N�:j]Bk�M/���l�h�r�����nV`4,c��g8k H�X��_�����%��]OR,��pv0�)^c�&m^;��W��5�M�3p)c���}w7K��Z��X{���
�'lw���,��b4S�ݔ^8�n(P+��SO^�Xz^��(�|��������e�����ry�%Y�R*�{]����?ԉ��!�W��ه˃x���v	vjh�`����9m	Q?ÿ}�MO����%ʂ�V�y'�q���/_4�l,�����ƴ�ł��N���IC���\������8�!gO��m������1�M����|w��t9��z�`��S7���>q�6���4��z�����\KhJ�E�щ�T��8���O�eZQ���-���0�4ؿ�j�.��ϔW�:���	]��X�({:;+/H��Ѯ4�;�����)�T��:����u��]N.p�����#���@��/>;|�!㣏�K�j��H�5�H�`ؖ ^�X��,��#��<�j�zt�w�o�󺟍���"�)��Gx��o�Ng�B6�U� z���:k��?K����_�|?���1hiGǆ�4tD���2G[��[7L�(�g�����k�1hT�^d�NC]�^PB �}������)J� �4���
�U�,��ק���SdfHn�R�ʟr �3����AIBo�a����>jX��n'Ԯ�}oz�?5��<�fY��1(V��G����`w��j��J~Х��Gx'��?|w��6(eyQ���h,`M���˯���(Z<�1����a���^�1.=��z	O�64Uo޾v�Iq#�/����+��Y����e�Ð,FKȌ�z�� ܝ���U�&(���5���F8}?K����P���Ƌ����r�e�y��+����/t9&{l����C�Z|�.
�L�gg$��L��k�bͬ��q��`���Q C/ךn|�p�͛Y�3΍��W�7�D��ᇶ�!X녰��o$ ���h��zq3$�U%�t�w�=��\9S=��T��+ ���,L�R͠c���:L�V�����ÏR�j�E�F���ִ7
��cQ�w�����q���e9�e��w��t<i;'3�X�VG)��=�.��eJ� P:�<�������Sk��i�U��7�1lq3�Q~���YfA:�+���C�v}W���f��E;2��
�a�k����k+��~�0=��穣����Y�B�v��Y �?��E�ږe.f�3��˰��s
y�����X8�&��Y��E/Y�Z[��c�6~<��a���C;4�aO����xá��-��0�[à|f���<Jh�e�c���~CS:��ͰK�ϑ���)�,k�H�XC��Z[�x�'ʘ"Z2��?�T|m�B�v�b-x�og��[�n�0\1�q�-����Ě8�B��XiBaU�ĉ��f�Ӌ�7�"2���|�x�O����]<v�Q������Ӽ��$�bl�S��8�cבgR��\�(�����N �>a$����4oV���	~8��O��������u�[���ۋ�Qxz9C�>�p�n"��φ��m��%����5F���1מ�e_�Vi�u��C��hD��#�>��EK�(=�O�h�/'@KH�g�I���#���|v�ͯ?;|�_�`_'�َ�,G�	�Y��y!����+�)��Sx�[F/�-�W�� ��+�⪚��J���^XXp�#t�hO�Rp�;ް���F�G��םJ�Zb��Ad����׳��xV��L�ҥ��^��N+l� �����$���>�����<*�bA�IO�&ˀx��U��3�Uo]!�
��}i��3��E�3O:��C��qb�[�o�6c���?H	�S�~��{�/2e�i�s���?���Ãm+��3����,~�,D�<��r�.���C��4��Q��E*�K�2F}j(�Z5-թaP:�L���W�i��IO%��a��4��:�Yo�B�$����ƼQ�r]x��Gw,|�K�4�5?O�`:�;JN��L�2l7[��1���	R�ȎS�͸_q0)�Y[�"7K3�#�J�{�EWr(��2]���I`T�+�(�k��cK��z�5��ʣt��yJ�9��
ܮ~O3]�b�M�j��6�h�mX�a�C�Si`B�6|���i[+4�k֐5���ywTڳqv4`�8y[��3q!Ƴ�Y���S�9k���pgi'����Y[�W�eM�����_6��������:��gx����c������ȴ��R���S����s5֖��X�?4_o��E�����orB�����C�xX>���r��QJ��rN�U��Q̮6�غY�e�E�V������L!�#��b��A��XMY�ia�~��?���Ì��-��Y��K�/���!��@���IQ<;|��w3q�r�=���A�j[�F�
���]-���X�sU`ţt?����j�K�Ǥ��9�p�x���vG����ݳ,=X��c����~?�t�j'�"j�Me	��	�jC'(�w�?k�B��[*����ꨎ$Z�TWu\�{���)ϡ���gŋ�:�y����#_3�_[�;Jps�0:QN��5
��aTY�<�$����>�� .m7�L�'[���A[(���۝��Џ`s�.�8���_qߏ�/0<8��y�q-~/G0�8+<���N�[��"�����	�%�L&�ɵHsݲ�p�/� �}n�3Z�au���.����T��@��F�{�z�<Jc������[J	�Pf���]H��qxf�9�m ���WP|j�1��:X����}#���z���������Y���g�=K�Na[{���ε(ިce��@Z����Sr�m������Ⱦ1ؚ@>@���B]�U��Ϻ�Z�.�  ?^8Y��W!�-=��rVgR������?�o~��xi� K_���`��ެ[�ar���n1����$��N���mȆf�wEe��@{�)�����!�gL:!�e�cU�"ة`�3ģ�'�	�5��]%���_0g��?�^��'�`�-�yl���w)cwZl/K�͛���/��`�OǓ̡�9�M�F0&�3!�h/W�����|`Xi��7�fS �,3uLq>J�&�Qi[�1�9�Y_�Y��^C17Eƥ�����9�<ke`�����,��Im}x[���8���y�Qј[��!�������}7��$��pVo/Z�¹�	!8F�ˑ��'(kvE��Y��|.z�Fr����(�`wu>�`$�0K �i�XØ��g�TSL�{��ꆜ_g%��NU0�#��Acv,/�Z��2���A��^���/@0���I�xgH�e{&d^C�p�Q�X�40
~�_9��:��)V�׏,��
��j3�tTzϢ�����Dx[�c2}�Ys	�Y��f�����:�I�o��R �j��5�������R���~��o�w�w��?������K��뜬M=��E�P\p�^�{~���c~�w�g}J����<���Vڎ�f؟��A�E)��4_ԥ2W�Gu _|�c0姗��y���ȫ)��u�f�������e�x`h�������cB�� ��HY:�i�	���R�AꈰJx�a~t�3��"��$�ᡕz�,��⛔յq/8C�zDf_Os.N�1�0D��S� {e{^B��޻p��F'p�닱R�ݐ����W �6�,M�^ �_��QС��p�90�e=-zYʠs|!�N{ՀL�ͤ	���*n��^e8u,=�Is���f�[��̭GwϜ�ۻ��ܯ��mR[)�}{��y���Q{>{�	8��oBh?��n���P����'�ͫ	�'�6`|s�����w`���F],X�͞�k��G�X���8C@�j�d�(��r��~�&n���>l0/UN�=^pW�
:���)��O����%D���l�E'�fA�+1�;OS����������۝h�徑�x��г\qf�ڤ��萲�:�x*���L2BF1��7��}�Hkؾ&'YF�kB�����c4���hpS=o��U�Pe�F������-����=�=����j#��A���27o��Y�o� `�Z=K�a�[��Q=i�#ZC+k�=X�{(�Xy�1-�+� 5���*~'8� ����^0�.^̺�ӷ^լ؜�ƽt��,@��6<��2Fx���d�2�x�����~��yc�����_����ËV�VA�,�U�ᰗ-������e�"�4m,� �L�Z��1����L�Gi���1��`勢7�0�����~y����"��܋ ����}d����GK1�P( ӛ�^>�����1�"�|}�ů������M��B��fd�d�m����F�.�a6ۮ7S��
=�axhh��UV��U�Ը*	��W�p-�8��zh�{xI1Erӈj #t
�cl�d4*D��-ͺ甬��"����|Iq~U{�<4���d��Ͳ����J���&���ߗ%N�Q�&Q�j��S1V��ҳ��%x
��kRСu5���{M����L���b��@�ce�����&�a�$0o9�痖r�\m��e���S�e48V?��c]�׆{=%��e�Ni�E"�m�5�㩇J�������󇬀�̐�a7{>jw/^6��t�O����ʤ��l]�?�]
ړ��G3I�]5����W����v$H{��Ұ]y��0�!�~��ˬGv%XC�aϰ��pS�y
(e��WZp, ���5���Qtg��)���Oi��+K���>��ү�f���}h�$u�~�ϛ�^�5�����R4u�\�j��{��,��Iz�՞^ס���g	��I&e� 3�,�(��-��%nd0k��(z�&��Zِ�rPPuL3�gOP�(�r�@��lx�.�+<��kkˮ`�M��<:Q�S��*���t�E)��\�eT9Ѿ��}�z)���|R9��:�. �V���c�/���h�WT���u�^!����	"�`ld˛�WZ�IC����g��/���Ľ��t�tV�ׇo�,���OX(z�$gr�T�7**-f�	�y�:V{�v�S���U{�K_�'{��'�����ċ=�<�+�drcW�\'��u�n�$��'�����~�v�ET��l��"�Rb��>_NV�-�lI����r5�!�h/LV.��,'���2Hp_�ö�+��GOf׀��-���*�pԫ.�Z�*9�*k��(���=&����iF��n0�u�SFi���;���:Cx����� ηֳ�އ��1!Lӌ�+�!���0��h��T|���)�*q����R����̌k���HC?�bp�`�2z^o�v[>�g���(!� ��p�%OS�l���0W>3��s��� [;`3~#�U� ���`*��U3��"t�=O��P�A�}5,`4dr+��VV9
�=��E��;���A���z�|���i��=�(wH�i�X��)M��aη̟��"�-_�y�w�G�" w���-B���r�"8���L��<e�����H؞z�Z�f��|��Lk�`"ᤗ���'�-x�4g�%�
ݳ�v��z[/�z-����nk��(?#L�~���Z6�g��|J����`�.e'hF^�vB��^�ӫ�\N���`�cR΢?a��ҁ��e�R<����$xį����i,�Qzz��e;뛽J	y��%�m�t�a�rՂ������q~)��)B��+�r<�J��7?����ɰv�fiQ����4�zš��T���T�Qb����usp�!�:Ӯ×���5�\ڵ!�� ��������e��O�̄��Q�Rn�j�[Kہ��b"�`F�)j��#�ae$Fy�5J��O�(k�d�5.�a�j"��9������l-8(J9Z�u�/�L�n�dT��V`�xE�7�Iw�`)��$�(�Ewt�Ԝ¬����G_{��\g�bKPb���){m#������NV���Cm�����ݼ�n�����p,Ǫ�-�Ii%�RXmw�ҟ���-� W	��-���&��JQ�˄�f�m�S��K�[����e�p���{s���4��p��_�������"L�}�yZ��W��-i��v��}�:�׷ށm�$�l��B�ԣ�i��� �^E���u{��5\x�m!&�X��r����pJW~��8bl|��T���g�����~v�UW�T/20J�0���}Vg�/��ڴ"�83i�ޒ���)`c�*_��kq�J/���ih�4,�Fo��E+�F��S�OnWy��׹e�&%qa���l�<;H� w:���g̸5�r��>i�l���J�9��~xz�Ch��̸���6�g����l2ʇ��a4� ]�C 3��.F��S%�Ф�ɓ������d�鎃��0�ِ���4�0���ڂ��i�I+ǌ������>�|nNۆ�?�״��S�B��-�����Y�ꤷɊ�	8�1!�\JC�FA��<�#�@+�#�tT"�N�|��+%�O����ه,�iΟ���"ja�'1�wr�6<4C����w2�Ά���L2�9�`?h%����Z���M���T�����C=�0ŗB%-
7����!�ٳ.|�h��俆HSqM�/��$�Wq�9"_��%��;=n�׫އ�tM�J_6�9[/Q���@�%�L]LZ՗<�c�c���uq(��f[��<ZG�R��K_��fsU��]��>��lxWp3��zSɊ�v7x��UC����Y�G��QxM�����U��r�$߰^���s���aA���j2[��GX����l�E2��u���x|�R*jsS��?L�6�.���S2^��W/R��X��}�������~\�V�|��D��nh�ڀ��4ZdS{�k�Q[Ѯ_�71�zGᕾ£2�(����]\��2�)��m�5�:/��@Z��@4y����j�1�!}���r�8���g'7�l|�nch��|*P��V�k� �Vy4�iYra%z�3�[Y�ze��bxgضD����Q[���la�<Jq(
�ȫx�X(_,lcp��-�+���t��gñ�Y�����(���rR�K	Zý+Ԏ7��?§pmݟc��ܕ�b)�:.��)��W�l�u�j9;l赬�z�t�S0�n� �$*�C�]����q'�2^�C���4)�������d1�{���%���s��9|½\��\�����a�b�YIm����U��'���`uV��?<�v99T��pp�~�R��v�8���'PF���Wٔ1�M/���E���*��}��2�_�S���z}9>����������os�i�ňFퟜ|��+��z��ӟ~���VK;���hRdL����\���So���>�����-fF32-~�
�ʇ3��U~ߔ��v���3օ��{#�CR�hurۄ�]��Nuɣ7H�vo��������F�3�5>{����F<\�|ȫ5�n~I/k�cԉ��#���J6���J��Izg�Ti���+��㨱_N�9!8�&g��x����R�^T�R���9&��c��pY�0|�ȧd�2�z�S`\>����u�Ժ$��j$�+���z�U4D�o.��Y%L��l���K��֭�4�� �	����￨�N�i%毬��h�����)NmP���iL���l�%�G1)}�����ӫ�ϳ�XTP��aڸ5n���i!H+>[�ق�V����:�^������P̖gFqFX7t��	UK0pbWËOG�-vu�r��KG�{8��^�J>-�a!��8��B���WD�֊4,��ʷ�G��OQI܆���(��ZV�Q�k̆4/�|Sg��\tZ���4
N��*��M	���t,WBh<�1���Y��-��ge'��i�J0����HƂ�?��y����9YW�]
�9�=)f�������l[�5(��D�=���|Xg,LL���Y��o�S���_�3?0Cgz�pM9�w�ߥ|ќ�����gH��I(������j���R�]�S:w>Q�<�:/�Y�L��ݢ�U�+�Q뫇o}��Խzh�r�^�;���2����(SwpF���`Yu%guڿ�'��
ͤ��i,E˰rJ����{C�6%��k�hA-�b�a��K�g��,�5.�Y��C:�\SP9����t���΢'âӆ�
܃�A�*l��ٺ�����(���#�Dq���XA��� 8\q�Ȟ�����TL����]���ވ�}��Ôc�{�`����#�>58A���q���v�&���3%��ҙc�[�����n��(�]糟U�y�Y������l��)0z�����E��%`��k�ʡ7ݏZ?�6+N���;��n���𸌧�JZ�wթ��*S9o<s�">:��A���D��uB?|���׿�E���GQ��D���p���n��|���[�q�`<Z�r�J��agk�K�E��+L�G�\m�].7\oX�F�)(}�R5�\�z�N�/m-@X#+���0��<-�s-�$����X쇿/Y4���$ƀ1Ʉ�I9B�+�^����̰ŦYE���S�x%f	Z�^�8�؋��4�����h90����,�Bc,Ef�q^=MȘ�x�����t�hc�+��Ę���J����g	��!���hhϊ���n֟�h���;J�y�_���_}�26�_��Y�����&l0�0Q>	��n2΁�A��Ǥuˮ&��o��]/��?������.^����O1�K������f26>�S��=��Ō��y�襎_ǤK� ���$�^QWKM���y��?�a,`�\EJ�x8_:�/{�Qg(�t�m���m�#�뭘~3��OYH/E+�a�uB֐�U~Y����B��زnf�lX�p�`��L\s�z:�N4`v%e�u*�����N�r�:�Dk�f�
��Otj�M0� �t���5��Gx����*t��)����pO8�ϰQxJ�� �ה�5����WنDȪc`�x�:`�)�f���E3�El�t@�J�DP�'Õ|�(S���_Q������`���߲���77�l��dzپj� q���Na�L��,�p������:*X�/K��IPP	K�<�L"�o0Rz�zD�Q\x�e����=��N*|,KJ��������ed�ѷ�۞,3��=kU�y���<�m�e-\([�l4%���	��Oꆂ�2��,I�M;7V�Y�:(�^̤��`:��-�9
Q0�8�z�z����xi���+���.L�Wt���ǳmŏ�6>�Y��� �%m�3?-���A�^pS~����N����T���ʷ0�
��|���2Ǽ/\e�%e�:��N��c��H���ۍt %���;�~���[ܟ}*�|�?/��g�<��|�/[���o��� ��1�.����w���"��ۛ��M�����㽴���!��i?��z��i/���'e'�ZNh���o��ޢ>a�x�Y�M�!�X�W�x��0ɂSY�O��U��j�j�����i4�a�k�e}Q��k:˭ك~��ÝW�7:dB��͕�z^P���ֵ&;xZ4\���	7
�2��%��5C����b����d��ԍ���U,��b�|�53��5K+�N��eE�k{xYz���H��&���La�>���	�4��0���L��f[��
� @�8fB��	����n��2�	����p��p$�L/��1�[̈́������}0J�F_ĢJ���{��v!>��AX.% i�3�5.�:/V���0��;w�Jha���_�����֎�'��<M�7[�vF���Lō�J!��3��Q��2��+B���Z).��\
��A.5�ex�d��y�jV��U��#�sq�C���)�B�&?�k�N�c�w��-][n�Ќ�fW�?~��А ��E��sC^�ﲀ%��@ �$]�r��az���,�X�U���p[�1���oj
Bg=�pYĵ�\3� uDC�P�ip�}fA�E�U��(��o�P\��P��Ux�:KX��=zPC��L���k�jCs�[_�J��cˑ@�&��+�E{���l�0��rƼ�C�O?���-|�5��y�0ц�{���׷M��M�}���ܐ�e.��(+�K4Y��S��1�Ro������y�������m8Ń��)6���N(!�R�I��F	S�J�7m�GHY��R����{�ٻp��t^
�f�#V�w�0�=/��j����(�y�L���(��ye����zN��e7��(���%�h���I	.
�8�� ���]�-|!��|Ǌ7������K����h���/c�~�S޽�q�?,A2���|ɣx�/N���k��z����Ȕ�t��u��^d�ز�{��-W�E��aY6�B����*�yY�n&���|�gqa���(g��S�bm�\��O��븸��G����}"��N/�_�؃��Nq��c���,HW9mHf���R��2��J~=���2��d�Q�W}���z���z�wo�/j�\;��`O]�k����]�c��o��Cyr݋����VW�$G�yW���YzX��f���)/U/���U�OO�����٧Ƌ�c�8ف�F��j����Cz�N�T��*c����r�vA��W����x�o;7Nq��xG-�>N���&\�ZZ�D:{�[�b�/m���z����jג�\�`�P��DЊ�7Jk�c.?��e��1T�L!�����H�3+��o�*)_#b�	o���+��1=q��
��8�;�+P�8����G!����3�-�F�� [Ew5���!S7�x-��J`�{����䓫ƟC�����c�)}��f���_�O����G��Sii��,�o�O#�J�%�4��Y3:# ��� ��o���!�ogY�ڿۢ�@2��e��.S9� ݣ�eAH��`S����7�:ʖ		`�����w,���=��m��
6���XC��ߕsz��@�`�Nt1�D'��)��O�~����Q�Rߒ��f�S6��η�%�j
��:=)ኙz��"�5\�Вo3��D�1���"S�����2=����;�`��Z���)�j���X���U������O)�w�Nn�6�����A���m�t������H����7�R�2�˷$���L8�I]���öm����~r�w������h��k�1����"}��^o��ZTԦ޳�{~cW���>�aC�&� Y��ɡ�YX7_�/��݇+`�>��k�������M�͠V���9�8F0�ɺ,��G�,_J��G�XM2_2�z�ۂ�~V����G�K� LuS����Z��[��F/�(��¹���Q֓��]��h���E�]�O�@u3m3��U��E[[F�Ъc��^�f/)�c��~9JfyN����>Lh�����Ϩ¬�(�i[.�2���y/�̀n�$��r�@g�G�Ў���e���-���D����?[����N~ʱެ���V�Qtuccf��|i_?x����,�Io�ᕀ�1%�\W�9E����s-D��C�-Λ�z�J�v��EY�D`_Vo����T�'y�'���+�	;觇��+ޛ��<��(?K�G0��{Ǜ���&��,�{��*|_���jZ��|�iFV~z���R"����!��[��Z��'�W���z��5ș^a���uH��V�r~����>��7���x����6ry|��%����ڲ(�G�2yӁ�b`NI�ȣ�s��f�0��,�-|�`D����4gG�-���B�E�7u:@����j�u�n��M:�R�p��3r���~�o���u�p=x1V���BC�4�4DaAL
k�%�%&&~Vx�,CD��S�#��,�Ҙ��榗S��R�u2*�q�4\O��~V�C-�\��$D(WC�5�h��n�#��,ajvS?��s<�&%̶�B�Y����Y�^F	������"�ɬ0nO{T^g������tٝ���,���a,6����.±ЫM�_��N�ba��m��<m���(�g�
��!i�l���?oCb����|�¯C5��͚b8f���a�����Պre�'f�{@��f�4)�fx�z���U�,0�8	�L�6\�(R̏��7�r��ᷲ�eɩ4O+�v�ѐ��v�(�2��͔�����A�^��K
pp���gm\>5�j�����M����H�e�q?Oѹ����o�
LJP���z?h��y��/,�Y��V�Pap�9X�%aX��(�����w!�n?d��o��ml�n�y�)��:���	'V����V��y�߷�W��V�?�!�Ѫ�2�ki�x�L������ig���sZ���]rC;�e	�X��i�V��T�Bg��L։�.��M�[�~Y��Qx�Č��r�S��+@�cm{�y>��wNlћ�h��it�����]�:�����"	�"�0<�4d�!��]�*�K�!���)1�wy~>�5�I!d�U�M�L��j�[jh��Z|��)����C��R'��k�|)�X<w��(`���ٕ�QyZ`�L��e"��O��AS��Zf;���V�`���	�2d�d8�[�XuO�|���Iѹ���)��2�\�=��`⮰~���F"��8�t���T��o�/�����Q�_$�ś��仙��4��V1B��p?��i�4I���}�i�0��8x�@֤��k�|�,��+�UY*�>�[�0+�2��������ao��N
筶�|C��-C  @ IDAT{{���Q�N'���:G�=L��3p���_f���y~_g�	|��uԒ|J�\��>�7����d<ЬҨK�����{a���c9��&���������`�;��l�ʯ�t�+�T������m���W��/ �H}��P0Ǭ���/�R/�꜈���8j��BX�l�9�<Dܻי8�.�m���"��䏕2��ۀ������	w�-[<��-3�'��tx�����t���P\����kV�J�2�#���q�:+�1`_���4��׿���D���?��p���h��3����+x�p�2Wf��/���L���@��`�G^'aw��2���*��cF�O?]:�����-6��4Í�!c�Z�YV,R����S���U��c�6��_��Nf�X�8��G#a)���,͐��jf͙
\���ef�S��P�������s��JCx�G��������iG��3i�f�~��O>m�A=��9��c��r�
��,`��T�V��Dd��3%��D��Y���D�x�n�_�����Yݒ��o�%���dK1{nE�����׺3��x��~���Z���᷿���7��6��b:�7����B�ij?��-���Y��w�s�Ǐ��9�w�+Yj���f�<�|��X���@��j�ך0s|z�a�:.�,C�6ǲR:�5-F����q5��)�+}݈�P+ߣ�{f��bP�b|���ơj�&ɤ6x;֮'����SN�5�V�6�z�17�
!ł%x	` .���(*���-�sE��L��Ҁ����@�E��8y�"4�N��c^� mG�hh���N@p+v�����ԛ/,��&�K��I�p��1�V�+@�$��ꧼ�u/3�%#1�\�w4����DUf���TR�F�	��{r���?O�yi�!x����q�9{?$1��L�=����f�����g�z��:u��S���R���	ϣ�/���F��N���BnjdpP�
��
~�w��e~��3t]/Gq��l�
8�=�e?V�Q�����|K��k}������+���O�S�Ҝ:ݳ�u˫�@�da���%�~�������p�>嘿s,B�;�F9L`�k���^��T.��]iM��9�z���+�A�'G������91�a��	�=X���+�ш;�3���Ǉ�\�"Ռ<Y�u���#}%�~P*;�����f��+��}�����<�)�f�_z��~���������i�9�`t|҄�Q�j��}�
����|'k?% u�;$��S�o���^���h�_�;�(1!�c�O4�^�J����A*k��O`���*��7����fף
�[�V8����ݓ���9z�����aV�L�T�����.��[����z����{���G�P���wm䝊�ظ;�M"[(�(A�B�u�J�l?M�u�����s�z����xY��P�Q�uQ�����4=�Yѷ��d 0VBJ��.J�~Z��Ptb�D8�6����W��%ӊ��3	BB���ȡ�����(cZA� `9�!��Y�zc�z�{�T�jP(�]Ϗ�Ӑ_#��@�,,
eC��+m˒ ^�f����4��igMs𧬯�����o�VYV=kd��� Q�i|��au��,�+}��%R�7��e���,������~�LT�Y��/���(v�?J�E[`� ��¤;��:XD)�9��F�]���҆�)ۆÕ�#�gՓ8�l^�VB�0��1n����5��z[�mx[�e�(�L�\>7�����p$�����R��	X��`�[]9	~�]�)]:/�0po�TR��6��|N�s/]�n>N/u��yY�1H�)#e2���I0�4%��E!���2���~��o�5Ac�(��:�|=Y���/�~�3L'S��bɕ�v�*ޗr�D��~��H���΢�:���[
�!@�ા�_�9��g)_f8�j��l�U��װ���X�KO��Fw��u��8C�c������(~X-�]VwK��%���\n����R��ܺ���-l��^<eW/�~�zZ�O]Gq��/��W��������Tb5"�:����`����yWb�y�ZQ�'\i�������me���.��wW�]Ź8V�+!�)�ű"���=�7�M�+��Ƥ=F;���J�����S=�]<O��pTٌEzb���s_�X)L�����R^�(M!k��?��ˋ��;� J��)��^�܍�M�'�))]�G����W���TZ_�(~��N|�GE?���r}�g�[9P�����Z�c�;��SWC84��уq�z�܋�`L�z�P���|�P}SA��ΖpW�<�뫥��g�*�ҍ�м�«�UV�5��ƭ֭괶�Q�i��%ua��V��*\�t��^�!̽�"�!�t�k���&`�&��1`��~�.�?<����Y/�G�~��|N��P&)`Ȯ�*?3MK1��g�� כ�*>eGo�i�����~++%�0���m�NN�1݇Y-��<ςc8O���j�5�X�(�'
6���4_B�����g��,qQO�7A`Y��a�˞u�@L64~l�{��RJ=^c��OP���Wu�}y4�8�[sk��������M����`*��aD��5%�~d�RT�E�5C}����GB��$��-��(�GshY����`���q��F�_%��h�}kf���|�l�X�Z�,; ;��a<Y�2u����Q���܀)V�Y�t3S���|y���ހ��-8�A�G�:�\�P��ې�{g:��,Y�"�����o�o�>V
��n�;�S�����	.�74�΢����J�z�p0�pD�W:��K��w�l�t��Q�[�?F�S�uF�̾��2�U;^�;|eP?H�I1)Le7��Ce���ˊ^V:�|`DUk.�Sp�efZ{H!�t(NGQ+L�V;�ڐ�P������:}���f��';8����u=F羕֫�(�޴���=�k=!
����}��َ-��BD�3Q ��d��v����(a�1�rX�͞��1E��*���u���M^��e�3�N��(fQ�Ck届+�����P7��w)`�G���N]Ǫ����N�_�_%�U}Oˢ�:
>�u?7�R<
Ǌ������]���`�}ְڊ/�y��`���V鄿P��U���=�r�M; �@�L.�Xd�U�dԄF����tx)_T}�-�����F�ï0�B�rh��Mo
���l��&� t\A�Y�Қ<{F/��,>�C�t���5\�_ŗ��d̒3a�̴YH�ʜ\^�6���|�O��)�#%�hƑ��X�o�ݛϋn���eW��Y4ȭJ=�E��0����E�]`���H���q�Q��G?P���*�Ńw� j�&����dם��~�{@�B�\���aI����1c�c�*6s���޹=����[	�M����#/i]�{����0���^������qr���x���"]��z3�>�
�����nʊ��q�$�_0��H,]�,��)߶*���ȟ�q�M�עo1�*�JBְ�a��o��#V���Pbv��E
����/s �O-&�ে��=L��:R
O6��¸�w����J>��b���ë���M+�6�h�%XТ��Z+���ޫѝ^�8�̆��~9�|-47��@u0Jf�_k(y��w��b����e*��|P����S��'D���8��
կ���\`*c1������^��G�n�P�ǌ|�Vѡ���\�'��_� ~_�	)��W1\�����w ���i�?�|�Ԫ;��PUkY�wt�0�y��c���c��%ت�f�Q�Ks��s�&%̒�7+��𩼎�w{4��[o�1�Wh����s{�1�ʐ����b�1�-�����-���N�onB�9�m�MJ��٪4�I�"d5�ax��.xF��$m�!<���N@0Fp�Zmʹk��($):�7��}A��fV��lE��t���;V�|��hS��%�\����R�r ��hA�/�C�(E�G畆j����Ix�W6���c����Y;w����E����(�-��#�C1�v�E�n=[���H�v�2:��x��ٗO��S[�שS�Ҟ�!��c�My�Ǫ��	�(��P'�`
<P�x��0ނ}�[��;i���َ	_�	���,��{�|Dz�ߕ�����-�.N)K|��x�7�z-��o=�:p/�ee��ޮC,+E��X)�ub-��덎��>V��fb�.�ds��
�s�3ч{G�=h_��d=yNp	HY,\mJP�]��y��ֈR��@ɞ�Y�6��O�ՑM��Q�t�J7K�>�Є�!���ܕ�����z���w慯+�z�>����X�_��=Kr�|��2L�Ǩ����N@��<���Y�A*����x���{�Z�[/��vO���WF�j͔�����/�̒hf�V4A���L������̀4H��jS�-��.��S�-�^|�f Y�݈��W�t��#/�Q���9ș�YEB�{M}�����lY�f�B�I�6��iJ���d��)A�f9�lb���}k��m����C{̒��F}��զ��GM_Mſ|�^B�O)3$Ec���㶍9+sZ��J���u۰�y��~<��/���ӆ=�j�fT6����� �k ��0@��- G)9+C��>jc�?���~���4��$����|B*�L�if�G�����u��|NY��=!l���,`')`��d�9u����z
��Z?�g3�*~�35V��SNO�ޙ�A����|��(�c��&y\o/��,:G-x�<�����N����*�-E�a`L����E��ey�0�f��(��V�KQ��>V��ynX�`�����	�Wm���e㧕O=�o�@�Q�X�Ϊg
�;�XE�aj��9F��SJ��-����Y���Oz_0NKgY�JB�l�Mo\��wp���W+ǮxYvd����9�wJ�Z�	~N�Q���,��`�5�i꡺��3�'�a)!��/�Ҙ���9��p�ЄD� e<O+_�����L}�5�I�Ճ)��h
1��b��9K7D_��t5$o,h\���5�L���n�-���Q��'�_o�:u��eG����&��\>_Y���j<>Y�	�_����/57%p��#r��<M���k7�M��v��_+��jh��}���'ڝ��Y�(iv|0���zf}�T�ҳ�z͓�U�1.L�W��!�p�ꐢ�v���V�|���	��s�>澄ĝ�����~�	*�w��=L�ni�L:�o�].	�u�i�:���:����:����eBx��=��c�p
�
$dgy��qg�������"�����$ɘ2����~��W��qRW�t��ׇ�UttK�s)4Z[�1�i���,d��g6פٻo2�tr����������]���N��No
����;F��vO�/48��Y��#<;�hsd��߽�:�נ����<؛���[!�d�u��+א���̌��n�6�xDC�����YC
�ҟW�{��������`G���\Kb����G�3ԓU	�&�
JPu����R�޻Fc�N��E��v��`���-:�� !������K-kp-��i=����W_�Ԅ��|r�h��
�٬KSr�Y!�/��Ys-?�,z�/������p�����{1�����$�g9��j(�6x��칯���Yv�ZH0$E��qq����{�aP�pV�a`,��?��{0J[�/��uѾKq����r&H(�O)���a+�����T������P��~S�OM˭��_���iP
/��VC_s��cj���{1����4z)�|t��(b�	K"+�^�q�^��Zs�R߬�9�g|���+��v�����-����f�F8_�+ey� �+G�.�O�6tc�7�ސ�a+��b1�n(�zUk��|�G���M.��`��X�&%0)r�����a�(R���w�~0�a2�e�L*��eC篮F#)�S?SW���YrB�M=���_���U��et!�hp%B���b�HN[@]K!w.k�d���W6��I�b��C��r�*�Qf�~�8�b D'����߫�������� � �C�
�]S6���Ktz�}W��S���p�Q��Q�am�����){���<]iͺ��0+�똥N�>yϺ6�P��%+��s�}�<����כ$s��)`���/�F�OZOy�ޥ��8ܨm;YV���u6�����
}l�7k�3�NK��Y���,11H����_� ����`�R�s���c�=��[�=�%%��G����ݞ�
#	u&�u?7o��i����N�k��0{�� g���߄ߋ�v�r��:��g8|A���NZt3;h���c���%��q� �Jr�����
����7�������6�����~��95׊,�
3���:��"g���8��n:�-oJێi�/�l��.o}�ob�)���0{�&�_�;����D�=xfgȰ@,���� � ����8�2�
�σ��=͟�Hkk\��a�����І&���t�MB�����)A�7���~;É���Q��j��"xOn{Ყ�_��jhq��
�U�%�[LS�i�E�ޝS��<[/�<���+1���8�Q���Y����W_}�l�Ŵ^��j��G-%�4�ΫǮgr�֭�-2g5`ӝ�ʗ#�3��"�Y5=�9�Ճp�8�8Lg�j}��Ԋ������ru=�s�OYz�̾G9ϋ|�rt��p�G�6�w���ӌK���	-�2z#k�]�呂�4�`K��Y[�K�zv�w���Y+*�U�`�(4��&��pɒ	5�ݭ���>ɐg9����J��]ؙ0�JQ8�B��ޕ6����hh�x�*Ryg�}�p߅R�LHIە5Eg��w��D���>����|�i�(K@Bö�m%�侩?��>n/�.+m1$�B�t���'Sp�xk�3#k�'���D+�Ugiכ��0qJ _[Z*Ǆ(M�g��ɕ���Y��Q�����a�4��U��?��dؔ6��{�K`m�*��5�k?��eN�ô���(�,bƗR�`g���]i�zWޔ������A������H�*��41�k���h�%:�,d��:�GA:�(�< �{��9f؆Bc���ڗ�8�6-�{C4�%Z���V��Jp�_��?!�:6r4T=�{7B�[���Ȣʡ���Ű���bv�`��=���:f`7�i�%��O뢸�4�8xu0�r7ֻ֞lf������4�+��ً,��P���o����x/��nT��W��"e�ř��Y��U�fx�	H�f�F�Ã���5
X����?OC�f��|��sƆE�@1s��x�nT�����ە��L�������m%f��U�{����a��Cy��o��nO����%�-X�N߽x�U\������l$X���C0-�"��(&���Wfd�e|���f�zm\{�p�T�s}٢��L���Ѩ�1��&XQ�����.y�c��,^ƀ\<�y0�Hߎ"��h���u�Uz�*�]��j^����"�ǺE�u����"����x��[Y�L�IgI�<@���\��y�[w��o���sE���*��U��]�d��*@_6LIˡ��6i��ü�[9���!�=�����(�n~'�n��Гvw�yG�ƨ�qC��xL�(Xi��t�zo&�)`S8F�i^3�jX3�XC�����a�S��=]�,�KP-�2k�Bp5�R0�) ��5��3�(<��I��e֨��k�����e�@�T�#(,��
6�׃��­�7θ�%��rVe���Q��K��$�����:�~�ʎu=��.e1;�V��l�R�����u�R{�5���"<���Qj�$�hwx��ZO�c�E]ͪEIRUʲ���blhLP?�he���_ߦ���Ь���dc-�+���Ǫ5g��i96�̧/8[��EJ��fkR�� 3�_Cz����(i�������0��5�z`nqY�j�z���3D����?w�b|1<S��\���aR�(_W�'�zuwf͙�s��p}�0%q`ZӦ�b�R�шm�Xlp?��*��t,��0�w]�p4��.��
�5<����c���a)'f��MP�}i+�dO��Z|cB��£���n�4m�\���[8�ꈠ���]�R��/�@�~��~Ĭ �ƙ�9�N��^��ʙ2�~T�f�>f�S��Jۮ���ә��,�|b��N��i�{���Ż6��v�D��4��^�2�����#%ʚs�R�����uȲ�������Wu֮�'�,�R9�bf�/�Q��G�jN��F(�,7ꐽ{���>��]vi�S���t����1�6>���:�;9��|Jc���=���p�҃6��K���&��������a�[��:��
��{;���j��'0�N_vY;az��P���:b�|���97����9?�}�������E�|%5�2�Y*�2��Z�o�cxP�7>���So�:��tR���l�SVc٬`����{+EIH˛�u��s��_��=�P��� �,��{�%�Q���pn�O�}�X�	��c�����>�_�z����ۿ����!�w� ���b5~�ˁQ%�z)_,L̎[<��q�FEZ�_���v\�Yp]|�����[�b��z�'Y�.eq�;�8��f���j�1q�1"=��VY���������W�w�>iP��"���y6��S�^e�z��~�-qe��->�$���e=_�ޝ�34�q(i)h0���������k�g�{d{������t�U���sp?x����X:�^ˋyOS��))
�gʚe�L�!
�YRWR�n�t����i���[�bf�ys��c�O/�d:E�i~m�&�>V9��~7M������c�\�V��X��=���7�W>��B��}�J����H;��Jr�L'��}/�^]���X#yf���_�s��ز,K���Z����6��F���Z�5I��L$�@ ��HbZ <��A��%$��.	���0-��Y���n(��Ո
<Ym���ʩ�0i�����[�n�z�) �[r�WA}H%�-T >����Q�P�͕��Wu*t��;
�U{6�6v8�%-/1
�j��I?岌hZ��G�7���K��y:�H�fY��פ<⁪�����M�v9N���k��Q�誼	��Y��j���w�?���4y��Q1��vQ�v��9U�m@���9���U���_Q.�I�Q�i�ĳZ!z�dڸ��w����Y��N41��`����.���4���Jl��H���\���T�.�8�i���z0bf����)��SV<�.m߅S��ҥB;���[ʐ���h��ww��E�v*������C��'\�cD��<��Qi�(��&D=�,i3f�:U������qf���#��Y����=����(8U��&)XY�!�G��}��,�-Z�G��=�b�H��j���ZW���	~��?�7H�g���y�����>�H훖���4���]��߸7_��a�c���jto�Ц� ���ӣ�����wh=7��8�^�~��V�;'�i[��
�O�����y�;^ܢ`�1����z�~ �б~�,��M5H����Oy�6U+f���6S��-}W�{Y&D���}
�c-�pط�ap���|�p����z��Op��<�?U_|>8:��(���b,n��B|�>����,���J�7�L<~@��Jk�;;/�\+�_�g��]
j����#�R:GF3� (9�RȻ����q�OxM��X	V�&��O��,L��f�)����}p:~��L���P�N�H�Ϗƶ`X0?򶣛�%�w�w���r]~�ƝAul�!u��(���]����ӓS�	��-o�"��q��^�'1�G�cW@X��T�������-�hj�������<ĳ��H.�(���L"�)�M2z��E ӫ�އ��t�i���1�=�P�	�+qĤx���2İ���C�(�0q�X�k��� �]���No����-v�Y)�+��'�x����?����U�)$:ym�`<i�5�y0�sĢaR[�p�2�i|n�[�W;Ҷ��U��)#�(��S�rOK�/5`2P;�ơ߇ ��)4z��!P!#��k�[HN����:=�p�h5S�6Dh��o��w���a��Z�=1��;�Y���j$�����L��g��,l��}uA�2N�goU��	�[Z�^�$��#�pkQ<�?����zWR��tg�rI��NS���b��iA��08}+�
�.ƈ{qI�����iz�{�/A����;���W �`]wN��ZXRkm'g�Fk$s��\Ь]i?9!� K�Ҁ��۪;�`]���tm}ă���!N��[T�Qa�x�!\�p7���c����x q�OI��y[w�x��޽|�4B���!6����m6[v���q��~��&�}6ܰ��ZO����x� _~r4�p״��:�Pd�0��7���O�ߍ�/8�Ҿ�?z��~��||��x��֫u��W�k��>���;C϶#y�S�h(���m�����7CK:��lC�O�f�q%p��t�qD��D�����@i�T-��;xG�}$�L7�B�m/톫r!ɻ:��Um��U�����������^�jY��H}^��L���a1�,����W��ҭ�*��%�$�zho۫�3��l��^���~���3�5�t�wD ��#h��p��*Ȫ*�+��J���'BG=\}���K}�Q�Tȭ���ʶ�E��� QB�ߵw�W���4m�XQ���7#`3��#x��j�Y'�:�(6�i�T/�T��»���ެu�Z�-L2�7EG����]�ftZQK n�r*���<m�ā�mG�h4ݽ�=V3�!P�Ãm�j�b��J��c���%��n3L�i�k��=�4^w����<�b�`A[rҐ�m �e��: ��>LT��<��֐|���V��6p��H\�K����M� q��%���MƂ�-o�3�8�_��KA+-;��xŢ�(�'pgjK���̊_�$o�W��`t�f"�/�� �}4�Bj<�Lu��{�9������ ��T�IԖAm��(Җ��e�e`��@�t�x�_��pu��"��n.R��;qH���p��V��0�5�Ԧ�"(��S��^�G;C[�8�K�ȟ�B���\��L\�'�P��t�^�SJH0a�8�D�XD`
j��vZܸ����-Q���3�9�\�G���bĪVk+<q���S�>�����Zc�4�s:�JJ �ۗB�4�蘒.��zP�P��0��@��OAFtN-$����C�ދ�.�,a�����U�,�Y^a���S�W���,��4?��n��2H�'�:K��= "�m�K�D�T�cZzV�z2SPʉ�kxUj1�CЂ��6^�;|��|�~�x�^X��M`��j1�_���.�c �f_�2xI�{xgh&mR�#�p��?<�/��K��5j;�/���y��z��o����������<>����q�?���1����}˻�=��&P�?1)M��_L�'Oۦ��W����@��9F2k�>@ [a{�E�0W�g���A����!��Je�~+o���[�AY�V<��D­�L7�&�����%�IC�.Ap�M�G�Qn9 �rxf��k�V%$}��4F������J�i�K�����	����3�K~�@����`��$B&�����(1s�!(j�%b4�>9#�
4�7��4DzOD}�(���p�ڒȵE���9�	9�_�����'{�mM�V�Y��ӵ�D�őTɏw�U��%��h�1�!]ᨑ�)����)'m�����h�T��G8)T�0:ͧpV�]˛o�e�1;��2$b�����D`$�$|�Q��(���k���8�^,(h�A5}5�L�e��F�?I�@'���NC��Њ(vJ�iς��pA���H�|��o��Ӯ���l1�'�<n`�.�(m��Ee�I�;���t,�r�f�I�j�	OyI�`LR�Trj���t�:�*#P�!eJ� .�n�ؾ�/"��0a����T)ੱ�]��w�1i!��"�9}n�S�R[�p���Y��2O!|��Q0���&핔���ţ9�Kю |�|���6$x7�bG�R�d/̄#v%��U�@�<��t�� .<����tN�����]$p��&m51��M^jV���0i*#uS��A`㚝,�&��.��R��� �j
��4�9��=W�Cl"ϐ��4�i*DZU�G(,g���Yx�,�������g�%�%��Q�����*�8�F�]`?zvԝ�E�;6�JM��)��+���@35��$�JJ%�� L� �<�^��>�"F�:n]d�(<�7���+	S�� 2%}�#�Q�Уi/2u�L�Ρ��}Rh/aA��&�F�t�b���"Fxu���k�O��O{׮-��N���w��-���[�hN{>��y�{㶣�k������KqS��G�9yTv�S�8)Z�.u���ө��T�c�̠���:�ʛ�oi)�D}�d�eԷm�>�*v���̆���	�H����I�� uO��Q���^�ǁ{x��r�2�#?<��w���}��b��|�hX�鏞sc��/��S�X4���/F�kl�ӎ�s�n�8��iq�]�Z��W\ۇ�y���0�1f�?���N�)c58	H��VlI���WD"��\e&���A�v���¼�ϓN�2�z�>Q(�����&�X6�Nƚ���w$���J��6|%0��S�S�DL�Q��RP�"�C��,F�j����%�w?,�K`>�N"s�b0(#�L�.�Q�� m��ȝ�!x��<+����I_B��������� �ܬ��k�O!��NHZƵn(EV�.2���# @�P���W5F�-Qd�1}��e�Y��D<�c�r�>�QN�$b˒��Hg���ip"��x�F�R��`����.���Մ� ��PW�<�L�O��`(��f|�Ь -��PB�i*X�X��`Ж�}"������a~tF�z��aEK��g�h&t��#K R���:TX�'��~����%�H[Љ��4��CkӔ�>��[5r�T�)-��m+��F�������Aja��NK�:H���Nhm�+5��^�$���A�Ep�U��j2m�]]����2j�4x���~���(��S0�����b� 6@u��j��� �&�{��ZXB�/��y��i_��[�25?�:?�ތro��"�ؚ�W�{�e���%j�l�Һ�G�Sh*ܸ�G�d�6b�l�p����d\���<��:��X�v�p��+6fG���Fkoo���Y�C���2��_`��^�.�I�j]����;?m�0qG�tv�8�Mr�^� W�h]?�L=n|G�!S��������Гu1da�ۉ]���kzү��h#��|_M�u��k��\o�j�����=fmG��=��R�`V��1�XB?�I+%���C�{�3��FZ�(]����6h�׽�?�� �G{ni�����8���=�k{׾�[��k�ϋ{?�ky޽����ᥝBW�J1��EY��S!X;KO릝3�5b҅�V�%�;t��h�հgp�`�A}v^Aӥ�GW�ߢ�ϑ�:<c� }�(Wco;;:8�6ڸ�9zʯY�50>=�wj7/�������'��/�6���}���"\۶R�|�`��}x�������oh��'�4>�iɷ�]!���p$~W�h�� Ȉ�(!�@n^	�oK�eX�h		��O"sӰ� _�N��xzwoD$������+��F���YH�6lG`<�G���Z)s���J��b�0S����[�)i81����ŝ�!{jN^)���hi|`)H�����$N��~$C,:�����;�����:M�r��˴��#��b�K���Y5�����v�����C���E	^#|ZxUd�򙪲�5i �`�G�Y�rĨ������r�������	3��4yk0?�+�MP���4 �TH����C�x.�Q�ʅ_��%#�k�oݹ�֕��$(x�u�R��G�u�E2 5%�V6��'h0u ���K�Ϋ��_�/�D[�y\̺r�z*�j	`֏4%.�W�H��C��_�>b#S��\'x��T�%�(�-e��a���@ٴ[��كP��6K8I_���)΄�b?bJ�\���'�QȨ]q�Qq:hZ�xI^��I^��]���	��k5�-;Z'���b7O���*�����C��OI�B�|��Y��b�e������#�w������O]?�6tG�@�zsA
RxP�e� xd�2X�},����b�]XPQ���i+v`ְ�j�VY�JcV"Yl=.bT�� �0�՟���	A:RHDлD0r��>��ɦ���8�$��=�Y�q�
��@��n���=͓Ǜ��Lu��SS�Ȇ�{��yv'���
�_��tH�=q�o:�SN�L�d�1�H|�I�,��Ua,`����{o��)��7L*�{����^���ЛG�Pӭw���O˫?�[<Ϝ���0n{�}����<�;.إ��y�;�-���(-���k�}N�N�&+j��!�I:""$?y�� }�.p�Qu��eRM�V����߁8�)�f���&�+˸N�O-��T;�P��fgN�;��x�ٝ�!�uU5sC�e�����L��<^m;�a�/���;�[�C)^=�ڞ*���m��R���gx0��ωc���蛔đ<т�C������rW
#�����}_�������#�� P��a��R�f��#�&��\�2�B�8l (���FQڍW�������� ���0��-��)�!"7���(�ؙF˅�����/�'%>�YnN�v S���k��!|�p���w0)g:b�T�\d�
`Tq��~��hԀ�2��c2J�;~�]äj�Bģ���+���$8j�!�r��آ��i��Id�\����=�ЈMcx=�
��D��O6�����D���3�N"���J��ޫ0{
�18���N���o���l*6�ī{���{_Ի�t͜r��S_�4#�GnaFvtN����t�vv�Q��Y~>��dX60�)�Et��4�<�F�qibGi���B�:u~�!wr�1B�t�j�\�X���%|���tS�ӎ�L�~�}q�]�J+v�����<���M�u�ܭ��.@�� \ �v"��j9r�c^V�>~���k�*�2=F��J�_��<e���^���������N�AJ�{ZaW��C`e��~r��`����@_C�����NG��K��:�C1I	:���O��<��=<�v��p��]����"B�
Ya�G�ݫo���k���C�>�k�����r�1��[�0h�)��$��؆�ߜ"�th�V�h�o>ĸy��-�S�j
Ĭ�T���@[��o}�����Y��S
^n�B�8� q�L�x��4�@�i�	ڥ&'�	���jn�-��#�
@v���wg�}��E�4�6f��O����W��yӛ����J0]�x*8ȯ/���z{����!�-N���);k�'3�ʮ,S�6Z�G�l��=�$pyJs������ЄAՙ�@���|k��G��L@�cXu�v� �?,������jX��Ñ@~�w�Q\�i�V�7�ܾii��8��7~�oW� �w�	���4�h�D�|~V��4��O���A��)>$�k�#��~��U���
�¿��e��ٳ����:��hw��Ϭ;���?�U�1��cYI��W���M��V�0�]� [�ako�̓�	�E~!���@૬�p)ķ�����_�1�����:��*\�L���<��� :v`<E�0��vꥁA�Ҵ�����p<U�0m+�F���_
�����
7N�����o:�(��?���s�4},�U2����w���zc��A����,�!����  @ IDAT(�p>[ǩgt��H�}�\&[~L\:΢l�̀ ��m(�8�=Ezکh��j�hS��Q���S�νG&�4�"SU�a|��e�4�f.Zt�C�\��oO��Q��@s��s����@�Ax
@�����ԦH������X\�Ku��Hz�����UWN��Ƀ>i�p�|�MA����H�U��5r�*��EV�d���h��a*:���t�J�E��9�y1?���%]�#W��|�����4���B�ځ����:_渜DX�Q���'$�Вn.�^����E�0/�xR���$�Y?W0����a^i�L85�m�Hj��'P#~钗08|o��i՘��ޢ�i�I�eN�D(؁�T�����,��1AZq�	>�:]��vc���vϞ>D �dˮu�U:_�е���%p@㧸�8�X���F�(H� ����Yᇮ���7#i@�������;��@�77���wO=����0q�2`5bG�J��9d�w��}ܙE�a�n^`�:"]��}	��Y����h�Cw�Gx�-<9G_'n+��[��A��q����ҙ�=|�=A�z���V2����Zc����e�"V�C�k}��ڽ��~�Սn�l MYo
�qG5��0���)<A�#�e�-.y�������{�N���������.#0j� i��&�&\��udN]�#^p"m��q��Q����E�hI��I���>���iZ�I��GIwދ/�ضY���_�G�{{��#�q6᧽�4.Y�Ż��3�|ǿ�-�m�|ǿ��o.����t����=l=�|	��.��[۸����<
�"�ڤ�]�VJ�.��o�/�����5Խ�ecs�լ�h�ϻ���Uڜ;*��w�!�j;|r�p�[~���9��hpO�k��8F�����Auq�4w�s�"�*S��ާD��~ÒQ�>$ן�1�O��I��W�B��^�тS��#R�w��ixդ^�!}��<ڽ������^��:�<� �L6�s�P��2��}�G5�B����г$��.	�p��t
�ѻ���f�{��v
����Eo�:d�A��L�����<Fp��]�=Y�ZB R��a!�� v���VGvt2NA�Aq�y���E�INǘggv�JA�ߓi��tJF)\�EʙS����c4�gG'�D�%��Fӷ���S���x/�.]�x�+s)2Y��}J'�j8m6t����'8�c��g����.����`z1�d+j�2�Ε�n�k�˚�>C���1em��⽰)lF S�`4醛��4D9�Ӱd������!)?����� 2�+0�`{%5��D�idq]�f�z�t���"��s9���Q����e�$��H�Hi��v��t���K��w��<��꒩)]�h��9A��nb�����(
_h�t]���^S�E�5�	e
y�0a`H�O�����1d���0��4��X�����W���{�4�W.j<!�z �v��CN��D�2�ߡ���W? �Mi��
<�p�%2�5��G���G��Q��S���N#b�=���C�#�i�C^��݃�|�!�m ,|@�c��*ӟq �Gxm�P�a����`�ڥC:c����[���x��N}j-������ѽx����d�ԍ8�nl�<�v�8+9�{Ys |m!���3���U��46�뀇 |���S��M�:�	p�r��T�.�d�-E;�44K*E����`���l����n9+����Cxw`H�F�T�R{��4�*�=��]����<��ڻ�P�-�¸F�j� �p�����+h�	�p��rZ�����K��Gkk^�4`�]�QT�>�w��4}���i_�X��oy��]�����ӾO{�����ڗ�ų�œ�g�A�iG�Vp]��ڠɴ۳r���W��@�n�G�ĕOZ�6X2O�3��>��T�׼������K�[�6��� m��>#/���L��WpQ��>����i�+@r�}s�"c�ay�����SH>��p�u���`�
a����*q�wۉ3<�C]������#��8I����|�������Xw𴸾�4�(vk "IB�ډ�=��Ř6	H���'�}M���/�������-C�>I��MO�\�@���Q+�>�ߙ���.�8��8��
�<����>�9�ma~� �m�$Ҿ�O����<�ga�>�a�@�9f���Ѹ��Su�N?�h��8��ʬ	zW[9�TS� �7e�&���}4W�:�c0���S�ɹ��1ƽ@ ������T3�\��h\�F�=�50+��yΐ�S
�N�
��=�d�i�+���ػS�%oma�sZF��B	�P�Οp�U	вz��{�Z׿T�?���m"4F��|��&㗔���J
u$ߒ$�F@�g3�]")��S/�K��� |.�itjg^�"s(�t�e|�Q*=j}���W9��H�W���f<�Uvr�P�VG���q+�E�z���)��M�czj��<�k���B#e��u��|5_�:DTK���yZ��E�[<dS[���Gx4~��	�� t@4�
�sL9,�.t��D�+ݓGh��?���{����o�W�ܼ㜑�5H@T$M�u���ٍ��2��Ԃ�7���N�v������4���Q�
ӏ+0��\�-g�9������w�L�.�k�S/j�d��@3�W;�ͬ��g;;�2)�E�MM� �m�y4��׺��9@/�<�=���p�_|N��mb���YQ�C�"U`������h�� 0$�9GRAK|��i�ֹ����x�M�:\�w��ZgzT!����*N��!�E���d��l5n��\(7K�M ���b�r.����6=�iH�kk�c���\�
ϣ^��{ʧ �^��>8��4e~�hu��zI��q���^����*-����qZX���}������<�ߵo���^�Ñ��XyLg�(\IM���<y&� 3m�n-x�����֓Wx<���>^��q��E��
຃�6e���y��apYmB�~�e�쓨p�����B�-���!���Π�t�1��e�&1��_�Mƾ
���۲Q�*���O�O�ѯ!����X*�IhT���eL�c�ʼ�}�����vm;��)��,]�$�RT�O���7Ja�U7u���3Ҁ���5���F2�E�ֿ������h�g�J�X�WIS���G��
�,+�.!�C�r�+�d̖����=H�wy�O�h���E���N7A�������ná�����k{w���n�)�i���Kw*t��XAM��i�����)���imz'0�wl�����?��;F�+�h���r�%:8����/��o.���i��{�c�ߩ���M����v���QKӎ�k3��ӿw����o�o/�a��F�%\1eC!<���V(�z�NJ:�յ�����M���/�U:���O2ճ�{�����~|���A�x~�qN1Im�b$�A~�X��ď�[]W�I�f�r���`q�/L��H��I[:�4�4�-�B}���Qi	�P'�ϰg��7�4��&+�<L����M�ΈzP��kh��� �]�����փ��|���$����I{;�y�]���~DxG��~ړ�4nU�/��q�#��+�>e��� f�U~��F)�W!��?�#F�t���Bɴ����#�>Z��g���WO�'��*NB�:*δ�X�-Y˔{�1�H��Y����E���xJ�8_��Շ�lX���*�T/��\�C��>M;y�L�fTJ����j��Xpd���LC����fc�h+��{�G��\C�ۂֳ�A�e*D�}���Z[\z��(�]�B�E��ɍ���`�9�H�Y|Z��|�^��[C�u�F�b���i�7W�]2�:@h��&G_K�;7ԷS>�O�Պ�1uׅ؄A�Ҷ��&i����������cD�Q��F��Y(t5�j����� }:��,���<I:�AhH����@7�e��G♎m�����/^TmA1i�n��k�_��8�3W�
/��q"V����h���w-�>�w\�1}�ܾ��x-���hq>�����{5�L�s5N�.8l��{�c<-q�~�ױ���2�˴��ȩA��]�i�
��j%�g�M.�8�o�dP��g�/� �B��T���+�A���xƒ��[�������!�^gh��=I����(!pM1Uy���>+��0z~�Uƴ�k�8��d���AL����������<��OBePI@��a2��U2
wlq �;pd�2�r%�u��a2��#~�7�����1S��U��O�ly�?���$rM�]���.)�x�,=l�k�G��@��R�������`a!]2���ǧ�a>��F]^�I�̯�e�����!����MaZ���do��L� =vL*�W�s�h��?f~�݇�؏�d�Si����(� �t�I��S��=����=~�}���|��p�[�P�Lx��_���NB{�u�
gk�}N��3�\�iKl��i(�	�oS�t(t_�|�}��_o9g��(~��Uw���ea䑥�thv�(8�c�\�cnm����۾[$9��Vd�^ P~� ����<#^7O����޾Q@=�NP%3\�S�)*T�Hģ���^���
*4���{��E�����ع��6�Ə�������|苂����^��@�4�25��	K��o��򦾀D��ɢ�%I��b�;�PzPq��mP�LĖ��V>��4M��Pb8~���������e;��7��f"�EB���V�����U���[�Ɏz�7U։F��T�b�!i��>\_���)��G���WU6̖^�!a
�|M6�g�U�>�Ʉʦ������+�L����I4ZGh�#��"�T@Y�B�A���g؎y�1�%$-����	�wd�C?G���E��aS�������;@��eZGH����^As����x	͑� V� �8��J�b��W��b}H��M|�th��-Ӧh�s
�U�g��m�S�|�A*8c���LM� D���4�XO��~���o~�M��œ�ᴢ�-05�P�s��S�0b;`�	��`���I-��$+�yH�W��֓WVLڕe��1�D��ՎJb��y�	���֥�����ٟ��׼�{An�8�G��;�z����7�ǰG8�}�~�j�vn)�>{��޷����ϲ�F��b}�ײN\�zl�3(��"N�>͖�y
�3!1c��Lg�I_�P댏���E�޼�\���3K4��LK�|�X�H2@wK���=�B7|F��@O�u m3E�a��h��Q�����i���Y!Y���%U�/����S�={���{mg�WQ8��B;�����3<�A�������i��T�mW!͕�W�H6Wd���7Z�1��i�`�<�-����Q�����"�-���<���L�F�t�Q&�i!#�Qd��8��nl������-���J1�פ=d�h}A}�����wF��_��}> �t8�yvö����d��̛����08���9%V��I����`��k��:�!��ZY�����B��sqt�5O�@eZ��L	l��B�C;����l!�E+�[�Ht���0'�.�w��+RV9;��Ԯc�iB����3���F���`L�4y���a!���$�~�ʱC��sd������`�N瘷5?vj��Z	�:���SMŊ��*�ZA^q���V�[��V������t�\�ܭ?�CM�S���!\Mo��.3	 ����(0�0%��+'ߩ����g���D��M�-�bD�J ��S' *��O� 5����	�����YZx@'|ֽ~�c�F���z�:BH��^��h�$n����]�}�F����ى6D��m:��������ѓG�/�z����L���ϻ��v��c��ZN4;f"���p8Z>S��Uf��UW���4��:Z.��0��>d�:��۹;�g�:�$v�Y�p��ֱ��>��?�¤#t�Z���Y�'���G�u�I>F[��I���o�����ʾ���gؠة��ӭ���/��M���.k{k�A�v4�Ǵ5hg� ���ũ:�8�0ykB���I�$lfps�|����x����<y=~��z��n3������`�"��*L�X��bo��բL��Y�W5~���_���ݷ���ՙ.�g����qz�Ц w.O4]@�?� ��(P���=��x��* �V��+���m��^���Ԃg�W���C���:y��Ix��u��m��l�~?}���>���.|�<�H���w���ƿm�Ҍ�ѧaX[������ȥ��a<�g��l
G܋�m�ҳ��ҕ3�!;���0��ʤr�6�mQ@ҙ���������)?��?�雞}J4�����}�hr̞�^�,i�����RW%�@&�`�j������0�3���/�Ou�c\`��-��{w�w�q��J(�Fi��r7.	HG"�ғu.���r$O)��eߦ6W��d�{&�>S���N�;u�(�"���_���K���+	�hr��MA��@@n�X
�>���FV*T2��ދ�g�a��L�h�Vp	�̎������uNU)R�b7N��Z�5�a� 4ާ0'�q9���
�l�lr��X��.Y����B@���e�j}n!���e�p�4�B�etՏ[ph?4��n(�ڭMtn7�~��9�wԨ�E���4 �O�U{荺Q�V�+Û�#XfŒ��4�:���`�o�:o(�@5W¬�xs��%�`d�A��f�"�I�)^2�iGjG�=�4�Х��+���͓^l�1�}��DnȺ�	jS� ���Z7��xo�?�r���{��)�އhM�?�3�����b�e��c!p�J?L���>�0�i�`y�`��<��]���z׉<.I��4�Lݤ��;#�VR��g���}K���PTiOa'7���C���>^�s?��N�iy��*\C?2,?MgF���
 ���I��\�wO`r*��׏ �LB�Ti�w���/w�~�{��AV$����C����#��(�]�D�`�M.#YW9�w�S$2m}b��Sj��1���8�uJ�i�kh�C�ϡ�#4c����V�4�i�g�z�V����A��ח{�f��^hp%���G�O�i<�JM�Lg�����د�0MrB�1� 6����5E� b���6^�8������o����h�h�(�i?'���4����u>��Y��������l3^�%j�h{����.ܠp�%���~<d?�Y��R�T�p/M�>B ���ݗ/��씡�a5�?�>�#�m�M���u^Ol�IGw!�eY�����R�G�c���$l�J��#V"�N�{��k�u(����P�
&BE��~�M=��d:�%Hxڎ1��?�+l�<�}V"y}������q�j�}�oR�?�O��8�����_[�[����۵��8��SQ�'��+��;<��ie�R&��U�[W?O����3ؗFv�p#�tlkR|�E�1��S�,����w���������)�1h��b��R�M��!oq��TL^�,�ob�Sh�Z�k4a�EX�������h4b�x�
��\�I^�=�Q��Ϫ�g�Z���jҦ���Q�U��#�vL����$���*i4U*!L�?��>-pz��n�äE:�aa�(
PD�
 1L	2��a&����� P�n[�e��D�ţ ���0O���J������>�*�����G�2�"'���ϭzD��%S�?��^�y�p6
_���2�� �hA��|ʰ�	���4}�#ˌr�t���pe{�p�0���۽Er���K�+!���^�T�N�S��hVM�g`�j�T�{ 
��Tbm5�h���2�Q�Y����d�zOX��5�'���2Ƽ�Ď��a�� ���H]+ R<5d�,I�e��,�v ��16��#
��g={���o�����l�)D:�`yP��A��w�ק�J:В����������ۿ<d�؃+�h���v�(���2*pf��ܥ\=A!p��f�@�4��B�>A�26�2+"�z����#:��1�X?����Pe�e�AXB��_2��,uh[է��M�����^�gW�g/�w�����w�y�}�l�#Z4%���K����3B�&? ,�- 4���B��*�#�H�M���C%��ܶ��bt���E�ii�_٧�k_B߿����?�{�+���E�E�NZ��O�0VW���q S��+]w_0��#\IƩ>0
�jg&�t�X6В�P!����s��=I�)�v�;ݟ��}�������#�թK��X7ؿ�ta�wj���h0����Nش7�\G{��o�
�bϩ�C��L�\�bx��>L����. ��V���vkj�Ԫ���6%F(8�b�O��؄��K�֗V��m��k���6�ѸP�0�l2(�/�����~I�sHZ�</+���6Z�f�Kq4�'Q��m���]�%N=J�?/8.��wI�>��G��ƶ��5���%�MK�:~����7��\����k���E�}�Sރ.1��9��y�H7�����L�����P��Ȕ~�8�.������v���/ͿiCȄ�B����C�.���'*x%�%��\4[6 [�xu:� -���>�DaN����m�iu1�"�]"��ԡx��ȳx}
�W�l;%'�:l{�<ч�s]آrC�����2EVIßm�t��Qr M���Ҕ%�~�Pvy��(�f�`f�P��'6~�-�h�f�a!rS�yh^}O-$�U�URd�F��̣�UPq���aW
@Ņظz�/X�.��&��F��P���Sx �0�e�c�WpI��r��K/��0C���	�����Bt�;�MC�S���}���#jp6`sQ0F��T�NI���sSH�t�(�ה�l�C�|�����dF�<e�Nc��7�:@=^����P~�܍�e���P��l*"�n�(�Q0R+e�)m�D�04�9C�u������2��!ґS^�e��SKG��
��
�F��AYwU\�;OR���U]Y3uX��!~yo�&^��
��ӯ�W�9*����X�֫��Ѹ	���!�?e�F=Is�'5��Fe�7z�o��@���q�y��GU�1;�>�Yg�E!X2?g��BB��s��Վ+`Ҡ�2ū{ w�����U������������sZVmȪJ(1��dQ���2���{����ў��tvz�cՉL�!�O/ah�*G[C��j�kh�is�v��-�ƻxf�-�����,�[� ������M�������C: ���6; �}X��-��w�A[����Lj_Bc��i��]Bu��?�lj��� #tp(���?D�V��W/��S��͸�\�m{���{eG��m�\AU�v��k��(;;���Q8b�ir�ۺ���t)|dO�h�b%�=�u� L�@�mo�S����d`AJ���b��5��c�=� �8@�]e�St#o�k��,'l 4�`P���޿������<���6J�!tQE���v���!��0�E���l�����g���ԼyYU�&)����!U�� X
���������%8����Q0ԣ��]�����+����w>���k�z�v������u<~�3���}{�7���G�]���%oWp��	.QKߓ���p9а� >�uJ�� %}�����DA�x��<u�3b���b˕c�A��h+j��b�3��GO0�������%t
w`�H]x5�L�0���2)XpO>i�ɯ�gG����FL��<VN)�Ps3�o�#i��-U^��4�$�� A�<��i.1y ��:�̅x_ԅӿZ�	HH=1�9�O�? :E�x6�^�q#N�ƺ\:�%���� =�<;�R�Y0Ӱ�&s[6�ZW5��R�R:�a{����hP��X��I?�|_�#Sx<)�Y(��Jɖ�����x慎Q����p��x�a�{��i:��	�lr���ʳ�:�� /�"�S����d%
���a�X�1�=/JkC��ѩv7h��~)|�0U�H��t�G&{�t��M�i(�uj �)���ьf�D��w:D�Z*�e�+��Hlj�ʷS��t%p��e�360ƼD��2C�	!DFY-�1��B��::�Z]9�"�3f���u�:��p����_"\'1�  ��f�z.���xMyč��� �h�"��}\mP4=W��ʆm�f��N����}�a{7B��_���n�� �J����rG{��nF�m�)�Q��-ׯ���*��lN�h��r�|���M�VInl����k�b�C]e�C4jW�h�Z�#�Z�Yڥ��tW0`�@iV[�I�*�{BK.O�m��5�x�'�g� %芟^#�[
^�H�-���z%0��Y��]|c�b����y�7��bK�W:H^2d��Q���;�����?�۟��%��j�vd�*tN����OMP����Z0�jɧu�*?��|�!��;>��"��&T�Kڲ��iE��r�)E@R���A���C���fe�ww��y�fj	�e�����d�zŗ��u�����uuu��y�[���fԖNڎ@�Y��_�6,�	����UR�4�S�Nכoh쐡���%��#/���!���U'�+���u_�qَ�p�����V[D`#������c�����7�k;o����]۷�����[X�;~my�����n<������A��C��$H!������L�pM���R>$�D�V8���#��	���s�f���ndt_�Y�g�����{��rH��a�][�� o$��y���L3н�{�]���?3�aG��o��Ǹ�q���m�UR V4�C�mk3��f@���c�A��HH�ȩ*�vfN��X�f��;h��l��ӎ��;:��|���G�E��fF� _�C��$p�&����V�q��c�̓Y#42�M�J���$#�+5�����#i��*;c�P��[�Ќ +Sj��vtbL����8�`f\���I�Z�/~DBK;�"�Q��r�t�-L
�ڦ),�"�M��>d��W?~�{����seyb_5��Y�	�k��g�j!�p��
_��)E��k���)S�p�BB��@���_�&A��ܩGWEEc�+�q	c?î�8�Z��:}��(��V3�t;�0�ĪV���x�q�҆b'�"�$0�F��2F�ȩY�Y�*�Eq���L��T҇�@W?����QDn}�/)w($ϩg�'O㤮D������M���S})��T�r�P�
U�2i�����!v0
W��Gh�= �鴜�+�E3�������"�iDm����C2+���d���5hwq�4��32 �f��1�[|h�M�fu�N>I'��
���Y�u9d��� ��,N��&���J�v�QXi�p.
N2M�-�5qU��h8L�d4f���](e���y��U�c+�i�l�%��0�q�#�jP��ԯ.n(�Z*2	S�2��\�'���yv�i�ĕ���x��=TG��ʯ�L�m�6��K�YɗN� ܒ�²�X�2��'��Ew�(��!�==w�Dr����䅶��c�>c�4݀�lգ�HW�k��m���BL��[���&$�Oӄ��GlKJ����W;W���P��y�G�FC��+�oҷ5Y�"Ϸ)@B3^�,�6}f�4t�+���t�b�b=f�"5��W�8@b	a�3�.R1�}�1�g���#!�������w
��o���0�+��7M��4��ޏ�m��}������ߴx&���������v�q�g�N�<,ֻ}�L���)�J+�\�ޟ��5l��9�Ѐ�z_����Tn� 5��du�%��:A�M[r0$�Ќeͬ��<u�L[q��mLT���>�&x��3�����&��qk6�GU�R���� D�H��* O��A�J� -��d�HO�d�{#�7q+>���m���u��(�L��+��6��7�\�I��`�����L�h��
"�<��l^�CbTF��S2���"��dRf�~����qG�>@F���rm�@�c��Źh�����;yG�X��~VH;Ʊf��T;�*x��x��o�G=O�j��FԮ] 0��*}#\�>lv��ǿv}��;b÷	:��i���g�e�nu��&L�U��@H؈.A�!�U#C|%����+�8��8����Q>��[�Yx�&�dG$0�I:�+6=�a����#m;�h(4�w����27�g=j�k��C��cT�f�LI��*�R�i'�((���݆d������\��c�M�]�d�����)�ʤ����[�
�%DB,�d<^���?p2jd��~skb�q��;pFB���C_���A֑�6@j�r������y(��1T|��f�::����V}9�`�}�v���<�	S�j%i�aG?��-�)��[�Z��y	�
�j�\�p���E���7؞a�������c��4$�����W�
��Pj�d�b$���җ�"$+x��0it�ЕQ˾g�95����}�V�l��άsӡ�I//��4�>�E�˗�P��hWJ��H���Vv����1���b�(��+��tVZ��2_Tg������t'��ԥ#,��@&�
r�d(W��eF��)tK����Eީ�Y����*(Fˉ��>F�
42mT��<��2y�Y�~��+Ʈ�R�lT5}������[��.��փ��k�4���C�t540�(,?�Y+�v9�4�">�����r��/��DT��]$;[`�y��eԵ���)�-��;;��%��N;��4^�/3(k-����ݫWYW���3w�Y�
�:�7��N&5��Ǜ�ml-?�hGZ��:t�K�E*?=F<������#oτ�X9�9�]�3?-���-���	.-O�3���a
9��<��iߴ4�_���,f�U�/ @뿃�Qq?%t�^
�
(����K�����h�ԓ�`���wW�~���ݗL�/1x��Kk�����m�����^y���?v����O/ :�ͯE_<ٽz�W4����U��)/w`��?G_<� V�l� ~l[���PT�`�v�-����[�RA�4��'ЦZ?��+y&�3��U[C��l�3?ZRH�M���
��xl�g��ݍNڼ�AƔog ��$�˯��Ѐ��|q�mF�����1�� >v3b���pec�`0nnD�LEfSs�6%X� 8Ҡ�$(x)�iSLԎC$4�@,�v*.��w�}�͊���'~���:�fF�
����y�{��Z���9�^[����M��چ(�im� �i�0՜h'N��$s�Z�$E����c:��g�U���V;/=ٟ2�D?M�2�YT�׮B$]�kJ�$��e����zҎ��!{�����,��N�|3�j�ڑ"�����c�%LOphǯ�	�ө
#e�!�9���YL;�<RV��~�J��8y�����S`�s�B��i<B�($�]�UXK�:g��0�vj��K�:�o�J��IJ|�]�3��*�Ԉ�A�,�����-͆�-��$�"�j��R�a�v
�;�<�<G��K�`�x�,U��-� %�h��3p��$�\[�2��.�|�%�xo%�N� $��+���Z@=������s�Gx07ywU��}7]�&���u2.aXB�����/��FB�w��:�f���]�.Nq�{];B���~i@T�I0��)��u>�AK"La�ѥS(%n�����Qgi�i+ЦXu���p�ʎp�*��A���U���G7'�N�k�z��
6N�h�B���IY��e4��ؚG�ҕ��9�):�hͩ��U:���J� /�sL1��L�it<��`�_8��]�gA����U@"�f�v�;���p ���A��Zn�X�!I �>��4��b��
����-�%q�����	+|]�Wq@����
xv���]���{�іI�I�*�n��X�=�DbH��5m�Nཟ�^�g[\�MPj���o�����������)�]�8�������QG�.��Q�u�"�Z��d��vƷM�(�Zz%�YzЌ%Z0f�Tt��s����2�'��:�U���g��g�Md�=O_~�4+�q���g�c�G*p!�Gڞ}�<�ٺ_�E�+�q&��M����۷�����3��!+�5�e�	Y�풅8���?���?�^S����7r,j'�@��rq��E��N~��:�M���ƶ���o��S����S"Y!���N)��2��2I� Ty"�"�Жea(��������_�7�!6�E��@�r�6�N@��#�E*R5��~� O�u%]��301�@�"�,��!�GKg�v��%�H�d�_��Ʋo�mu����!��}��n
�Z\j�n&�i@��!�,~�40V���h�a딬�=��:�9B;�JP3��*��լ1sF���r���U:H��0R��/�܎��)�]G�t�j��őo��$W���,Ԓ�3�Q��.�j��&Q�V��� ;(�������b��ܤ�%�

����i�Es�sz�*�ecr肤��4�s%H"V��t������7�ߕ�|�w��mU"s�Ѡ�������F���*G�Z6T�l��a�3h3��s��<#��_���t@Yތ����.Р\8��}# 2)W�����SvB���|51(��iArB\� �e�� C߀���h@(Z�	�4�T�Zh�W��ug*��j u��t�Ǥ3Y���v�K�hx���L�����I�0�#��m�eꙶ�M���憫�بW�	�ntu�������.'���h�1���&m?Z��`����C@�m�iA�Sah����圞rJ���OC`�m�f��w.�|��2U \�.A�)W4QԯU�>lE���r����-Fꫦ���� O���|��u�7�^fʵt ��m*�(�|�=�������T(tE��h)�d�� X�ỳҶ��$h[am��9��T@��N�����&ֲx�T;v�Q�^�ÓV���,Q���M;E|�4��A��98���e`��L�غQ�4C���C���߳Zt��&��x
CSj�J��[;9��aX^y��ȳq$��;�۽�zO��q�\�ޮ&�}W�����������~.�������C����]��Ĩ'�X�։��W����P���}��_]azQ[*h��$�oT&P{��]��5g^�=0o6�-�D��D�U�sU���v�*Xt3@ [aaї8F��k�(��Sg��Tc���ݻ����kv�xL_ACD�qWy�3�A%�~3��D�+�fym�%P^x���]`��|8}�ǧ�E�$����q��4k%�(��24�ʚ�;��\m1%�_�W��T�ͧ�P��8������B7e�c��Dd����d����@��֫�a��{y��#����a!�me+��d�,��_�#�PᎾ��S�8*�Z����pI5y�S�Z���6:!�F�=܇������߽����m�~��%���`�c7���)�i�1�'���a.�ŕ$sd$��)<��"�H�����{|Y�U$`#Q]����;A�z�4Wl,l82+�/���U�!�|U�z�f���yة�C˭�c�%37��.@�rT�LC�Ɛ��>]� ^h��q3����9ժ�+!5W��ڸ��[���ا4:��u��Z�O`4a��9DTq�JP�K���z0����Wz��С&Ɲ 9b�V���VJ�`��D|������g+�&S��v1�mr�tf-'�7�DF��1�,ª�vC�B!�4�����!N/7��f��¤Z��? �h�C�|�m�;2#���X��7CEoDڄq�Grj!n�+B�	�=��lqi�\�+��v�&���bI���t{C��P ��6\N�` ?ƥ ��Ro�2�3� \�66��Z]�_�ڙ�#���+�u]���|o�h_UZ�zs  @ IDAT%!��R�
`�XS���c�C'���	����9i�‸���SsS��,܇�%:gJ��/(S8��oϻd��h��Q�:����#��O�+a96�ң�&��1k�XUx�7��bl2-���4g]H;һ�w1'P+���4jJ��T��x�?BP4L�yq(4Y��)xB��(�%4�+���UM��2>g+��jI��0;+���� ��=:�w�c\��w*�m�n����`G�M߹*�Z_�Y�ǒ��[��ۜ[t�,^�h뀣:5��Ҧ���Yz��;0�W@�B�q�����5i���Uk׻�k�����c���v��������x:����dM=9T���w��v����C�SW��
)�L��C2Og�p����b�3n��v_�������B�p�i��s������9���"|qj������Wd0 n����fY$���:��]���{�ж]��^�F��������4T�HQ�����J����他K�4���M�������Ն�>�q�c	u$K�{���!1` .���^3 �`����?�rim��rt��d �2|�IRB����I��5f��2���!���x,tr��-�S��:n�!�٨zQ i�F|���n2�m)\}!"�q��'!6H4�J~"DCl����<�#����	�1���?�����	S2LNh�s�d�IS�	"�>�\��H\D��"�k�AG�vAﾪb��Iy�#

����YE#�՞T�MG��;H�t2�nګ��#�L���|��F�����0�����)��0m�Ǹp�m%iQV�ذ�Y夶";P�z����{�������fcwm�y4 1����G#]ImM���E�G����3
�ddM���_��Z��亂� �����*ՊH
�������#�%����W5&i�NH-��
��#y��^���:�]�k��^�W�0���#��ى0E�h7gY}'��	9ʜ���`B����+ݩ�p4xJ+K�Am~ˈ��Ey�F����Ǌ�N��d�w� p ���h�ċ'B���QS��iR<�����\��V����`c�ȅyҐFy2]H{B0΍�+j���W[BuzaQ<0���ˈ5�)��v!�`ii_S�_�����C�|���]A'�µH�u�z=\�Nqn|���s�]�\Zu�B^�RP^hO��I>�fz�Ln���&NU�i������t�XI��ց�$S�L���~�v�{�O�7����D/�
��,2�P[���2�����g��t:�����Ll`�5:�.\�5��C�o��7��U3vt�αi��i��r�G�ήX���4'�$��/����<{�m�ꂂڽ����\q6��@!!_m��|L��}Nk6<w+�£������8(ap4_�|�?�ԡ�o.���L12�!�y6�s*I�
�G��Ȍ �J۶&)�!d�`��t���C�gN"�+Ҧ�����Ȱz&��=�ǽ����[�c��;~�]oi��[x���������g�o��3i�si�o[�D��>خAl�`�GJ� Zē<��E�05ȘbP?j8��'\��<��j���.��i���}���/_d����u4c�� 0�MCH�g�?�\�2�f}_����^�/+���~t����>������;?d���l\P������q��=�ٽx��>�klܽ�\*�S���(�i��ҏ;Wj��k�!�
c���p�̵�e=X�4'�G]�߼�'���������~�>*���%\�v����]�.eVε�=�a��n�;6�1�rs�|Pp��O�(j�`A IG*D^zi+�6�w|Y����������.�ڈ��bR �n����H���{�d~lx5�[m5p"I�������.�u߽z��G�{���ѭ���b��U]\��S�nM��i�a~
VJ��ޏ��{>��0:F���a���d(��jW:1�TF4���Ǐ��v^�c�>#�%��	+/����4B$6F$ _������,6;
�2�h4e)�&qG98��a��Sr�`1K�
K����WV�)�Y��x�:���ش��S !
_6R�� �o{� ]���+�>�G�%��Z����]\( 8, �-;��4��=�پ%B��)i�pC�=7`�F������hK��|������/yvT�V-�0D{I����M2��!(��6����Y�^gd�!��\ӱ�)�@?�E��`��@�\]e�6�N/�O:�n�u��Q�X��r�$��>�\u�h��ݗ�:�tD�� ��M�+���(���1e�(��C���Nܩi�7i�f��F�/Gׇ|w�f'�'ZX5?��n
2iAo�'�K�e�_)@Ux+���W�O&���i��r���EG�Gt�`���4x�k'>����f����!e�����%`sCia��kۜ�f��B��Vs���5�#�g�Hj�t�<˩������%��BRH9�� ����Fl�)h�:��&8�����fzN��o�
\Li�i����I�zbҕ�5��E	�f��'Y$'L�:�������r��9��ߜ�g���Q�;[�"?�{۶�^f�c����Ή��A>]�U�����OOy	 ʫ�ލ����~< V����?���r��I
l�(\8ēa�j�uS_��nH�g��9�}Ks�����O�!��7׺�c��|SNi�,���-�h�ƨv�>�6f^���`�?��0����J��cr���RS�	 t`U'_h����U��Z�,"�y�v��P���	�?��X���p(�O�)rQ�	B�%��|x�C��V5-RPre���a	X�_r� ���$�K8+�TVM���mP�)��+��S�V-�mB�[�~k���7�NhK�ch>�헶w�X��齝���c{�F�Z�
�㩗s�:��입VF�ը�[;�].h���}��z�+�{���H� f�_M8������2��k�MG���j��̄�,c�q�q���G�p^���?���ﺉt�V�����-#�I�gؔz�_SLG�od�Y
.RG	av(�Ua	�\����QWQ���+xA��E���mm�$}�d􎟕yV�h�~�v��7o���`��ۘ��_)[&�شIrS]����qUA������6ސ�P�[i�������D7��t�J��
�W!����5�ڒi�딉��l�*�(O6XV��j��,��<�V��J\*`H�9*�NȖwb�?*�'̋H����QxO�����S�����Z��]��D~����!�[�V|�y��}w��%��Eo2�u��j`��[�"DC0���o�C�vz�>W���������AUa��]�?|���8&�f<j�ՆJ����Y�x7�xZ��0�V?�^xW�/��V܈s�]F3M	���#B��3jj�T��o��wo߽�vp�
\�ha�<|�*�M�7V�h�$�O�O++���uV�:R>`Z� ��F{��?N��C^|�E��&x�h_��K{��������~��2-#|9e
�15���ļ`���mA��ضL�!���![����O~�q˕���L�(��U����HrttWsD���ɪiڛ�i�s;m������F(�����G8>����
�P9��K�pV)�Ӿ�l��;�UR�2p��Z�I����!'�;>���P$X�-�,��5�p�b��q����Im���=�,0<�C��Rl
YP��S��*DyH;�-P(����YWi/P��#;hy��xH��/���0n"$b:�|�����h}�/�n�o$���g6Ó��+h�۾$~{���u��4���� �i<�}��~����3?_��I����|��� AAܲ^�I�vX�uDcı*�xJw�dZ�j�,�ڥa�c*�zkk+���㇇ъ=ʀ��oF{E[*wLj��[�jj�t"�Q#��Է����M��>8#�w
m+��M�{l�>tkL�?�p�m<ъ�V�>WcW�}1@p�*z�$Oʭ!?pV���)Wz�x_qD}�l�Ү��e!�A���4p��RFޫVӞ���� +��JJ���=M��K�/�ΰ���ŋ�B�͗Z�	:�l�bE���a*��W�[$���\,����!�9(� [9��é��H��W�!+����$~��e̦�Ujz��p�LO`\�G�� r���[�L�a��0^��za�R��nu��}9�(#v����z���h���u��6!D%H�NQa�� ��="%K��#>�0�r�omeT[���L�����r瘮���E��������䣡�,�&��Z�iG8@nj�޼����Q�`@�@0��)��R�U
Vͦ�� ��+�f:C|�k��ik�f�d
�/k��t�=�\/�Vl��	��E%�)��W��Vy����"4�R~W *�E}Ng31��(p���\�F�V�3F�$W�	$�%u3"��@�V2e�Q;L���Dǹ��2YQl�fhL��IM�ً��w���7h>@$m³��$[v
v ➼��W�V��L'K@�!����a�*��l�DbL��fhYhvi�q�h0X8�|����2�+��F����q�j���0MRߙ�i���S�{h�N�rt���°�S�~����E!!�[�+�bYsN�7�]R������4���8=�
�|�|l����v��	��܉ee��y�Р�厮3�]�%L�� J~2�)ԫv|
��Rf�jGm�L����\���g���t��q��Q�8A���ʌ���ll�u��	vq�J�)CO3y��VAۊ��.�CL;f)�2k�!�4�3�r1kz.D��]�,�di�)_�
���6�N.�pu�#,��#���lb5���ږ7�g�L<��~#  =�gc��E��IBoKI�ߘ�4���ʙ4�8u�W<KG��4�M�Pt�?������k4�k�wx���4̫OP��58�cw�m׍$�����G��HM������v������*5�RJM$%R�g����RY��������"�  xdZ|m��n�Q��ﱘ��.�E}Y{�V�O�� �����,�::�$݋�w����$DL�26����'wf��t������N�YAo�4AƳJ�!��`m�~��B9
��0����n��I�c��d�h�a*?Ⱥ��}T��Wx������j��' ��(M4aV��m#h�=��_�W������/��0�,����J�nW��o}�|�q2%�E��y�<'oT�����|�����or~;��O�Ѿ�Ǵ7@A�f��(����K"� J�� ��"�=,��k���[�e��0��i��fR��c�UvZ���꿒s�Nf���$�����s�U8v�v���V�<̹�i~/bԯ;ne|R���3��5&}ӎ��9+
Ӡ�Q��+�5
`@�l�=�6���l'Ql���VJ�N!�#���4L�f�߈�1FVL�����]r�J 5��u�F�|ql���{���ϥ0~^�;�]���#c�����(a��!��5���xY�^�`=�S�L�J�=�f�1�"��/$8��YZ>x5a�Cp�6F��ځ�p.k���rVs���a���"8)(��lo#Ĺ�r���Z߄
Z0]DG=S9��)��������Y"��=OQ�&�h}%��^-F�x�@~�<fΎ*{-�@�]=���1BVQ6��oR
���I��YI���������ײ|�Za���|U���V�=ɡ���"�L�Sl)���h��3�˲g��l�Lp�����$[�ѝ0Y8f^�(�[���bG1�:m�[���X�;�Z2+��X�k����|Y�i�m�p4��bh���}�X�,��Ot���ެd�M/^�S�ދ� �|U�q��V�kgx1n�Z�U��͛,5/S�m��v��(�T/ڿ�py���/
&n5��_�1�b�@R��[�'��)�Y\Q;A��d8v�&�TN=q��kSu�m�����g�}dj������m��?�@2y�?ܻg�s4�2�%a.}l)���<��Y��Se���L��ϳ�ܾ��!VN�h�uO[<9Z���J��G0����dxx*7� >E���d``�5R�}��:�%�M�L��|����3~����IQ�uʞ6�SQN��f�8J�����3�V��O/�^��n��	Щ[�=S�q�M�t��{�R%�?��^эҁG�E���x�(f�+����6Ͻ��w���hb�jE�V`c��棘�[�)Ń�e0�Q���i����BY����M}��G�P�|��ʠz�����$Sm[��r�I��X�	��S����S�~��Rm��fx�B�E���g6	.Q�]�r�D��L{W�1FDk�!�������oR����Sե�kX�w<kk�	`p	�?K�������~������lq��F����Zy��Lh��,�um�'b(x��]VHuG'��p�W���	L�B�2aF{�T��8�V�L&���H	�8���[�4��hI%'^_{Šhi�F\�{��0��L��]��ʥ��ӈ�ٔ��� !w��G9�˒�n�%#��4��鄳�F�*}��MVG�q�L1q6Z<�z��ʥL�U�i؞�{c��t(�/�{����jg@�kh�H-6���M��7cZѹyv?�h�tJ�Qw�N���Y	j
����������zԙ���A�:W�i�[��s�.�'�-�7���V;7��'���>�F�p)��⇫-�g50%2�d�xT����:!-��Ǽ N�q���ɽ���U#����k)-�>8\�ߨ�,�J�n	��آ������y&x�Z	�y�݊9N�:;�z��U#�����Z�}&�vS<�z��`!�Y}�u�b��g�l���-�x��e�O+!���V��|��p�*��K>a�艂�#���<�W
МW8u�w�`�s��M��"��|�c�������P1p�����$H��S�.Ep��>��tac�
��İ���e1e��1�^?�s;K,�ש��f�����B��V݆;�m.8	�}l�;g�,�y��󍂵��mP��+l�B�`u����˔�y8`1��e܂��dM?�������d"P�'wV2󓊶���W[�p�r��@�dRQ�����Z�Q:�m����ܙi�(`�pS�f�j��ʧ�c�	�h�v�L��)H��R^ؐ���m�l!R�������ژհ2�杛���,��4�V���+�mҼ|u�� ����|��j?���Rp�L��ږO��߲�R���G�������Sߥ���X���۝0�6<�]/�~8������xG���A#�[0���j���~UF��V%��\��׀\2c)`���u���{j�2E�H'�Q�.�,`"�=�O�aW����)�k��B{胶�R5pM�J��)�������!���-2���|i���G��h�[�E�l��>��{������Q=�o�OṬ��|B�d��:�A�ZA6��ԯ��];�FPk�����*<?�x�2��3�E�qiC���<C�{�>��/�%(lW���q��!��Ooo�O�����4Ztm@��Y��{[6���6���I����6R}ԴރǦM2�Ձg)u�La�� ��梒�	ٵ+`����F�O'Z�}��*�ʮ����":��v$k�Μ5Ƶ��X�>1�VW9��tU~k�˜�UD��J�b�:����"�:��������zN��JYm�����W�>������^\
����C��%�Y������q��R������;wm,<��sr���~���Y�Jͧ�I
�N�۹y߼u�y��Y��)��~�䛏
� Ng��1\h���ZnXu�/������~�H[Ey�N�<���|Y�]k���x�у�o�����tW���]�Ͼ��p��OZYu!�|��ݙ\�2�}���!,@��w�ՙ�X#�F1�L�-%e?i*�^D��k[����W4��D7;M�!�	.�E�Ír�3�b�FXt)�YJ��,cW�K0}w��g��D;NK�%��#�0�s��7-�O�0ܞ����ę6�0�Q�����7��*C�b ���̧���{� �[x~{i�0)X��Q&����l����w�[��ܓ�Dm��`΃1�#��^϶����X&(�Ng��qNMa{Qβ��!g�v5e=>j
�a�S��C�gs����G7:�1��C�� &Y��F���8j�rb'��?���}�<l�a�+�N���?�v�Ŵ&��(T����!���=���0�Sۥ@��n���on��匁S��	DD��?~��w�n�9���<ܾ�s�ڴ|��D�a��h���d:ի\����2�e'��A�b��ӦhX�m�j|u|���ـ��xu������^��S�kW~����M�?�EQJ��'|���0�%EW�o����.��τ�x�4}���g�&m�i��N�;�:�{�Z��b�q�#�G�]#��l�u���Ѝ���/2]��X�ɹ6~>JV0�>�Eʋ�R^g;��W7�ǒO�DiG����~W�/�\�:-+�
�/�Ǵ��L�Œ�S�dR�`C��,��>������`8-���W�2�G������ߕ:��|� q���V"����p�i�_{?|)|P.XΟFg��k�rSrZ�h��J0�r*�>�|���f�d�p�W�z~����{N�Q OG'�zCi����~�a~~���^;���h+���[��X���6D�[���U<|�:Ր.ֱ`\L`�|i
��u��l�ٞ#���P������N1�@g5z�4á���:i�5i bJF[K�EDc��NH~�h�x1��3f���N��8x���4L?K��zW�G�myҬ)�E՚�hY�X�?O##OL�m��+�j
��2N�����x��:`Z�\S�!���[sM����d��>��J�1q���>��p�J+6�:J�7��]S�b��U������d�N�3���0gEg�Q�*cj:炙)B)?W#���+�ڻ�������/�l�؍q��(�FN,��Z��gdY���Y*ߝ��Bӆ|Vi��Y����6�������O?�Ҏ@)K1�Y�[Oe�{|���1j��>��5��7�7n~�u����==���03�	�'�j'8>�� �p��^������A�f10-��{2�:}Ã-BN��oZg��cpx����3J�9��}��aamc2�;��x��٬�D/k���Qt5S�e��z.�w�F3	���$�d��Dӑ�QYς�N�T?���tuu��<����~�o��D���3��=����l��$���o��[��o}\�(e��WSً@��5��G) ΅��?���mJ��.�B��e){4�y��1.�0۞̦H���d�&�P�˜�?���M��:�����]l��Na��t�m6�~��|M��0�8F���8��3����[�/
O귦����P�����t�����:�1(�Xo\��EK���E���ahY]����᫿v\K>-�}ޅ3��N�Կ.�$`�߳�T����_��р�<�x��4��i
qS7�w<̽����X�ǂ�ϛ�
��.�(k�SX��e���;���m#���,i/��j|�m�s��9�#��/�C�-� G�AË�F�<�0�
B���)�
mU*kj���i�!�Bahy^��ޣ��4Jӳ�O��X��oԻmyQ j��Q(`���!
$�fs���>��K!����t�n���yʘ�6[�ӓ��z 8�_	vJ���Sذ�)�>�]�i�r�i�d5�d_̑�▏��$��utrf�_���Ԭ�}�̻�2��O9.5}���>�u�p�ƍYUL��7���	9��yF�'�^�Eb$��=y1����A
�GA���8�%[�R!��_��y�	K�wi��q]��,�)8\�H�?�J���3:�w����������GVk 0U�R�ƨ�agxs������ �ǟ��/���E���[���ʚ�@(=��͞1:M:�
�ϟ�I�0�& ��p�p��Q#���u3u-D�<!?�n��+0k����
ѹ����WcO�T*�� R��6����@�!{�nȝ�M��p�.���м� �Wȑf��ꌔ:��hc_��Ѧa�Bd�2B�p���U��z�ӝ[1��9��i��'9s����g��Ǜ	�<��ȡF�I�f�W���ԋY}�v�|ɳY��1��u1�s��EQ�pd�o9���8\�b0Lt�\��c>�]v��Չ��N4���T֡W���V��_����Sq+)rO)-u�1�������#���YS4'�ҶYߌ��Ͻ�����ph���ɧ�G��;Zxopլ�����F��Q�kC��	���c����������/�����*fП����D�M1��092�xF���D4�4��㘇O�bC�p�BA���(��-�hےs����)�'�`V��1�W?��%Y���<���!�,�GY�ޥhP$=i�������ՏR�v��ʻ?W��������#�$k� ��&� 5�~mS�ڤdpG�j�!A��^SGՍ?歍(�|�8�^,ޭ�?j�����wa�k1��EB�h��������ϳ��)K�)�g���J�v�k�Z��#^�+��7�F֖כ>��A� �NT�ҕ��P��A'�X�{n���w�B��{m?�Kmz�������p���/X��#��T_�h#��S��0s{���ٿ��2
8�լ��?��Ӵ�Ub,�`셕��bP�͂��D^�Oݦڜ�A��dy�*]>t$+����r}�l<N������W?���ng������&vg���)gx<���a:�i����ÍkW���/e
X��Z���o��O�������&ZK���,z�e�_�ՠ��,nf���H�.?0�����{���|�Km���'r�
]�%:�3}�<�՚cş���7M��7瑆 >vE�|��r��'�L�B�/b�p��$��
@
8�4+��-B��?�0M����0��,C]`\�
�������O��_he��y>�N~1<������W�Ň�᫔�{�\!X˰ꬾC����l�a>IOs%���N��|<I;ʳ��)��v��Ǉ��_������3�^�5�+_���iۢ8k�x���/N�1CҠ'�����|Ƈ��E9�w��ժ|>h�$�k[���?�*q��gz�𚠋\����t�����~y�9V�+t�=��n�f��e M��?m+���=#��rt`�B^�I���6Ɵ?�v]x�N0�T,�jS��Ջ���lE��(d���6b_�Q�M���b�e6,�E���V� ���=����|��~>1����Fp{r��0> ��̷ʷ7Cl=�V�i�:��J�P<�:'�)`}(e�S1i������r^�� ��N���ߡ�x�ۙVH�����0Fs1�r���cF�[�ȩ2�E�/:>&��G�܌�R&i�6���0�!`R������ّ<�Ϫb��#�ߍ�[,3T��?=|���Ͽ|}�9߯�9'9��pq�a3-W�pFXY(��	E|oL��cb�6�ub Fs*nl�dN�m;֯�p�=���~�˭�p����>�+'�!eZ�(!�a�	f+MY�XX�^�����s���g='S�l�'���}��{1�a��+�Nw�����v�=�,@8�5�t#(Ϸ)���z��i�SB�0�x�O8�H�mx�$��? D����KXv�����y��Un�/�>��:���5������)�/�q��i)5s�W���$\YJM����Șb�~Ts9%�Ƶ����A� �6&hF��~A8��yJ9�u>J�X��V��N1�*��8lm��<���1k'C���]�{?E� �O�[��ht���$�����K1��-¡��������xG)_��b�>1d���O���������/9��/_��p����S��l�ܑ;V~Y�9x�&|�`Ã ױG�63е1�cb(`�:��qm�F�Ó���FW���W�g�wOS��o�d�.��	�o�Y�}ӂ}}�`~��K�ͦ��C�������SJ9�g�?��e�oˍh�T�ݔW£����bf�#�1<�����c5X�o�F{�}&��-L�~�ig�O*�D��M���Ƀbh���)�_j�WݗrT;nx��|��W\b�{���8S���bԯ䏗�ì�X��x ��a�n
�^8�1���	)�>��jp�%�:R�o4���c���k�F�Yg�*�@S��U;��u�z� �����������S������9GinZ7Q�y�`���7sRk}�������O_�Y����>o�� ]M���^��t��ٚ��+� ��/�<𗯿O&��I�Ϧ�����1ᴺ,c�^X����ʧ_��n����mq&�߮����j��~�V���}�y�G������)m����I��e6�[���x!��9g$�{5�5�jisK�_��E��<FFH��Uo����1;H}كiAH ?aD9Xs��&ҙ��:���k�/�Iߧ��@[�b��'�Ja@6��w:X�	D=���[
�=E���L;&g�t�N�:#�P<�r`)ܟ��\V=�V�K)���7+�bB��+{Z����z����v�v`q�����ӏ�����ѵ�ex���2�1"�P�<���O��WSt'�o}�؊�ۍ@����/����x���s1%�ϙ^���0B���W��\]Q�~���,^_��Xg�&jds���t�v�O�H{w�����X<�/�����p4Uu%%�b�c��U^-W�f�>��k��a~�q�=��ocVE")�(�L	ӫ97�43fU��d��x+�^G�F�i�#|�g5`�z�h�b�;��SDMYU�_RFg��4>���z+o�s�����?�.�n#�p��������:i){O«�g-�f��.\?>ugRН��$�ܓV�=zf*��E������COm�Mh��{��_h���]BeY����~8s @鿟I��w'��6��q�#l�hϟ��=K��
Ǆ�Cn��[�%����N_�OU�r�5���=����~n����1�_�=<܉��5�O_�M���s������A�|�s��]�\þ�MR��6�У�R���鬫/ko�����
,�G�;?VJ΃��8V�Qi4���p«sg~���]:�ۢ�Y�����ܾ��(�7۩�Y���մ���~�,�BJ?�՝���w�e�b10�zY���~�G_� �y��7
�|f����sy'>˽�־���Ý�i�d�r~)�U}�<M1N)�� _Y�!,�uX��j�T���M�0�Zq]1)���D����� <�J���������,��_V�ZY��_����̾q���,�>ScL��&���˿��o�=����������}�ot�&pO�)����V�	O�.3�7p��蜢:
`��Ū�n��e����-6\�?=�8x�V��hj|m�Tfðȯ8p�]����O>9���������|��k��R�k��|l��.������!�4���3�K{�-u7Xz�%���(a�k0@�?M�:Y[��?k���o�
����XT�BJ_�՞b��gk#�\���}����e'�4xӿw�J
5�e:KH�S�1�OY�b�T���Rl{����/�
��oW���ma�Q7��k�b�m:oe��D3�v�0	J�B���c�\�8�G�%j� ��� ���T�Ç�^g�⯋k�)�p�,�ʛ:Izw
�Z�3֯����Q9�& hlSYd}��KQ[q�~ o7m�z���k>"[x/f`4xg�1��)B"x��<G��	B�`��,R�Y����KЗ���Hb{�f[��;̯bC�Q��=��։��M/$���z�&G��4�u9�s����o��"�����͙��F�ά|�2�'��Y��a�0�T����7���hW�a_J���qN⚿���H_�W�=�;S?d���;�X�7-�ȷ�T�p2��t��w}�6~��v[��3��b���'�������+M!aF✋A2m��<X@����0��
�f�,b@�))6N��m�ʱs,\:zS�4�Y42�m�}���Z�'�_���#�Nm�s��������, �`�Z>�呂�	!N��8�O���>�asA47��]�P���,k�N��":���q�M;�J��Mۤ���$���X�9��Bʆ�`�j�i���Y}#&����<��=�}�(3kH�&���Ӎ�k����i)R���ӥ�4w�3��i'���T��F`�r����BD�<Sg���Mo=�|��vg	���y��]Vڙ֢�5�2��&��6�^Q:g������-��zОd��z<�G�?���� ����N���V���w��RR9�'��)�2rV$?&Њ�c%|R9� PY/����S����E�=q��r�L=N1�����ˢ"ֳW�FU�~�S0��:�����KW�)���jԿ���l�a�+��fV�����9��ʰ����q����m<�J����Qm<֮���5B0XXb(Fc�	fp��_6�<��vDJ��ŋ�}hL�Z�x>��������|zk�1]eŝ��'h�g@!�G5x�Й��;�o94o)�)A���%��$�k!k��j\4���3�Q!��R����7�C� `gB,qJ;�*����L�V�����^��s�OS�����~�Q�R.� �B�u�c�fF��޸q���^�s/x�zQF��Tw�md�fU7��	A�f"p��*|����m*ݨl���q�Z>O��c�3&�U��9��`��E}���.hz)��ύIx_��o�Qc���j�-�ޯ8b�D��&�-/��7w޹ߕ"���~�y9y�n��i��{�r<�E{�س��:��-
�b���zV!&�EG�Y�fJ.�왹��fa�:f�y�Y˽�:M �g�� >u*��}�t-�����0�U�����J�o} ���4Ԫ�BG�UL�N�X�zo�@�FM�͘�u�IJ��|:���2k����C��v����v�� ��p�5��u�~�>�z�*9��E{�<m�ȗ��̈��F�7?� ��M[�°0����yk`�g�M��2S�cv���í3M{%��(1�}�Χ����N�2�)!s�Q�28V�n8C5ZRyfv��ʹ��Yپ��Ct��K9�=݊�L�5�t����QY>q�r�m>�8�o_��W>|��&r)�Ͼ8\��Q�E��eǵ�^
�(�!x,<am:|�o݁�������6��"ڤ�D�kX�OD;�YB7Z�rBa.b-��׷	��)?'��]
����I̞q����t~�)���r ��'Y�*�mx��w�}����R�l�0A���I�E�g���fӷ(��|��3ϩr[�;FU%j/B������K�ӈ���Ch�M���١Y��/��R�	����p��).�ףǭ(M� ��Yw�������j���;����o��6,�de�g���M�����M?6uc7�J����~�7&̟K�_�P�!�2^j9����C��Y�B`Cէ=��j �se�og~V7J1�>������ F��?�B�"�d�֦����y�t�ijKFΤ8���� �P�]+ �A�&�����>kP0֫�g��/�4M�<xǗ���"�Ņ /[���4�٨ror5��O���UK�&�WSoR��;:�Ό��s@kY|�����;M��������j� �n4jݐ1SUw�f9�����X�A9S��D�ƪ!�sH��F� ��2���M��
�p���g���QJ���ơe+����Ž�k���t[�|����Y4@�,8�*�k��\
��:���?^�f�²�7���(��c���6�����س�K��	���i�چr[���z�_m���Y�z��ׇ멵%^�����c%}t�G���C�6<Mc�`0�3�	�,�`Y%7�;��׼Ii�-��X�ӹp��N*aY��x��U���6��o�Z��<���a3PS�)T�u��\4/^��y~��/9�5Fl�  @ IDAT�C�.�[��}�`R&�̆����آ!�y)����b�S,T;��Yσo�𿽘��e7�}y��V�__Z�;�[�����MHpDtH��8�o9�|&q�>�ő�6S�y����כ2^H Z0�>�R�q��:�G!+<�=¨���h�,AJ�t*���q!ݮ���P�Z���1D+[��Z����L�޷Zx?
X#d
ؘ�G��*3��@_�N6�BY}�{���,��{ܥ����$Tl�h��^4_[H�{� g�?'�;(�����?��I
��f�b��a�Ѧ���<��`�c�.%�ݾ�w�xV	�t�W\��,F�*K��'7�̼_8��1��}�b�c&�*)K�g�#�|F��ھOwv�w|�XGO&�4���/j��,h�q1g/\Iٺ9�RY?s�����Q������qD)�+��f�6w8��5G���
����E�$xZ��~G��m)t�DM�ݵ�6g�٧k���y�3��Q��(�u��U�T�ڙ�9��|���	�-ſN	��;c)bY;�5�ʵ�����	
�x�Z1'J�-P��"��"�"6����Eco����� B=��]_�1��(�;{��%D^;�y���ՏS&��`_DGϟ���R��!�c�ڂ�-7��B���G3�����_w��M�_S��S����Y=N�sH��:c�+����B�Ť�������~5��SjY�Lѿ	>#t���J���@����r�g���ń"�+�_h{��L�8�҂����g�m֣�c�� ^��c�k��
c��W�qdG�F[o�wp���ƚL��j�����6R.)��8t�Y��d��,+�9��b����Vwa�1�J������>�j��_@��p~����A�������(����;�̀�J`��X�(2ng��pp
�W��mm�iS�A�_V{¼�>�ˆsr�+�)�K sȯ��g��25�Q>.�omc#X�5g��z
t2�ϔD��e2۽0<L��/]��Wc�S6��J�����N+E��o9��L�aPGAVVO�%a���QȢ5u[�kla�((��'Yk��9�'|����(qɄ��ף{S�|��{Y�l�LY���b����J���J?��h*k��Iu�$�N��).U�@���A�s7�:fc����f��gCo����~�͵h���c�/~H>N&,����&��)�ڇ�S�.�����.lfK����и?�����$^y��5�x^M?��bl׏��<�{ģ�&VT�
�-�VDU
dڰ?{�O�
�14ak�y)�T�"�b�tӎgS��w؄�|#̖e`L ��t�ɽ�ǂ�}:Lq�$P{��S�AL2����B{�-I��Ƥ\�S�jiܹ�!�2⧴I�u-���S�O�V�l�&Y�չǌ�^!�s��.���1��x�)�o����l#�s�:8�тKG#�q8�j+(0��Y �!�kt\ÿ�-T�E�B��2�g���Y���s(�X�ڲ�Q���8��s��cU����,
���ߗ����\�W.m�3m�q&u#I��E���_����.,�8RCZ�t֡�A,��l �l{^�vpK '�N&��N{����X<z�*N�S�d����0�����l#WL&�<�Y=d�X�9YW_~n�|��ᛯ�/n�:K��wC���!��W�L�3��<��tg��/Xܹ��V�7�����^̅�%`�% ����7!l�j�`�݉G���TH|�(�Mv���7%��"��~	xm��[u5����^��)K�% �C�~��j�n=�-�;�~xG@�#p�ь��+����� NM�88!Qm_K�2�U7+����z[�ߧ|K9ʗ-*t�s.e��pA;�W[�)]h ��l�Oo���脉�kф�}�tx)>Z�����}�7=$T�¤L��Δ��hZ����@���9����,!�}ʩ�|]����>���i+��䩄�>~��Z�W����,���l��f�,�`�����a
�T֋��.���C�k �g�־`��wG)1,aV�W��^8����y�X��CSW�:;�o�4�,�(R�|��h���4�ۿ~;���;���:|<�,�tUu�fa�(�Pt�r�4�~xʑ��.���و$����l�;���r��W�r�����o�����/�m��^��C2-P���#>���^ŋB���/w�5˄~2:R�t��q��sNA9��h/��5��trڠ�U�Q�f�S;i#%�&�4�cKn|�lV�"�d[f��6a͡в�ٷ�ĉ��b��۬�A��+%�%�>P=��S}�gP��A��5A��Եdho0���#��}���t47�a�j�Qz�O)��o�O[�����������s�]��oO�us�-^gc\ʻ��oyT���aRn2Qd���u�vkĚ80�R��Ciy"�o_���ZvC��b�E����J�SA��h��3����5��q)_ū��),�/�w��g�m�s���=����B�� {��ŕ`OTF��C�^״@q#r���
�"��
�N��E�gB'�B�'	ZS$'#v���a��Qg�N����yO���Ɯ�,�?VL%�W��v"�T0�j*�����������{oT���G������S��W	,y�Z���7D�CTW
���La�'n^�=���,ᅱ�	C
�8ï���wp��o�=mM2��F~�鞫ڔ,���/\�=9�@=�I���c��l�S̉*^��ōi�J��f]�+��~����0v<F�Ց0��ʂ�+��Y���Õv���Z�g�O����.�&�ڤ�C���D�@xU����}�3ʓ��/a9SG)a�X�08�+��'���#��b��(@�Lŀg��A��S���8ڿ{�XE�_��8���c��V�N�Yq�͑���T��n���
S�]ɷ���a��l]S�Rm���~ݣw|J�&��n��PT�\Ԏ�U�˦8��,�W�O���Z��Δ�:�\��Rf��������-��C+F�;.�fI�
WH����]a�Cx�r�(�Sܪ�j�	�xS�>)'1n&���g|r�C�:���۬�e�U�l�qϨ����go���YS����K����_Ӡ�[� �a����M.�`�B���?��Q&ݨ)^�?s)`�@lEmG{�"��N��ld��Ӷ��M9����4�Q~�G�9d�����w��(���N2�Z`��TV0ӹ�Lϲ�?���u����B�G��w�ڒ$���5���"~R��$E�3�,�\�Z}nqzt���Tv����n����\F>����)�� V��
���Ĵ�>pA�/J0��M���ǟ�>��AC�[�JƐ����)�%��(uŮA�?p��"l=�����o�myo�T�v�!��;Y�b�,%���7�V[n�B�����2����sXO�o���A<c�7t��߅���B+�z7�z�O��O�f�'b�O��CA���0BV�w9�ˠ�>�Lz���q�wSJLJG3�t�B���Lg%��7-�d!n�J�⭆�}A�w���Ёa�W��z.n����Z��+p��dVJ_�*gK�����!��AVU�a�g�-|���m*�1Z�爝�qdJK�4��9���$0%�O�7V�F���m�pu�E�yQ0��q�A� i���WF���jY^�� c��NA�AR`*�rF�0.��c��`C`�B9�3��~Ϟ/p^�5m��7��,���Xy"Z�#�
�-'�]�B�1�,�+��4�Ⱥ�f_���p]�^�9�i��i���0J�:ңv [8vb��r(ƵW�#*6��e5`���@5���TʫM��A1�D ,�L������G�L�Y(b���D���(���Xݠ���o}k�2�S�z9Em_�C�/�4�<��`u�W,�8]�0%�O�������&�ˊj�c���Z��}��ʧ��&<`F��#����A3������Fu�#԰4jj�E�3t�����(,O��K)��XKi`ٳ=̫��Zq�&|YemH|��}^%X�����eS�����JN��Ʋ��)�ߊ�$��g!���ҕr^C�#b0�E���	�U/�����w7�+^a�b��t*�V��O��^T�p7�+t��5Q� ����\3��	L��C�z�Ry���f��œ�zX�q���_���a�µ�
�,�PY��a>�L�%+�0�ϔ�z����T{Rjb(��gmA�3*�Zim:��o�T~��}�>bd!�~3~��k�=4�쵲�S��)�Z���������ύU�:��f)|h��(\Nu�u#ژ�b���>�2��g��וg#f��g~��^�/_�h0F.���p?0��`��3����ٟ���)Ȼ�mm�Q�N�!+�;�)�取2U������H쯥n{��]~�X����k'��]�*�J"����/���5"Gj���.��#�1
�@��|L���{��W�xr��>�,۫�=n�S��~�[�#�ު�+'z	�H���8ݼ�.|o����L��+�B�{��/?}M&�lqz���@7xܪ�D�O��PZ���U���?�Kǧ��H�F�Na}�^�t�8��:� ��BHCd��8!��K�Q��� ��2��Q�ri�j-��w��t0��%F$��$����2{�p	
9o�8]�m�˪k�}�ؠX���+��W�%rVr06�se�A8���x?�T�o�,'�\D�%X$Xy):/�p����D�k��`��.�Z�X:~\��V�пi5�\c��>�H1����l�Wv��`�Xn�Z`�v�״����6SI�!@y,���Y��4���0����`a2���*l���;���9�ho`���Ɯc����"Q�uw
�R*����b�����C��	���	�,���j�
^����е�|V;����dm�8����1���|T]��2����]1��3��U4p�k���0)Yl�Y�,���8�&�	�Q`���NT���3fc_��0%���ʫ�����6XV�E�T��X[Px������	���B�>|�5�&��i�~�Sy�ߟ~0|E/���m�1�3����s2�pu1�du0���Yc�6�c%��_w��Q�e�1��x�܃�;\��X �=� ��iB�>��W_�d�V���ch�Óôg`P>��C���ѵ�4~+�����V���>C�Eb՛4�',(q��V�R��p偤LY���3��;�?Wܳg�T`B������%�j_�O�c� ���Ϛ�V@��o������=&��M��'�GQ�_Za
?ܔ�1�����P�v����J�]½��cC�)`c��w�N�I}�r�G�.'[8Z�l+����,ާO�<َ!XֶQ�Wc�o�h��;��z��ҌP�������
'�d'O�i��i��������b<��Ԯ��9�e�����՟%��o�55Y]N4s�m´�1��P�j4�
X0�����C�j�5��&z٥ľ���l�a�[�>B�[����� '�Ff�~�+7`V�p����Poq��X�OL� ��N��&���Z���~+�gi&L�	p>���?�59l����P|�"nuE�{5����bb��h@��� N%�)`�f2YÝ�1d}����隈g����p/�>�����5���0x!�vi���{� [~����M\��������_������/�Á�Vw���#�J)�|`���&��<0y�g��~1;��^��R�|1?4�*�zŪ����۴�JP˛������;&�>
�ș:f��w�7�B����ރ,W]�e�� |f˅^bj�OV{K��9՟)��ø�$tu��rZ���>L1*�|&���)`�Py@*����^�$-�Eث�5J�*L�}����N&Mp���T?S!R���K��^��8�d��{����jg�y"3��d	�W,AyLw`�h�;>?'[ql>{meg�1׾	�l`+q���*��+~`TL͵����;��^O[F���LzN�ډ�����r&�m��:p��0O(�p�\Q��a,�A&�Q\�v����On,	�5�o�E,��-��ۤ��ڞ���o*��*#�S�ԥ�Pӭ����ń��e�# %�)R�v��X�i+��,:0�xU;=�����V�^k�Y4�9(�k�Y�G���^}��M]� �T�X4�:�'�?h����\.�H#'mY2n	 ��?Y�E
�!/ūgڳ4�m@J��t%�oq��+�+ %�mS��]#��r���ͱ�/�	3���~`F���t�5�VM���s�\�x-J预Q�X�N�GgaL(v�k�E�H#�Ok�^���^��Ee��p�_�E}�"�lգ:p��bOW����y7��ن� �����?��#���'�Q�X�:�<�뱅 );�8��vZ�a�ӼN�`��U����i���R;���{f�!�;�~�����^"��w9�]_}�g���^���.C��5��耼��̖��Xue�֧���vChR^������×�c�dЊ��6�rí�
�)�ǳ�9�H�`X��f��|4��런�Nh�߄y+g\^���H��6����`��o_����w���������x7q��~,z�Rmt�.��K���K{ӫf Y�z^�vt�pR�W�*����>*-�) �M���ʬ.��zY'ާ�����M���C���@<�X��߼�|����U�����b�Q��_q5҂Y�w��W&�l�o��K��7�I�a}�������B���D:�ZY�àQ�<��g��L��H�>�T�Ө�LZ������WQ	>�F���N��	.���Gf�ޡ� ���G:8sQ��
�3JS�
���W悦����L�y(�S�������ض� _�z����͡��~-:�vL@/�*upԭW��W��*3�C#PY.Җ��o��`�ߤ�� ��V�eY��W���M����r�?��}Nc>�!`M]N�m�M�t��)��4��;F��Oc�c�#�w�L��h��Ђ2]S�-ւc��:��}�m�i�B�kXW������&\?� �<tM�apнf�O����A��aɫ�([��G��j��f�<e����購*s:��"�]��~di;�g�ʙ~>��c�.���Qz}e��������4��]g�����󹔼WY�X�^��������瘥-(��j�w,�Y2����EuWG8d�>!�wV't�0N�F5��F���S����W.�o_J%���fꭸ��&-\�Ԛ��5؄�)��)�'�}�Rt\,2����U?���D#(�?��xR�2�5��*�@�\��,.7w�3oϦ��a|�o�����ڵm^FfD=䐯e�tZ���
��K;����p��oK?�t�JS��~�Y�L{���6:J������L��,EUU�w�˩8�����G\<��H({�9Ks��QUi)K��~/K}J>����<��»U����x���%>�s���͆�h��i^�hH~Q�R�z��tJ�,�V|�6*O�̙��ƕ�B������oС����sW�aH�Ki4���/��mY��ą?m3m(��:�t�Z��0Mn�wSA�20w+\�B݄	c~l���7_�%��W�y?�n�Џ=�)p`��-������-c�{C��r}�o��
VM��4j�?F0s�	ɪا�M�^�a���0�u�i�E�4̦��\N�ƛR�����w;���M���Pbi���Bb+�z-�T8��X�K�05��As_����B\]��&����o��`�`��_��w�Ѐ.q�s/N������6Z_�B;`�����N��|J��I����Y?zW����u���9W�{���V�����+m�y�U�I?u)>��J�]VN�z\0��p��Zʏ� ���̅��D�������`[��@-�U�>
���I���s�?
��r���9�~W���}�7L���]���!ia��Q��Ì6�^0.�ʅ�)�_�����%��E��im;��
1q�[>��jw��F h��Tn���ޗ֥ݴ�p8�B͏���º��^�e��߶�DC�`h�M0�ϲ��`	p���0�7�[˹��8d�#�l�9SD�"$
=@lQF��曕8�����`1kϴ[�(q�](0(�C��q��;(�⓷�\%��S��n����Ꝡ���ǈ!�v0����e�h��)���i��^�=�8c?��S~+����G��^mg^�e5K�o�iϦ�8�gZ��m���y'Y�*�ReO�smG�������2�����yL��ih��*����5���AG�ܻ����W���!�v�*ъj�>˲�T�?� ���~�M�Y9�j;��
�ɬ]/]>|����Z�k��ٴ��3��W�p}�?��dx���]����PU����>v��+���賺��~|�#�A~e��շ��]}��?�����'j� ���?׉,|Y�(�e�w��;G��D���-�s�.���6(����J�Q}Ѱ~�=�"�p��Ct1��F�6:>�te�������_K~vP`�W{����� �;����G������_�ڨ�M���(����pRp)�a�\�fi��G�	�r)�.³�Kɟ�U�g(d��R����=�2Ur�'v�S>�k�i��Q���p7����^�ߛqQ��01���\�����Wv�ε�Zrc+V/���z��zX���'XL'�I�=�3޳ޞ���{��rh[���|6��V�2��W̛�ӏ3�1c�?XI皊y�B&���g�@��	�~��)~ş����xV�q�)y[���{���{A}~���8�� ��������:�����;�w8'ǉ\�-p��X���7{~D\�ˈ�[i��rv�z�oK,��N��;��]��y��¶�N��=H�c9�'�D��$�<="�zT�k�iǞ� f0��
"K+�-bO�E�s'x�D�}���fG�O��.Vغ��,�<)~͡�)c�+k�Fga��S\,��Ji�ؖ7�e��9����{kivl�z�����!�(Y�f,!V\%�N��
6^���4�c�	���
��~�4hؾ�^�Ya"������X>�������!;}0�����b[e��)�z�ߟ�ٛ��Np�ؾs��^>\�l����\z�^A	�U\���"E�l�ގ;9q�ޛv������rs���ӭ4[+���ʶ���(�a���F��Yن��+��(�Tp��gΦ�
J�̆��U6c����c�>����)�O�����2b���)ĳ	d�_��7:؞���n@ݽlU���}������ݙ�hvm������ڟ#�+���Ca<Y���o^�z�򳛇p�<�o��(�?�4N�U�%����?���?�H�,�p���`h#�h�f�J~�bͲ�bw}��~[\n����^\�/3��k03te}w�� U�JC;��<��/�H؞�Õ_�yZ���+x) ���΅�h���^��vY-S�C_��������/8�|�*��X�����O5���EV�S�K0�)��2�g�Tb�@/l�aʿG=w*	�⏅�U�A8�~[M�mceS���~���,���U��z��b���������G)yVN�b}�|�L�^�T
/A}�ϫp�`sJ�(��G���� �R�����]\4B�Z�X�S]�;��Rgnڤ۴���2u �r��Z�T=PiuӚ�	I�8
�ߕV�E���MKᅧ+W��t#ߺ��I�}��|��}��N��z��|v���W���X��o�urm�������_���!�<e�Y�#�_i&�y��x�c�w���5e�c�3�[pϥ�Uף%˺ɉF�����g��H�Д�4#(T��g��2?�X��Sex^Q=Oh1��^a�.a{�[���b *���Λ���{��	_w)&�O��o�Z��qV	[\���nUd��h��Z��<�N��w��4�ـ����½@�v���c��q%���As���y~�P	��_a�}u=��lo�`��_ǐN�⭔[�mu��j �#ejM�UBiw���+��MHa�>o�7A1�
�k�(ʞ�z��M��,���DN#� ����d�ږ�p)`��޽z�%�S?�!���o1+Sm	�~<F�gj�"��7���,h'R欆Z{U%�:GM^g�)V� ����jv�	Gޫ�j�������=�P*e�+\�q�r������y���k�/?���;ۃ*�������]�;v(<]ho��7������9���J�.;��@��$c���_�=Ӵ�=/��?�������?>��a��5��qXw���t���(_V@��ֱA����O�c\ �'g���O����#��?k�MY�b��[�n>����o:���_�6ʯ]ﵛ���~�f�,7�B}���D�����OR�RN���:�<v�zV�K	��ׯ>���>V�zၲ΂8��F�QX��&E�z����n�����çr�C���o�8|n��]h��v��ҩ�Mw�Q8�b�_�I�7�pȯ��N����>9\��n���?�x���?�����6�9V�����y������͎���� ���V��y���?v^l'dy��'�n>��o_~��Z/���&_�:A[1�@�@� eH{��.�z�2[��Jy�n��;��볕æ�L}Z1l�e	EԦ������*�lQ�-�c�*��J�
뿸�'�0�S��w��O#���>F��})z9��؆�u8�X�.����H�r�Z�O/������=ȏ	�-�OY�Y7V��ۑB7�_��|S���m3��r4y��}���l�Km�������xD@�WO4<��u��G7�>�jy����_���?G�N�(�p�=Q�X٠i�ʋ1��e�����M>``���\�X�Q���᏿KQ�\��������u����ׇ흦��A�۪�_0p-�[�(�\ӯR?����a�����G(F�ǯ6�t�N/��`���`,��[����@F��j�!/��׾\���d���F6��t�؀�����u1�64}�� ���ـ����R���$�F� ü�ۋ~��y�#nwo�}q�I��&ӹ��G0NО����[��/����^(Ԭ���?�)8�N�g���[�{!S�qC�SqJ)�@��D6yN��	W���]+?D!��rŘh}�3�m�����D�b=���=��PX�yǩ�i(�U�����n�M^�7Q��q�4OS���O_��=K+|�}"ͻ�~��]���c�}@}Ҹ����"b��͆�C�h)<q�)V�%L����4'��6aC�t)��v�?q"kCJ�MY,��@�@�� d�4J��X�ް��&7�=��V�\��.�ۢ�ӆ��M�&l�u�c.�5�<o�����`A�3���t��On���O��������)�1�n���voj��H9���%� Q���hM������$����d-�rp.kх�[@\�$�������_|Z+΄k���������:T>!����u-e�,ƫ�o0l��T<��]��,a���e��iGn��ow:xΧ0|�r��nn~�A�/-H���?��G�O[�g�¹��O>�y���%�n>LX����hR��Kx���ne�)#u��f���\��CE�xEqO!��`X<!�
���Au��Bh�p*����FG��|>�%i�~���H��k�]N�	��RRX�.D��?�t��on>��|���V�����~��M4�ΑS���V���n�퍏>l��2��򣄍 WB���3,/���ܵ�����|�8�]��t~���M[	� �������]����f~3y7o}M]���4����:����?��F�cP,(T�[h��ɻ���;o��\�q��E,~��Q�J�C�,��Ŀ�[C�u)�V��������?J+I��5Qq�t���۠�����,F���M)6�ejk�.-����߼Y9`G5Mw�&����!�'�����z����N�����||(�����p?F�`fE��ݪ/|��'����o�r��������֗��]��y��O3��MU�P���s�"u5���>�[5���������W�~�q�͎Żw���	ngy���"���.e����E-
Ze���n=��D�\�w�x���	�ߋ��w��G�������ٙQҵ�qǨ�5`���_�ߋVyh,�AD�3N�M�0�:u���z���B(`�ō`�d��]h$�����_X-�����}��O;ބ�N�<�,�cUH�{8`��W�̵ ��o�~m�x;x���Kܐ~�>ř�V>[n�d��}���Ҭ"e�*Q�k������ȫ��<�|v\l�<{>�iW���A��xQM/W��Ѫ�N���A�v�@N�>�tҮ�n]��rGQ�[�+���RJ� ��>�m�m�t��.$a
.=@��~Y���*g�o�N�E���*�i)���&��w�;�3��p�UB��V~x=�j��\7�������/��*��wꨧ��ý��i��[>���[[���MA4�²뜶�{G�3
V
�(b���]�콚L;N��r]��S�����{���I!+?����q�JJR�*ۙ���~�J���yVxeͰB� a�;���F��}��:V	�M�c����(G�}�.��x��a��K����gu �L�Qx4���)���:��bmlUX�]���w�U�h_��qhe��0�O��{���ۭ�>Jyi���br���M��X®4�h:S>�����2~�U{!�����t�Hݖ�A��L�u:�Ƣw������>ِR�#b:~X���O���~���}�$�;J�����:o��b�i�w��K�9JI���z!�B��8�U��YJ���0U��S����8�y�ii.P��g:�T{a1���{E��dJ�`/S�������s#ɟ�����b�l
>����OYE�P?I	c�6]g��:X�uy��k�-�r���3���*A�l��
ӕ>|bz��3ܠ�_�&���6u��YQ�5�n�΂�Zl��	�V��5}���2%(�"8YGg3�(�q��\��h;�nJ�f}����7�����"_���);��sx]}3YV�߿ױ`Y}��c=*� @��#���v?|�.6`��ʕ5��r;�}��N��;W�ƍ+_~��7G�_�Y���R�P����;��`�qۗ?�\^��$�9e��^��L�o�=�o3�<E[C�e�l����{�B�����;8�/?�����߿/ږ~ޕn��>ټ�D�)�IfhX}�)����7#���G��o�̂5Т-l**�+�3Y�"*:�@��\pQ!�����@��\(O�=��C����<&d2�U���͏R�����v\�J�7��l�#/��:I/����w_@���ĵ�gZЀ"n� 
��y)��U�	W�+�^���5��h+�=�%����g��c����o��)k�fH�/�.TXD��I.�<a��{^�ŭ��Wx9V
�hf�k�߳>ה�ނa����E�>�#�����d���i�5�x�Þ?��e"E�(Sc���/���3�'��x#��4M�e%���>k��C�SX^������t����Q��_er�$�o��fg�|1>����2���6�}��m�7�}��I�,�5aR�*|��~j����p|�8���!b�g4+�0�W�\��1I�6�4�Q�J�.�?j�˦N9���o�o�!ۦ�f���Y�nT���G#L�5��Hq����5�)�s�*5V��9��/�gd?��M�s��a��7~|	J�F�b�bE��K�Ք���fN��s)VY�&����wy�u��[���L���.+�=�d�����5����O�: 	)N����w�޽�&j�=j�N����}X�(`������vZ}�~��[�3�|��{4|)gvrb����]��q򾚥M{R�(�;����>uX����X�l�ڻw�D�o�v�'Hυ��yM�����S(z�ZD��b�U�΢;SP�����:��Kw������ڏ�G�xwxz�)�t�i�gf�ά��R�.\��~���]��*���Qt��X�(�dZ46\ ��la�?8�ʖ3@I�%,]38�a%7}9��"���5mfB��؈�X�>�;EIߛm��di��F���;#����~x����G7?7��X�(bh����-R.m���E�j����]S�Y�*]����?��ߦQM�R�m"̏q�!�iO
�լ�7��R�_�h����x��Xw�q���'Y���^���vR����p)k�l�����A�)'�|<+.��HFǗ���S����u/��'���޺���%�\�(!��$��M�畻�{���;%���&z���UN1��Q�������[��!�a�2�#�E@����F�.�H�U�-p��d�����R��{�/*�+�~�A� ��>e��������o��*�d5_+le�թ�U��9-PvH�4��b+őV��L�3������
��	���6��<+��}~�ǔ��n������ޯ�&����R�*jW�-��Rm�U2!��@�� T�*��D?���,S�8+�I>o�+�=���V����Rނu�oB���+�q~`�L{��&��I�ʅ���^=�O���6���>Nq�s���_���Ó�g���f6��q�`����������$�!_��ֿx�{t`��Ǎ޿����W1�u�য়||������?�����q&��|��)7�R`�cK�w(0�2�S�i�A�L��6�������L�����|`���L ���)[2p@~�4�����W�~�����ty�r�*q%��^��`И������(���/�M�a���M�=guL P�XY�޽��H�����g�4%��'�ԝ��q�����|b��)K���1V��?�D8չ�/���v��Ʀ�.��P��/�BAsh7�!��������m�/}�2L�w����e��SH�����Q�kN�	��J�YtQ�R����j��� 7<�E08��l{o�(]D�1�M��L�6��,�����9�_H�����7���}�b��>Y��J�G�ՠ�<��,'��/�Lk'J���5�?�}Ѫv�T~�����w
����U�b�H%��愂���U�~|�0U��*���(�s��U����)'�hl�����dm<ۃ�<�b+�}jt��^���C��*��pS��K�Uek�{5��l�]�=�x������>�O�_k7�;y����/L�q���/�j����ch�O[��V���]�Or��w�_��h��z���rf��Y.�y���{}�r��k�>����g+_����;4��#��s,�*�#C��k�-���=0Gc|�X�}.\p����"m�0w�e�FA�~����^E��&ޗ>P�y9uG1�5r����U������~a��������'夙6݊��o�>��2wQ�}�UJ��䫗�����]��N�[+C�h1J��<�wϮU����ƚ<��8�����Tpubl� ^�{%WZ�ۋ�������_�N�ۻ���c
(�^Ъ�q.���r٣�%��d�BV���˫	�{�p���qW��w�
�
Y�!����5	w�$��)���o���B��D�0тa�q�+�(i�D����.0(g~���	���KuR��p������O;���k����r��m��.I���h	����X|.K���']9|��sp�,P[f�8�t\�t���#�cf�	��a������ʋ	�aF�Ü*�t��@��3��G�+󣜯�f�j�̋����1�BcQ���M�R�yT���.k���qEN�*�3�*�ܦ�^e�;jZ��ֲ�@`�˿��U~jMѾ�������M�g��p��;������~�S�pF����D�lZ����Ȍ�[ui����ݟ�������'f�Bq��6N�ǳ�����YC��J�9t6鬠dqK����:���"q���X>�k�]LR[���u�c�
�6�$�Od�8����v������бU��?"�������$�MI�˚��T���ǚ�դ�	��@^=e���W�C�h�-�v����7����R֕��7�ž��O�<��ʆǬ�	JSShX>h����<wVJ�Q�  @ IDAT!}:P���p�'B⺲����|s�쪏��z�s�8:b�SW����!�0�
ؑ��NX�()c-�#��/�+m<>C��^4���~�!{ɖ �y���[�ڗ@:�����Z3X��='w�|�T�4a8�a��c��X���b��a�fz�Z��M�^�z����h ����.^�)�+���_~�9?��-`��*��0���Z�O��l��u�iC4-O�P��q�Ȣ7��?e��n/R�v:�N��J[��� 闬���Ac�^c������ր��G�1��^���(�R��a[`w��k������@�|�_�W�L}ig�h�ra�]��8��?���E�Hܿjy,�����&劷z�dXD��>pWq�([���D�Q�Rܮ@�x.w�q!B؞�C*0�ھK���z{zy�LB4P�<O�U�D���5����7X�{����+x/~@�t��@= y�}���q�^���Ȋ���	�FK�yջ-��๼��=	W��D��*p�t��R,8V�����=}�d[��;�Ni{N{���������@5:�k��y������Pw`�d�>��1�|��ߊ�h��m�`�	~�3/�I�0�[�f2�v1au���S���1�31��m�F������1��Oڶ���ºfY�*�d�O�w'!�"����h�Y����'�l�6'����6���y~;�/cw�]W�$��� Ip߫XU�����#�|���9������uz��Z�⾂ @��O�{`�H�}���KdddDdddf����>�D��BX�Z�@��
\@�JIj���0
���>LNϹ�(b1z־z/rJ�t�a��^a6��1=UÎo��΢u)�=��uR�����W+E��Fb5�հĽ/���?���3�k���d�;e�Kbuq��;�r%?Cq�����'y���ì\,��}�l�a)`��󦀽L�x��qt�q&�峆Ƀ�^fhFUq0��k�
�!y!k E�⒈�Ug��L�:0̗p�`����2�6%L�*� �2Y���~8pG�)���X�� SG���$��5���Iu�G�b���0c����{?˞T@me����.��0�W�Á��q[�l}�P��Je�c�3DEPn"��1�?�>�F�F(e�a$���Ǵ��K�������̒�gSV'�p��^e�-�J�� �^����4�!r�_�AW]��`kL�,���N_�ñ������~�/~:��]U��Z�숞�Ic>M�?��<�[0y�Ur��^�(ͺfh"i�H�
���%�;׮u$��Q����)���3���eX,����d�.�bi���S��k�^���6
:��~z������SG���?���pE���ZV��cE���o[��q�P�ʡ4���ñ�F�p�D[��(ǽQd�l!�:(c@��]@C=��F^w�v8V)C����z�+ທ�|�g}/�n�G�o���X��6T�護+�ԩ��]��}8����D��]��!e���7��� Lh8beȓ�!~�6���D�K#�Jwފh��:
Ť����Ig�!~ާ�9�p��JûI��)�������`�/%�ʹ�Z�eW�ݗ]��ڽ�o^��+u��@����Ľ���*����(`�0�W-L��%N$��c� ��,�4���R�{��>o?�_=�s��~�0�ܥ���w��@��s'������/�8V���X��!m{��٦�{Y��.���j�P�t�~Y��ể�؀��`�C�d�:�PHr3�A��y�'�	���°���z@�k3dci�˗^6t�0ƹ�`|���*��+�ےf�%�1��n�c*�ˮl���A?J/O%�LSy����71�̫�)4N�̀��Q 5Y�Y$|�&9�R(�c��'��0�1��&4L���ŏD
��?���'���X�����C�T�e�>^c��a
��N��Gy��I�t/K��v���<	1E�?��B@��%��d���wc���%�}>f��e�3dJ������B#l��ɇ�<tE���E?x$��m �$w�"�^��a�I�� $P/7�w�2��]�h�)S������T���:���c�DW��cf�%
(N���!���!UC�fd��L���f���(`�!�r�),z[B�B+�S����V7Br��
��ߖb(<eA��á~(ÆEa���*4
X��h���i��U��7gEih��G��z�:V����=�����
�=�M�-�W8�W��o�.�򱭗��)��)�:8�&6��dk�Y�K=£�ɓ:#����N�Hʑ�f�Ni��k� ��a,�q��<?�
�,����9�[�f^���U�U'lQk7�tS��[����M@�f?��X���m͐<�Y�-;���8v��~=/ڙ�}E��k����"�D��p�o�����K?�Ϟ�0�>�tZ����gU�����z�Ғ׺��"̣WN]�	�S�����r9H��E��YZ��p��f�m\�"�u�<�.�a�o�W�E��G�A��Q�_ѕ�
�����9N#2ٞ�8��o_/A��b�1�v�m��w/��#�m��X��z�����9/~�E>�$�,�T���qb#a%�\=���U�m�����T˄۾����ӷ����y�!8�Ƿi��6䊻�R��<v魔{�ݧ�v�}�S���C�0��"a�	i��as�t�}W'+;����ug���bWZ,����)1
G���P̬���94�*�R�Ӭ���������9�1!
X+N����ޗ�+��Q�6��?�b�-e�I�^ʺ` ���R��Y����$��:)��w�h;��h1�0۟���w:�2K�EL����|;�)y���B۷��Na	�1X��l���U޼x���[���54&)���y%?~`�1���a>E�T����P
�Y�Em�{C���.4㍕��E�.\���X~hY0)}�U<y��Rp��e��zi���˗�sxZCh�[%�O��&ҕ�����!�*�(bk�au�B�9� X��U�d4��6C�/�ao�f}Z'�p7���������oF�����?�0���X�X'P7�2�t��=�G���0���ѽ���/.e�/"Ï��F����(q��\oIa9�[�`Y��
|�m\%��8'pߦt����Km�vB����~Q�w�3%���X��={G�7��!p�~,�vZkd����|��8)��ь$�)�g�ʹ�+�g�qėo�{�o���E�Ƃ�u:f�Xm&���H�x?��ᛔ������ڌvc��4���8ʗ�&�T��13�@�?��nVI�i �h�4ojký�/^<���O�|�͟�
uڎ���.��U��>�D���_�0ql�d]2��ZT�RO�J{=y�j͝�S��?�j{G-�{��e��k�`V;�p�!~8�t��|�7+�A��(�� *<�=�����ڢr��7�rx�X#�
��!��M\�u���쮻�^���v1������H�Ed##����SY ;��D��Jʽ�V�j�<��E	M�c�gZ%!��BF�����vZ�S(K��[e��m��~W�y @`j�t�f����C�����z��4ƞ��D��J�ۜ��J��?��g�'�����S���)�6��𦠻�?��$<(��kU�)�z*��d�;w����>L8/<�4'����䱾�]p�W����D�Icy}E��XE�=m_��;���/���8w�$]?������߯4�w'�%��P�S��L�F���%ƣ��U�МbC������B�/�l'�&~i�@��6+_��M�%;L%�l�E�z�B��o��,��B��W��d�2��bk?�f���aiZ44���=��´�t��%*�>�2���9�v�o3�.�}^�}YWt O}:($�A�{=���"�he
:��0����7B�0��*�cɋ�>{��e��0��mY�?K�����_Q� ���T����(�#Sd.]�o>g�fm����V�����J~fCh��n���ݶ���'-G�a���M1��~��'��0��$�)_�|V�e�l���8i���B��aʔ;X���c�}CW˟�Z�@������)�{��I��,Q�I��@x?��v�6t�}��(a�P��0�^U:x��z���딬W�������Zc��X)S3l�Jf)��p�z�`G	�D�+J�t�'�;�t�G� S6d����ӣ������y霫sp���dk�;y�ҥ3T�������6ڢ�ɉ)xq�"X�����`:�T���>zuz��B���
�׈�k��VJ��]�)nK�P)�I�@Ie	5�L�|��Z/��O����Z)2_��{ְ��`�������&��hrГǏZ$���O-&l�Z�x'#��]ǂ��G�н!���נ�y��[J�3\/����*f�Pe���V�纡ެ�8傯<�U���Q�&�Xְ��,ޣc����x9�^�	ڈ�;]W�u�ʚX�W�o�]�.jS��c[o����ےu?/�O�uxᜯ��Q-����k�\�	|����u�	�}�S�bM)׹�Sb���9�W�?6�����;]�G��)`; �7��2��7!v~����oUV���Sc��E�*E/G��4y���U9"��w�SGdˡOeB��
v�u����!�9�]�*�.n�K�Na�����y�l���o`,�?����nEY��|X�`���6����'�9������aܯ4��;<M�-��ij��Dܥ�q�S�Ή)�-�ַ����v@�����U�+�]:�H?��>M�q_>>O���?�GG�� oR��4�Op����U�nN4����8������z	�/��r��y����y�|�Ϸf���6Rv��8�t�W�^��{�z��Zɜ�K�`nTe�6k����q�q���u���<��\{�����Ö�nĞ�{���41�Y��?��iW&4dA1�@�r�R��_|�Zw6������}��w����0�)���l(��%�h(����mCd1S�X����U����3˫ن)^��s��f��'ܿ1=�e	.޾8C��{�E����K�U��є����Ϻb�˥E���c䫮O"�������3N����Gy1L}�fӶߡ<نfާ�^��2�l}H�L�{�ऌ���h#T�#v�"�A���ϖ9�l���LH\��Ke5T�b��)]C��;�x�.�~�V�3�Xy�Q=\����2M�����7)�?�X�*�����ʊ8�Ce9!X�ZWul�_$��*�z�]	�_kf�����͹�"e�_i�x����O�|��	�����kY<1S_ֆ=}8>~V���u����e1T����N͊�L��@dwN|�ѵ�P]��E� 	�	��
������4�W�Ȧ���"/���"�e���[+X��<��qt����}2K}�kr�&�|�g$�u@�7��QC~?���z�nf���ς}DQ�O�!��[K���_�r8�ḡ����:R�ZJ�v:�u�
��eV�?f�:���*?K�����#�������ɡL�/:l�8+0E��xg����)D�$�Ks�sW��4��լT��KN�Ts�������y�f���z�����O�%#�1��=x:N3�>�/��	�)��΄�pz��i��{��w�Ixm�1Ō�p�l�J+T�be��A<����È7�?�1<#��ů���k��-D��~��આ���W�zM�z��#�Q���f(�9��ve6Fb} �4��DGp�������SV��r�tc+�6��Md�'e��4���A��n&�ݧ���N�zZF�*�G�Ŝ��넚<���(֧���-\�X߽Ā��w�M&���{�f��i���.΄g>���n@��ӏ=Iˡ^���W���O@<���l��󤕧g�bb=Ztw?.J�	��5�c=�hq�I�4;����Z���#e!�w�v���m���R����U�O�+�����]2ܬ9��a�M�ƺ��n�캅��)�&W��	S]�0��D�������
ob��KYbD�"�l��b�ڨ��D ��şI��B���%�Y��m73�b�x��9b��0V��.�ڭ�q�:���?7���1d��w-H�m��)/̛b�B��0����ἝBs�z���9�3\�9$��(|_|O��o���`�+�]˺]��{3�c_��@m�5��r���Oh�>RF�#�2��X? Z��_�:=o�Re�|ŢY[|�O�`If����=V/C��3xe{G� ZJ������k��(}`&T)��T��qM�%(q07m��['|����A���yO�L	<���w��b�#���I��t��,uO����պzoZL�i��8uk����u: ���W �|u�0'��J!�� _��3�쾳u��L֮Mm?
б�K�d�6�dG;n��͒��I;�. M��83�J�E
,ƲpD	<�Pe����Z|uW\t���[=�,,��7�	�f�P�54bHq��&��<�Kx�YD��gY�����[$���_<21��h;K	OA�pV�����d���C E�j���f0�r��uŃgϮ0��P����L-��C�Ƣ��n~r/�
ꬾ(a3+?H�l[8_�`d�5�kB�o!�͇��L�+�z)_���IM�!+��}~RE�����aL���]E�Ȗ��QbV��+�p;lz\*6.B(Lc�%4�АI+�Б�ۧuFl̥�׌w�֐�j�"�5�r�~�:�ʰ`�4���~����g:�̧/J��Y9쾬\��]���h��E|w���~�f�0���� g���+�
ׇ�O��wH���W��u����~�T'��y�Ğ�JV������������7?S���}j��*�ͥ����[�aD�����"%J:A�����=��P�������H�I��,KP��W�?¶�Q0|۠`
��hǁ���l	����_n�����K���u����L�ț��r�i��~����JGd��];��]H�T�S�옺\�w肷��B�Tm�c--���0��˭t�n��s�ٰ��x񼭁�%\��(CB�0!lbR���LwR�.϶<g�Gl�!;
��I��%�@�ey�9�W���D�@�Q���6'���W����c�fU����������<�x�A/�($ Y�
0�d:
X�zg+�"�a$��
xc�W�k.����ٿ��[p�^I;�������J@�6'(�p����W�G3��^�k3�k�?�ʝǔ2J���W�e7���g�!���Vf��F�%ؖ� @�x��*��'�P�LjpR��0~���,sO[Y�]�W�{�fk�e]d����.�ai=�G{Q��(���u2d��ю�&��w]��5��`��w�d�.�f�EN;|���뚭l���g�j[-��~6���,����|�޴v���n`m0��A@��2`��k�m�j�E��7<�~�i���̭v7w��N�@W8����N�W����PV(S�+;SY�U0��аFݼyk�n�K�ŝ��^f���y�o�����k��w�����|��,�����4��%�Ϝ�)~���r3Ͱ���R��̶�Wd7
4�J^f1�p��x��<j����:\��\
��_1�^}W����򠍚�bk6÷���
g�4־PxiA�䫵ҢD�}�%���?ex[{������G2�w�~�|��W�S��I�4%�<���*����n��4Cl��p7�+P�)�?Ƚ�qx8�$�p�٘��zGU|����X~҂�z���VZ�)8طE�bH�pp1��UH���G�N�ՇR�[����W(�nE�
_�*GA+T��(��2�m��}�����@9��4��� C��y�&Bw+�|PwA�1R�ջ]�x�t���uq�vIKg��{'��۸=MB��G~�}��:�)���6�y�~ ����~��o�\�,��p��kC)���VGQ��4i���.x��~�vZ�I-(�ӱ��s������i����xc�4��#[��Ĺ��]�o/Y6t�6
&T1�-��a��̣�$&��B�h�)�yCa��m<�W#A1��L��E��?��k
���M9ԃs�UN�|��Y��g}�9�W�%��E�(��"��eW�YCXY�!�e��Ug�Y,JA@���);��^_`)y�a�>i9�7�g)7ÂVT[�Z��f��lQ��f�H8[��+xaE!��	�'�k��d��0l'�Of�I~>��L)IA��o�P�P�[Y�j�/�6&��y�=�8ƻz�Gi��F|����;\,�QS�@�8�ř}�7�Xt�]�c<�Raɒ�)J�:���rz�=+�3k���&!p��!Yå)�]u��PR����K=�u���HH�"��B�&�+��"� ��u�|�ۄ��ָ{��eR~lف���Q�ɫ�E��5�._M���0���B3�͔�]^|%-�B��L"�3��#����,��w�wS`ӽF�B6\����ͽ�x����"z�4���z)E��[{���|�kK�<	�f7S/�������F���[ �/����~��v��f�C���}U�xV�.�����y?I��r)������J��ꨭ������T~eG���X�0�nK_�3�_����&Y��m��OR����Yj(�{� ,`�%{S������v���j`}B��������AXr�w�>,11N�,��y���aZ���%���� �{���p�	�㴫���i9���j���U���xR�,<oU�k!�g�<��ԩi��5�3D����������h�u���A��W�e�K�����S�m���l�sf��Rn���u�g�k(�*��rJ=6N�x�(oj�o�ԓ��p��4�K��"!�/���\��d�	��8Z���\^%	���b^���ƥv�3U0qݹ�cI%�	�4���iC�1�(�3��+�����L�li!K��k5P5�\`�q*M�z[ۼ'ت�	\���
�1�]�C��]�v��-����<��:T�Jm1o+��)dA'��f�M���1�*T���1���Ճr/
L� S.��,nB�^�ꁧ��^O��pƧH�=�{ֺ�E�B#�m�q�\��D������u��[iH�]�V���ml��DO�,z[�4Lu��Ζ ���>v�z��L��-��kG�W��׹z�mC�b���g_Gf��H>$L�tf���I
�9��1���=�zSf ������c`쵚�Y1A�S�>l�X<��8�D#�����Z&@+Z^�7�ߧ�8���
�h��9�waz�W+���x0h��8�x&%�0�����A3�m���$�!��}ݹ{�}$YS^��=���k�e}i�U��$�n��f9ܳ674��E&�06ԉ�D[{YѮ��m�mI��"r�.���o���s�n�\���'CϪ 9.'�6�.ޥf2*1_�K)L��tኯˁ�}�m�c>9O�S�1�W�l�+��]3^��u�\�	+
����k
7�+�dfK*>b�SZݬՐ��P������V����e;,�$l�"�|���ײ��~Zud!XC�gR	�o��a6]?������఍S�ݢ�W�x�" 4�R�o�����\�֬�x}.��$��vV�/�Y��Q�H0{^~�<>�|���,m�o��xP]�D��[��X��g������ffF�֫:��Yk��R�XU����z"#����_�������/h��v�Wu�R��0cT+��3�ޱ�/��^J�X��rxv�┧���)��W��l_�0_.����k���G�>�S=����/7?=~�E���#��w��9_�d�ÌfC�H�Z�\�z�	!_�%���[��i|�U�:��q�Km���L���?�T����"'ѓ��N������<w���%E���	��Z�Gm�l�{��}�h��m���V�4��QO&8�C�2�l��]rr:{��s����+��Z_K���E�k�~#*FI�D��{*h���6��8%�q�3�x�0���:����H�
�1lfݏ�����g7{5�s��ʨ�T	���)�J� ��@���/�yr������~�\�ɞ�]�X֦��F0���RBz���P�I(d���}���h���E����*Ly�]Et��J���iZ��ޟ\�V�p�]���y�s��`���Sxw�V��G�Ѽܬ�y�}��l3ƁB&�W�����p���z=����W)�8�A	,��i���u/�	(�X��%8��!Ȉ�|�ܣ|�7��z����t���Ð�RS�#6s��)lx>�\�B�sт<D�=�34H��4D[g-�`�c�${�Q�S�Y���6֏��:D1E��ٮqr¦���^��>�GըЇ�Y�^6}���8cͤ��q�И<���u���cu����:� Z�Teq�x�w��J_���ۄ#K�g��tr�*�Wsz��$�8�=,x��r	)��x;��;���%�vD����_��]�������'��+fB$&���*���M<{ږBy#f9�	cD/;j�����^)8�;�`Ǚ�^��Ǐ��_�~��̼�㜥���w��g�P�_L�ڒ'���l�����J�$� �P������0�38��6���
�jdx��HV%q(d��gX.ED-<��k�ڛm�}k��Q�_�f�e|n����0ka����{��!=5j��U��|����G�)Ѕ��;�xo��	 ��Q���岁�?����,�\P�bYj�^uh�ٹ��}�N�F�+���ƕϬ.u{��	��l�L�������ʡ����|����v���\�v�K�/3 �n��f��:/�>��a�����kB��Ouu�]�^�0a��G�;k����|�62�>��P� \���smYɂl�
�`Klml�Х��*��2%�
�i�"�#�˓��-��S��4q�����ro���@�uz^e]ɏ�\=\�G�/��W�~��p����Wt��U�c�O��C84�\�Χ$�z^�]���ձ���E�/�LS'ɂ���a�kf$�d��S��Ʃ��>B����b&��g����_g��£Y��T$��.���^C���=�Mp���,���ϟC�ƚ��}0�Ί��Qw��7�f��je�	�<��x'%>�J��'�t�}��� � >����ޙ�5��Him����8�zA��Jd�?D�#d	ZL����}�v1��*���ښ���ć,o�i�(d!}�8�Cd�D��e��d���zl3�&x)a� J{���c�Ì8��g,H�;�Ѕ$��Ǆ���n������Oqܟ��9=Ds�箥���� ��~�DL���
ٯ7�u�|���.oW������ޭ|��SZקm��1���l�<�f2�;oC��)=��A�|�a��[`fƸ�/F5���>`BSh$���ϻ� ���j�ދ��˹��:]���S}�%0�/rM@\i��Yl<^d�]k�ԨjD�]גK�T�	�r�>.��X'�z��/J� %;����fp-�a��K�*���rl��0ʔ-O�����&]x{�����Ǳ�/������F^���b]Ѭ��6�
m@=��w1S�8>��(&��n֌�z�	��ȅ��쵠jm/�U+�O�o˓�F|�,k�^#G۵`j~s��AB�p���ݻ;���;�RB�$�d�9	.V7{ENϳ4ߥ�!����)7����8�mHm��{L���Ҭ��߲�5�Ca�q���&�t%�xG(�o��=M�|ym�Ň�L�5
����0��f<��������,a*�A{B�u���>.�x߼y}�W�����/��6R0�7=��?�\���bR�W:|Vٔ@@���>���.�N�h:���a8�n�HV�G�$V/	@�g�y�UVIJ�G��o��!�iǒv��m?k-���ͯ7���ެ6�
��֋4��^oj�g��߼y�R�n��/��w�5��*�z$X?d�Bs7���Q��2��	�axfe0t�����㧯�e�V�my�f�E����ﺥ���\�p�^^�5u��Q���HE��_�1$t3�>	�z�ϺV�E+�tխs��/���N��-�(��D	�)��װ}iV��d��,\����Ney��.Ǳ��_���S�xg(.�C��-W[=��s �����g�����Sjj��X��(��6������w�w�a�%����l�u���(��X���=E帵Y�,|�מ�M�%��S�2iCSй���[;!W�U<��+�����aCuݷ���R��+.YW8�6v!���LHLL�#2JUkm`�
�=;���[e���6{�Y�R�.\(�2�¬7Bfp��?�@�]�'%��Uc�m���o��0�:h���F�Zz ��I½F����-~�c
��W���,�j�	!�JNoIȾk2cK��Ͷ01��r/�o�D�t��	��i�����wE���HK�(�m��n�]V�	����Z��!�]�Q��K�MЁ`���ݥ��[�d�Xy���k�"���R�b��ׇ����Q����o(&���0��0�U�v�	��F�G���
�}�c}s%,l�|)���+)�5����j����̴���[��R�#gb�S��d*gŞ*�qĈ:���-K%73XùT��:�� �QRj]�J�����1�z%�sSCܖ�4��ڜ�T�JY�@��T9ϚSؕP�^f0F�`�����f���i2�i��✇����au���,%a�^t[zh\�*��Ao���U�:}�ZX ?��~���6q~5��/�cI�'5+sm�#�ؽS���[q�!+��7n�W�U��1\J�}E8f�X;��x��L���i����Y�1C��&���������T����,n�#V���J�e�ȫ���z��Zg�0zy�J����ȧ�8�&\F!(��Rh��sz�vґG�A�.�`�l�Q
Y8�4]jI��)����᫯�la֛#D	pul��0�����З2R��e�"���}g'Y���Dp]	��:�gh�>.'��� @���h���
����F
��buhz$�]qZ3+�|'k�W_}��*��N�@Q2\y^5Q�y�W�	��wP�3�C�r��C�i\���H��`h׬>��X����whGq�qY���-��7_�c��6�<�
�>z�G���m��Z|gxO������������0
~�FƉ���m�w'����ދ�?./��E�Y��%�e���M!��a=���+�l�S�rW�ȇ���2v����vF`�$�
n�����j�
Ƥa����{�g5�4ڿ�B�8tג/�+��Y�)�nR��jT�=����Y��s�������%��e.<�|��|AM��=+}\�R*)�'��6�����u���]s�����Ӆ�@!$;�Ử���Ë��F�V��tL��ҋ��W����|�m�-�C�vOր#�_��:cB���~vuW��C���m��FpS�j���� b��Y0���@u�!����V
L�=��^a5����j�슑�s�A�k��?=�{V/=T@UP6:|#�Ӵ��<�@!\?��.� Ƙ�ۮ=�_��A����#�b�Д�b�Ґz6�2����S�f8h`
]c1Z�2e�ڡ(��y^?��E���\1��,�Ϗ���p��4�Ҝ�^�r_�� ��X\w�vq�\�]�w#���w>{\iz�Al{%}ջ6�q�r�1�E�G�<�q��Me���3W._�X5�s����":ӳ%t�=�dpn�2$�9' _�p�Ɍ`���E/�ڵ�s�~������Q�IMe/!t����ǘ�^��M>=q��qB�$�cV�V�1��)7�������
{�JB�a$fsÙ{ьu��i��P�!���y��TG����W"g�6��n�D(oCW��i�h~/�cS���X���F�ebΧ�]�rg��PeFT�h� �j:"��,�C�	�xL��S���������v#���~_�Ja�j﷿�]on�I��-׮�����5��B`VVR��E�o6x���Q�P��ן��jh�c�G�V3��^Ĉ��<a�/�f&�l]�P7��%��@f��N�b����ל��Z?�@~U���ݏvS�"�a������)f���S��KOh�7��^��2����e��w��fە�tRS����a�p�~��Ejs~6�;��r0i�����ٓ')}�����J&X��u�aՐR��}yws�΅��XY,�i�p�(� %�7��|��& ��M�`�{W��a�^)n�*�����A^M1fU�$k��r����o����͟6?=|��4�Z<7_�3������Ғ��h}̺�!_���<,b{���+<�3�խ�S�gȧ<�����gh��V���������>��������o�T��<On�X�C�!���d�&��^�c,f�S�x~}���X	�ä<=kǔ'��{քҁ�l�@�:G���
.1������3r*�cֿIE29�9r�4(�-��,���JV}%��x}j�J��i����mv6������V�X�"_|���B�S��2��� �X��^+K�(4I�֝kc$����7)^������͏�ؔ����ˬ��?&�O/�:)c�S�(`$��J>hh�����-hU���E�:G:�U�����B�831��&È?�	�:C��3�����I\8��L�?j__��	Iy��k#w�9�Nl�����5�Ȅ��j2��]!�����6�Rqа�IL��i�tT�z3�>fczM,��e��p��
�SM���\g��)m��m��*�0r:���Y>QkՐ��%�0����vm�K��{ç�#B9��ٙg�[ƨL0��:)ag����G� T�`��Ғ�?كw�Iǔ�����g�ZC݅��O?*x�&��R��ʿ����8�I�t"�{�h�:N���ݷ]	&��a�U@�|1�Jn=O��,AW/�Fr�_���|���"��	��	��5���ZC����+a�`3\�K�� 
? ��Õ��:-#�:s��I@w��P����X��	�����T��?ւg�G�a��5��� G��]P��Ԙ��!V������.2MC`����#�T�#�^�!ߡ�ĺ�YK�ʑx����_�)�/�5eM �ɤ�w�6zs|�P���E��]�I�bB�*�i>33*�;��gx�r���S�c�?�t�ꅆ��6>�pPu� �����/����cF�&��� �JE+�"�ݤ�^Q^���䰞8e���sL�I�c�Zluc,nwn��X>$z�|�(x]�J�G�K
�b�����������p��Ø��,�߷x�?=�<J���`�{��٘��&#=|xs��s����͜�������:O�ۊ�zS�����-�[8�{J׬�U�sZ�԰$(�:��#S�Y���|���~~u����]�jNCoY���Z����7G�6fd�l�Ge����Z�E����_����1<h�p����㼫 ,�KiW�����v�@���	Fk�}�����כ���a��)/�^mb �«設m�,��M��?���%t�,wP���EJ���*��
c��6�pJ�̌@ȫ=�2�JJ�ƈ�k�������}j�+��F9HZ��o��������"������ov
5<��	3Ei)~�Z9�t�q�y�c���Ք�Box�Æ����脯N�3�El&4�����7�����q�eZ�ah�u�?嫏)��_o�?|V�6]�;��km�v���ѹ��(ֲV.�)eR�C��a��)��BYȬsY�-m�C�����7����]��)M�`�$���^�C��D��F�j�Ѵ:_��E_�2�Ǒ"f�Va~��O;��X�G��d�kYu�*W��X��Z<�w�E��v0�{�ąm�o)��e�������u/^r�!�{_|1���7��/��o�,ڧ�S���c��G1�s�}�{�rfd�'�]�YP���H&���SD��+A<g�h�N[�(�`����,*���=�R�
��>�	���1����AT  @ IDAT<k�d·mb�X���/-f�C����Iw>�й�p��>TF��!�T��^e \t�{)L=���׵Z�����f��v�N��p�c�,^��f���q��x� �`�4��R���0n�eᆁx����z�7}��+�ީ!��Ͳ"�߽~�yؐó��в��ݼ�פaXWƔ�K1�	]J5�ߐؘ�%� �Z��^��Ow��J���^54=a��|b4�tf��	��[E�b��p��v��X�X1���#>m�p�10�TL����63�\i�mm��0V
���f���3�@�h��
���F��,N���{�� ��`��g��R�N9�SY'Ts�.��u0(?����?~���(`����׿�����fV�=C�W�𬏥T~���YUư���z�?4��fC��ɟ��RE�M�꿺���Z���^��wY�&�� ~)4�Y�{�v.+A������O����?����ZZߏv=+�o���6�m��/fؓ�1�8�	.</ڀ=4�ѪG�!�A\W�1��'͌d���w�G	3S�Q4Υt���_׹����<���2fڻ�"���䥔����(�3ms����t�.�E�?\��P����Ĳ�c�I����?~�����0rV��,|��_�W7��_;��0|<�C���;JP�6��)ozܲt���WH��3\���e��9�L�[	y+�ğ�]��7��u����כ�������nVh�u5c��tXn}�~s��6{)��o���fG?�.�Vlu�^� &���F	c/F̠YmO�)��l,L�ȩŅ笞ܶE��o	��3l�+Es�Ko����G��b�@C��@�� ��I�w:�^�
~b.��Rk�g	�S�#Q�)�e�z�~�6�~҂�ϲ�ܺ�B��(���hw9�,�˂H�z�"��~���,��[m[���R�4�/���h��כ�����yn���(�蟓�aM�Ҳ��͉>�}h�j�_	W�:z)K�|-�������OS����)��Ik̭��N�p|��E;o��\�>��u$<R�0a��;�q����ͭvm���t���+�)t�R��X�ԟ΅�i{]��OXʖ�U�S��ߎ?�g}�C�W�ы������on��ӖOj������pw��o���&�|8y>2�{JN�!a#���Į�zӌ?��^=��KJ�XÈ╸}5Hҝ�NET)u�k����#�O�
X���1��f!����SOqkL`Za�0�\���b��}���(���F�Y�TX��9�I�.Ѵ��g�@S�����E��p�&��SX�kt��@��x]E�~��`ʛ��UC���̈́��qq���[���6G��x�m_��~E��t����6w+z�S���D�|Xl�c����~뙌�)µ��̼���}ڍa0�jo��Mí�����d�	�������lim�[p��zRE��Oco�m��Y����c��X�)*a��:e��0��As~��ת�'�����o.à�o9$$t,��GiI��E]��v��n��������N��M��u��ȑ��Kļx�y�-���[�PǢ�����P�(o6��:�	�h��5X>�|	>�[��a�c}�rs�۟�fx���Z�az��{tP�j�f~���M�xU#��������c1��YL~���u���3�z�2s�b��R�(�K�%��?�C]1Q%Q��: R4)���f�[�F{o ?�����m��3R�X�=Ⱥ`}1t(n&�FX4����Z��̃G�gH�N��Wc���(�9��a�K|�]CS��ۀ4�e��y[�|C)lf�m�tTo���Zk�|e�l��X���3\���������4��Ѣ!�k�^M��ng6o<�b�d�����Nu8ʗJ�-�ǈBt�I���O��h��G�f�.TZ��Q�XPl�^��	n��yR>{:T6p�i֙f�BC��*/BԽN���V���&�+3��)A�}��E�%�z_��@�V��*��~<a���|ލ�W�JE���|B�q���nf��0Ьp�Ef�K�J��@Z������_t�������D	���O�}�`�C���Yg�r�E�6K��x�"��l��o�xɃ�,�� �yf���PsK�����Y�ds6��zL�B/�CZx����f��zY}����*�Om�Z��JX�z�2�|��&-���/g�+Yn�5$�#H���C�W����M���i�7
X �������>�iYlw����8n���p��-T�hD��?�0+�Q6eg�:�Pg,�����\a(h&޼~+�v�r��6 ��1��D����[�����]��#�/gm����0<@��H�nL׎*Чן�����-?�Ri,_�n�+�=�eR�D8&PQ��!�&a/Fluq��=��c���?x��y��7A�>i��^cp�j���SQo���X�y�Qe(��P��������E�U���Gt��ٽ[����=�U���'ֳ���	�e���$Q���=~J��o;����,���rf?�b�Yc̊�;�/�>R�"DV����k�f|b�iS��:�����;�b[�m9P�u�鉤`�>�c&}�K$3�]��e����>ƥ��<�΍[9�$��?��z��C����7{�)��c{��� �tf"aj���{�}��B2�u��Nzя�+�]� �]8��H��� ��Ճ�֖E�>��Bx�������5�^?�G(��jx�3������X7��s=�6ȣ��߽���4�ėa�(1�㔵�/RJ�G��Mf�,�kճ^'�������x��b5(m�#��S����(T�f�2��Ũ��̓���?n���?�Qz5L�8������8�!_�ӳF����d4�҇SD=|"f�7��I��I=�G)�O_6+�Uտ�1�K�:vS��e�p��[^����u��nfKZ�� ���������Y��n�Xc�R
��\Bo�4�	u�%){?�ۥ�����:�B�����IV��y|����x��`���4A ��M��ϥ�m���t�m��c�5/�oZ��2����zux���%��%`/���1�Z6@��x���?tr��胆�^5��Y6Y�f����Oi�¥���г�[�5>�zU��c�O!@ˌ2��E��^ '&3�L�*�iO芋\V\�W��څ=$�~:��P��q4�X�a��VB]gj �m���f�<��Fy�QeS�Q��p�������-ؤk�U�`}W�ݠ�p��y����T�z���U�����S��yKj<�|���,�W����tCw��CK�|����OG{�"���x���x����c� ��꘽i��O����`\j��{Y���Y��D�h�Z���	���o:��$��,x6�&K��~���˜�E�G���Uu婍�3�v�������+>���?l�������_��:��Ҏ�K��,gk�?㉃25
�Il:�]w���A;B�kJωc�J��|f|�J���(.��U=.��Չ��XT+X���#���:�����I3�˾��f�V8�Wi荏��K7j�wǼ;S��#�S�P03���P�f�P������n�BM�H�ba*�ߏ"�]jcM�T{��W�k���WC�3k��[V4~wﴵ��k)
��x�j�O�!?�U�E��L3�#kI�8滅�����_5wn���-�z=ǎ,=�}� �o{�4�q|�v�|~���]����b���"z.�{�wɬ|>=͗)�w!���g'頰p9�������}�?e�b���`x��bކ#�V�-��p�t���Y��,�����`ޖeW�]	�u?�تwF�3�2��ݲ��f�L�[�����������9+KX��M`W����{��:z���N����k�֧��`�v9=v���I9xV/�~N�?�ix�����O0Cy���1���q2��p��$0��O�0+�γѶ��~�FD�@ue�[S騥�5tp|�<��&ң|�^�R�Z�����/�gZa�~ç�I،�!{8)��5�``��_g��TY��q���m�'����`>�<V��m,�V��wZ�L
uU)C���)O0������~���~�,^[��Y
�+4b���Y��|3gM���YX�+����h���ċ�6����\�z|�^�T^m�r67.������K��8��~�5��_%l	�7!�63(S�Y�!��a��ꃈf�TO:	cIq1Z��|(<%���G��6O�/�7�:|���yʔ��f���p�T�x/: ����Qՙ}���,4V�ױ"'�F�r�hج����8�봰����J��E�N�|��E#�51��������wn��gm�Nf�N�9��y�M�ӟ�mQ�+/��B,$�::��&�� W=W�p�:����*�S]�5��*A�V��YOڥx�FNVn�$0yJFD�rT���jG���<�t��b@���"G�g��.d�[��Ŝ��O����3���48��i+)�cݧpt�Q�+�i3�%���&�$�R�S���^�x���Mz@����N[� OAwx�,����~|����?T��+������k`
4�_p��L�~��K��7���7��b�/��7��E3������C`��!�q�ul[smksh�|g���zF<��uů�m`O������y�g:��Uqt�-�����u�M��FC� ����x��_�Ͽ�p|*������v���C�b?���׭��Y��Lj-�`�[XHUB���~����Q�ʳ�YD?��k�I�z,0F�0��X�zOc���@�^>��-)0f��l`(�e	��I`\�|�����l�7�4��?}Sɑ�(�Z�_����9![�F�崯�kl��$ ���g���pR�yP�D����������Xa�z�۷�l�³���bl���Y�}J��O��'@W���6�y�}y޶�U݊3^[�4��Эa��f@�l��aƯH��_�b��Q|j���c�^�T�|V��0eF���� ;8�2%��_z�D��}�5a,�K�ܮf�&��%����l����	f �f�MaT�W1��z�	˽f�+\���	�e������~�=b2�SV�-G@N�~��·rR�,�`/;B���ML���ݳ/��%!? �D����q�3*N2xu�e1�|R�X�ݖ>eY�q���$��Ջa%�k
�U�u�p�,F{{?���A�Y�o�:ţe��Bk>���kY+��h��/���^Š���6kR6/���e5��Fg���g����� ��V�A�-�ɱ� �|?��M���r��Rv�Î����oR���2���h������x~L{?�@-�x6�1R(L����xN�R���u���˕�uW��}�g<6�wz�W���i�$++����a5��ي�����Y��1��T�*t׳�\A�3	��՗Y��E/�+���}�VF���LkyQ�o�m�d�~YGٌ�cCNM,�x!^/^o�U��f~>�|��C�ޱ�ĵ|U�/�<���T����,��Ä�aFB��冇�����Ti�/��������M�Ҏ
�ݫ3�8jŘ�f���K}YJ���/6���򏳨������,Yw�5�J���W�iG�l�������~?�v�I��Ű)9�2���sC�*���\S��>���Sd�,d���k?�?�Fյ�rT�����u�o��o鎜�vKޥ ������\�����[���)��������k��:�i�C���LP�ǖ=H�ئ~&�4����m,�N�x���c/J�a����������f�6C�/�a�e��pOV�i��a�$V�׵�)�/j�,p�	o����:ώ�+��a�_'�+��t��/��|�o���a���|]^+�f#�M��0�a�v����F�|�t�k_.��k�:ǃt0���92SVψ[�ĤS��l�>��h�4�a��p�X��T3�1|�e���R6�`ֆ�tr7K��_|m�w
ع�_��tєC-�0�Y��������"���E�q0]�6�W�Q�z��#��O}�n	��G��v�1O���PȾ-�P����1�
;��a���]��XlaV[��r#�Ӿz��h�כB�!�tn:���4j�iɍ��0�w��k�˺V�V���C����?�Q���uTL���]�u]��ٻ��n��z��+�>�1DНǕF��o��
'��8x����,SҀ?�z?��o(C��w:���s��Q��x�������d F���d�g5��<AS>hc2��=�w^�/�N)eb���<����X�w��v2������s	�s����½����<Y��w����o�I����`𯙙�@'�';5|L�z�Af�<=o==${�.���]&�/L톐�+{
��fq��>����<�f[3/��sEYe-8QṘ	S����N����|1����m�`�򇶳�嚹ܵ|ǔ>�%Z�̪��pұ�!�4�C4>g�3���:����?Z��������tŔ�
3�����~��Κ�qnݯgx9��R�`��x�)Z�����qz��C���/���<��̄ Z�β8,HN8}�VI�>�:�*G-}r#k_����2%�l��~��Rɢ53Q��lC����SXq~Lx��f�r��'�z��+	=F�C��[���T���=�n���=% ���L~�-~H�[Knf�Cⱺ@f������s�s��1�|~g��uqr~���͓h'V�����"kⳬ`,���n���,Z:��.K��E�uPrװ��e��6���$2ҋ���\V���-�r���zy-�m�Lty.�Td�+aJ�X��>����0�߶V�D�������a#+\������	��o~H���đG�->^�z�E틀�h�b�f�����%�Ļp�dYm/T�\d�G5&Xq��;����r��	D�,�Գ��X�)*۬�Q��ID�v�$�����Y�'Ͻ(���{��0�dk�,,B��<ʉ>�&�p����Y��ߘNY�|�@A4V��&����:�g��}���~�Ƈ0���p�r���O���jmx�Jf�ϐm�"31P<Y��ɒ�&._��|y��o�������φ�|h�7���W��Wǁ����Q^/��Z�Dy�Q4�-�p�-Y=C�=�g
\>'������������n=�_2n�͡��V�^��ϩZ��?謰H�_f���3�[]����¥֩���ۿy�����/"0%�*R!�<k�p8���N�S�Q���:�5(`w��H�p~:��{1+5#� �&�U��i��h=���W�C�'P���l�W���i�,��Hq"n�����4�sws�k�\�ح��m���_6��y}|Xx�z�Ґy�tj�12c�|yfy �7���B9��_}����P�<���]*��oWV���^]fI�	1�&�.;,��巋�n�"9�a�b�ۊ�P���ճp����>���,M�Q@'�,������֛��Eʴ�E�uq`Ä�\��{�̰co���k��	m�
ޙi�я*�!e3~�d�H��(�A���RB���r��`+,���Y&����0�K��cci��(�A8tկ��/$4f����),/%=
X���ef)"FKe�ad�Ae��0���a��֐�:�����bf����^n��V���o�vs�L�FZ��N��j/�������^��2���^e��o|ߋ1��d8u��W��kdʒ�蓄���7�?|�}��pAxW&����0�Y�h���W٬	�%C��s-�p=PnרϦDXQ�r���Ļ�V7�ߥ�F���0�nON�bƖ���6�G���X�5�F����3��U��2�=�ʿ({D�8��0
O���'k��'��G�'dI}��ʛ�6V��F�g)�?5$6��<|*aA`�
F����G	;�P��Y�O0�#"k�۽
֥wш���sq�_[��G+�=cmH	:��lt��iGG	�)�_�Q������zs԰b~b�ԜcݡuD�_p#za���b)���!�%,�q�/q�K��vtr)����ϯ��~��:�ў�Y��ǃ��G�@[{߯�,!s�:y>����ϛ�����j�%wh*��^Ёu��4dG���UN8�L�q@�|WYM)y��=���Ҫ\X�� 婊E|Xu0,�r.i�����[��U�X�����-zʱtʯd�3\5tnag�fg��P���;��6�!���������l�\<��n�S��cw��ƒ�$
Ua��E���lx�N�Y���>�����_l�n�B�ʓd ��=|?܃��W�ze�c�Y���Q�NJ�+�N���X�2�7c�������
_����*��]o�=k��K���/��~�U��v��b��t���*l�P�������A�5;[�&®��!>f�ȌTg�R���Xy��@�u���'�M�0I��o_Yk�]j+���.g�P��򵛝�������ْ��S��IBc�	y*q�DL�n)9�
	�r)"
�F3�S-�9?�Fe�W
!J	$���9���Ө��'��c�1D��}��b�?W�5T���4����ې�f�5��w����N1.��p�ey�{��nj��M�4C�LVB3Ѥ�s��z��N� RZ��.��	���O�@�v�\q&޼��.v�[H>]��>mӞ���Mj��O�
���N��m#M���F��s��- >�D�x�c�Ҿ_zi�kp�I�b��d��*㮜�u�;�ա��WH/v��U�B���ߣ��$����Q)�,� ���P%�\�ɣFRoR�������Uf=Y^�#�a僔����>�ˮq�-��)�����7/�9L#'h8z��G�!��:cE�T�ee���,��5H�lu����Ka��嗭�t��r80N����Dﴶdhk�Q* \(�^�O�zR}��
^wۃ��'�"D�yC�6,�I���"~'�E;�r�S�)~x��4V��ӌ����s1��_�~+�M8�r�n��j�>^�p���Qu�1����u�Ѝ!C��B=�����$�D�}W~�h��
����+�oue�,Y��|�ΕA�,�Z����n�8�5�����S� r�[��`�Z�(�������qJ�U�J�S�uH�R���3�6 ھ$�f�����ůC�5Y��HB־��6Sj��a1�m�~	��׃�Ged���G�����`>_�5��b�@*,�t��%��?�zU0�x~��LK���$��PY�g��;}��@��2�� W�~�w���	����)�������me�� .�oc]���ৄ��:,�����+��pЭ�Ԃ�k�L����
�Ǌ�����ژ�����^��f��{闆ʮ���r)���Z[��6��)|������"��Ŏk���W~R�z���a��n��N�N=�DR&�Fǫ�7�Z��V���Z�W�HyZl���t��������Ӓ��"N�%n�7�ï�����.��J��z���ҝ[76��՗��������"�)�%[�ٰ�����'WZ��Z��7[T�V�XG�"�:��q숗R9N��ɺ��aѝ2��D�
K9��� ���ǞɵJ^�1�=�o#��&�8=���u�N�5�1^m�KC����x��A�*�xT��s~3���oR�4AJ'Y�E�a0�Y�z4̳3�0�v*���cW*`�V�P�)t7��zBa���C�6	�����Dc�[��0lh�&3��=�U���q��9aG����)L�ѣ<����4������f#����l���W�
?�C����k �'՚�0P&�ٗ��Ma��m���ű�U��>?��g�Z��u�e�y*̖HHD� �xú]�y�^�>	��~A�^�#�Փ?�yʲ�
~��X��)�N4���E�!��P��pB�I��-4zs(Ji�0Т�u��U�{�l��xb:���,�;̾ag���� (o�%����o��aC�<�,3�603~�ɭ�(^5���h�k��5�Q)����%*FL��'��ԉw5��֒���}]8���/k]��0��B#{�7I#�Q�yk`������=+\��}H�a�Bde�k[8Ð:4��0�~��&10V�Sd˿�"��9��K���F�4�p�&�C�j���VP�0���.�x)P�m�ײ�]��^�Y��M8����uȧ�t���I�e"�e�Z0I͜5��_����/sJ�(!�0��0S�\�3^ºͺk\{�ڀQ�.�$����l�YT=����`�b=W���fKa	�A&LX*�,[��b����r�����}���E3���1��LB���*qBЫ/0j_��p&��S>����$V���I4�#;�S��GAs	����C�!��"=��q1��*.m�:	�F��9<)�����ׅ=�9�R�"��-�+e�6z>E-z��h�5�.���L3rϵOe��o�B����0������Űri':(��V��������V�o6�\$�*^G�1;�/��;E��ګ�`T������Sm�Z[������R�;Y&�vֽ_��7c53X�g�.�Y��n�-�*�SU���}�wu�I8�pa�V�S�W��jѡ�F^F�c�N�+Ԭ�YB��%�"���7�jYJ�t%�YX�|��N]�K�����#~���|�`U�¼�>���C]m���	�q�O2,�B�Ϩq����f��ۿ����|'o��͢M����w�ݬ�ݸu/����F��%�S�f�ӻ�6��}�RV��U`��"��E���F=a��BVu���p������ �i;��F�`�ֵ�-Kc&p����	Xso���ex�A�wJ�p$-p���l�^�BY�Y���h��[�kէ���1�n+��Fh�pJW����)����>�kb:��z���9(���$����L��77B��0O���͊P�V)g�6.����TF�^�2��u���*�i�!��?<�'�M����o�+�6�	�G�X��@B"|�[�s	�A�ѝ�P1��
�=i���;�/@��CYד����PC ��L�M���&�琚�+~����6u�-L}Y��qG	�1��r�>�1OKu��������J@�a�P.i��"M����T�)��)G߼7�-��C��,e<�'l��Ǘ��iR�n��
�.��Aa�u��%yW"ʺz��}���M��wD��,�`��i5Q�C5�-M���0�`?�w���|h�w&���=��4v4kޙࡰP"�7PF#�q�x���@�UZ̲t�A����ù,��W�j�4*�ԕ�buO@cg7B���Ga�7\j/,s~�"�cB��b�3���琞��W�_�f�j�~/G�%$ϵT�A0Q�������Q�H?
�K�(�R�	Jt���|�%X��pѝ%��s�N�(�w�0C$�a�G�s�$���C�@CGʭ`%<B	��UؖQ��W��3S�)��5Zq(;�V쁨�uL�ũV�>���M	��?����Z�]&ꬭ��D��7��ɹج/�A��T>)�#lJh	� ��}+,aA	����h_v�;[e�m�Ug,)�%I}8��m��C�� �)YC�f�4�~������3�NEf��p6%� �2tg���,Ъ�I?�R����?9@�a)\(\�6Zu	�� �=ic�S�cV��%uJ�X�_>�<m��g���yX��߽=��k\*d�1�򜌷Y��(�"��Wg���j��Ҙ���{a��W:��S��Mk�iaV����ee��g��(��\�U���gʠ����@���Kr��a�FaBa�J_%�)˲���u.�	7�]��uo��_|��$Z�il���
Oa���\m�w�k�r�_�V��Gee,yy��-�M�p�/�v�h�Ӕ|��mDO��ru�l��r��&��7|�#G�+�� �q��34��K�nב���g�L#"�B� oK����Mf_J�L��@�w���	��E$���*$>[���"|�\���V�V�ш�\cx�9&��$���h1?C�n��M���Ů�4�;er�`�SYvb6i���w�%�L�&�uDt!l98���1�̜��f+���έ����_�;�nsx�I���bU��zp�nJ*S;��!_EL�o��d�C�`N��8-S�p�9� S�0�B-� �bu`��)���窥��P���a��|��zrLϿx�0ԸkI������E�@�UA~��J)��#�<� p���0po�Sdu'��~Y$��X*{)�EH�$��Uq�qj��^)�a��%�}7a4g�jzq��8d�~��B'u�1��S�H���й��G�1)3h�.$8���K܊���I����7(��4lq6�a��I�|S[h�����
��U >���]�#�FP��|1�`$"����8�2��H+mRWa��t�b�J�/K �7�-g������E���0Z���I��mh�ަ~��w���:� �Ӱ߽����U?U[I-��k0��(%��U����(��.\{�X{&;�+m�$�U�hO|�p�������?�ci��")nغ�y�7OU݋�3�����ԩ��U"j��&�9��������u���(o� `[e�q�Xz�!mbl��4���$s`����^��Ǭ`����v3�7ڼ�d䂗���o�b�k&�q��Njt�;~�ż�Ǒ�g��d���$,y�s�s����}mo�<Č�k����8J���Y}Ħ}'�/��}V�������Y>Uå�6�������3��3hz茧�a�+嵽%��]	a�A�����:���`�YČ�,:c_�u�|�"˷_��R��\;xU�����w�����_|�S������ӕ'/��f?��Yq��=�P#N�k[8gp��y��(�ҿ�^��k��a�g���:ެ�p\������}o�y��X�����w��c[J�>��!S�\��|a�v�mwyi49�G| h)��{ë(.����e�+tn���jѯ���u��?�I�s~������9�۸����Yg����,��Q�2��\���e1}�}�O�[|�
��_Yp�����?iS���[�e��7ob��7�y�Δ^מ�ʕ�Ѭ @����/��8����ܜV���G�8o�!���J�4���J�k��j��y� �8J&>e�(h�BP�@�ՠNFN61e���¡{�m����?�g�f5��|ʯ��(}t�/J'�J�Hp��)SΗ�4|��w������8�}��+�+���G�F�X������{�C��M�|��3?��py'��x�಼��0�F;VM5Q�Fir{e�jX�`p�n4{�X:�Ɯ��~���A���q,�������]�CDy&xY�!(r��1��"�i@�:3���3�����\�y���������c�&�L$6���0^���$�P�2.V�N���C[��lJҴb&���O���\�5,cK�E?m��P�6՟�Zc�T�A�C�۠+8Q�˷6{�ɣtt�#r.���$u�s�c9���:4ӂ��	X+��㍃c����n���	\�P�m��MAՓǇ>��������5�x�v���f���L�i~���toqz|E���æ��`;���'m�B��k�.6t�J�P':���K�&��'��ۋv����Q�v!:��s�ϕ�m�:�_�ˉ���D崅�l��?:9
�1�$�����{ToZa��01/��N�y��W�[�����Om�j�S�j!Jl�-������\E%"]��C&x���1�� �,�Y@N�:Y#���r!�x��|��5�u��8E�`'����H�6Ei�?dr�VF+S�'�9'Q��Oo� �L�MWbg/P��!�^�{�r�_�g�����^_���'��u���D;�U�}�[��x�8�mr����|�\'�cύ��F���U�6�@>Ϧ�'�����C^��9��c�5� ��b--}�_���;��pG��/�)}+G������	xy�
�
�M>{�2��d��Hi�I�I;)�r��Rg�1�ʸ����ż��r���L�mu�p^�#�����.���'7�����ʾ��W�z�e��6�C~�� iۍ2��܄�w��y����_��c~��9�*��Bo�W�*�O��������	ߥ|�}>{�彩G�%^�KAp��hd�t����$�+I?��f���g���l+f\A$���u�G�d�C�.����=V��֥����x
�$��6�7�5���,F���b�]�fc��Ug&�4Щ�!���+KxN����8:�E�8p�޻�����G������Kx<C�����	$�����g�*�G�\tP>{XbVV	��b�!��5=��$wn��xE#���U_�7�z��%�_�������s��?������{T<z�I�/��B��tt���Մ��~f@D-wp�����0r���Ϫu&9�ڀ�_�I�v�`�O�)w�{�HI�с���<�$K�a�nd����Q�t4σ#e&LkN�?�ʁ����+.����� Ce.
��5;��N����H��[ ꨏ�D��r�HA��GtЄ
�2�6�:�f"�������d|$M�Ε*+`!�l�ji.�����]��l.%N�\(쟴����$�,�;�����ӣ ���㧙0)�!�5�`�VsF�L��Kg��+ҕ�MK}9��{���>�r%��i��ŪL� �bc�A:�9Y�K@ e�/Æ��������ᅍ�'�47^,R�+��r����eE�v�&�u�c�ހ����%�$!�>�*�G����F{�ש�f|��b1��{AI7Ў8�N�u��r�Y@5�r�h:���Ύ*j;XW�:�j7��Ki3�S/��+�Z���OR����jc�mmV�P�ʑ0ag*�aO.��nyDTR�L{��9�̠.L�u?���w7�Y��D6G�h��&�	�_:�8�B4}�9��%����Ue��xCo����<b�D�[l� ^�8I�v��Z��RW���CV��O�ʕ	Pm;��*f�~+���W���Gl��������3_HMo&_G0�Jٟ"r�/bS�vV?�zxz���`Q��ɷ=���/����~��:_��kb|'�?���qu��MP�O�&{���>�I�Z�Ț~� Z!�׵��p�Ε���r���A����y2��?����k�+V7�6���_��/��ww}z%��\��;��I��rC�+�W�ydH0����p@���C!�֦�@�_T�?,6(��*���	oF�l���G��3|��:���y�FV{G���.�W��r��h�8Q���g��/�V��'���c9�g�m>4��N
I"�g�A%���7���%��э�������K�)}���[�`.��P�Ci$GFx�2=r�b�竗�'p�w���덣 r9�aT�|[���k?�;>�K2�d���#3�YFU��J��7{��C�� ;�� �P����N�Àa���#�A���JM��!O.��t )&����_2��JS�:�m{��*.w:`��kW�8�7�hP�$��Ƹ�m�� ���ݾaEfİ̀G+��6hemal�cPIi|ʗmP��n?	�BƄ���(��)��
���&��#�rC443IS։HGG]��0��%�L"Z�`���+V5G��
0!s�`�������zǁ�a�k69�"'L�� ��	��y�Z�τC��߅A�U4(]�#����~@.lrĨ9���c��Cyڰ:���F^��W��;�X�e§Qo��KHlA:ڪ(�2Z(pd(˾\�����]�gBں��A�\�XIo��+�쏗��uKF�ޅ� ���z-WFm�0���Ȕ��.Y��\�ȡ,�l�OyT^����E���b�y v�Q�8�N�G|�������x�s�,���'!^�`�A^��ړ����K_I���n��P�Wis�.7�l��5i��Jl�ŅfnH�P1�c׹�?��:7!+<}�7J�8�Ӥ�l��ݕ�ƫ�xq�6qߺҏ�>z�54� \�z��:d��M[n�.����l8�&���t^�*cmݴ�H�Nd��/r�����O  @ IDAT�p�x�'�C�ݲ'��~�g����s��E_�z�/#e�E��>�]R�~�JV[�O˺=AKZ��cu����io�cV�#����>���oL�g?���d��%�����_|O�=���r}��!d�>D��
K�]�_�/�؝~����	�q梍[���D9G�<F��;�c@�q��ܣ��苲��@��ĸ��څ�U� �3���`���mup�9����͖Y��¬L�,��x�8:=�@:G�U�*7��Hӟ���/O����z�7J�U���VZu0�>c�ɪ`��+��c�+6㥺��#v�]�{\N����s9Ox�����y�������/p��q��CA��/�º�n�	�!�1�%���q��������\g"e�`UC��C6"���'l�i_�q�J�N���u�ȑ_��,��|�`{e�s�r�z�T��H�>��Șc&���K�6�<���u�������;8���G���8�Y�3v���c�D�,D4aS t֢��P��|3��"泚7y�B�t�v���X�XѾm�/�*C�	'������J�(NƂ�r�Ib����{)���`�-(v��+J/�����y��"�c����ɍ���BT	�=����J'�9Y�4���:Gm�L��'6�Z\e��&hV�DD*���PQ������*�Hشp�ɾ���b$�E����z���V��h��������1��I����5��N��[Z�i���iu�v1-=�(te�>����"s�bd�<�[�4�v���"m��y�9��R��f���!��[����,�����\���E�?�W�����n�y���9�:����r���[L���[n�x"=�;����+��
��N�"�:�&�Y��=|�\5�e�ON�ù��b�J�^�Ѯ:~?��嗬t��|I�
%����g�U�?�W�� ��ȣAoT�Ǉ!�^�aCG۬��LGv���#�99Z&:��[��&I�K�7�O����>��}���W����ot���΢���cV����>��0��;G ���J�z"�-e�2��`2���?��f�������/���O,}�S�c\���ͩ�����(g'����s���eK��O��|N!�C��>���?�B��پ�3�����G����8^<r�+�z��oQt䌸���.�=^5؊+h�QvO�Y ����7��ҶS�MF��=X���6VZ����ڱ�H}=�����^�3�|�O�����+��\�K�s��!LG^;��2�b܇���b�q�A�\�pl��#�۠?b��/��s>�yޒ����6y1C+;�wK���SDQ�	�O�H����ᤧ̾��!&��aV������=�q��{u|G����3]ϰ�+a~�D��Y�S.�.��\e◧�B��g���Ѣ��xN�0�​2�����?c���8�N����*J.~���jܬvev���<���I�B�"FU�$6���,{�w�Co����N����tp�8�e^D(_�4N_X�lыlV~��T���� �pL����RC/Z?�L�S�����R!}�Ȑ^�� f�����x�(J�3�Vx��T����^�������T��;rV^%s������
?���4+�꿩���J��)�T7�3h�����j��QC�J䵥8慁L�eY�����(�:�r�*&/�<7��������=DW�$ԋ?��R�E/&.�Ȧ|V�	� ���D_�'X^�MMy˖F�p?�T�%b0?�#���f�N��4�V�͒��a�f[��]���t�!��5NOz*m"]-�=i��4�j�]�?v�6�v���&�n5Q��77�̳�Z���z�y������>�4�k���]$��/5<&�&��=�+�w���g�y�G}>u0���Mo���c�زr.�rmվ6b������FK糛�}�h�s�K�u��g17�\�t �Z���1�`���o�d`�.�"�[,�Q>ڧ��9a��Zu�*�P�Ĕ8_����_�:�����ax?g�=_��q���v#?��H�RH_/1sK:��JE�u������U(�l�"�r�0�S�M����yMէ�z�-]TR9�����8ay��+_��"C B��ɧ���c�W^���=ek`s���(Q��)-���	'��Y�«��flC+M/��	KxOp�>�Y�����������I�Cm�32&��3C��� F>����0l|���˗O�+�n�P����,ϧ?��L��9�_�5w~���?�JaO��n	oP�ҡ�!5�QL�lM�Y+e�L�Ty�~:��
����oⱺĲ��)����O�r�?���矝������ς<���׼����/����#�������f ����E���wQ�ځ<��H׻�|w�
��5�]�g��jtB�!�v�ji�Y �ʝs+6o�mL�aܴ�-4�m�݉{J2�aw�~�Cʜ���-$+��=Bg��!s`�C+��-]�إ���>�#Y-Z�R	گ��z��o��ɗ"��?c�@�5���P<r��v�*��b.�SW��
#��h%�Z1JHaC���o��r��5�A"]}D (�v��y�#e��Ʌ
U�F�j�*O)�-��GlE�0Ql�u(|�ʖ��|_1�+)��j�u��y�8�9_�Gi�>�GG!P�/Ћum%,�(�vI�/��h%�f�ʤ��X��X���X@1�ܷ��F� '���|W^�����s�rð��ؼ�.1&�)cNz�>�<�6�47x4j�#we��x�l�J�����x]�(�u
����9�s,��+]a��s6[9����Lۧ��jP�/���E��|�<��3n�q\��=��/.�%<���+j\���}�-��_/�'lF��ض2�#."�m`sV)lw	���*W��k�Ӑ<#���7�>������={V�>�M��鲼*������Cu��÷6�6!�M�ӈ�\���"g�A4��C�}"���%쇬~��2~�>0�>��k�"��:oe���ў�3�D�yK��V�F�p�Pz?� H9�Y��+_I�ʨ/��9�l���n\�X�+F�ȫTi+�����4@	�=2"��^3�j��ý�c^�����;��P�D��H`o|~�3ޏ?��e܏�e�҄.�"Tn�g�"�R��#O�S�D�U�����+>X�;W�X	�+M���WZ������_���������K��н`.����n�!�ΖSe�\�$�0"���h�/��+.�^s���_���şO��o�����<�#6 �b���-�|��~�&��1x�+�c�<��ZF)z�i��lV��0�L��uvN0E��ؖ"���ˎF,�Û2��L*�,VZy��N3�w��2o�=��NO�Y2�u�8���ge�lX1*;��B����	�;n���#W.��u�G�NRh./�L���*�-);A�WO���M��\zA]��\�����.�0iyt��	�pM�$�H�9Ma)U6������)e�4!R��CL�\Cڅr���tn�/8� ���1�<�?R$,�l���Wk/���
�i��HGf�I���g ��2Aw��QohP>X̪�9V"W��[�z�%>�ml�T`�l�dN�k�m`C�i�8>ș�� Q-��ks�7o?��N��/
�j����	�G�9vEE[�o��I�ٙ�:�'�7A�U�8Hض6�	M%�OXW0�� #D��x�aM�⣻�K?��L�nVx?m@��z��t���k,f��_H�?���'�)�v���O��_�W��0����t�"�ݮ!r"����a��2��/!q�.묮=h��ʕs9�{}������ԅ�G:���2k���9ֵ(S���ͩ\s4�ȦB0��P��7�-¥$/�,^8����{��=�%����k���|��c�"=�+]3CI���M+ 
��Y^	���[w�-=L9�R��{�r� c?M�׿�Q4�#G��w0�+�s�a�t(Q0�U��'�Ӑ[��l�!%�a �{u�/٤����cx�2�@���%fz�~'��/7���X�NFq2�+ɋ�õҵYX酒�(���m�w4����+�U���q }[.����_�����������l�g��_C=�hr�� �X��&�E��ɤΔ0�^�|��K���c�;>W󻯾:��8}��/���5����	��|w[<��R��(̤�HU�cG���d�)r�P�4�����E���`[�a�gLq��Y$�鯙��IYi��iA��DM��`a�?ԛ>��Ҫ���� ��Vf�d	�=iy�\�K/X�v��B�Z+�#i��f�Mn;�Ef3��uF���<�E�{�������e�a�bx	�Jf��r�x;	9�ڧ�����CZ��AR� �O�̓g�\WũX �xhI�2i���&Gm9Y�ŉԡ���7�l��K�ȕ|J�SMaI2jU��PJ��N]��RH
��
��mŃ�W�eĥe�X<I��$eړi�8↛�Pg���G\s�t�Oh�O�fN� G�q��X6�����8��2�b1���lЩJ��U�Y�fT�T�m:��.�G}���[~����܇�b��#^����_j�l]�ؠ����?�����t"�/�\'�K���Ψ׹�n`��S��N:x\��8��0�)}�Fye��s����-�cê8�!䐳�u�}-I>�.��>����nEDf�1�]}����Rk"
�_yml���g�Xhe#@���+[X}|��k���w[}�{������B���=��Зi����CW��!Đ�&�%S�W^�̧q�HV�^��i�m�	��(>��̇������M�\������Gyqh��G�]V��$2k�ȩ�?F����}�t�떨G�"y�����C�u���׻�����V�[��S���'�>;eҠ�z��UX� �,*8N1�8`�WéJ�.���4��V�������	�/��+�na�|��\Ȭ|�*R1V���^����Q�~��דe�`?n{�`����~�3�G��',Y�����r�:�$m�H0���=\G0�?;6�����6N����/?��W���W|�n_���o����2��s<�#� �3�Kw��"�ҕoқ�KEfO��e�9��	�O8	�E�;@��e�L�pl7bes�2�L�\(�L�������
���Ea�������ZK�l�[g.l�5x��'�C�ǊR��d3��>�>鷱v�#&>��I�#6P@لq�d&e'���L��-8z�?�u_���k���!��\4�7��� �?5��Es�����RVǣ��X:����=,=�&%k�Y*��F�-Y'��$ILڄ��B�XZ+kO�t�W�LURl�5� ��o(n)�����[�ށ_mkF�8y�&�^\J`�c`kc��0G�Ί@%k? C	�m����
	�R�� �S~V6�>�� h�	��ɩZcI����rk���<������F���pa�����˽�I#Py��)�D�S�	�KJq��S=�z4�xݿ�-���=�ok?�&��d�/�5-j�sBA^�Ͳ�׀[�h�ZypI���M����q��'������ب�cڿY����)UW�I�v�H�w��ȧl@�.�W܌kK_�p�u]th�(��:~u�GS�j����}c�'-����k;�8;�Ď�iUd4%֢D�M���YiS�|��o���4�+:]KF�a��0���<&?�T*��{�$[}[����M�3򩇛�9��m�\�0�~�I˯�]����0�
����.��-��l��,��y�~+Q��f�#VX�E�DK'x�FE�g�:��1�qU��g�1���P��$�G�5��%M*s�@��a�T���f-��0	�m�yΟ5��7�#e&����P�GC�:_"�
�����dH�ps�"�֨���x������ϳ]־�7���Vq�_�������o�yG�K�o9��0�8�� ڙ	K��6�	oufm�$�t0�;�"v��j�#�4v����Dm�B�!�d�L�w�='���+�s�C�P U���l)(�̿�tz�ir�D��z!Ϣ��7F��uJ���M�T8Pm�Ka/��K��G?�>�w�[Φ��ǖ���@3&�@H�]��:#��GS�	��%�u�LU���"���j?5?�2E�"�b!��u�WP%�<�!�3<����S���v�(s��ŋ�"���M�x����cڶ!X+� I����V�G��x8����X�� �U�j:EB@�)%�v�S#>m��<iZ�Y�}�q�C���;�F\���r7?pk�4��>Yp�*f��+�iG=���T�bVW2ns�����>��d��{��3�JCeS�r����Θ��*��i ��]eI[��ہ��k�����.�[�'v��&�z�{�|�H�X�p��3�!�=��]E��e��c��G)��ʬ��~K���#�3�{�n�g�]�'�@��Q-�=�K3�JM ~���r���*�C�~�$N��ƹ�)���ߛ?��M�0��}�͹�jO?؞o���5���,䍓�82VFΎQ�$��Y�A =��W\a��{lv����W��5���~�д8�6����x�,���mWx�|u��]ڥ�W��w�-_0ȵV�v�ssr�d��!y,�!�6����~ k#X�ښ�VS0��{�T��.ʞ	;�v����RF"H6�H��i���V�&��Z�#1�
5j�M��tD�	ӡ��T����WQ��kc�;֙9�*��V��v����b9�L�u����_c��f�<�'��h+�S�\�a�YM���N�@���t\˜Ǚ��i�8^�c+ڭ�8S:Н�x���|�C��mI�P�����4{�%^�[�QQB���A��V��<�|�lݘ�0YIK`N�M���Vj��0'�B$��t��[o�{x�El'�5�YM�,+ג-2X	��9x����c$m'���8TC�S��b)1�G��c����FJ<&���o&��ߔ�[�.8�"�0Q%����u�J$f��X2��@�-k���o��m��OX����h� f��qS����BÊZ��!l�	0���� �"�J�V���bZ�lpȧ[�XOB���uӶ���eR�O�\�9w�0��*c@���He]�ԉ?W��������2��D�����-�M�ǋ4�c�9oB���x'�����]JT#���ٕ�Ę�� pnl��Յ����~�~��'����S�i�n���_�P��q��r�����h�xF��z\o��Q7�~q�"����<�j�1y�l��%��ZP�ro��e�?{uz�':7�q���������x�b��#+Y�z�3�CX����7qƟ�xC���F�&�8E�̢�+s>~\y�G�4dE)�t���'����#U��I��z�{S�J3*���8�5�z�fa�+�MyZ�Ǣ˿�Q*��&L��oG���`X�DCC�{��p��@�_ �r�,���q�˅ӆ���˨�~�F*⌤�sN1d��T�,~���va����pi����w�3h|A&��g�_@:P�$e�y��簷	<�kC(�:���*"��B�����N���~z�#�?��4_��G|������N���<�ƶ�|�v�Ǎ�&�E���@�RA�ڽ�:ˁЙ\��R��\�����Q�i�N�gP/��C��#��ӶO�(g�!�J�,���2�	��R�� +�+������vi��,EJ�sb�:b敽z���sn���e���.{��1-:y�-��8(p� y	'�y��M���*��	qm�HY~5,��a�ߐ�Cyn������=B��(Q�+OV@�����j]Dp��)��K�E���T�8�-NI+պ.�Si�`꣋�(p����2�v�*�Ƅp����BR@ dI��;c�vi_2�amS���)�bW|qj3p�6��	����aX��U^U��V�3�,ٶ��B��,/L$�u��Y��K�#���͉�[��G�M�Z�	���G������q5R��iL&:��3e6>껒�=b\̽��Y^�� ^'V���(o��0i?a��`�~H��ֱ�xK���^��d��_���)_����FqPm)WO�_��c���aV� M�6]�%�x
�>e�8��}�'px�?|ci+�O�����xC�����K<�H^s�}���00�'���1���8�����G���M��/}&������yA{k��i�qd�uƐ�2_h��,� ��/�e�{�z�a�+ӝ���"qQZj�o���i������� �~�Nc�/b}����.���{�`�I�K��C8�*b�X�p�eŬѕ8�O�a�$A�X"e�~�t
�Y�u
)`F�h��Ph9�vR�������x5jZ�H�����L���]#����Ggn�����\8B4�]��	����j���u*�.!�����`x���ד�>=}�����n↥d�r��/� 9_�a�e�g�f`'�����GǖG���f�K�7���@2��H����3 L�<��F,tB�͎���ShPMIHW,9I�rl�]r��QX#�f��(;L(-.�C��:�BnQ+�PY�/�#���>`^����\9hǤ�o���5����L���`SV�\��no8�lr���1B�k�סS\���waRn��q��#�X+ �ڤ/�����G�2��bŔ�/l�V��B���mBG��%���K���س�'t�=��5��¬ �8aSиv.v~��$Bf�rTV@�0��-�U�Ė��ڭeI���~֟��?P�!�^�T��-�
ۨ�S�/���zq'�R�k�|j�B�U��>�)o��XKޓ��EJ[pHg!�����`S�x��a�d�g���'��~�x�2�W��o2/��E�Y�S�����n�Fb$(��3�i��0�g#<H�ڄ�QO�7����e����3�e����`V���I$��/��{�P�.� �0"ٶ���ڞH(�>d�����ig^��x�ёD�+��jy�m��v�_?�+�/��mĲ��c�mH����`�t�݉�IZ��FVEN����袽��|��u�F���!�:2OqV�)k��H�	��B�������kkۂ�\#���QER�#��U��/�E'�YVl�]yD�I� �J��9$)ƈ6��Q]Cp�hpU�8���������S`�Q|�^�Ã�q�xg3�v�@
�*�.E+���G�~��x_>�>����rBC���7t_���v�9����m��X�#�������?��!d���_�C~���r��Y:�W��^�|�=���-t�GW��gƦ��S�"_�Is�1(�g�n#-�����ʿ�Ib�Ħ�QLk��ʓڅk�� %��Ng��-(�=�f�o����9���H29NpX4�$-~�����8���X�**���S,����}���I���&�)�ALV1�j�M�����N�o�z��J4Cgii���D1�֦x�N�j�F��	��0�!e�+cSѿ2�e�E�p.
M��=���R��EUꝜ�'�]�u�Z�
k��/t+H����_��/�X�#y��җ�!�"�Bbc�,ik���6�� ���6�G��D��U喓�1��U�Y1̜�8�|����[��8�!"�8Ҹf� .N���xU�RY$���8ߋ@[�fn{���YM������J$#\2���p��e�W��G
ƌv�:��FGϠ��F����)Y[���#��ί)Iw ���>�ݐҸ��{�y��..Y���v?�w���Y�)�`�qL��k\�7+���E,�'�L�"|�1_���ؖ�፺���d�Dz��u�Ix��.=t(�!�/&�|##y-r������8K��ʧc�e���dB�z���ܸ�/:Ҭ�{�g���eb�+#����N�﫤,t9Ƕ�A�YE�8a0r\���`A{�MI��F�\y*w�&dյU�6����tB^ʋ�*v��<j�@�`�7���]��&�3�}l'���Ȍ��~�O�N���SI1<�tYJ�<���O`x�B6A�D�Vw`ٛ�0�^gV$�Rd���i���x�|��r��e�w.{��N�QeY'�C�k��0��yg,�*����x	�NX��3��A7U��V:��4/ �� 6c	xΝd�iI��o���MN��FI��I�б�L�!��Tӭ��v��'��
��hlp�[��)���L�U����^��Q��&D9���y/*�c�MS;BF6e�K�y	/l*�:�-���g�/K(�V{NYN��V�chYJ
��B`ŕ��H���
�t*����Z�&Y�R`��w�*�8�K���$G�bWz{�)�b�����2u*��0��~�>��\]��0��8clF�#���~�U�=��eY9�]hU��Ҿ`~�It����c������WpCqN��%��6�����F�g�Gr�r�!3aJC�A�yS'L92�f�t�
��ط\��.s0s�+��嗊����sK��Ż)�ȫ�r�xy(�����, )W?���t����P��u���3*��\b��'��r���ǃدh�ۘ�%�����`#�Hm�8��K,���_�ꔸ0(}	)��N�E����� I�~��(�s�T�a](י��`�"[c��s�Rze�b�ѧז��-�I�~����! ^�Y�cm�,�lmy�OrE��$�
���)^,fbaZ��� �F�Q�կ�&��Y�͵0.��N $i���&�(K��9`{QS��/�/�q9#�΅/�se떲��a\����f}���+sǃ��U���_AL��[���Z&F�+b����lhȥ�:"vT���\n�᭳?�WS��^�!�QX6��yp�]fc��4�����G����8�#��C�u��`{?���gy�}���e�x�#�	nq�⌁�{�0��#2��FH8�S��q"-^��<�[+��R���6�����02�'���0�e2*9�)u�����Y�����1���I�U!ek����+|�aC&!��@a�N�#r0 ��q��d���g=��8�!4��`l֠��-"e2��@���F� ��VQ�%��L�drs��Y'�%�8����WJ�;u���:���$-���V���S8K�+�^���¢��Y�a���S:�k�j�K`�'�Vy0Rف��8���C#7Z�k�M�0�t���4#i�� I�a�1_������+�w��o['Iy�e:�%�(��1ds�#_�-�ĕ�B	��<�I*��#|1-V���#	j�P�s������ǒ\�!�
��ٸ�)]�H��1�I׶2����4!e���ӫR��c��6�MVy4�qI��a_q^u����V�(!}ȄAG���w��
�A�]�:u��^���e���B*t�5rV���:)U/_��/�����b��=<K��yU����`�+_�;��K%�-4���SV�%���{��&˙ǔ�y�J O~U�����ol��s�|�Y�4���f���c�$:���Ȳ�TC�uOPdz��� �@�W��;{h��a�P���'��C.ܑJ�"u歡Ja8T�]����<�|���l�T�
?xS�Rb���>��3_#�Z|�l�@Sno��PB�<'���d5�F�0!A0o(j���^P��+G�A�r���;���y�/'�Q0�8��c�=�)�	t���L���6���t���q�d�c�)�A�2+�wO����ݴ�.���M�B���ҕM�������d�¦�X�۹6޲��*{-\�'q�끹�|�dj���*s��@!�ӆ��k�v*��]������i���ShHG9� ӌ������F���� 3��L�RD_���FBq���]�O�V)C✂���`�W�R�S˒.�4�舗`�]zȻ��-�@�x�D�F�i��P�{^���Hk�ܴX"H�$W@������z#���v��Y�RS�#R0#���n�&��`���b:�ԉ���Sfb�)��n�aU%���ΒE��%�X��T4R�x/�Z$�p(ʴKs���(ٽ�Z�R���S���Lj�_QV�A}�wiE�:H$-_#�4�9�pl�n�Q�$��(X�a���0�Tu�f>�dQl�N/��N���N��
����ɴ��L:>��B��8v�-��p��%n^�
���J�*�#o���:#%b0�Ϋ�t�'u��B�>�.ļx�'�Y�;~0������?z�E�7YQ�	T& ��qH&Zɂj�Px�CkWe�n@�<ؑG��n�|}4�D�K��K�}�J��F��ӱ��N�ѕ~���Җ��۶�=��w%��U+�z��/�U��稬��,UA3��ϸ& W��5�AĆ���
��ԣ*ъ-�gE��l��_��AP󮄱9�z�】�b��AV���sV�Q�҈��`�Pƽ�PVu�lv�:4��m�X3O���*7}��RUj]~�	n�bB���6>�@3FWpv�3��Z�M�2�@�x�@^q"̊YyR�-��SvL
�X�M�aO�!��;�8�c����q��2�h�)�TV��n�!��l�I��|�g+a��56P�PY��#,�i�g{Er���H#eH���o�)P�%�~p��Sk�e�(��RNb�ih-�!\�{n�1��[aFF�nZY1� &��5\�'Tsͦl2��
�x�N��=��Zm���f�pL����0��?r-�R�r b�����v7�&��d�S�sQ6ͯ{�����M�J�<�W�,��z���E���%fV!�DD#���m6Pae:�,�Ԗ����Yn�˘�(��Y=�ˮ��We=�Vy��2t�(��,�u�I	c�K���L��6�i_5U��1$:?L��D��&&	U�pm�r)����'5���A(Gi4L���F -��w�9�y=��:c�k:'�f��\g�=q���gO����Q��/&ܾ�|�ggU>����@��oY�PpHnT�<�FA,���Z�"34�����{��kXD�sʕ�]%���
�0�� lgv��F8�����;65V����n���b�.L'�/! @忎��359����"�����Ag�����/D�IH�&�9���5��2
9�b�-��@s�O�W���ء����D�qg�o{I�ʍ���LC����Gxgv��� �f-�,h-!���0W�N�r��$���f���1���5�Yq͇Xt�@�	���7LZ�cX2Ď3���`��x�bJ �UXm�Z��2[N0N��I�B�!R��C}���Mq���Bb���L��@^$��m�i$���2leK���S��4��{��W(��i�iVh�M0rO�xS����ت�_� ��6�Ej�w�٧/�%S:�0�C�xqI��Km�/�^䏔ϫ��!���Z��8g��/�i��b�5i|!S�d����M��N�6.��Aӄ�b�l��'K~���Ʈ���޴y!���sS�QuIG.��K�!�`N\o�/��r�d�M�|Jq�������G�Ny�²������֚�ta7����Zq�g��5�-�����F�>����ߌ��ȳd�t�قKSإ�'�d�7G[���`�4ȍ떲��н�`k����_T���s>����S?T~�V����=�yvz���q�x��rPf�6�P3�����`4n��*{c)���/6�	EA�c�_�{]�<iW� ৫�{�>�W>s�&+L��n�Y����S���7�QzdzE�lD�!�jmq�I�����t˽�2�.�FT�x�Z���E-DdP�R;�[��pK��:i�qV��Ug���靼4t���c�}���^�,jq�Fg�Cuc�Ѓ���9�=ҕ�h�5g�`�D9<�/`�a���+�od���R���ITV ��ף<�O�!�hP��I]P�yg�V��%�v���Y�Z/�*�(����\��\z��6��m)Ru_�0�Y^�������v�/٦b�4Z�&�`�ca�6���
D�D��F�\Tc�e�2tZ0�G�M���G|���*�������$�;��L��6x�[&U���Mȟ *��;�}4��[gz`&>�aT�J�>����+&Xv0�&+[%-+]�y`P�B�ca$:�>:Ya�xqdaz��-���R��k�@�=|h� `�Z�8'2�[<2�N���o�SqO\�N��k�7u��؄��xK|;�-B��
��c��l��G��B��R-��0
Z�!ⵕ
�e/Z+��Vd�l�\�� 
#�T�Դ��TP)�-C���/Dj"�'ߙ���7��c�����������)_�q��5�O/�f�?`�W��������H0b���W��q�R@�bɖ��R�rme���4�,
�T�8=�������V�J}`�/��B�{����c$G���&Z�ڐ%����'J����s��uEk��P!m61)sбq�]3�Ҝi�Ͳ����j�!\S�q�c�������(�q&%�Ik��n�\��]�z�:R��������p��|�xߘ�N:(�@�6Jc�b̑���RQ9�d��:|i,͡m4���MV������ԉ"@��n%�=��%F�m���m�lx�[R�2�"������n4&q��O���>qUh��ӎg8d��6ٵ�����J~�Y�oGi?q�3؇8�>m�Ʊ85�6��Z2m����ƣ�u-YT5��.�]�N�2��7��v��j��L���Yf�9��g����,92O�e~�J<}fhLl����Q�~ܖ��~�^A�󶒠��B�=7�r�A��}I�AW��a�����0[:�M���j�zrD̸^*���cxO��tb�)��;__�e��t��v������l���6h�D�R�M��o��Δ��#�Вu�+Mf
J����\GR�	�BZ���_�8�)^r֣�9�k��鮲��5Tۺu�X ,t�����2�!��xs����}����O�4���ĩ�c�g����ї��1��)4QI{�wNn��6K���JêY�rK�okp�E�g� ���)^�Qaq�q��B��`������x:�����@�"Hf�P0#���8+�ƫ.Jz;B�e4�so0f�aئ�8 ��z�:8.Q���<�H*���I��0m��'�-XZ��2�#a���/״�#�������?s�`�ԟf勸�xKq뤕lq�����g�Qި���%D�Bu;J��=�m�����=��F�����ơ#�BN4e�@qV�X���GT�	Xk��*v�M�P\��\����:�042H�O��G�.ف��X��.�C�c�$�c�z��H)�:"3�;�0Ғt�GleY��rЃ(�t��2��u��.0b1�JL���IO|�$G�c��/NY`?� `#�D��#ސXMt?�;J��Q>A/��3�3�� ��,���X�c�c��޹2}��f#�_�Ba#y���#�IO�y��C��{�������my�ns䱗��_���:������S`���������M�/%�<J��K����2�?.�cU����%y2�3/�׊�v����pi���!H����H%�\�5��^C鏾�e�H�
���+�7�p��<��˾0�˿}w���oy�'y��J�<�{�÷�|uz�7��RP�]QB�<�#+��&�P�G���Z��ʌ:�<��_�}��@_<[{����s�+�u聪M�y���>��5��#�U���CVd�e�H֤�NR�p
CU�H��x��f�XX%�Y=I��p��$_�bQ�J`Hc�v;h�Pк�Jg�%<d&(���v���@�B��e��M�����o���Η�ݾd�2��8����g����O�?���yyŧ��ݾJ�����4���/��J��C��z8��V����kSn,���_'5%��q�(MX|C? �vж�p��x�4��5�9/���@"I��	=�K�~j}�cKs���> vr(��{��r�����P�?ۿ6��I��0��dH�{,��%�X�$��w��݅�.�<� ]îk�'<�&�v�� �!%�NhYF�=�������X�e�  @ IDAT(�qdT����و�U�t?����<�;���?|�{�X�#�U?�&;��oʏ��N�m�/_Bh�-zK���Q.�̧l�<��ŉ<�[?8�e�>h��d�����f��R`��8����LjH%��u���`]�bc�69����G�st���H�RԩSde��pTC<��)�>�q%9J8��f�hYp�ڲmS&غv���ʥl�F��(<K��Z:���Ʈ�y	��w���O�L�ĈG�����/__��+��~�����;}���N^�&_r�*��|�tyS�+6������\�޳ų�]mi���Y	f��Uvev&Ε�Cq]ɺÑ����(C��]ĕ���[��B��׼��߅v�F�8r�oНoa���8b:a�+G�,#i 8oaIi��+�_���Q�u�"U5T)�Q�(��n�Ǽ��y-�oY�s��eXŋ�^��Q�ⴹ�񁛆-g�vlu4��j�)��B�Y�������'?W����oO���8��aYT�h����_A�B>�����f`�2a9|�L��uT�Q�0��w� �7�Wʑ[ٽ��Nqt�R����[��4K���t*��6{��H��6�����ᑘ��_bN�����྿�˙��g�7Z�b.���,��m���s��6�����.N�b'�c����͛m�p�ZmR��=�u��1�p{��P�Nد����R�#[ ���J���):XޢJ��qL]�k������o�;]�(}�őH��C~�AV��:�?a����� ��oQ�:�iiOV:��eT��?��S$i�h栖P5�Y����`�x�Cp�\�ߙ�o��N�Lت�2�^ ,���A�8z�U�#3�K�pl��A{M\jf��)n�B�	{�H�.�p�t3w0�U��ɁM!Nq�x��5�7���ʜC��_�B��V�*&�<]=�.��ɛ���.�:a<�c��+���X�z͵�U"����O������_��u}�����7�����7��__ް/�k�Û'�;���xX�AO�c�_m�X��f)� [�#sV�X�z�cFc^�����[�v�x=�u���T>%�����-�����7,4���$���O��C�0�q�X�j��R��	Z��8a3���4�v�:a����T|����tw��C�^���T����Wt�T��#\�I��mB�e�>�;<���\r�b(
A�	��X4:墀�8_>�u�S�����;I~ǳ�?����?������;=�����x�f	��Qܡ�߲�ӝ�'FyK���'{������v�ԥ9�F~T$U�v��/0�C��'�;`*GPd�j��3[.!�ٌ'����V��ua�����
�e���s��'Ζe<��~�MeQw��5y+������7-v@6B�U�W�Om�i�S�. Ǯ��LnG="0�%"Y�΁kE�Ji����W�1��(VÖ�ȏ��AJ|(_��ŷ����{o�4�%�3����I����\H��:0�g��3���HGrCcb�&ؚ�^�e�Әi��&���%����6> r${�q��8��-�GZoUN���-���Q�����>z�g��w�M{r^<έr�`၍��wv� ��2oU���5qz�Ħt�$5��l$�@!tp���hX���1��4�!���y�^��EN��s}�&����*:a�h9��a�J�7ߟ�����o\c?�����݀��)�]��	��0�p��ӹ�Z�Wbb+y,ybs�۽QZ��� 2O� �S0�_@�Ֆ�|A�=�*�'M������\)��=nW��^���ن%�W8a>1���͛�H�V���Z�0@�p����d����ڌL��th�[�Ch��8�G *�ڀ����}�o~E�2}Ń�
.{��z-������lR���L�N̦���D�k��G~6�s>�������~����߰�͂�����������G߄��i��e��"���`�"�LHBI-ఓb�d[0�-�:'j: ���_�h������[V�_�$�R] ��&/x[0)J�$����v�N2�e/lw�O�:��K���`�K^���G��K�RfE�V(��jTo��U�'���a�D6�e(^y8�w�7:��%2#�eʲ��r��	��/,��_LP�,��?A�ަ��I���8o��["��m�}�S�s/�*<�ߡl�1e#��Ǻ�}Yw��;uq�+���#����䅹ܛy�9�eGڗu����^��v�����>�M���0��G�[��^X���j��oa�m� �H��#���m��@�~Sl��,ի^j{(�]_/ˆ�^)s{�p���"!8ɓ�k��Ԅ���ܕ�M��*Ѿ��G����o�>=}��7��>~r��g<]�Q��ʅM�>n��1���oNO�؜�j�~|z���|d�mA^�	�t��\y�\�s��%�{��y�.���
�;������XRZ�J-��3����/<���1�+����.DA�
�_ᑏ$�i8t���Sۃ��WdŶ#��a���Udk,M�tf�KO/��kV����J��ŋ5�G��9��p�!�c�|��#�w�+��r (%8:������47`�p��E���Ek.5�SS�A�3\��~������ߝ~��?��������eϫ���?�G� �U�v�[��^젷��m,e����T{�S�XZƊk7O�
>�`9Z�Y�N�)�48��m�X "l�����Kj�9����������[��8�=��,Z��I�m=.;J*}xWə(m�h38�:m�@,�b��%}<�L����nL'��-���䱸%�>v1��d�<е�@{ $~(�Y^�{B)�{��SE�u&e�%��o�L;�?�Sj,����z�S���K�Z�X
�j���9���&�x�h�J^ʣ�����IO<��Ҷ3)����CJe�.<lp�5����,����VC��2#{Id�������}��e���G�	D��M�O�!���
�]�1�Qӱ���NGJd�ټ�rw	�H�Sw���	/*/�nm��E���_����V������L�+8����
������0+��ќ?$ˏ�^�p�S���ԧP��}��������W/��>��%�(�ľ��J���6������y���N�>�r48�n�ޤ�~��o�޿d��%N��B>��mA:d��1oo���s���2��~!������K���O􀅨�k|��|��]ˊ����%���Q4\��
��H�������{;��V�	�pj��'HY~�	 ����t
I�[��Q�e|\��'x�,�ad1�3%��?��O��R#�,!Vvxied��F�h��~�)�?5�����2������������/_~�Q��{�C�>��eX�>�,�
�-+_��K����!5 ^�Mg7��˦�,\k�d��kf_��rA,�V����3M������T���'F�s��-��L,S�|}�2v�i����*�
Z}�W��c2�*�v�ŏ�΄���`g�8ȼ���y)<8cK���z�<q)�`� ��Y��DkG���|�ٲ��ԅށ�.�2Ӌ��_i렸<��4L'������_������ļAR�#ȅ��J8�{��ty�|UoQ�OzN?1�K�� ��S^�Q�.:�7?�}��-��a�1��?����Paٔ�����{m�0��]{�!���f;�����'#M�9ɷrSzO��c�ipJ[gي����'�x��e|D�t��(ee������Hm����>�E��U6�l��P^ɤ��
�<Is���L��8���˴������� �kex�˂��Z���C���_`]\�n�Sg�Mw>�"�E��o�w���|�5����x����>=����>�5�v0"W����C6��}�5>�׺f�a>H���3������ώ}��?���)]�F.4����a��c��/��z�|��w廾��n�2/.��C[�c�*ƛO_�!�N��+v��׼�Ǔ�;�����#���- ��~��/W��C?�����_���K�=��eUGI�"!
m�#]&��"�/6޹��/!n�Ru�nX��y�1�~׳������y䌌8E~$1#�:�5�2���[�����tO��Wu�W�<z����t���_�����s~u�X��C�lV�x��'�8�������6�as�R��Ѧ���5�v�	D؄ؚ���1H[0m�[�7�ڎd��*�\��m�a��īB��@6+�^/�)V�B�%���X�)3� �d��+y�T�m��vx�h!�ӡN[���	4�v��: ꢷ,�7/ e�`��~�ޫڭ���֎+,���Ű��|���=d���"�j�%2A�"e�Z�������>Ń?�@V����V憟�	-n䘚��#m�
��	��r��76Ծ�^�z�M_ZGz�/�/䇈�m����uP-��->���S�Z��#�t�ָx��K ip�Αòv����
�s��S��(�t
��,;˟H'LG��~:*\�Sѫ_d�`լ�Ŭ^�Tlj��sp�ӆ9@�L�$��ٲa���V��iV�(��{B��c3�:?��"S�c懶��ڃ��[w�ٺ�(1���J��7����Ͼ8=���?���k��"�"ߒ m���P�5�5���ts����u�F�|T��n:]R�~�=�uq�Y%Ιp*�ў���,n1�b����#|i�����n�B5�w��ϰ�㓽+�G�����
����x��䀸��E^q��g��<�}{�G)_�����>�t_��W�*f�˔�&�@�6���`w8O�Y���8N����~xz���q�tĖ�ZE�	�y�*�+�+��{���;H��o����}χo�}�3� z���Q�����ߜ~����|�����}q�Y��8`l ��ro����;֊~�9�<4;�9m��&�]��	�JNZ�|�-�0v⤧���X�/�&�j*�&�r;�H�VҚ�R��*��i�t�� �Ge�x�_G�D����t�/1@��ұ�P��mz���Sl#��ot��/Y),|k�t����~��e�t-Q�Y"�&eT�^!�PD�T;� �ѷ�$���+�������c�e��(�5��I�h����X��J����R�����~*����$6˟��y�_@�r)���X��z��sʷΛʝ��wh�of+&]{��C@�#�)?������+s�2�������\�	Ȕ��m�&�����i���`H�@tPC����3�!�-I;3kbs�,y� 6��0k>�
$N���W<eȕ-�7���s�yN�+Fzj\��\���KV�|���4}�~�����W��Y�x���\s}䇿�/��隧a7<s�K���d�;�B�`eXb.�<@SP�(�E�h����ǵ�+	�_��yE	�t�,S9ü�@	(�:�)^�[�*�Û�~�#�W,P�y�
�X^� ��㡕z�6��L6�A�-��4��^���6,N��1�S�h�*]ޖl��"�_��0�<
�
Gǈ$�b~�ɏt>˦�7��灎��nm��e@_o����<~C�l�����W����ק_��������_���J���;�=`H_�������Vw�|��w[i5V%j�1��`����4����K�5��R'Co�ۧгS-0�;�de� �T��(�Y,A�����ȉKFz���KGڑg�\
W�.Fؠ9r�ݖ�%QE71�|Z(�To������cq���{z�7��Z���0��
Ȯ��jX̛P���:U���W�9�XU�P����l۬ܽ�*�з�e��@$ZĖ���T��Ps.j���&�m�����8ھ ��@E�A4����}���5q�䘖O��|d��Ė�{�
X�I�k��VI�ԍ�i��ky���u�;8+֞������n���[�d*BO�G���5�h������y`G�������<�3N��w$5�Qv��̫�J)�d���塼M�5E�SeH'Q����t��,}c�E���F=$<��Wqې�RWiM��R��:��Ѧ^z � ��<�����~��|�莺+���a��ő/�~z�������>���M�ON��S0V\ta���
��
��!��h��|e�9i���c��Ca-���8Ҫ�wi����\��K�5>��$I]��cN�ڕ��o�
M��p¢�P�Q6:���{��%��*�{����}�+��AB9�e��G�>e��)�)+N0�//��Y��T00(R*K�4kJ,��x�����3 o�k �Ig~�ͳ���}�_��Y�^�wA_��U��H:����+�^ ��i��ἸU�|����_|}�����8��o~�+��K�H}����}$d��w�������>~��M,_��������-DL�4�7�$�X��6�zL��`��<z��٩�׊v�I�v���a���G��s��e��L�t��"_:낊�2�v���aA(Q���ȳ�J2{?�ij�Q��Ioho��"���J�đ�ЎVp����JiQ�W���9!��)�]p�u�`Rng��䱘�N����� �3B��,2��ch��yD�# �0�� L�Չ���^���Ğ�T�R�"�w{����Sc8�6����\y'?qJGq�V���,X�^�XY��W���=U�+B�&��ꛪ�M?k�~�ʡ_JKU�=cQ������r�2�t�#�R�۪��{��R"�*#��Aώ)�W�U�ɤP�^�*�iƢxbS�ꚫ����f�\-���%]��ՑRvx�� ��p�8T�B�����\�����˱�k��cl墳�E?�{���ɢr�N2ׄ����a��/|��z�!m��F���&�ag�%�H^^MW��>z��)cb���@���۳�t�"����E�����[��7/x�����ߜ���7���_������~��G�'����G����y��՝���=�t�m��8<qL��ڋ4���f����U��5�����&�4���X�u�\�2<T'|W�ڻ?���՝Fq2�x��6߮�C��g������3c��ￋ#uC���H6��8��x{�%9�$=3�L�P����#��������ث%G���u�1����7u���DU�CZ����Y���5�=<\��{̓�:��uyp�j��cV�p�S�l� ���U	tθ�@�d�|�)@�{u�ߌ"��ŏc�k��~l�0�H~}��Kh�,�݀��|݄����s�=�d����7��������n�_n;����@�̷0>��W�g/���#��K�1V�\2���6;��㜰�q���9�Rjv��	R��<(��R�%hR�_�'���H�8��Fe�>	�R$�9�h�:������N�.�K�eG�N��ݲ����w�u���3�^��F����jQV����.g�ت^)�F���WiR�6v���*����X��P[��#�|�)�)��s��:�#HT��# �C���C��k8����6�����E��8���f`k�'`EJ�C��0݉���arC@;��X���_ͺ�q���]�ud/��A��őW{�����J���t��/}v�/[F��s��H:�;��^�������XXvA��̪�~����УUsaV^CN�vx���x�o��^摝P���i[�c�
>���"��A|4�ʶ�/G�^����0�v�E��4�&n&`A���Z��T��=u�h���o@�GR���zN�õ�oC~�n�w�{>�B���^��O?ݼy��2rK��}d���߱��?��6���� M�L���9.6E!�I2�(d��9�G��\�3i"&�	X?8˃���_ �1y��/���Zݽ`���K �"�w��|����۟��,�<�O?��	�go��,����~�x��$�>@���H����߼ň8a�黿z�1W4-��-9��2�1,�M��1����g�wk6i"E�����j�z �n��d���{��0�$�&k@t�� �����������x��n~�����C������7���3`/_����� Y?�y�{BL��ڵ�	���!�j���Շ�vF�-�����(㛀8�Wz�F	k׈[q��۰�-A1��T���$P���"n�h�e�Kx�F �b�~B��!zbwص��7��?�������^����M]*(̎Y7�s�t��7�B�+���n�-	�ڃ��rr��x�V'r�^��6�a�>�pb2�_�g�Iw�x/��Ӿ]v��J<�f�1�����o��h��fl��1��v�cr��[�A��q�e=�[3d9������2��1uA/`�����EI���N=��)�]�:��D���O�#o���×��t�����Ə����c����蛺:��ľ�9��Vu�e���9'|�Ó��b:�H�S�3+�$h^s\'�]k�9��{A���s�]w���|D�d�+r>�[�w^�J�����w"�x���g^��F����7����_yG�_������_���_�ɢ����7��B	X�}3qb��ռ,
��k��'Jk���>���}�hd����S��j�05����τn�9���Q��t1)&\.Je��8T�߄|�B��$`��?������7wo~�����=+`>���K�Q��W/n^�zE��n�X�������2�L 0�1*�Z���9Q�l����Ӹ�L���� 3X��	J`�'�ЃHP ���[�ˋS���Od��]_�=+_>|�m�|����-0��z��7�����@���2&��l_Gb��~M�v�[Z���K��v��.>���ц�ʯ���O��=�,E�4*wP�!'�]W��6��t����G�c5ek�A�l�Ҭ��������%~d����/��=�s9>{/��Y�7y��9Q��ս�x4O��Q^���nυ��ñFR8���.���z�rq��+�:�H����{H#N�v�c��Ks���}��7s�1�]����x���1�]Ni'V���g��<^3�>��3'|�i�Y!?yF��c���ߴ��c��@ʵ��+2i>���}z��;v��w��c{ʂ��5�e}���Bo��]�X��yc�K��l�X�����꣇Fd��X`p��#��U\�9�m������#�%�6#��_��M7���Y!ew�w�!�^��5�\S�)�6���>P�?ik]��bA�3?�����>d��cC�Cd;�X���Ǣ����[�Z�x���$a_�f�(T�Κ>���E�b��f���&{�2�<?�����q��/�����vc^ ��P�n���cK�\@C�s�JW����?\�����s8,��������`~��/n�2x�n~�۟n~�+�����&\�_���������o���;�,�6�a2G�.����@:�����$�"�VF����$�BB�d��m��Eq�XW��;�f�o��N6�o��J�;l��I�����������?�����y]�Wo7���7/���k'��H�oX��g�|W�A{��t�Rqw����)7˂���6[Z��?�Ʀȡ����+8�,���p2�.��hX�_}�XbNbZ�'h���h'c�O�X�H�X��5|h>vΑ忮�gS갱	�'NK�t�~t�\�W%�(�gXk=E@��r���ӖD7��ԿC��XraPLK�"r�����1��tH�0�3�?"O���o�򞴗��h��}�=N����ζ>���9��_��������A���Ѣ�QZ43N�rw�
��k{f�R�c߱��

J�0.�;�feH��XN�I��Sm\��xw颁(��j!L�����j��|��=� B�t[����`mS���"�yS��{L����:�����6�v���m3#׾v?ii�l:�:%��>ʮ\!\��ܩ�/H�[V����a��(�z�z��^ϟ������0V�>s�E�<������ݼx�5��Ǜ���s�?�������v��뻛��5I�a�����_q[�oF�������%w��J
(��,�6�+T���A�$�c�;zX��|�%�_�w�Ý�5Ѳ6��cw����'�|yg�����C���$�o�G*A��U�������y������Mn'z����H��W����sb� �@�%�w_̧k��ֵwdcp�q�-Z��,%�"Ac�攣�N(q�ۡ����L�:w��I�U�-T�X��=�����n�����g���o;������?߼�%^Y��_&[����

�/e�|�^��o1P��O[u0�ԧ���{��V��,�*��D5Cq�jȊVO�Rj��^[Q�*6�<!9�-�e��w����r`*�nx*��X�$p����m	]��]�:G>�kGvK�IkL@�nJ��G��"w슘S��R��ܘ�v�P䛄~�q��1611>u��tSq�L�����hG��>Z��u|z��e�>~�=�iÍ�ѳ�;�Z�u�Z�5om|܆�����(v�;�3�96������<�7LFYWs~�h���L��q����S�4O���1�-�P-�m�c�(	�ǆ�?�ж%�����҆�B�X��A�c�����U�g7�S�½v����a�˼H��J�m�2��5��C�rǇ�}��b���r-�Hb��2�8�����h��$Q�mOg`�-�5�j�%�q����Iw�
�_��u�śܦ�5��e�_��_7oH��)����� ��᧟o���/7���'���[M�^r���_��x��4��cR&G+�U.�-i��U0�D������[dhwb�sBV���;�77ٓD���y�	���F���\?�����W>ׅ�;_Fjt�j�_����/$c�6�����/:{��*1����('��0j�G���|��B�U�3[/H~��<�\ B���<�vGp}�Da��Q�@'�sߌ���eeJG�2���7��_o���?��I��D��	�}c�G�_s��._9��M����u���z���{���mKo;�����?x�O��9_�
h}��(-'�Oۃ�r�V��2�
��5U@�s<��|qNnme�E��1z*���˃
��/F�ి~��G�-븲�=POE'�^Ћ�Ԛ����a�_�˿�\���)�2�׸w,KQ�g������ݯm��=�?%�̈Pʈa6β�@��9s�$��Zg��)���$���Șzp_)mN�_"z7z�~�,���tT���fy��3rl�6��G����Ɓ]����14�sji���9�Co�������4�����z�?�7x�ݚ�3zw:���i_�N?�����b�e2�e��d^S'q���yf�h�z�y-9y8v��Mlx��Ŗ<���#����:��� ��IТ���#��B�r� ]�������K:��%�yK�<3A�5��o��k��xߺ�­����v)r�wy�����e�r�g�9��X��_y��]�z.	�|���R�FY#��8�J��y��$PM�����ަtL:.�ʟ_T�	����X��[L�̩�cil�5*�qc,�Y��!w��c!$�2��w�~�u����2Q�җ���@%3��u���b�m�kXjL2G�QQc}΁#�:���/^����Ky��9_p�6�:��_H������o����*�W��|ǫ$n}����mG��ŷɼ��SC~�o��'��a~�B���yFVm��	��G{��֔O\rb�Ta=�8�8r�$2J4��v�+`� �Wڴ��SC���j5�W��V����Y�e��{�7𙨫/�muNd�"�P{��^u�~P�{ڤ�lc�t�� =݈��od�'�U\��*�^`X@1�y����Wl�>�m���T��6��I �O�J����`c̸�y�]�#���1uĭ�>]��h�	=;I*�l���Wş��pY~�~I�L��a�������Sv�z��!ե=�f.��9��ϸO=4{-n�>�]���=+��Kg(��� 6��`#'\�����\�ʽuA� J�;�ϖ��v{�C\�Z���t.��<vFg�Ȳ���!
\�4�S;~���ۯ3�๛��r�*Rٳ���\{�}+���ZԬT� B#@D�!2湤+6|�}D}^������q=�|��]y��{~e����M5�[�\�v��7�V��l2��Vϟ��֥d��$��Z���	� ��WF�^w�,�[��k�ga�R�ç�4+h$`򘀙|e��g�_�����r�x�����q���g,���W&5<3v�?�x��x��޽��>�o�4���3��m���ֱn��6�U��ױ.����xχKv���%��\y!��m������Ш��*�p���$���3^���=mz�� 0�<�Ƥ��4d��:��� ��!��S�1���w f�m�8���;�	xn!�z��8)C�`�=8�Y�9h`lk�����D�{�| ��G�)���pm]�m;X�I���T[��jeKa�����H�j{h�n�IwҔV������|%Y�����e��ꏭ��!�!�C{ m�ࡕ����(C`G8o��Iq!w:�7�9��-7�;ng,G�^�����E��:�UC�<?Kܶ������`��
>�
z�fB�N�'�1%C�D����M��ݨ/�1��C7���L���ǋ{Z��}����������g�ط=��~���7qn3o"(h�N�9���S>�9k�m�2�.�wm'F��;�ʾ.�?u�avw��]��,�*�y�3�`�x�$z��-�D��j��OY ���e$I@iILL�R���e8��5��W�'S��lȖ�>��9����)'Ux'.�\�5qܒV.�>y<ً���5}�[y���ڨ�V��_�7����Ѽ����r��"��g��6
;���ݰ�xU{�[jz�Zv�5c���+%.{�1���S���#t�{��3xѬ�*3��`���e���m�6���}�;p3Q������Oe���X5�p��W/��e����+��X4��$:&]�1mj��>�Ձ�R"6�0�pnu<	�K�oYi��8k-�2���q�m;��� � @�W��3��H���/�����fP\���/��z�
��?��=&�"p���`�+KΙ-f��S9�`[�٬��f6����;�y�ˉ��@C�B
�
'1���2��`�b�c��|O&�/v(�1T��*��~�@��K�ե5�wu?-J��ZB{��]�:�����B�6���~�MC66�?:�je�U-�V1C�Q�n>ܧ�E��:l�]	O��>��|�:�8o�Qp�_�}�[��v�"��_���FB?v�a��F�sҦuv��1}��´/����m,ړoyyű�8H=��q(Fc%:�ݍ��?.��J��y��m�S��mS�2��n`Sﴵ�j>,�v�]94©�<q,�.wcK�z��s�:ؔ��s�f�����b~m~<����c��a��kZ��:b��ɉ����pR�}V��N���nYT�5549�͵�$�*�9&3w�#��|��viy7i�8$VC:hp^ǥIn��DX;�F��rK`^�P�9���,6���+mr��8�SL��D��ק<�S��q���p|��l&��Þƞ����ay�p�4�^���WZ}T�:U��E�g_����v�;_F~�ìp���-�w<�n�m;�X��y�h��7}��+t&_ނ�"c@����5	(p1�M��9�	&�D����ӑkB���-���e��>��_&`������H��=���۔w�K}c�-~�7��/�=ɥ����^}w�ҟ�ʟ�<�����Cy��`��>,�F���
�X�@�m�	ȪC������Տ>õ�A�J���9��VG\S�o+S��nW	2ر�y;NX>ɟ*�N�c} OQ>:��ʉMS�7��e��?$`��k	g?!X����X�!	��R��'I�� �;�JcŒ�);�&��w{o���q�B���c�/�.�Z���x���Wz��.3��a������S?&�ڮ�y�׼��u�zw�k�/�w}O�R�c�ߢQ��N=���čS��Oå8����:Bu=���2"�z/����y�贆&�\	7���ڗw����]���D�����l�mӿfN�,+C|���K�/���*��wy�Bq.r�I�R���<�G*<)^���=(�1��K˯�$�L}�)F:G�����E�|SP�-纯ͤS~��kW�x�������@)����+(L���[�*a���^��5�Ď��JQޜ@|��������o�݉$�ލ��i�A5��u]����u>���蓏@}��u�$`1�=I�{�c{��$[�X*zGM��	�[V����M�u�� w��X��Ή��,�N(ؤ1��Ǵ`"��j$Q���T9�GqV��D��$MJ�<�G?M��P�W�35_5������{p��L���O��2�Ws����G0�Mm�1w9[���713!bF9�s���ӭ�M��c�~g�j̕��c���Dw:���$1�V����/&�1�E�X�\5.ג�t�'�i���;۫H�[b㴩�E��+w%4�����+F6�Q7��@	��,����V�Χ!��Fï��Ü<������Z�T����~�~��^ �)��yH
i̯�:zǭ�iЗ��w ��=b�j|��W���~��ZЗ�B6�&^�<���_'�1��`�mxJvǩu�@�x��� ����T�DO��	)���#l��ue<�ڑ�(�m�A嫤C��n�M�c0c+�Tù{�b���m#���+���`�b�P�F��}8\�p���.�/�f��hĜ�v�L��&o7A^6��ʒ�1Ҧ�� e�b�,��4_0���.�p��ɤƟ,z�Ő\�Y�Ɋ�(h�E�GQr=�pd+����M���ڬ̹M�����_�Եd�J<�$'�pE�WZ�b�z��IH�#�z�#^<�u��K|�oJ��������oɰ�x{�>��=_���jR^���$f�����=��xW��!o�8�'�=�2���
m�dZ��Ϭ�#��-�g�5��!<���dp�^{܎$ �}����ک��o{x��7�j�3+7�f�mn9r��@�#����X��Hb6p�F�+qNTlD%���p2�q�'����E�!�!�(�{0 ?���%+��a>L�;�vh��D�vh��ׇ~'1��+΄rz���9�qw���nh�ʉ30�g�_��dv�РG�	��yS�����Y�q,�~D��.n���O����2�+���~�FY�ݔ�V����v;��Lߦ�S�����qj�q���H���KN�;���#���w�[K�	�`�h�S��%�@M�U{�2�Z��d'�ǱyO��O=4����eM�O=6�1�ݝ�V?��1�/��4[�%.Ud,����O�Ѫ�Ʀ�3���XVƪ��Z�׀�<I7��F����m���������d�=�������nt^ văFdMp`# Uj3�MXrĹ\�놫+�A@|~�{�F����nކ��B��%�s{��5�~�6Z�}
T��<`�}���qMZ>.Np^��9�!<^�+�g�� j��3�ܩ��5�����/������u��k{�1ZM�ё.���� �`;��8� $�|�	�ڮ-�?�m�O��E-Y� �0F��o�-�%	�`r���	��w�^�α��8�i�oR��WV�\�2	��t~��{�(B�=�0�N��p�#W���b�>x��-�.Y%;Ѓb�Ë�m�n� h>'��70I6Dy��_I�^k&C����q�HV��u�ަ$��G�7�u�}��G���Y��!�|�o!�O�Ua`�<k��D#����霓�˔�X_C�!!R�%Ìn�lJ��S��[ҹ��+l~+�̺IXf�[�e�+w��U��O/`�Ol@��.Q4G������0.ntG��!֠�^����f�< uV���ix �X����dQX���A�0-	5aD\�V��h�%Хw\��q����^�p���/y�C���C�QfE�D  @ IDAT��T)���b=�i�1��t6i��U?*������P��~9�1~�c�ԥS�F&*`����tdd���~jyF���۪��16_�jp����׿���v���F+�������C�?�;������+;v�*_Ƒg{|�⊿5��Lka�ڻ��y�R�Ѕv1Mԍzq[�4�O-�sKƗ��_Wǟ��=�Gv���f�$���3�Z��ے��G�\E�$�����-�,V�3��Z��2�=���gQ�:^��ˑ�hpdb�|^Q��YMcj��J�ḵC9�<Bd$7�Q$o��:�/,������=�,dp]���V;cD�ד���B�11��c>&�l!�,溃H�M��y��/-x�;l�y}59��Ѧ<p��7:���}H�u�>��U�9�B~��_�vi��|p��~}P����N?�w�N�ߊ\_���e�Ё4�:�n닃Ёn��7�
�n��	W�r��Q.[�ì<�`����Y$��L��>���./M�E��2u^)A&�����k���EH�����N�8�1�S:�����h����f���s�xP�o��/�s�=;���DN��C�1�Z�eW�} p��D�M3�sr��:m���g뮎.�4mJٱS�1��q)N>�Z_�&�SD�i���ei�WĨ2������Gm�C=�%ch{�ڝ�E�$�O���3%t�;Icx��n�k�*��Zl�6ᕪ�񷪆ZD��XtT�R�2�3^O�>����:�7�)ʟ� ���UP���u��؞�@���n��1~L]+FQ�9��]��q����k�U�I��u\ƿ]����m���Ў܁[����O}���k G�xۏ��c�C.�Y�B�=�ʔ⌧�w9�����?���Qa��;q=6O=��;������i�?N����
��%�P����\C<\F�z�-/?�{��e�\C<K<�N�y^��Ÿ6���y��-_��B�=���v��՝'I6�T��c�o3Z��!S��V:Y]�a���(���G4����t5G_�M�>��y�ce�|m֧O�����p5�~���u`�pmЦ�L�[r `���ج � �-Z�Ng�'r�F
lx�mR�'����W���K���[W�E�]�C�	��Г�������g���sF��T${[Y�_��i�Z;�Mcc�JQa�X�h�J��$�����<��u���	�$�i
�\Y��w�$��y��d������d��2dK�ZU�Z���b�O|��+-�Цv�B�nʪ#���˵�z�`!9"	25�4�;~���.�M�
�y�*}mV.~+~���y�T��F)p �-�2�~�� E_�d<%W�Y���	�lÖ���C'�����!/mm��BJC+b*�8-�_~����_p�i5VFgAٍ7�Ľm�Y�� �E�h���r�ʊ��Qi���j��!X3M=�mRO,���D��$����1Oj��ًo,9�э�@e�\1}���i���C3���!�R��nXA�1)9,x�q�(p��^e�Z��lUٛyj��G���Io\�I��E7�Ӟ�R�C>a'T��-&@'b�}�9q�dx�}���Z+�m��,���>�R[�hl+�"�%�O�����]	<��?�o	[��B�EWs+��U��D[cY�tC[/���Q�����鵣g�_m{��[�~��o?޿�ݙ�o��+7��ᖋ̫ׯo�����Ϟ��>�E5�}p�TH�c�e'�R��f����4S����g�8\�߾��s�vV� �o��:���8z9��$}���I� �d�9	� ��E�&a�&p�M}��J��ҏ'��u��2y]�R�<�h�J���f�b�BF��Z�X�-w�&_��"!o�Ũ��s͌��9ω���o���D��`��[���]��r��(���qH�	7�,S�N� 5��&�r�o��t���(�!�I]�cD��Z�~{�����d�
#��4��F��; ���h���R�kG�Ýpm�?vi�Dꁓ��~}o�U���k��:����?������1���w�����ߔ"����]On�2/�������5����6ir�]��v�[?�HʕOiF�2�E9�����%
�#i�+k��G��R�+>sMq�7Q�#'v;��6(�Òm���t��������_ɗFĎ�16.��˅F�rF0�گ�p"[�zK�&z2%�"]Yÿvة$�u�Aⱐ:U���"�+6ۢ�-��L���2rC�×X%��*y��}�vn}!����-�e?�y=�<���6V�W���Pׯ�h<%Y�V������9���R��p/��o�s�.��5Ih_�i�j�R�fȨs\2����D^h�a�����Ƭ�W�l�V���^%��J}�;_�`9�h�0�3��u����*DBb��=2+X2�T�A,��9��>"�����0��z,���|u�Ǫ	U�G����^� y.Y�Z9 �eu�;�/8G�0c��=/%��o����o���Y����O7_?�?o����p[��;s���[�y�a9mh��sN9���A�G�+�^���6�k]��^���m�E���3#�sJO|�O|������Sg<vL@glb�<+t:)ҵn[�!��L�.J�k��)��pr�u�L�L�nY9���\���k�<&�lW�|[�_HJ�몥y	���4�k��y�����AV�n�[�+_���|�Yy��uLY+0$ ���=8��goY��Gc��^`�:|z��E�%�5�tԀ�l�$��u&a�k@�=>�G�(��&a�U6jVj�z��nOw�ʌ���@R�x���	]XPϳ��~2;���o�a�����O7o��͏��{ws������o������{י]c�b�ȡΏ�ה�B˲����7v��޹��&��lh��'|�R���L]�����މ٘?F��`��M�6"�i_՝� �PN��C��+AG�m�:�5| ��m^#�:'�̋PV@�K'��YZ��d��>;�r5bJ::0��/�8���ʛ���)��F(��a=a'g��.#�X�A����8�Gc)}�
�O��u�?�<���\�_Ҟ8N�m]���yL���	�����'e}�\����0��yl4=省�"N���]�ԫ�<��¯j|��>�cC����0F����t�]��]1Z>JV����f�k��<-���䌼�>����
��F�sE�G�C�@�?�-�&<��`�O^r|�7��Yy��o�C����~�V�˛Oo�u��'�f����|1zW��s=�<�_�����ߣ�}���e��P�:MX�X�k �jg!��Ny��;u��CB�����J��͹���F�4���FiFoe����f�:���E���k+��k&��Mf�&O!�l�� �t�5�D�r��$&	�_���{���G��%�j�N����ݺ����fu��T���\�u/P��ؒ$\���d� ܝ{�����%qB"4�.%��JQs�V'�V3��X��hO@��&'�gc���E����ɦ~Pk�5��Ձ�}->�u˯��Z�oo����n��?��@�J�/���q��_���7�@r����0?�i�"��������V�����R�"\&S�ׄ��.���wƎ������w�����d�ԫ��t�[�˿�HU��t �QD_�����i��!�A(�|ِ>z�Mj�1K��n��/Hv�����G����W>�v��/4{e�_���l��6��P~�K�&w�`�X}8M�#Ov�K�ˏIZ?��ZՐ&�����)�,�]�7���\��X-�mڜ��Q���4��2���^C�`E�c[ɉ��t��OL�ch#ܘhsc��96N�G���%���`G=�Y�8f�Ί#FyaV��U�%�귎�Ӷo�V3v_���W!����]�˴�<�o=�	�,��P�o�c�VT<����|ͷ��ɞ���9wP~���o_�����ׯy������-/Y�/���ɷЖ;Xs9s!_Ch{��6��m�o�Q�X�I�z4R���9�i:�KY*���6�wW��i����,>�I�F.4�#_a����dс�Uyə�3V?s-��;�w���|� ����s�4yo�
p�v�˥Inf#�F�oyX-�]]��
S3���?jA�b��Q��ek�b-���Mwb��	�b��\&}l�OquO[��S��I]IʐRv=;�FwI�5r�:P.X�a��[hI�g�����6�4̊_po�_q�����O����<��`s_?���>T��;3k�T�ð�ׄU���֠���k`'}�>y��'F{N��[�;������N
�BU���P?��H��XI!�}�n~��2�22T1�*���1ȷj��xe���O������n�&��Uz��.��@�b�0�.M$�=���.ťH�����I�sͳ��.\ k-�f-[R0�V���/�	-�RO{q�X�N����!�ktD��9HcF�ŕnN�x��ë�eӡb��;��gp'_�2�-��Ŕ9䟼;��G��nȃ���������;$tl�اX-�hO�L�9>�ơ%b�ң���)!Ep�W^E8& 騻1ΫZ�S��{y�^�ҫ�G���hWX0��=*����7�������;�tL�|��?-h���y�'�I�g��績��w���5�C6xt������{�� �6�T�BR�#]mY�(]0�O���:���L΅5e�	�����,��C�0��V���oq��o]�"�qf���/�?���w/��'�n>,�,����&����j"4o��`ȅ�l8�fc��4�\E�b_�:�<���§
72T
�2t�W�R�ؗ�ɶ6�5 z�{���[¯�C��Vm��U��F|[�(�+(~k$���`}�r��_�V~��υ�ۈ�yP��o��y��O7�9�~��w7��_�����Y6���[�����r�-���	�����%.��l�*d�{p�Ӷ:����o��2w���sR�6���_�5���E��w2H"	�c.�B���w�=�'d��t>E��,��9��|��~�)��J��'�Je�ƎT��BGJ�iG?5	���=���3NE�>�� RT�	n�(l�t���@��ӊ�ܶX�CQ
a[U�Cx䏒5I����R�⢜�����$I�;�2K[J��v����a>��s�;thjHǳ�Gګ}���9��zK]������%d8����[g�îx^Iϖ��@V�����!"�Z�&an�	I4�*�j���*Ǯ�F�H��z�Թ����ܴ�9�_��ЕL����5�c��0�6.�UWƼpM�n�o��r��k6�V��u���!�k�I��x{iJ|B��q�݅���֏�_������/B:�=���`����4��74�u�Zm����b'2K.�=0�#ϊ?ڑ��y��`3�]�^|3�9����!t�J����C)UYh���U��ZI��Ļ�x��{^�OM�f)�����  4�r@�ի��
A���72���d�d�Ĵ:p�մp![�*y����36ȝ6<��r�#�������^�<	�I$\��.����g,���[���۽�C�a��t�?ː|��8y�-.�B�f�$���_W�Ͳ���GL��~�,K���$������d�0;�N�`;��CE�VXzɽ�>�$
�C��TK�+~ ��$V�'��s���{���!0$�`����ǰ�
p�!(if<䰸?lIg���'�"<|�t��}-X:��_�-)�8�ퟸb)�*'�
4�k�l��ݒ�~卯���X��4��E�/�����H��4�B�`Y6�>�����.�#3����N��o��^	{y�y!g$2�d<*��ڮ���*��6V��R��q�Z��z4����IH|�8ˉ�`�T�� m����m<Tw)u��> W����+]�Y�ߣ��hS異ӎ��6ܹ(��ײ��x��{����W��3��{�d���˯ӓx��|>J_rs-���]�e\Po��o��gsF�Un�[�Y���:;��@J�1!	�;㑾s	��݂3��|���)Әz�Ԁ�����"$�9>@Hpo���k�s���۸�Bh0$��D�[�J6�>���5�P���3�9^;a�	H���_m��GK	%��i-�t�T��񁫧�G�,5�*e5�җ��1�:x�H^�K^`3�����C��؆R�]YD�����FG@Q�j�	�[����9�m�O���	f��b<~|����-N�Gɏ?����'~���~M���zo{�e�2��һ%N��-��76��B�\1�ኒ:rA�N�A�tNZʳ����v�����P}���{�9&�r}8�J��f�צ_��?|
3�2{��ϹM[љeh\����HR��+�z���^��Kvv��� 0�)K�e�z�w��trFsw��Y�Ц�zy�/Hʣ�R|QIʉ��Ն��>�
��N��ث��_�
o0+�I��/�S�̩��P����m����R�2.���Ա���/��D_��rƇ����_.�_3-��B����a����XR�0\���!ҹ�D8�����mIr�uз1t�Z���1x�[@��Wt<����8>3�h~ c�z<�f����F��w]z����\C���˯��y����O���#�l�J�=����3�H3����69S��mǫ�y,�,��2�_��m��6���P���:�=�%�s]k`�d�\4���xa9�D�<!%���l� ����>
cl��6x}��/�Q��S�$:WV#���#�5B/�T��E?�_����tq8�*C{:<�r� �?��nY� ��X������f,���Q�99ѓѿ ���6�H`V�$OYT赥(}<Ћ&�����B<M٧���EW1N\�s�p�#��ׇ%_�t�н�����|byO�e��w<��R<<��zii�,�',cvq�9��7��]�m�\j;	���_����+�1?
�x=4��J��=*�v_ȥ]�2dAщ�r�4c�;��v����THv 2�B1���U���ܞ }�f� oȵ��b�HhbU�����Z]�pnRl��U�)�W���&fh����,��F�������R�+�����K�џ��TZ�O��:�׻�# �>eIw��e�䩶bB�nt��i�&����yO����S�hѾǠ�N��Sh��C��Y�؂.y�6q��!���ꑺ[����'��q��G�vc���sY���׋�zܦ�j?�I�\��r���e�+/ Ѻ{�����oo^"�#���Y�[^�<߾�g���k	�R�;
��7Fڛ3�:�ie�R}�I��X�	��{.TF �.�d��Ҟ��#�n6m�&BJ�@�tc�b_���DPxM���)y,:8�C��&�Ҵ�w?|[C�hKU�ӆ//� �&��[��.2����M�nn?�(,���b٭�R�%po��ݖ�r;ӄa�_�d�g�T�&AQ֒�t�&�,-.�3��;�T���@��P0�%�!$4z�j��ʖ+��pGO���>��j/�Aׯ,k3+(�G����������9��6�t���������|���ӌ���H��G�;:�Pb�����ډgSc|쒗mo�5� گ\�"����Nb�ӣ;eTΣ��KCo�K��GROZ ՒA�V}����0�����	 
n5Н�_�J_��<�Bz0���%Pxڵcl,xⷓ3{��#����7(�x�ByF�X�{�؀�x��Gn�Y��>w�O-~�R�[�4�|������o�K��T��<b��-���m�$�t���:�*O\�ieM��_==ϕ�}���0Cdl^2V�J��P:i�E��m��h-��V܁G���!��s�D�]1�䈜����T���Nd���8�y����5�b�w���5-��{�_>õ>UG�����eڽ"����_O�� �)�����4߳�n^��_n��x����8&`^K>z-��}V���rN��jG=6�w�b��@]���#�ϼ��L��ִ<᫕���h�NtV~�Rڇ�;�k���}�%-ϸ�/`7~p	ps�C�>���%}*H���&�1��Pߦ�<�KͨU2�͏]s�1/\%������%W�e+���& f񱖺������P'(�`�P"�`n�a��]֥[hS�HV��ͬ;����������c�N!B�Vn�>��X�kr�Ƿܣ�� |��K����O-_��~�������8?r�(���܆��u�eu��-�t�,s��84�(�1:A��ˋ���'c�V����ǀ�3�7�c�D�?�ӆ�#w��Os��s1!��x'��
����S��;f�  �~�Ϙ�L��#;����J���G��[�K@�ݨ�IIyGqL24�O��,�P7%��a(z:���{�-��DL��C��\����UwEվ.;*7��Sj��e�W[�d��.��vm7���t�_~F~m�9((n��x�T�jS�j(����eq��B��@���l���ј�W�A���|n��f��eC���n���y��@(r�4-U��<�
qqQ�@ [Ү�`0,"�|�O�ڿ�6~��-E�~�tt��#z����S�-�?��� �M-��Es��)�<f���p��g^��ùo�w��;'�<���00�3`\Kh�!�C>��Z�Q�����w�-ĩ��u�Ѯ/�c����]�i�O܂,�]�h�F%RR�Lmgڍ����2ܯ��6y�5j��7��4�k� m9W#�]oI
9�l�Y]
X� ��k( �Lΐ�a&I��r�;�Y��˔������e�GIS���u��6M��U�=�ҤLz��SW�UC�@�4xq^�ĺ��<f�(j�����n=��kVňI�����A��]�ӍG��ཀ~0���/4��ۯ��Qo7z ���- �ɠ�s�&<6�r�Q�o|�3:d9�J�c���/Q��z��/b�Y�B�V������W�#�2̏�7�țzC͌Wl�dT����2�sR��W� ���6��v��/�Evѭp�0?�8>yCs�O�C,�������QǧI�X�K�юNd&n�%F���O���}#O��cR@E-dI��1�!�����~�V��'�/�c�(�7v�;u�ʉ_���"��_�$�x +~�:v��}(���Ѹ:� ��=���A�G�����2 �p�C  ��ι���9K�C�ܔ��m|�����"�A!�j�l/z��u���,�a�_v#��@��	?N�V�J�x�o����y�K�i�)[��p-���6���[Q��W�v(C�����<d�S��m��O��p���wP�(z=f��=�˳�^<E�?�G�����z}��_�a��|^;g#���x۱O����&03�풁��g{�O^�(�M+�F$��D����z���U�� �Ms�np�a�r�-p����(��m��I�]�K��z�_E$��1W �f ��*��<��M�1��	���WYy�����u�Ր�v�a���d���Q%���%��I�aO]�5�EV��*]�I�«\-Q��^�Y��,��O�罨G�>�W;
_�4��-���O-�^*l�QXb_0&|�n���m�P�6�#�����7���E> y�Z�H:z��fK�e�1 i�5>��Z�P^�8:����̗��{�7i�v�n �CL �$�fl�D.�s��C��>�z%/�)�"NJ3s� �6������	�eW´���b�Ъ!���=�r�q��מ�s��GG�`�8����o���@43����DyEEi�����. tb�@�T#��Q����U�yDE�d4̡]h+l��qk���iYy��j+wm���6��!tft(�]ʴ1�cS�ذ������6�.�*�/��Vsfd�#����.u+\"=��y �٩&���Tޘ���ꩆ82~��lǄe�B<��T��[��w�Ey��۸B�&慝Ȉh���<{�a��[ʷ��e� 7�[�z�qCC�@��U����[�����Z\��������|dr%��}��u�k��s&�5[Щ����)mז�C�*�e~���C��\΀�VM���<���˳���Q��,��ӫ<����>��\P =&"'�v_���S{L(c�]>��.'d����K`�$`�֟����o(���$�ַ|�M
6�;_�$Q�׿�e�l�s����+��\�[C��EV�P��ڊ��0�J�_uā�{�"��:(�5��:�Bs蕸p������]x�ז�Ԃ���R��Y�͍��em@�� ���3����率�3nP"����Zu���E�:!��˝���G�q����_�c{���E�89Ú���l�V,6�Gu��'��";�;�p8���MK^�ĺϾ���:�EW��결�E�l�à8F�˱bc��߿hN;F����=K?��G�";W���q)�LI��^E��c]t�gwEWCjmefE+� +�B����#��$v�kbdS���9|�z�
]�B������a�����n��(��Kwlz<���J,wlO�:�H����9\�"|�0I"/t�[���d�\�g΍��ً��]'���ۊ��ˉy�9������XH\CLǵ�b��?������-5����xZ���������M���[��wS�̅]�2Jxl�f�v�e���h����=//yN��wi���A¥;V?���!t����M�r�b5,��RFC%�A9 |l�X�����Leԑ�,����Wꒃ�ȜZ|�(K�\�<U"{έ������ΝԂ�qF������Y��!~�dZJ"�;Ċ����3.F��s���]_Z��G��D^�QN�뀙-� �X�"%��_q�,Wj�d�[cCz�"bY���/ �����`Ac�&he��ړe&F�*�r��T��&�z�EVV�¦���r�X��r��mLW�k����tŦ]��*J��M\!rlz1�#�I�	��=y�
�׆
T�>L��
】��
vKС��LL,��(��Q=�1ֻ��o�����ʚ��N���_�Ǿ���
.��8~p=�H�j�\��~p�䕤2ʗ}�,x�ʪ<etsn- �����8V�� )��<�.�ұ�0zѦ۝��2�ֲ�@�QI��"�4�a�E�8�mq�W:ن���JOo�a��Pe����E�ɀz(N"ˌ�J���[q����~xĴc'����Y���\�x���>J�>4�ZڛpW@t�Y)O���Ws>�:���cst/[�e�q� ������[�M\�}�ܲ����9�u*s�c'�1,e�:��#1���Z`�R��i���x�9���<���� �Ҷ��0r�k?Ub#���yw������&Mɍ����iK�q�n�U�ۀ>�Rޑ{�AN{] ��/_��*O���!X�[�%�X���]�v�'b�*@yn�(֤����wFd����!���O��;�9�,T�7�ڏn嚄�P�w
�>���o�*s����\�}��OI�\���"Wd"���s+c�x�n�a��Pq�oUڏu��^ݜ,�O1^l,:�����R�mR� �	{k�va�3i0�'����R �������(�.�{e����>*0NJ0t���f�������g���z���g��3`�����3W�|(��O��:wL�f��H-�8�lb�l�A$�HH���:YG���|�~��h���Ȋȇ�M�����BN�;�' ��;3�Z��"�Ǵ�=ji�
��SE���]�h��p���o��S�QE4�W[9����'q<ǘ=9h�4�R�E�Zz>����R[R/V���'�Y�y�,��s��*�G�:&�/�|�{�H�e���]x��y/+�OB6�SDE�G�SШ�uby��Z3��P��`\T�)��g����JA�NDte7e5�v/�����Ľ;$�����9��Ωs��Ո>�+��:�#���!O��?>���͎����6�a�t9��H"Pʒ��6�浪�����ǼX�:��wi����s�kæDgzp�6ʖ�Ϯd;�Hq�L�|?g/E�Y0���L=��*瞎8�+�x�Kl���3��+=�Q�JNW���Ԧ���5d(�b\B�vT�g�&"׆����Ⅹ�z����c�zu�h3x��k��Ԟ�{~�4+8�R;�;2�����g�X7J<8�����V��sW�a���2l��z�䎞�b�1yd2���bm�εcwLGئ8���A��/���K�`�!0�Q��� �XȒ�2+�}��В���K`k�G�#�*�@v�"���E��^2��<��Rٖ(�Y��S�}V�b�S8��r�7���Ռ�@��;��-��ZT�.1�.�Z���Z}��Eǉ+��9&��~�!��;����z�
�E���5����W�bK�GnE�-n���>t����S1-q�%&r��'>(�ǌȷ���hZ��m�_�"2��jøK?�B�Ieq�����-]Yu�"�����o�]��^�K�0�R���|ZXS
�y-��x-�1Wb����[BLm��0��/�L7~��W��,t|e���-�u����5t����Y������F�R0-b��C^��X�ȓ���e�V5�N��R�q�1�d�樂f�/�4�����z%��$2��]~�=2
Ou���H�`��N�|.l�V�ȡw�v)l�����b�ah�K� o}Y���b��F��t0��F���4oi���.бkt/)ĸ8s	��&a	��@��hn7&���u<��|�Z~��E�������Q������B7��DpX/	����a�����w�غK_3w��"�T��U�dG�fL�!ֶ���Rg�sN����+&�m�ܘۤ��� �ؐ��|q
�9� �0�Y2�~"���O&���p��\���tS���!��hu�"RZ�!��W7�d�&�+?.�&� �,;�h[j��tL@��7;�B�
�<��tL�Y�=���������ޱ����<��F@aʴTF���Hzm6�E��q�cgn5��)�>}$��!WzN�p����[G���Q![;$�:^؝,�z�ꈐ� @������Q�>H �Bc;%ʖ΁]�
�Q@�8�.�BX�^*�尖����fc"��7iT'Kآ"���(Ɣ�[��f���l���/�c��/MļYub�
�c凉%�=6���eB"wtD�=p �[�Q˛�g�T%_�O#!�;�x��F�'^�����1c���fL�qu�ze�z� #�ȴ��N�l�&�xHkrB���0�cf�F���{0��?Ys�I]�	��{���ӺI���{��FE�.���'�ɘ�l���$�*�C{rYG�V��î�b�P,"!���`������K�� ,Q��jOlnQ����l,^r��:Q@���]�޵�yw��J��PV3�����
�,8��s�[h*��bg��i���w�5��	
D�P������Z*����(j��`�-�5F6ѐ�B?�
�]e��]h���g��� ����1�MI�2oSQi�.���	Q�}���M����=����%�p���:s	�Lal�Wb�mr�/4�࠿�UX��u
�	�A�2u������b7��M	�vU���Y*A��8�H�z���]|I��羹 H����I�������)*�Oy#�F����(A��~'�G� �:l��D�k_y�����,�ٍ\�m+�@HL��ht@�;9)p�������i��@�y5a��'�=a�2˖��X���`�Z{�	�*��[|&
ԑ(��O�ʖ��t�b�{�ڦ�#+$(�f��@�'[����J4n���f�%��aL��%��E���I�!Y4=8� �����t�豳�K��1^�un�,�ĕս��Ki�����[ 6��Y������s�[����$���q���fE$&n���	(��C�MF7�	a�:cU"s�]�����c5C�[H�jFe�~��	��iO<�, ��V}�=��aMW���^ɐ\>,qr�T6�!R~���cm�^P�I�E/jr�ò�`)�i2������C�<#,
�9i��B���ǿ�� K����|����n��9��k"��%���8U�rkǪb��� �����0�C�^A�O�μX�S��I>6D���:F��p'n�Kie8��~�\O�ܹ��1$ˤwݎkg�@k��Z׷˱lhe�ŇV��KM>�OQƺ���)��v�f�gB�4��Y��)t�W��*gO�ǌo�Ր�/��G�`w���k��.�h�O�'�������{�&_���qV)���Wq�����y)��A��6jC�٢�!;�J�xuꙷ,a"����<�<�6��ߏ�~�y��g���[�\�{<�v�������!��IȞ�:
�y���{p�q?Y�/��tgh�D��P���ǯU&|h�`�ҪE�\������Gl��AG�>�Η�;���A�^?��ܔ�Q�i��m��"v�i��	r�w�F]�OK[���rۥ��aYt����T�,g<sg��~�t�e�9ρ91��E���R{t�~�l4M��F@&�![VJ.���.���]��Y����Q��G�_j���klt��*�e�2�JӸ5�.^/E���>�fJ��W�}E+�<�����1�Α$�9F�/3Ig
G��p\c��&�E�v߳:j�3v�C�˿ew����4�V�����v`ֳ�O�D�c)"��ѕY
�gZJ�?�w�H��H�B&��y̲��y�ӟD�A��r���<�`̡��Պ�g�]F�<=���/q�>���g��T�;�F-��(�-���AV^W{��7��EV�,qD/��;�J�Ly�����~�n�6�r��l���EFϱ�{�Y��'s�0�v��]ٍ���h�:�˿Ԣ��96�\�i#H���ǘ;��L��s��Ǐ�}:+=��,%*cdWO�l��r��}�����Q�_�16�O�o�g���K��U��^�}P����qz�I��#G�]O{R��
QN�z~)�{�fXVm��yt��֒}������\˵M�h�X�濘��1�C�?�&]�[=�:Go�����Ӯ�V!姭Ψ�}��{��	�w�ADiCJ��w���mf�����0�6�ӫ;~��o�PW�6l�'oz�{>�z��
����<�L�J@��h^�Y3L������Ƿ7��	�������x�<G����D!����d�*��/�z)1�psR��|6c�'|��p��� ��zB�2�Y��6Ґ*�[��x�I���	��PBڮ$92y�F��\'F��Ȇx�{Y��4�VWD_��ZpíOS�n�(E,��Mߍ1��k|�r�m�6���!c�r�q8�U��C'�>��_�D6�>J7��Dӹ��)ó��qX���ԡ�&��F�!ι9c-6��==��(��OT�����$_������àz��޶sQq�u�@�s� �/`i�G�˱��k��Z�شZtT%H�ֻ�H�-n�'a�$%�ա���<n�9��v�Aڇ��Q�,`�w���'R��#]�;ϥ�hl���M9d"���R\,��ƽq��R?��tr$:�? �&�u�PYK�XȤ���V��8��숽���&�ig��.�������Ԟư��$q��S�^F��j��SВ���Q���JC�s��C��Mpb���ڸ"�G@�Z��EIP�K�DZ%���U��,���	n�Ӧ���D��e�yѥ����~Ss�b-�=	laO�kad8>�@�g�w�T1b3� 
ӷ����И�C<���o$�O�l��-r��]C���ݰd��3�`\>�OΡ&GYp�\,s�� έ&3 �O�ј[ b�-	ܭ���#��EO��.��2g���'�snpnj��5��׬�Y��P�uޥ��t��?�t���3�#ex>�y���ޱ����[�/�	]	�������wd��a���~���[Qo����dq��߁��o9�?�ѡ�<����޳:����j�&����vl>���M�D{;���9C�����%�z`�o�  @ IDAT��)��=W~RS������� ��Y��׃XU�����Cl'�c_�� �n�AH��n�g��^��KQJ�"��#Qq�����!�r��3Xi/�k�4^�� ��R�2F ք�h�h�/��C�>������zdN�a}ɧQQ~AؓAA������L��R�}p@�h�R9��7�܆c�6H������(������5i�J>�@�o���c��GV��2]x�]�;o���e����;����44���п�\���K�����O��	p���cG����s~#Z��4�dŊ�<�-�0D�\��~�f��kY���|�x�%�R߱��0�*H>,)�2�!\�=�)���s����r�L��?+5��_���÷������󭱜c"��Ġ6�:(mK��նڿ�Z��7�Vጝ�f��wF��I�a5n����/&�� )��*:� ���9fV����E;�Kr%UWj��wJi�*ͼ� |٤��:mB�c)�fT�mVָ�8%�*w�*���(+����*^��g�PhPۮ�l���8G	:/�n<�M}��ĸ�Os�FF���,�>z��M�p,�.(���y�}��՗^��m+�R6��w�K���F���ZK��c���46gi	��-@P�S�IW�>s�t|����t�
XWȼ�u��폎� ��O'"2��D�g�o�~��&_.2��8���c����	K�2bz�Ķ���~{w�/ٸ(�gf��W7���*yρ���L�}������L��$�$� !������_>�|x��{ŭ�[�@^w�쎗�)Փ�_��ǁ�8�)�ߣr�p˷�L�H�|�,6£�ޚ�ȓj�6 �|{ Y	�$`X�{3Y�|S���-�~8�k'��di�%;�Djڵ�}�)siv�V��-��o=��hd,J$�'��<��:2۶�
�6�KO�hX����ףCH�۾	���)��%�	ߘ*S�I���}��*?'�ŵ�U���kcb[�B-����vw!E��֡j0�jN�'��,�p�~x�����C�+��=�8z���� �2�b%�?�k���ǂ�����Pe�~���]_C���������/�p�E�M|�C��+]�U�a��Cqu[7M�r�s�Gq��N�ؖ�!��bw؜"Ha�?mg�I���`��ɛ�������ؕ ���/�X ;�=WOw,�IR��{d���Yi���wss3sss�#<Zx.��èR�)8�2u��TX/ա�GJ�üS6BEE�hg���3y��%F̊�t:Sq<�&\'��R���ę:<ɟ4U.^�SF����D\�
�Gn��G�I]oWa
gOgP��݋����5q��<��1�<1r�,����8a�á3�l����Gx-Z*���2���"E�x6��`-|<���[:&ə��Ɖ/�Q~�77Sם`ܛQꊱ˻E[�OUe#\�렡a|��t�&�u�#��##��8�s�{҃[�r���1v�.[�׉��ȧ��5�f�A�'���7��F�\4�k��	��ɮGc|b@�ƣ�,*3H9�<��02ӈ��:���dF��M_�3��"�a|�~���ƽ�g�g���ݜ�D�t���ɺڝ�@`�q�����y�^�-�����6��M��o�'�,�^��Xص�a$���%Ӗz���:c����˼dt���E�����e�lc�7�c��哞d�"�N銝�Is$��g��Ae/+�A.;st:�56�a�D�v|fD��z�d�4�i�<��'7��+
(k�	so�C��	��VJ�Ц&	���S����G.2�
�E�H����ki^���D�2zm�E\v�����@�t�@Yq�a"��S>����(8��k
Y�Z��L���c���uJ���uG�����=u6~�Od	&6�JY�E������V�ڡ�����t��5���Lʺ�*�
#!���(>|��8`�YV�� �a�:c ��i�dԏu�����t
츨Cw:"V,�3�WƢd��_��qM���4Q��U&$L�q�w�l�K��61P�V�� �\���pF%�A�D�ʈ��j|ʉg�J��]%Ϧ�AAc�+a:��G�6a0�^��U��h��_)4-���(��W:f�g�P��gg'���7F3���X��hY��,�#�\�
��7%�M�<��&�.y���٫x��s$��_<�~��<ư�8�����ʔǔ�ɍ̵��KF�Ki��c�{=,��,"My�rAy�	i�L��	���|��h*Wa�%��[��[�(�_􂴕?�H,�Ŭ
KP���Oі�/�\��!�!U����;�yH]��<��g�i���uD ��Ǳ5�Oݏ�<vP�n�q�P�������:
q&�����N��a�6KQT��Y�B@z�*٧���C�!ʌ���z�L��Ӵ�O�s�.g���Θ��2[���r*�KM"��t��������U5Z����_<�/�Q��Hyp'빶�A�N�sM���.��ܸ��u�����·Ŝ4.��b-�|��=�)��8��+��e�=S�[4|M}wg���T�j%���FȊc��� ��]�k�a&!�O�hu�������R�J��go0l�z�G �y��	�)+)l�[�ˆ��WB}-t�[���,`@�W�YNVU}���G �}R uW��R�I!x�w�Jo��|��CXAj���m{�@V���)����I�:���:Y��|4�������t=���%9?�����"w�&3��Ɵ5���nr��������V�|�݆�̬���ŋ)(�#��r�[��MN%�#��2�����p�`G_p��|-��e���zx�&�58�Y����EH��݂K��/����C�'䅢W�#�G�k#`�a��()�z��I=�ef�♯`��<�E�o�����Vp�N\�6�P#�p�jO��8m�uP���/�L�:�����ND���q�����G}r��<\�@�p���5�8z�C:�����yH����jX?����rJ\�g�Gp���[��8��O�^�ֿ��g��"�e`Sm:}��"�A*��=|6{K�4bB$�7�xmh�G˚���(E�Mӳt�!�I� W�U�4��Q����铷�｣��{����C��C�;f�
L(����t�����+	��+��i�G��7E0�*\
�z��`�\�ϳ�T��Y�ɑd�8������\�W9B��r`�s1]�h�b�qC�u�2c ��,��c�׆�m�ڥ�崤Z�g�OBWp�Zjjpɯ�Q��m�#m�%�jNٚ��ԥs�UXt0NW���1É�R�S�0u�5'�{�0�8ɬ��~�j�5c��1�����غ��w�+��ԋ���ag�La��⊩I`�Vq��BIA���t�W��8_����	�I4{�� +ͅ�*�0��u$+8�[Q����Pp�6�05��T�Zo��i#��uw�#��3�[�*�W��4!��Z�%�(GWF����&�E�*f~��C\	4�� ��	�",���T�;�4>a��$oPV!�2�.aӄ�ɘ��*a���N��RJZ����H�ȦaA�v����IQ	�t=�>�*D�;�T���1��F	��x�͓�U�hH+<�i:�vT,*w>�M���]�_�b�3����FA#`�x{s[���&=�P�z�t,p�a{s�[2��;�p���"]�6#A�/������hIU����b@u�U,�FUZ�W���Y��A���p�8,�A��k2/J�p�s��>"YKG?��N����r.���0�S������(��=X�W
»ś�y6��]�Y�e,�J#x�o�f��w��Ƚβ2�a�������(9�ɴ�0L��������2/�'ER������vc3�K�J�Ht%zBXV���Z����/�Q�^�\�v��
����Z}��V�V�iFt��f�,�uV:.��9��h��% dJ~q�Y��u�!I�cBm���G^I��U�d��I�������!�b��v}�k��b������:�l��@F����:�(ϑ��3?^s� ��`L��a���9G���kF����J����z�r��L�Ϭ�C�\��ׅC�y�m\�����ӏ��:b+��m����nǞ�ġ�*�t���V�#H@�hq>r�U'�>�N�^�\����들����͂ܑ��Gm���/����I-*�ķ�ѝ3��ҭ-�2\<3��xq]���2GI�EO���i��o(\Л�1<x�0�O$e�o5PflO:^"a��i^y��LQ��XT�,������W�/J����j�X�<S��6�����-����Ϙp��\�o���|�|꨹(����6M��� ��>�9�E��9x�Iɚ&��m��O"�5�c�$=m~p-��L	H4r]�j!K��ypD�Q�!��x/�1ʈvo�"�/���X�cz1=Bߘ�/ݬYh _DU��X�SY���[��hY�:^����+�l�^E旣fT "��-*�C�%
u���B�ŽjܘՏ�,	v�~�g�H4\`��;�ZH&zx�+���������˅�[���L�Y���p��@�]0uo���T�3���Ac��<��3����ˋ�������Z]ZbG���	�V�W��R<Ri^��C>��	�e���hpk��S�z'�8e�|�QTx�B��2�8zo�ڡ�o�'��ް�2��u�GQ�t$3�H�R{�8{Ze蟲�>�
'�`�#��^�����&)�?��ro�T�\�������U35C�a+�0�5�
���7���a�Wu:�"<|I��笼�u���!�*�-��)Np�		.�9a��^e�������s�������H�E%S����j]��G�e�yhb�_��O�E�1��KOc:q=||x��$#��ׇp�Y��Y�J[�C�se"*��K���!8�u��
��Y������W9�yU:��/p?�/#��N�cu�(cwY�÷�-6i����)Gg�̆���x3,�����C-����*=Eͣg���Q�r�O�Ti��цz�>6�i�0���!4�//:��` ��ڗk�����-m>|��2��{��Z<�M6[����`�rC��k=PV���\�#D���*P���t�P�5�
��F�ק�␑x=K �2����bJ���g�Ly�SX�k@�ұ�x��W7,��po6�bb��ap�f4y���4M?��JN>�6���iL�<-�RԮlByT\��0W��qUar+��JqTT'"x����ʉ�ܛg�oR���FT��'μ�+�F��#<&�LZ��A&��[����G��S��Z���;�4�߇�!��_�(��S�ቮ��ou�0;��0��/qN�+����Y]\��^x;��p��K�5��TM�A2=g�,��3��9u�=��]��g���p,����-���a���p�������a��!�
<�;o!F��;~%-�s�G�K^���׏.G�(�z6�p�q���������������<���l�W�>um��!���7��{��ڼ��g�+-XH��D�1Xu�N�d��t��NK�9%(�ـ�74�Q5i�v�����r9lo/���]�f���F�7����}�Ӑ�u��G\׬����6M֚#9�e�"�:l�ϾܠA�BN�p�E�W�.�q�����О?ҁIi��U�����q���:`W������� �㒌L��zCg��q$�9�пjVK������'4t:��6������q�M��{�����x����2L=Qw9jj��8H���:a;�,�͵qN��9u���k�x���22b3#�c�NZTx3�	�orL��̒g�)����ðI<�%In�a�P��4��f�ZZ�r����91̜%�b�Cˣ�]z.���k��$�m{!W���-`�9���I���抮�63o���iI�n�l�YW�o���ݧSz��͹3�9=<���X"�=� ����oڪMH���1oۢW]�:m�^I����%���ҕc��	�/��ɦ���=/c�|��<�U>��''��G:�T IlCTb{C4��� ��9S$��b;�k*�)�)o�룟���LI��D]�:��Jm,������W���p	��K�-�N9^1O�A0؅��1�u%��:����½�������ZR��r�xy�qùA�N������
Տ��u*H�#i������봑u$Z�(��ѫ�ȌR����9�X�LgB�5^�.E�@�h������m��c/������Ȯ���}��S�]W�|�P��F�C�D��t�m�j��
c&�0GS]�U�魰��P�}��4D����l������e3⋬�L����Qtdn��\1"{A�{N�i�]�����pyz>�t�H�c����lxr�;�z�|x��o���C7���z�J�� &���B�Ce��1ޫ7`A��,S�L��av�
G�V�����ߑ����19��y�S�Tk�
ne'>A�\r$_�n5Z�c�l������^��"i��N���'�i42|��[�)2,���Xp�C��vy��X�6����]���M:��C��׌V^�Ϗ�:���c�h����E�W�:#�8r�<6ӗ�p��(�g�s��W�§\�9S���':c���s���QV� ��Do�p��vnW�E��Axט�_�-v��.#b0���q�L'h��*OրZFb�~k��i�ā$���]]��9bA+q�m��:d�e	O�����Gy�!N�p�]�]wu��6F��Ĕc���⤑�iuqD�"�x.�㓙q�Xa�pD��!��;@U�7����aH�+T: &|�|*˖ʇ��3|6�f;[\78bE5�8��q	aJK[;1�h7�R�����=�ɯ~�� �H�t�I��p�#[��aH���K�2�ԣ�s�K��&v`�̀3 :]{8]����;����ptx0��逹I��eP�@&Œ��aZ'lZ��b�[Js�h4��n�Z��[<P�ҹ��������~�A:�]^^>~������&��0�AٯP���B��
�z�䰇ǹEo�ڞ�3y��a��N�R"��շe�"_�鰿�#y��
EV�Uf�>��ZK�y��)������k{�\r=��~z�	�)�^\�p0��b�K�cy��&N�����hÈ�ԝ�^v9b:aR�W�lT����:�<�,� L��T��Lml�M^�#\�Kd;M�W�͹�W㳾G�u��>=�ďʗ�i�u� CkO�߇�������"|pH������cɠ�����M� r��������Q.G�l0����踮���:e9����Ek#�	���%��b�6�l�ً���q����F����8CTJ�;f�����O�_��2���S������م9���;��'�Û�����c: ��kR���/�a�P�b����u]�w9���K��I%.�.1.����9k?���������#����ϑ�2��qݛ�c��K����Jcd�2��MQrk)B�������n�\!��GF���Őw8��f�����0?����`g�Z��<�џ��G�ĵ~Iy�~E>��F.���#L����H،Q|��7 ۤ/�Jfr)<�!�/���Ӻ�fs/�45��r��˧�����6T�O��nrn�Î�ꀩKWvb�c�Q.��^��6@���Ɯ_\�޳)�'�3�+��[�Ѝ>Ful��S~Ҫ2]�j$��T6�H�b��8k'��N��~�o�`2k[io���c����B�eK�X�ƩK�_���?�N�{Y��?y���1��1�L�#w�{t��6�Оz���}�� *����>��	�,�$�|�#��TE%(9�\9�Z
>2��2�Y��_��K;uȵ^�8��7��3�lF���-Ge�<��.��Ϟ�_>���������m��r:��X,2��+uƼW��l�����z�SZ,�����&���F��� ����\3�n�i�H��c�t�}�ԹK�l� |xΈ.��/cQC�1noP���u����a�,v`�9��=z>����Y��-�LaHfr����AIũ������j����`�q:,��jqy�BR�LgNcqE�����/�O�:c8_'g��������	�.}�BsŨֆ
�(�@��~�Xh[���U�:��2*ؘ&�TW���b!v�+�E���*e��
� �\3-i�dPU@#��_�+��"��DV�	��%���`oڑ䍛��	� ���pH�ϡg�m�{��244�c�T�P5_eՕ�M��f�#:_^���_��l��N5�iI;�$�ET�7*�������1J��`T��%Nْ7V|1���N	ݒ_w�6�ӹ��o�χ�S��\Ov��|��.������{�G㹿�9��\�fPki�������rȍ?u��I�bH��!;8��?2󏃇�6��p�p?2pV�0�#�W��8�h��<Ia6�H%uK����6uթ����ã +�{i�*Ov�|v�/:��L��o�ƪ���(b��Ù#yp�c�B)�(���.�d�DƵ�af�S$������+���Uc���e�C^�y0�W��?kQH���i:|��r�]S6w��u�Ĝ���{4Z� l2��h�ۜ��mP'�,L�#W����St{�Qۻ'tl���.n�qr��Z��UYJ6�2��ڜ/��^�!�`�7��[��̆��B��fX?���\�:jjShL�UP����d�@�%V~�ixx���'l�/���\�Q�zgϣ��M�I�	����s]��Ƨ�z_��-U���u}�>@���+���s� �V:����'��0��0���`��=S�m���d��.ڢ�����Ö�/�O�|�}�b����c}��Se�;H���[wU��j��]�q��A�a],��Ö-�^d�ֿt�ïKG�œa툸 ˑ\Nש��0bw8��B'CA���4#z� )#�ˊ�3Y.������o��ްf�9?HIيkrO��:�b`HaJ1���m
I��x��#d"�m"�4��b�����p���)�%�:bV�k��5~�����������?��~8�<'�Q��e�۾cZՆ�7�\g�d�pu�:/P��^��GFS�Ѭ p���$�`�9���|̦�*2S�F��c��p�^ǣp�hJ��N<�>�o$�K����+{9%a�A_�7��ô�ٯ%��=��B+Dm�F�H �C@���]�a�JI嶜. �^f3�moj�i=߸�a���G�t��6�׹�'���d�[�0����q�v����]z;4$8`+�/�3zic��g�����p���܏��BKN�`/�WԱ��9kQ?15yZ�S~�a��%��p�i�éL��v}���1:���¨�G�JR�� M�	S��]�Z�QZ2ſM]]"����&��⅐\̈́�H�0�6D�щ0��U����3tK��`4��=�K'�:���#hnj$�t�-�O�#��l��:M�'�k���g��#�,j�E$�t
gPu4�-�G��s�(W�)�WH�O(���	,x���(��
G��Xj�H,��'������_/��cԀ�:[L�l9�����0IȮ� |�t��͋"(����7L1�sH�%0mv�|2�*o���(#7��#cG���)�[�񓧙�<g]��f���������G0/�ر��l:���>�PXa<O�D�N��|"j���1����5GJ+e8��zTzgL�_��<��|�8���5� �W�\����ga�?�_2�'a�V� �P����V����6�	:໹�:5��Y5RG�w��[֎�l9�����s֓�M�63o�����ۗ���O���=�5�`��⺾��>���5���.k�Sٰ*	�,pH4�5��X�9����8�*�:{�Ħ���M~U� r�Ǣ��Ӗo0��A�Z.���O�_͒d�㔩��::�r�/�E��-v��S;:z6s����$�T�76	q�d�LkzA���f	5�C$VgO朊T8VJB;�Ԃ7�a���cfevM����C���W��SI`��)�����	sŇ{���p�~��#bg�9��N���vF-�Ȑ��<��mԦ-6�:W�"���>&�Ftq\)�o+W��w� 
�#%�?C�A;G�rs���a��c҉��L��'�j�O�`�q\�3A-0w�#�ǘ�gX�c\_`^{��k���2}e5�Ȑ�xX�s+��/P��U0L.��O�WϏ��^=����[1�v�ˊ�}KO[�m�^�m�P7#�� �^�@1��Kp��p�&r�o7��g�)?��� Mj�Q��?�w��k���9� ��?tΨ�~�K��֋0�n��' #ڵ��ҭ�&̪�Un�L����miŚ���� ��� S�w�͒"l���YII�뜪�S�=�W��:a�m�1B���JD���C��B���a���o�Q�|f4��HY_�8'{n����^I�qj�p|GG;4�\x�t�M�=�%j�CF5�!S����N+yb��7bu��sZ��`�s��t�|xK�_���4���IW8$L���,Rv�G	�6�#3
W^�}��9����t�n�B����h�^kW�a��8l�]q��R�,�	y���p@���s� ��M{@�c��?�|��[ ��	F���N�؉?�8�~1<{�rXи�1��O�9��������i��1Vn�i���xԤ�2�UM��FQ�GiS+�1ԛ�EX�i�Є�%J�.�_�x������"��� 	h����K�ò� 3���Y�QI�d�x��$���&�Â3:�ΐ�Ⳃ�-`��e5����{����e�~�������xgtvW���.�}�z�����W�_O��I��HM�2��vZ/Ӎ�VE"M�7�L9%n��Z��tX��ٍ��L�2��q����Af�� l��˘\	K�&^�|�s?Cd�y]�����W��gð��?l9�{�Ȗ;�oѻ�|
ȩ����������=z���.ƛ��2a@I��IgUh� �烒�� �*��e�����@�|]R�Ti� 8C�z�����r�(H�րq=;?M[�(S#@FT�#[��W���}�v��?ҳ���������6�ao��Q�;6�]�#�/w6����#�W�A�UB	�r�4 ��\e轏Uy��I�b�Ucc2��HB0��(=���o$���*ȹͽ�u/���L,�b8�����3��E{�u/nQ�cz��1�+�H�|�`��֨��z�'�U��9��4c(��ct�`a��l|\���~������f��/�oXW��Z���>���7�N?���>a��E���5�"PP����������wi��� �*�|��2���|���85EÒ����4z.���ܮEg��2��0���0լ����ص̼�D�uaP�2U�G�H<Gi�Wr���������\��z��t��3:�0��f��W3Tb���B��-���/���f��z�5�D�Q���M�h����4�yt6�+��k���+��/�<�S����Ʌ��"p��Jr�	��$eC�ɿ�)��q�HqH�t���}��1	�rN��ab�[�>��D4F�Xp(��j?�+S���5*�nhV�����t�<i{-�8��#]:[�4��ٛ�dԉ>���p|�|��?B8n�o�u#e�[�W�8W�R~-��`��aޣq���j-�~�ɻ��aVY�I�-_h�#d��F��CƋߒA�#8�%�}����O�+��PyJ^��$�kݯ�$�yN�_A�n���������ѯ��P����?䛴�!�nA�ɟ isc	u���z�V�3"M������:UTZS�i�չ���퉰�Y�Pg�b�_O��i�;�-�龈l����3�c���W_��ś�뷯�1FX���\ /c��Z���s��=s��y�����et�u�3� ��v�5��_q��9�)E�|Ie��0}�Q+KyfD,i�Md�Igf�R� j*�l)�M���N���34�����aΛ��o-J��_��m?�X����������_3�rL /�R����:�~�jS!U:�*�+�=�Â��F�8�EK岀�Wcd���0
N� 8�F�ȥ4*Z����U1x߉|�2����a�}ggxBE?�u����p@/p�ъ�x����ƹo�O#H��R�rL�&��;*h'�;ZҞF
�	��)Vfu�w���)�,�4���OU<�`U6�%�����`L9�K��%��5H�,b�R��We�zZ��h��Ea�DU�X�
�2{�+�n����d��|�'��Ux˳�V�%�qV���'+��ќFy���Ѱ��A:;�e]�b��z�Ou#�m��`j���^}�.X겙D����Г/�Ew���N�P�3�$뺬�y��������:��F�\�m!�	,1ʩ5��˳	8��Ø�ت�����t�u�#�[/��{�Sp��t�`�*�kt�E��h�ī����.TQ�)?hțS�m2љqJ�Ƽ78����"�&���+D�G.�h;�i��D��ǖTT8��!(�������\�z�9���b�_;��95Q�˿U�d B��#N'W"$�G︝�wFՐ��bb����xt���2�Rթ]ܴa�&�����A�(27?�����\dL�0,�l�����,�w�',����L�C��5ڢ�x����Q
��0���ν��"lo�糖��¼�A�8$�l-5˥4�+I���I�[�����ନG|O[���AF��y�PԓޏniC?}D��l��(;��Jo4����^Va9EXQ<T��ǏZT�Fuz�&� +�~�3(Kց�9r� P�|L$���xo���ˉ^�f�5��n��Fb{���gÿ�����o^O���fꜵ�N7^_Q����Ӟ5��Zq��e�����dԠ��L��I����z3^P�SA�xv�#�bή�.UR�5��9�vY!8�Ui5�6:�]�>��>��J� ��N�E|��Y���!^hJ;������WT0zFG����8岿�ҡi)��e�7�,�x�!@��N @��)\��B/�!�8G�$�ڙ[��@�@����ao�r�PY��r�`��ҩ"μ�d>���ŭ���&���y�G,��~BIò�b�_����|�K������?�������#�kE�z����35Ox�LK��Nw��0���)	���<$>q&����7�Ҧ_5�񠱕?$,����<�	��f��Y�����|�u])'��4&�w?AȽe�ռ���>���������~���>4)����}�$��C�
�T��1V�̃?eb~N9R�1�T��H��.z���]�K�H�6ӊ�������t�������}]�.�p�B�u���<��%�+�S{-�:_���]L�H���.��n�4E�<)�aRZ(�ɶ���y���B��?�+����A^x��X���CH��G�u.��/�GFp�p_��р�'N��_�R�m �.�r��9G��	��Η1��4��ru���-�	��&�ts/m��@�f�3i��13�b5�*�\�_10q	��`��9a�ߧ��[��}Ȍ�䃼�喺��*���r3��A^e�]�Z�{��O�`�bz��|,������鼁TyX��ꬂ�����
3i� F�K�Γ:�EY;��ϊrpz==w;ŌBܰ�?k��=u��/u�)��X�̧숏�K�d���aϻ��f��U�r*pN/�Cr��'9?�0�B�F8e-��W����e������:ڶ�=I� N��Q$6:�P,��s5L~���9�#8�a�F�)'ʰ�>"8� Y�'²���g
�е_��-a�M��#�L��Ί'<����״�~V�7����C}�a�>/������믇߰����}P�\�x]��8:�Ҥ;t͙:���70;;�Kvi8��v3����u�V��7���Xkx�[ Ai|e�����;Y�w蓿�/<o�9���ce�Ea�5��q2�:t^�9�d4��/��?�ﴀ���'��rx��C�J����%�f�.�֍������C�k8��B9��F
�a4�8
dU��7�<2��9�}N'c���2�D�4��RXЬ�q4�ŀnh�(�kn�ҹE����.�e6d� 4g��1���OÇ3F�xS�qH
��ǥ�n��"'�O�Ґ�KoO�JcD�J>�t�Q��2`%&d`� �(�#�ex�SN{�0Co�qfu���D*�x��x��T.r6�0=^M����[��������O�;�Д=�	��^Dx�~�ZoU�!Y*��3Ϣ����&�z�Z�Ę��z�+�J��ܠa���*�5Zy��^�AX�^:m<V��W|��tb�?a�S�xY;���pA������e$Z�  ��)ZF=?��=B�??,u)*Z*^�z����s
W�R1H�pG��T�4���W>e�r�s�+��m�7?%�Ga�GEN�������	<���q$g���'�$�/"3/����#/�I?�љ�n� w�;{P�7�8Qŗԍ�&0G�Bg��w�/yd��ў8�[9���vCõ��>��:25�rC��)�L���7���L�/�(�;o���<�O�S����@���Xyk3y�;�k�wp eĢ�t
C30� XC�zj�)31���ts�%��΄��r�H>]�{�G�O�D^��|�e�u���m�tX5��SR���"1��ţpL�E܎��T����u���D��\Tn�q��
��� թ�u��(�*cd��z�c�)��96��t��n�FT�jx��e83s6�P7o;�kf_���~���[v[8�!gM�itl墚��z�#/|X/���ml��I���GlQ��̞u�kg���O�,)9?��;�Z���Ɔ�� őTN�t�/O���O���0�'��!K�z�����;��-��0|�%3hsF����v��i܁��}�;������e��<M�`���x��8"`o�9Vf11��F�U�>�� X�9�,�[`Ąpj,��I�M���T��p���`=5h��bM(�\���޴S�¹AC`�P/WWx��F$��!I򅗗lp�_���{>�-�.	;GYnp��0.>�d7�����3��m�>����r)E��P��(l=�d��hhJ?����t:�eʬjV%N
mC"���NpI.r쟤b�T�83�|�
!r��[��V\"��|M�Ļ�Г���A?�����Ch�_�&��lDj-a�����JE�zdxyV_w�XIo���R��֊|)ǰ8yg��5����'�q(G;�O�'�%�ʶ��is��'���B��p��Ѳ�5�a0�d5���] w�G=D��A���Q"�n���?G��Ao�����qrWk;Hzw__P��u���G�2�`�I�|�Ӹ��q�0�v�5���ާ�+����;�~�c�|��a~�7[�`����c�H�Ӿ:g� ���V�7ВO�1�'�z�J�:���H�U�����d@�:�%o���ӡ�^q���jڵV�);u�p�>�|���.��y�TJ9��8tT��ﱄ���;�8�l���Ζh��<�:H����V�_#��\!�����]�
0����B:��H��4.�[b(G'�� ��V�������ΪW��=�$M>�uE/9���e��xKy�.��4�)*�t爍��i��T׺���w%��o����i���%��/�4ʿ��t��Y��)o��ZY�	�SR�z@�����	�~�"���#;�)p+� �t�%	�R��A�]�&��d6@�iG��$�K�Ns���b5�xv<�򻯇_��Û7O�=N�(iGl��[�V�|O�ͪs�F��%6�0ۗ��/Э���LwV��C�\��\���l&}�/�w�/��:��W���1B�T�y\:�Lg����1 uP~��~���*h�;G��_��
C��>��1:��u������[z�fV�*:85nT
N*#Cvmآ�¼  @ IDATq��V���e�"��*�^�XwQ�0�� �!p�ܰ^�SJ�zh��`�ס;��捝}o:|'��00>�wb�U.�(,��<n�Gp�=�b�l��Z�a��7�W�^���Iv���O0��Q;̉�p<\Y�Ș^94�bN���5�\�_�{i�}%)N#�<T�8B(��I�#�=�WryᙴV�4��^�<l��h��-J���~�C�v򓴅���"hR=4:�'�׷*�(+�&����S0%� �4�a��@v�����\7���Ȝ�LNqVm�K��SN;:�Q�6���(u�ڍ@B#V�9���6�Ŕ�<�[ ,��������Qyu\���Y/4�'{���Ax	M�3���Ņ.i�T>Z 7+v�g��;��E8�e��ӆ3�4�C�bК��td�X�C(�%��!�M�������2� /�m2�u�Ǝ,��G�1�5b��	�Ҕ�v�mس���z�4��rm����[V�kS�!�>
=o6�T[���&ɓ�o�1������v���M֯й��<��$`����8�%mK:�8vW|�7q���Ơ������C:Rt��e��u��s��R�>m~:#)[P�_�E��{��6`�;�,�NmZ^��"������x�OJ[q��O��]�<9��UǺ^�u�� [����x�^ݯ;:�����[���(�K���pb7�����d�����`�!��5��ږ�v�tv$��ږ �i�<�̶I�T���k�A�p�L?F�F��x�TƏ<�sA�����/g�r�n�~�y���8_������:4�I���up�ѡ�ԁ�2�����ëWoغ�	� Sx�VM{;c���e3T		m�,6�N�%N��u$/ZEX����͎ ga�|�B,�?�0�h�Z/�oy��.K+�u;Z�8]��O�#f��H�Kc�'4n�Ѓ
Z؃��%�!;�朧����X���"8����$N.��ق2���c�v�G�Ʃ���Q0	��}��	��p��c	a�+�H�����@@���9�>}~���U�j�j!5�d�s��cpb<^�(�����<l�W����?��� ;��\0�礑f�������Sv�,��M4D!>"!>�Bݏ���;5��:���4\�����U{�h����,:��N��|��	ݠ������!I��f<��������UxB璵	{���5Ð�a��z����C�P�|��Sh*Fp��� 9-��B�X���Pפ�Q)y���ccS  [cI�BcnB����Y�>��+�'����C"�c��9|�P/��F���WH�9L��`�'#V�ԫ�p��� ;�S/7/qLp���#��EYS�t�{�8�`�F�H��);;_��:<��Ο��.;���L	�&�C ���5�.�(gK��':5�|S�䧨cۨ{�6,����V�F{bc���/���|��յb�m��G��+��E�=�$_�G9�!�:,�!���-+��A�6��X�م�ph�Y��0�>�7��E���Cx�.��؃�&��T�u�r�&:��֪��ٙ�N#�|ltU�3�%�/kì�����EfQآy8���f�)�JZթL�S|)c��:(�:�e%a���ᥢ��r&�A��go����4=���u
S��w
+�i�Ӹ~����Ac�)��r��V��N�
��Tl�n씣V�'�̡9!Zl�����΍i
/�V{h�R�Ȓ���Uo����d�x���@[�T��w���)cѽ�^����g����7߂�u]?d E|��E�oH�5�83/���>{>���&����^�IN��*�T��wCp�f�� y��#^�z�w�
��/�����L����L�2R=�� ��)�H2�W�{�ZG�v񫎟�}{���,贇^Ǵf��(?�� ���%c�$��TŠ9d��x�[`K�G�z�w<;�dE��xù3�p"��j����"#_�'�����v����)Bz6<C�������(�H:͓C��0O��#g�0��P1�Lu�U��d5&?����-<l���L^�N1�l7[�Q9XG"L+k���BC�OA�V�3|�j�ˍ��d�M��A{C!���lq:���B�	��ƅ$Q.�* ����g���0����L��D�a8̏EC�FVc����v>*Q��ݘM��x��"�h�����,��s)��1��ƛ��?�^��ȁ��Tl~�����DX5fⳌ04�w��fer��-��*�PX��HnHm�O�ʸ� Uއ.�L���9Hg�<�"���������řmN�.��D��5�%_�3N����O-]1��6h�E��o/�/ԟ�c�{�\g�Y�^M?,�~�Q�[*�;�iy��k7��hg��F�ih"�l�dFr�l��,A���̺���~ZJ�����FL^�n���P��8�)���cY@_�z.������ �c}�R-և��d�F�<G�ÉZS�hz�nu�m��Yyu=��Ty�M�p���x�]Ǵt���*��h�P~q���t�\ܼ�î��넺�%��I����^�i�t8m ���c~�DTݲ�ԭ�@J�Nah��$+�鯄�[i%�����FƿpX_��azy�Ob���t���2���S廆��}�(�r��(�m�f���OhV�|� �� ~֝0�v�G�r���1�
����´O�7\<�v�l_к�+�����hD���Fw����V��'�w?�O�@�{�~�Nic�����'��ׯ�'�k���y����(�!$�O$�):H�Ć��̤�0
wŴ�>�9�o|q�
�MS��+O��l���$�䃮�	�Z�tJ�<:z���v-s�	�$�$�lGM�/f�I���ò�� ��vV�8`�x�����Y�3�(�N�3@V�v�*����"�̙f/)�n�W��z�Ǉ!~�+����7�pcv� ��<��H<�7�w�w}�������{^�H���טڣ�-�-��}�~�.�����|?��F����V$ӑ:2n�9����(
]�+�B�tE�U�P։W1L�u�`�q�8��84Fpġcf9�pR�(�cC��x���ada �C)R�(���	C��('���G������JT7Iߢ������g$a�~z����0���Ԁ�'��4,�>Wy�9��c�~DХ��� ��4us2�̆�F�7k��Ȩ��;��j5B��*e��U�呷�kB�ej���y'�_-3+}���]�k���/qc9T���Z&����I�2�w���<�Q�4V�JɅ::٨���Ya�+uR�D�mY������P�� �[�-���]W�>-����y�T�5�_wd�Bm�������J)�E���BD�b����5�ө��'�iS���KH���O<�6��1��O,����2QO22@Z��m�����ٌ�5:��
�.S���i�./yI�̩PG�j}nf#`��s�D?ec㦽yYe1�e�GY� 80���oYX �����ûN������M:Nٜ�-]�]TR�)��vz�p�m؜:��G;=�ٵ�L���G�nˉRC���	�ʺ�,��T�@E��'j��\p���r��l���YtX���&x:��S��Ї� ���t��S>|���9��P��[����q�ґJ�X�FG�%��?`2K���{qiG*	o�Ws�_��j���`�k�,���o}�q>��_���;�4���k9�c��T�s���u�;9Й���-uG�R�%}XĥL;�^`�%��)�휙-�3m+��p;"�x\}9�)��O^��r6{1%� �-ZXҵˈ�k�t��Y�Mፎ"_[%��ɚHDH�"�Cg~�{����ӱaJ@o�Þ�=�*������"��-9_�W�|~��d���u��9;��vf�8l�� R�9�ȯY��1'���H�o�6�
'��R�Ξ"�8O+���c��
���Gw�=������&���lM��$�V$��C���ǻݹ���=�WU<%Z�ӱ��@�d%�4��i�0m���n얷��%,h����t0��!9,a�͎�#+BU�d��s��0��a6t9i5ڊ�s��ƙ_�ϕgAKWL��6�K�0�r:�v���:w=]x�X�A���w-.
�{Dz51��OX`ė���/��_		@`l|t~=�0f�s��`��4�KK	UZ�MYy�meU�'LJ��Ս>ҰK~u����_[ܿ�DgOޑ�IX���dН��w��V+�H9"s���hu R�#�W��K�a8�����	5��1�1�����hY���cF.��Q%���4�0�f�V�ɶ�J��8#<:*.]�}���b���#�)_�1�Fa��	x%l�%�G�� 4��1�^�t ���jo�踺0�^g7Oe�ۄ�������_@;���a�~qu)El��ķ��i8�fo�u]�F�p��R<�8͟3wԭ�7����lm�_ӊY�s�֩e��׼���u3��W?�~J�:5�)My	^~��~��ƣt�K�i��S(��z/�c["��u���Mj� Z�p�kzt�a����=�����i���㨫r�4�3��uR�S�[��ڨ/?�%�'�� �3��ަ����G��:I}�9�S���+O�,��-z�*�zb@g�FՉO��2(���{G����*߲��_��}��N�M��/����5��Z�I"`<�m�/!D�**�����WG/n�qGn�&<ɐ�Pv`ε#t��-�ת簎��:⹲]F�n�.���=7(���F�/;hbG���5t��Q�ĸvX����3Y�$�!$������s��,���e� ��(�o$Wg�o
�5fG��XOp�G�q�������f$��p4�4B2�� �����nG�4<(!ڢ�]��7���)á�8�Xh��M"�3�V]�՛�|C�t���_x����q,�쉋������u
F���\R�gA�P�J���2��L��pK�ӎ���6{P�:���.yK��rګu���[WFn�ܑ���\r(Oe`|S���J�/�	������s��1���l��1�����1tDX!ݐď!H��ha���+P^r
�]��TJ~LTG���$_-B�M�ޥ?��:N�v"�J@�,�ú�����+Il�}����VV�,�.�PJ���yq�����t�b�l�z�a
t�w1Ʊ�(W�a��y��f� ����V����p��F�VA�-S�{�S�"ɟ���H��U���A'͑��N�.(�����8��NӾXrA^V,N��p�]��W�b�1����&���V��m8�	n���Y���f��<~����qZ i�+��|\��LሦΗ�ԕ6��l٭˭���ʎ�=r޼x�QEa2"K��m�jT�}���0�D{p_��4:}a 7��Ω�*Yl;�ˋW~4���N)�S�Ꞥ���V���/Q��/v]����ͻ0z��ty{�Jw�v�^��0Lz�!mu"�+gI�����<Ɛ�Iݛ��ƈ�#m=���:����eD!�kZ���H����	��AA����)et��&2�P����[�N'׈�/�s ��|˓Pf�:-�b~�_isͱ�%�����	@M�*�s:1G�g�:�Nݣl��5�3M��ҁ`9�N��񲍎�ŋv��z���_y�� �mjuҚ�#i[�>$�S����m�����&���:����*C�8�#�#�"�A�.8��~dZ�r�(�%_pD�E^郤=��UWv9x�i�ړ�V�lH���H�2�zx{���#���g��)!���� o�']X���+�,Xc{�qYj[���
3�hM�&�łt����1"Ʃ|��Z��DȂ�Ez��Ӏn9��<��M;7��9��)��FO��Xۈ{C�U��2M�?���A�����~�P���/!�^��{�m�y��^����
���!�+�s�x�L��7i���i�7R��*8=|6��ʻ 	��J5�_��nW~��_��f��4���%0��&3�y��W�- ��ńkdZ���\R�Ī�.H��o�,1p:WgJ^���E��ݰ���\q$l�l'qj�P����Os՛te<�a2��a�W�&������:���x�)'��q��BB0�	]���Z�-�`�%oFb4u����e
}�T�r���[<���ɲ��MǛn 	3N�>C�.����Z"� '��3�cOX?��O=ݘ?&W	K��֊�d��͋,�T+�g�7��#�>�~:8�-��(_ud�S(��i�y*!쑬�	�>�qg��E�N��S'Q�&�\=�G9av`=���Ё(yױ�\t첮NY
>)_���g'�C4��M@���?�<;����~�tk��6��+�������O4��<�ڑۼ�nۇQ�CU�'��)޽O�K](��OB��OP�nM�M��;L�^3��I�\ś��*��o��m�M�DG��lM�C��m��k)�C3��c��/�؞l���щ�h�[�~e`��m	=�j�Hg;B���4�E�PX�Rtʗw�&X
!#`
F�S�rL�Y?��8��R~T���A�OO�40ڄ���3�B�T�K�ܾ�QV����H+�6�qO:�)��W��WYO�<9��T)6���ܱ��oRҁ0����I���X�r��}#}`W'1ӎ|�Ag���<U��8�5yvjiG2�dv-��Sit{iG%3B�֞`������޷���8� ӑh7���0c���-�V���L=��{d{	��M֋���pdD#`n��2�rj푰	đ�
�漍o.�Ӌ����0`X�mx�r�l%}��0�r��I։��ی�)��5),.�J^��ԗ�&?Qlt�n�$�
��7K�y#�^��ۡ�0�uÞ(~�=B[A��7�W/x{��ܛMz��he�������|6/e�}��~����yh1A��^:3���Հ�¸)k$u'܄�Jg�GcՑ��6�=��N�9=׏��t��6Z"s�1!���8�a��0b�ƙ��: d$3"�ਟ��K��h��4�;O��NK�)�q�T?�b��� n��UO*��5y4��:QI/OA����'0�������n��M��68n	��-������!3�ۚS��&�m��	���P?��S�@����W�q�t���Խ�F{�,�C��1F]!���KF�C�=s*`��'��nws�6��c
n�����nh�cTʐj���@�����gy�L-S�����l�����iyGR
R2�݀Na�j1jO�F��:Jg6�i$Zy�#�v
E9�3��O��ݓd�3MK�zM0�%/�̆ذ��=o��7��<���>ca�����n;�#�}�G���~^����?��,��-:	`�2��0Nu���Q�uV(�D�c�������D�=��-�c������a�\>�@��y|8��8���]X���r�����w���u�>���:>�������Μ#����'����2�`g���tHRO�4C�-=�y6�h����D�$�+/�9H��a�/�<d$�o>n;B���پ-]em��CȠ��[���e]�,�A�jʼ��bk{�@vZ&*P�����5�@đt�r��:�����d:�|˩T���� 3_X\0ڵ��>/�I?H��r�ȗ��t�hH���k�(�H��{Q�O`��j�[�'
Ǡ����Yl�^��1���
��	�b�xa���Y<]<Q����a]TY�c�>!�ߩ@W�����%Ͼ��N���q]�aO2�;��;�� '��s޼x���Hޒ`��ޅә��]��M��V�=k�c� E��?`���������\�4��N��8����}<�^�&(f�M@�]�o��|����l]:E��s	6Z��!�>���md���P�}�
Q�e��06�*����.�I��-]���s�6���!��$M����WT�i��4e��L������
b�k��k�N��,�k�\nz�^�d�ϖ��R��k"��A�]n	&�p�,Q��!eD�ђ8'&&��x�#<HQ�T��7Hl�-��{陎��eUr���)���N�F���F���Hr}Z1B�BNל�.[`х�e����}ס�a��^e'=����r:j����9�[:v��'�l��+�E��� d�2+�p�5�Si���ٙ��7��l��F�OT�42�^�͏����+��o�t�SgC�	D^�z�ӹ�Ѵ.�.ld���#�	�Y@O�Z��o�2y_;�w�	���.H.����ϔHh�w�$��:xv/we}9	�
����|��t)O�R��,��+�,���-����_������5c�ПO� s7�Ζ�P{����s��"��Czڵ �/���,��R4~zzc
�@㑴a��ۣz��\4vZ��=�����u�?�Y�y�ΌQ��*/y�Rw8u�8�wO�t����9�ɹ�sW�?9-�WlR_�R���^�i/�N3�c�{��_ց9 .mX����X&�|��ԕqg1�N<��g�L'l�=�3C|_���.	���Q��<��3ټ�t�ܶ��`�]�=�<�����E��a 6G%��p)j�,/�\�CQhJw�;�G�!�=Dk�n�v�0����(A=�'�� ��-y�s�y5�^��/��2�f\�eģӤg;����!�tdǡ:+�C�NQ�s���#/�/��Upz�LI�'�k��1��N��
e\?��������F��B��#g���'�3b�v��RG��vࢁ�^�����d�����-so2j�u��/M�g��Hk+!�|��P=�`���k�یPi��/>���w���v��ßxM�t�3����+˯����Hs�|���Ȳs ڑ�k�f�؈�GYJU$���sJ�Mb�JX{n	��э֣�C"�8{�40�������-�SӴ��QY�\k�� ��9(W���k\�)�3�XFeI�.���(�O��KGD��{썘\@Ҏ·��`��!3��4�"���jx�|���!��}�{u�2*bS���x{s��}�N׈QՀЗU�Gݏ�DC]|M�Io�������=�z�H���k6$���E���Iri�Ӏxqny�qE��{�������;�4Y�I�?'\U�9���2���̷�ً瀺���,������L�"!�����_ud<��%4����z�nx�##L��S&�6A'��NuڐTX�W��Y��@�V񡗟2c�΢�>�iW`M�q$Ƚ�g}{W�Z�8�4^��ī#�;	�*'�K�,�V�؋R���0��)eQG�� N�g�#x�6��Ǔ��Y�����|�܆ܼ�n��c=u
��hS�esQ 6��7ZS'�0��Yt��fc{Z���B�3�+�) ��l[f	��'����\ƀ�e���w�N��x?���e-鸷�O�@T�DV�	�p�ǭ`�ݼ>"�]�g|_q��|sڼ=^2�4=���}���E��a�bT��4��W;d�G��kQ:@Y{��rc=��^�%�W|u�6�oN�ڱ �N��[|��7��lE>7���5G#���"�-7�v����m�Q��`�� ��Fft]��f��0�>�ַ�O��\{c'�?�[:��AԾg�9AT�P�P4z�9'dhGr(@�4+�1�~���0�		�a�H#YY7����d�TXT���p)�0�vpĦj0�9^Ƒ�l�*Uɴr��'�D�22=�� w��3��$�$-�,T��3xܙ2u!/F��*�lx�&��^��6��z��Ҹ:UiN�5nG��T�1 -r�d��(wQ���6î:bg,\=eS�?�4\��kz�n��d����1=�樝�t�eH i���1������Ǿ�(X�l�S� ni��t�66k�i|���Z��+\�P�ǰNO{��vL0O������Jٳ�0��׈��#:";���GeW����
�(��5�c#>M��d -}�`|�i8�h��
^�Fں,���'�3�L��Ux�-��`�>|���#pΆ\]iɚH���N��@G�VG
�-�I��vx��_�����_�0�C�y��i�׈��B�����^8=+F�.�f� �C�p�#�>�2�V2���\������9�-��jx��7��_|;��lo�zkw8w��	�3��K�_��`,~�a��~x��?�?�ȧKX�B.KE#_�ۆ�6:�m�{�<�X4���<T��y&��=�CG����-�� �z5t�����aa�>A��Br���Zn�uq^}c�F����:��zƈʅ{%Q�v���c���q5�w4̵���������V��d\!��]���@�𕛤l,\y����l�Ti:��6�Dy?@�4ܣ(HyU@#����ʻ"��GsK3�H��U�y��J`@G���76����L�M{�#��Y�]q+�[:4���Whc�&8y����R��.ys�^�ɐ���0�Mhɵ�dD=��!QI���7��������v�NH�;tl�љq��uj���+Ԕ�uG�ֹ�U{����z�y�y�6����DWO�z������Z!䋫#_�@xh�7�"u�����:'�G���y^�T)j�Y/��,𑰖�!��W�=Öe������6T�AVA�A&�_��5B���C	ɴr~<�(6�+��)L	�x�>Cw���2������3c��������N��Xd�"�:��s�􅊁p!A�AΉ&U��_˷R�����k��Ju���������K�SO��O$᜽|�4�(��BV�C�ɑ��wn1Vh�4R�5Q�|��YJR��,>�5iy���ʰ�X�"�W#��2y6H�$)DQH�D���[t5!X �qMbp"��܋�iD�h�:����~��������j�o��b~�B���00s�қe*?ejZ�X�D��e�S���-�i��7l�L7�u�����г�s�-y	Ў���Gh��O`
a"{2����L�nzNj��6(��C#���b*���.#_o�����a����hy����E�+ivT�^�&�� ���o6n�	:�����[�Y68���<�f[8NLWޱ}���v�q~�+�l���׿�~����%�p��E!���?����R)�ff�(����a��6cT�c�3%9!!��=d��S�)?i0 �F3R*y�K�t�G�%*ݙ�)�{���?�E�SN/���R�w��5��}6e�H!��b�Eg�L�mtϴ��<~���wt���b�oz9���Cl�z���=O9(��*�)g-��mfx�a�P�(sȄN�<w����k"�U�O�1�:#؈ߘ���u��l� ����e�o��`J���&�^�W�#]���Z\�)w;6��Y��ٔ�v�r��bg��x�)o:��~��[<��δA�g�y���BkT�r��k�A����;G�e �zd�k?�e+M���E|�����t�(��)�g�-�=�,��!���I7���G�H��
Q��n�ݩ�[W���䛛����[��軸< ��F;P9���E+�gd���{��@���W8�{�)��ً� ���K?���]#@�AiˍK	ě-a�6�g����IDJ�i<�2�@� /��`d"Q0�K�OC�)� [���x6`J/�
/��޺1�S�+n��6=Ɖ,���2(*���'��g�9�]�f���+f$��+�t��
tu�|��+_�x��5�`;���/��0���3�g56d-���CʧG�l�<�����=�JO��4���*�w���K�ٷ䑵Ƭ^�ǹ`Tfc�i+kbĄ���'����}�����(��Siԃjă$�����b���0A�`��0d�F#u9�1�RC#�4�� 3��ܘ�Ѭ�/�'8@O��f8x�:��&�<v���K��v�zꛉ��޲���96��n8�Z�O.2ft������Şm��b�|����ā�c*D��%K�#;�5šM����&u����O~��E�'�j��������z':��g����,�-'GD�T>U`9�#3���Ο� (yp�:_E��e�M�,��3�kF�L2��$UI�g��9��L��_��gZjM�KU�sc��eD��/�~#$KR#¯���� �Å�'��Oʋ{x���܂�t����O1���o���1؛��u�OOe�Yϙ�}!�)���wf��{�u�-�����yk^�/X\�˝<����d��؋4��1�t�C2ty橴�C�t�����uf�)�|�-��ޤ�G~�� ���-^f+w���O���0\s^V-j?g;Ѷ�4���u�N�l�G�E����ç�`�D�)��W���9�aߋ��6�������w��N�dVi�U9�x���F����2���(Q���M@3
?�Ѩ�7�ӆ	B�7{H�\�\� ցK���
�f&a�c���5�'�y7#�+� {8�����,פ�Ȁ
cǳH���L��#%1���*:��<�Ⱪ�!�����	s6����J"��0�T.v�93��%�fS\��� `/f�l�����]��M��K�7���5��m��o��܈�Q�����Ï���GI�y;`Y*��\�1�"��LA4�JA~��^~]��G'�4Ͷ[i644@���a�i������'n�jx^�L���
 xl���x~�.g<�nP6]�N4�x*�<�G�.LpX�%ґ�R�����l�Fj&#�i ��ځ�F��ɦ�m�d��,��������t�[n64/3�oq+*�~�Hfؼ���A8S��B��| q���7)<:��Iݷ9�����K����͌�ˎ;4٤������ �EB���F�Ŀ�`�v�)���?�|�/�7������Ǘ�3��@�ǟ~������|�_������X��(���դȿ�Q��[�ز���ѹ�A�UwxK�sx<d?�w�?�|�O�ss��{t[a��Rg�#]��P�.#�yO�lt|����:��6�1K���p{_���d``��"kG+l:D0�[��T7���g|��3^/^b����cdG�8S�c8���]:y_�r�öU��g0�I��Q>K]<�|^L��)�L:�f݄��x>���1��"��Ձ>��z7�3�̯�
�������)��p�����'��җR^����$�;�9@� @￸1���E���Ic[c֞��)��L�8�SV�!.���9��X��˳0	r��z~G��& ��蕜�w��Z;��̵ˍ��6fߛb�
13����5.eh�,ic�����Ww��Y��v_��B�=8(��C��� &u���\29/�dL���>�ϻ|L�&�4h���	�IE6 �:ʀP�Y10d���TT�ք�a�5S���z�]~&�V�t��'�+73���&�k�7f�T���0����1�W�E�qXΏ��H��i����p�Z��3�Qγ�����,y����=oa�i�F�}���e�C޼8�Wx;jig5�)�*7q�#�Д�(���@�o��xf����%eC&f#�׿f�^�_��M\{*Y���>�S���\҆���U��#�`��{�t�S�����j;�5��#�u _�o��D�w��B*S<���	��J����-4�1g�d�{��o�4�񋿿It��g2=���#�����^%��h[���z�Ob,�����љv���
˿�Of���ɬ�9��@�W����3"G,1����x#��.��=6�����|�w�y����܃6=K��ys�<���kE���'?дSr�������Iz�����dzÖ�z04Bp�����D�"(�֟zތ�F2%��.���]����ɕ æ���r�<4k�O�t�BcR�%�p��Ry��w����Y?��O��������s�zL��Y��ȣ��D��Y�
�������0d� fq�Q߶��dHa���"a�S��fM��5���H���;q�����
���	�N��{��O�	
�x�~�}x��ŷ�2[LYP̧��D�-�`�Rx����}��I��|�,>v6�����m�}�I�D33VA��bȂ�l�MF�S��!y��2 c���J��Ӧ�k�7���w�/�'�"/���\�w�eq���c���Lʃ�!�{��g �/��c��w� ��@���X]�$��␧|΀]��y;l۟���B��Aq���Ss� ���,� cf�ƜS�i�e��IW�U��Oc'_�>��?_��'a-TF����0���X��+�穤ͯ*5���~C�$q�2[❿d�?�B:�;�#+���2��ˏ?�"���z����ɰy�.�����WnH�[���^lAgX���h�$�� {�^a�0���>o?�ĕ� ��y����g�oF7�-��	iP�
L�K0����`�x�T)��&,�ش��m���ۦ:�m�(x&��ϛeY^$����wa���S0^y�6����u��ܧ�^`�xc�"���y/>4��@Yo�ӷJ�ؑ����ߖ��da��*a��S�:��e�K��:��)a��q��S��V�"���p�uW��B�dϘz�vu��Ǜ?�_�m���3��0cf�|�Gp1Ύ��	�e���r�����2��fZJ�v��v�v�K�u����y����~�aJh�7c/�uf�E/n]��B����!����AH�j�4��[�|2F��%�|�xyI{��o��]}�l~O��Հ���]�+��c%�0*�N���"�6��,D_�w��%.�e9��/�}��K��S�*��Ue�����ɍz�!^]�*��U�2kԔ��F��z����z"�kabܔa��H�>_E1�Gz����"��-g+�+ld��1ģ�4�r1Ķ��4RVʞ�̷8Q~���}����+Xh��7��Ʊ��N�fI�9z��Jc�������M�f�?�H���N�N�g��6%'��d��u�₃���4l�,�{���vq'c�Kbԙ`��R>�~CM;��}+h�k�t-O�����)� ��S3��G2��n�ⶈ^	�����qW�f�f���X�n�F�6�d.��@5�$s�?��/\Jt�6�I/ĶD��w�e���
�����2��X����QPFv�t���:�^��N��c�B���n�k^	I�m���Z��l�y壞�!�s����mM���]6�T����!���d$�$�k��B�^�	���?���4n�h.���,Q[4ְ�[��7B'��x���ӭ�I�-#{&p(���	x2��!q�M�	�5Yz�%a07���0�5�e���՞��+܆��VHg~��2C;3`��6"^x��H{֩dy�\�R�Zv��P�����s��**Q[_U6\�dmcG���s@�Q� ���/?챬��v��}3K)E5�ٖ,� �E�l�� 3��v�I����uH�x�A�a���7�0�0("����� ��c
[�)ȏ�o�
I���d�qw��7�?ޜ<}�y���0�]�X+����́�W]xA���i	S�I�X�Z^Sfޅ�S�)=�Mi=4<�F.�9y�Ω{�>��+eE)nΙ}�`�6J�1��_~`O,���lG��2m��o�=N���5��D��V���4���24I��f�k^E6��]�1��|^��_�@����3�'�>K�D˟�ɂyz��|���7�fz����V��l���2fߣ�F��[alO��{.�#�y:�!e�>��9���=娗���6�(R��P姜��bV]��r[�4Ml ڧ�㘽i�M}�I��L�94�֥,�'�0R�C2>�G7�81�r��SJ�N:i��W!
mxur�D���*�<_I(b\~�D���M�g�ґd�Lb+���L�����i,�\(e?���f���e��N�U�Ϙ�,~g���f���4�S!��2/KE��A���ي(e*�%�Y%�!�A��z-z�ZYX�P���e;��'���3H�;��T�oN��'t�y�=oH��R��g�L��:�&u�V�ȓ�V��4Iu� L�*��~F��V�R����C���wv�7y3���8h7W�,>����=L�Ae�c���8��Qw��|�v�,pClI�~g��  @ IDAT-�i��q�8�|��x�t��R� ���8���n��d�%�=��������;hB,�S��`�+O;�1�2g�ȟ�WX2P�m�.o��q�7�Y��Qg�/�3�"vD��F9QJ!���ӑqd�R3X�-��ig���4�o�u���l$�,�Aڢ�^P'�+e`��-s�N2���d:�[.�{�8��ȷ)��m�
0�2q.~�"�U߬�ݭ!�k��3x����ٙ;yK ��`��[�U�oF�(�-G!cX�$y���~�N�s��U�9��R���o=�w�{y�d>�����'໙ەO߷�r�Z��s�쳿�v��'|f:���H��dJ�_���Ыq�[ç����I?鏠��J�'�[��A�[ �u9�p)Ô��Ż"
*��c��_�P=�n��<:*ͅ��cʕ��`|���ʇ�i;��b�\M	?�M�H/l��c����S�`ڙ�Vg������u5�w�
���0}��`S���i�n��"=�~�<�� H���b��KR�@��z���!�n'���	���?���~<%<��4�xj����`F�W��D���QZf e@D�ۤ��Ӹt��L<���ss��P����8�>e}�?����ng���s��ӥ��ř��\�b=ʀ
�N�� �F��RfB�ԙq�ِ�#tfh�\x�Ԡ�(D8�ŎXb���#��뙴$����G��iYA�����~*��p��_[����y���0�F�>����
k��,L���5_���_q	�4E�4U������''���8ct���]�(��U���e����22,�r+��4Bl�pؗ;�Y���LG���p�!x�a峔%!�Ff�m���{hmGI�Us:�L����5�d��57{��uY*�t���eu5��2�J����*�)kO�?`�.Ǯh��r�@2h#��]^�>��wdQ�Rb�Q(us�+�Bo~Cѥ7������x���gͷx�	�k�=O�w�V#�J�:��i��I�ޖ�aSv�B�&l�'ަ�!q�j�7O�/�zʊ<yn >������.���<}�o`.��I:sbY��/�8�j�5��������7Y^����+��)�+Y]y^l3�m�m����^��ȓc�q3�6�.��u�ż���+G�v�#3�ޯa��F0Q�Sk�y��QR�ٷE_@�@������{Ό�w�[z���6K��W���0v(9�{��7����d�u�l�t�@�x��o�|×]0�33����{��㟼�n�۪9N%jݮ �bu�v4�/�-�uU'��!0�
#0:���4.�|��f�0�����,jP�M�A(-��}�m?�K��؎�N2��ϫ��V
�c2��f��&�[��ܸ��%�)��^iǷ>N�J��' 7��3�!�����ʅ3M��5����h*�wt
'�Ϩ5��	�ɳ?=V- �n%��ڊ:R���;��37�y�W*m��3ry_ٔH�L]�l�� Gu�AN�
�6~+|�NZV��'<�_�|6.��I���@�7I� ����Ӈ�8�I����qk�-��ԙ�(�T0��s2����"y�L��/K"��i�=�|�!0�U�t��Ci�rاLe��i��w�ق�#&#و�>kYy�U^�~]���:��R�t��bǯ�~���$��f�͆n�+��)q���}`����	��"̍�X��4��fi��#��q�[ڍ���pd�l�~�������@�Κz��7�������й�r�'��-{"P����
w?m��7"{���!�~�X���"S�A^>����r��{�>���9��.FD�	����B�S�xS"�Y�b�!{��6?te�Qm���v6�Q}�'�5�	�,��3�#�(e��l��"��D�8��L�����dv�rsv�%Eg�x�'_ڸ{O��d��oc{p���;f��7#;���=f��N�ӫ����"��װJ�g<^�C7d{��ڈ9��$q~�,v�x�������'1�����zlXUD��Q�}&b$Mx�nƵ�O
3��r�2�i	�?߰���)�3f)�`N�Y���M�a�3h���lC%ϔ��#-7�yv��2���X��-��q�zT��^�~���D����vh�hl�=7���c>Qv/sfL1W=���>n�u>��:���3
-<�0����N�����n�>%=�x��{oF���}u���')����M�3U�o����j@u:�l�z伥|0׎�@�g0eǂ��od��1���E�2�W�G��W'��}��Y�ifȚ�>�_~)��ӎNT�.���|(�>������8�G%	N�Jgׄ��i��c'ʔʅV��(��I�$<���������#]F/�" .-�DDI���+���2��B���(��Gq f�B5>7�LE�D%���u7}�3Ґ>>����5���7�2���j�S*�l:ƀ.�RM`=mG�%,R��S���l|�gysד�I#�x��\|�M��c̍�Oc^ڦր�r�	�D�����N�?q���B�~��Zxi��UY��?��wd���M�`�&�3���韲�Y"��p�9SϿ��#%�e���s�1�Ԑ���v�(��-fpvYv�C�
����H%2��t��SZ����
O��a���o2��ì�#�΂�<�-
Yy�d�������]��b�yj����$�ׯ+_������m���%�����af���ᐙ,ar�����7�ǅͷ��;t��8K̬�^�v�6drYh�M�ߏs��kۄ�J�?W�2�m�M�z'�D�U�LX��&�18a`tl��oҁ/���?����0��kő\�R@�6O��_��}3�9��ܤQ�_J78��t��C��F󖣑�����j}���ey�}�}����]x��Xp�C�7I���6�^2�������9�o�E4�*w�ʼ9>c��'���ᮞ�X�#�Sy����FX��O~���;��7����µM� ����o�z���aO�n�0'��þ��L�{.5��mE�Eo��-�C�#X�p(����?3�GN"� ��ԊT�f�ꚉ`(R�����	aV뼯I��'��v�M3S�_S�t�C�
��W�/0a>rt�����޼�{g|���]+�g��ӄWE%��I��PV��"����LL�1G>���l����;~SA�`R!9c #p�$)͙�6�&:���")p+>y&*�<�k�a�� �W�hC)�N7��v�U�$ע��<��*daB#�T޽Pɰ��92r�C#�Go�0#�T�=��zz�$��/e0��oAfm8D5z�9��h�4�9r���z���1�SU�L�/�y
��Բiy4`;J��d	~띳u9I�ve#/{�\��MN�W��W��o�2��JE�=���;�Q�P��g��S��S��6�
~@۽�L���m�|���������7���m~�ӟ2v�Ѥl�����ߑ��IΤ��o�	c��O���ᴜv�t�C�5��-O���D��1g"}��W���~���
ACׁ�I�C�M��ƥ��,ze�^6��n��_�� 3�������3��3A
�03��; �Xs�����
�+��<9���9se'������9	L�ҥK�� �s�yx�7P)�m�������t��UW�<@v��+���z��_|��ߙC̀Mغ#�� ���l�f�:/n�^�\E"��.��濲&>�b,>�{���U,ao!%�����Y�ª</������3ܼ/���yp��{��,C���l�6i��Y>�x��i�8#���o�e�\�
m&"EO�~�%_ 1��ǫ8���jg�"k�O���!�+�Sfj�t�y�4�/�ah��'���W��ոޚY� g�N�|��b��Ox����s�����Ձ���|�{�g�x3O�rS&f��-c�iX��9-CK%�a@��;�����{N7�X��٦��mv���>�j�fp�&6�Na��L-_�[�YFAY���G>��c^���l�.�W���iQq�?"}1���2"ld �v7��xg��ss�iE�k�c���^��H)����GX׍��)mȄ/�!>��RI�4a����1�&�
[:��!a76n��M�F������qz��I j��"����64@<i��z�$�Cd5�L��A���~�i��u�ƗF��`.��O�Gf�#/��*) �u��e�R�)u�ƋSܶ������#��4� �_w��<��+�Ż�	�K���8���5B�ȼ�˥*�lg��{ڌ9��`�Ջg�O�߼~�ls�U�:K�7_h�9�b��A��v�g�r���o�M�n�e}�l)���T߽}��OY�d/F�r��;��9W��Y�X��`D�C�3y�g�͠�P�~�X>���L;d��<�Їb x����r�z�@�!�^@eT���ʞ8axّP��)�Hc6���%E9X�*�l7ͻ�4\����0y�x_x��q3A��O��m��)�H�"r	m&�~������*[�W�ѳ|
��]��u��o;��g�j����S榩�,���pw���"3S�����l[�A Ղ4�j��`��ޫ	LT��N~"j SD�Ŧ�p�Q�덟��q쪮:�ڭ[~U��%�v��C�k�U�Җ2����q��O���C�Ϲ�dD&�NƠ�ON�1���ޠ��m�p�,�3ej~��P]e�M�M.H/g�������6���z�����@��½S2��;�Һ�Ȁ�� l�NQ�;�}���`��J&�y�*��4����V�Op�P+Fץ�����&�}������g�3	nt�n��UܷcZ�`3�ɡ^.x�����6�Rt3�_��ezp3b��H,,����w =��e3Î{�����s�qt#]R�,��N^d��TUIY��{<˳���ۆb�'-+�wqy_�,��?��M�sR�3X,ȵߦ��ґ��ޫ��a����9����#u;]��K�%���%�PYgyR\�Q7^UD����'�ؿ�{�g%�}��#�M������z��'�FE=���@;	�s��<�[\�Bt?�X�i�HY����OyG�x�Th�	�ٯ�\=��٪���u�җo��I�`���̘�������>�n��a �ɷ�m~`��+f��+��	{���>3�-�7�C+A�� XO������_k�=�����ϛ��Y�̄e����m8gѬP�����T0���h6��@ʟg];R�CϊФ�X?�˻������'.P3��qV����K]2�����6qh�	��z)���~���'��]�n���C�c=x�&KN��f�!�ȷ!��F�g�ɛ�.��d��H
{�1����6"dI�;sJG1;�^�Ɣ��٘��w�9��L9��!֟�����Y.���0'0��)㔑�3�q�J%B1s����¾�7O����why	�p?�&N�]�&����ٱD���s�i�Y�NÓi�e䀆�8z�����|!����2�����V_~{�98f@%1��ǟ̚�\.94�:���g�nv�+M�p��m��i�8Åd2'Du�L������3�k�L8mCN��W�G�[�)˙��;?��tM)r�	�p�ɨ���1��`�7(Y��j��	��ĵ��B�[289[��f<� �]O~��,���*�@TF_l���u̍�6v+�;��'_�^��R���ۖ�O߀R�{��5�?�?ޭq��x�I�<������MAax]^h`f��FF��aa�>0�ѤOŊ����4b������'����N��<���A��0�	��T�7zI7n6F�
S��ʐ<l��yF��B�R�/ B|�N��8���qw��ZO'q�g���ɭ2M�;��"JEt�ְ΄a�@Ŀ�Q�qe������v�u1$.����4T�k�A7�"_^ʑ{?A��)U�t�����A�檃:�,�X5{��:�t�d�B�����2su��>���8//ȸL̒.��H΁W�=�}�q��t8���f��>�|�����:��q���q����t�G$��V\J'�z&�>�i���j�ȍ`;���#KAo��R�R��H���4�f}ՠq0�t�,Z6�y�o���Bu ��fW����e�����2�mUqf�$��x�8e�V�Bm	�^s��$��_*f��p\+��W�+⁋��7`"+�3�T��4�	�b ��%x�g���[�_C��7�W���|�.��@L����Ac�(+���{����}����0�N{��W�j���q������E����%=h�z��V]��<K����'l�y����ε|p�����>5<8�u�ځ��C7�+�5 o)��K��\��%�����+�yT�c �R ל<r�!m�e�.�B���p�au�J0�D.�� s[m�[dI�z��r�،.�[鷼��*��eCtD˞�	�,�hX+֨<T߀ru�}!�X�{^4b;4g�Lu��0�?q���fp�mņ_6�^b|��X��2�F�
�i��l���9�A{���m;{$0�4�\�t#��3S��d^Fj�4.����X�����'Q[X��D�����D�����枵*�LA�9U;p�����[��f��PkM�<�R�a�8��=>�5�I�����nm�¶��	�-�מ�[>LU��A ��{F���)Y�U*'Ӆ.p�E�3e�ed���.;��ś�RQ*nԾ`�����0g|��f���l���K2چ�۸̨�0�� H��FZ��}�&U�IF%�"�g`��?��Un�vV���-�;�MT�d�%訹��(E��uкg�}���e�m���liGَ@���p9x�m�6������E��#�U�<��^�����E����{K6hKk(��qyԈ��9���拿��͗_�6o�9#�6Kz�I[��6�0�~�����>A�/T�>�Y@e�'p0��'����2�,#��΀Y*�@C�3mq�N��x�h(A&�����S��PWg]7�F�3���:Sy����������9:U7s��;��=1�����s2���`1���	��M�<�N�Y6#ל9���1�B�Ǒ���%�L���9/>ۋ�Ylh�@��h�V~�Y]p����1�e���G�ݔ� �@��٢��²�	�w�Oݴ�n�om��o�����G�1i�b8��2�#*�[��/dXKʆ����O��ND�-�y������P���i�p�2�K�g�o���ͬ�g�|���7]Ϣ_mD�gKUgA-5� �-8���������U@HUgl!�x�τ��+3���B[ �q�Au�=b;�>^�3 �<u����ː���P�W�58U�C���m��M�����,���^Jif4*R���+k��Ё�� ��鈃��QAf��F��6�(���_h��-�S�[y�����r+? �OɀkǷ���?r��g(�9�t�T/�l���^�}�4�{"v�L~���_Tl:;+{;ȡX#Q�,'��~�`�W�-��PHo�4:J^��ӯ1��£�:K���ٴ��v�>hn�o\���I�i1��'�o���d��wN�7f��ҙui�Y���f����1tƘnP�i,�u��/���]��r�,r��n�׈�I�:Z����2;�y<p�����C�4�Ҩ�����R���V����:{1�2R�m�6��5�WE+���)ڦ�<,��+�>�۱mT����ɺ��l	�ަ~~`���S�	������fc��ͼPg�����H�B�|0���Ӡ�Uh�*��!+��������� Pc:a�_�<��3N�w�˷)����%�r���K��0ͥ�l��ػ�<��p�F(��HפE>pI��̛��s�#�_p�o<O��.��5���d�I�,�s#z���(�e!;a�M�R>�}!�M�,�Q~���ut�|���P]Y�gn\3[������E�翗y�yKM',A#�8��W��}��B�y�튭!W�)�cxVG8��	�Cx���6�2ܐ�o���J���V�^�R���&� П�����n��<������G�(<f J�8\��� в�Қ��vʛx�'�C��F���9��##��]]�r�_�Oѿ�z�y�,ؓ�/����/��h��Y%>u
zy��n�߿�G ��;�g�*Zk��N�a�<�%�ɴ��)\�}�� �c�9q�KA(���k�s�f<�l�i9N��wVE��!e��}&Nԕ��0�td]Q���=���s�mFdJ��s��,p��8aF�-��њd�b����*�y-r�A*{^��`���03fW�,�D���;�.���Ե�ś�-#p��2���d_�y~�#��G������6�����	Jkשuf�8�q'3`�`�~���b�<��QYG������
��rlL+v2�xb)<aD't���F���7���?�r!���b)wC��/e�F�L��}q��<�'��Y��[���ķ��
/��On!=�VR�H���r�mCi�����0��递�2����t�X.�I�Y��n�t�x���6�-�rD��и�!B���(� 0i�f��5�Y���AK��#gv!g�@'6{h�1v&�<̢�E�l�r�[���O~�x,u��<L�,O��R@;L��Й�O��Tf�Q��Cģ�8\��v懫5��0|���@�,�;��Y�����X�+Nf����O��^�rF���|�[x"�Z���&
�!��>� {���,C� #�I�kɛ�7���z\���8oj�&�Y$���#q;7'neKO��²�a��5qo��\�r�'��z/��L����..�@�+��C�1k�L��J;BWG�_�s��Y7�˪ ��{�KW��)?���7'��C�^��5:X(�~U`�#��4����U����k���	%P�Kxq+k�Ǹ�K�W�����|l��AHg:����bn�/E݄Oq�o�)�8���;8"��,�����|�.�ɿ�����8aV8	zI�Ȃ���y��*��>ې	���Q1Ը',��'�
ý�Ϻ ��(����>T��$�i ��,.�j�p�l4���1|8�	��/�n�׿~E?���o?��e����57�g�Ƿ�:FG�u�7,o��+�����i�<�wW�(!�	 �&<휾�9g�����W�aY���7�{���ց���:`�O֩]��X`��Rh����m�sɞU�C��A�(F��]�%Hr2d(���ܻ����$� �g��Z�"C4ғ�7��2��9E4�����1�'dXg��;�S��[w9	#�O��?*R�(��ddR0�h���
���#�>O�_1:gyĥ��O�O%|����w?�ظ��eǝ�.����9�;lķ����pnWP�w}W�vH�&�e}&��ϙ,qH���.V����JhB_ᡁ����c:�p�w����#TZD,��>h��P�5v*���y~�SwF|���ydMKxdCl �	�"��@�T����*`�Ye��ȎO�F�7rt�$�i�=:K�=v*�9��jʃ Q�,����ۆ����v�h�ט�iALXER�KX>��Y�&�t	��_C*�<oy�����qx*�"'ՂӲ� g��?rV��q�lT�r�K�'j��U��2^�}-���ʮ�	Igj<��}o�ն�6^��VE���H1m���7�\������:3d~ҶH����w�N�M˥����S�I�H�5�alR�D�K8B'b�3D���6`��<	8��H�c;e ��w-#ÓC�-\�s����):���5����=w���8�z��
�.v�)F����P7/@梨�,F�7;!l-���1���S��-���yˊgb���9 0a�51)J+��X	�	r�B`�}�<T&�WO�8��*_�G"8�����+��iq�È^V������E��:x�!���S�F\�+�̀�I�R�ֿ�W*�i�R��ɋ]&/>`T��,�9������7?<c���<|p�1+`�@�P�4��ax9��O{��ՙ�����K���,����|F��wt��_�B=�Q�`�V!ܕ1��i�+O������sfz�͖P��v005�&��Ϡ�*���ڙ��,�}GY"�@�c�:S;�S B��`���^`I��f���#�����w�#�6�!q;2�W�"@�?�'���\�ãw�{���h����4�L�D����,>/e�h(���J���/�p�����,�^`|�����
�ʉ�_|*��'?n������-^m��ɼ|����pRc�sj��h�A��(_�#/N���)fĸ+ac��E�3~���#D���#A �Q��t#v�i��h�Y�љD^�MƯ2_8N��	�&}���5ݔϼG�3���G�&���O�Fը�����,5"�~�o[�����tZ�$��fR4<ӹS��>ڀm����Md�������y��dF<���
Ѵ���9K��m�
d��0��c7I+�d|�����|
4~�?�GzEۀ�*�<K9~�>MK[3��+�UT�P,�92���D��m���.oArr�mR���L�~ YJp��=�J�� ��XN��.H�k��zg}=�����1BZ�Gۢ{b�s���8J���g���?7���=��G�my�0H�D�i�5X-ƴmh�������w�$�;�PO�)��QWŁ[��/��&�ᶼ�l�����:�,6e�t��\�x��,YN\dFY��h��$L�3܎�0;���oz��Ϗ߾ڼ~�l���+Խ3�=�퐃���ep졮F�i��ݼ�5�wz��G���1�F��Y��<��^q�(��������
�EQm%aSB)�Ȼrm#����7h⛉*n�z׭��YB�-	G�LD8�H{��;��2�!|\��>�~F^�D��>�!�FQ�>*��^P6j���$��~��5�3����'�4�I��j7ʜ��=�lٱ>ʜ����cfV����x��p&��Gw�Kܻ�U6�9K~���T�/��qvɳ9ݓ}���C���ș/�Xƭc�������3g�N���=^��-��/�C8y%(3���:�Nf��rg��I��_Z�/��^Ύٺė�ȣ���+�	����~K{���'c2CZt��Ty<w����O�3e%�(����5�`�@
c!j�e���ϧ�D=(�C3�����Ng�T)*%������0�~�^������,�1KO�ң���Fx��l�'d�-�|�y���ޑV�3q̀�l��"O�f��Z��{�c���<A�w\��0����CW��c���/��[��Jc��fmp�@�
8BS��L��r[�L�W���ж�Jiƅ?qA+i�=I�nb�a�����&_����Q1�GŽ��tA,�q��\�+�"�+� H����ȁ	�Q����6:���a��0y����K:(��}9n$�LA�#+�v^nBv���]��[oB�?���#]yhd��F��,�E�$RvqKZ�Ǖ|��.e�`�=�2e��oÉ/�g1!Y�)�7�@I���@ҳ�c+����:ك���O�2;�M[.o�=�wG�^n>��_{抬�#g耧ϟn��{�����w����]�H}�h�G��-ƛysO^�Z�7�D�t��d��dO+w�5����MN Wo�SRh�<(��p��[���LyV.m�[�B��&�@dQC�;UG�Q�zL�L>�-Hgv\�rF�u��s���e�����gC�} 麗R�Ӗ�� �@o� K.���34�	P��l4$"��N7�yt�K9���]��f]#�.�i�2S��/���#;�$I�Xr4�� u�Tl-��2����|�iB�����ꩉ˻J~�e�K��V̟M>�G� ��T�F�!ݟ	Us\G���i� a�@#>\���#���ԣKW�l���,���1+N�S������-����<'�e�]f��`�X���if��E� ��^�eq�Ѽa=f�ΰO���>�Ç�B�`�g̊{�ӆ�f����1�ONM�����="�6���x�N@��/m1��r����%3ɗ<��-������x��!�� I�QfH�K�#xG�5�<v�gg�I8E�ʩ" Mt��%�I��"N����C�Bf ũԯ��Q��Pvw7�P���zqX"J��d�\�FOPf2[�v�*���Tx�2I�� ����&^o������Wߢ�}�;��^4� QJ��s�#��7�������BQt�PF�9��5&���\�\��J�&��t�߬$�̒w�D���OEU�4mq�z���P�O��Md�P�rQ�hiQb<�ۆ�����M��6���J؄��<R4�lN�q��s��,\�Nؔ��V�#]C�����Q�<��Bv��uǽ���������<G�n���ԙ���"�:�O��+�Z�S^y[���^���$dc*u�T:���(p�tK����V�Sj�(�kR~պK�$C6�"ct���!�
�s�l�紹;k�!�_�N���N99z�x>�zq���c��x������_=�ts��|PZ.\"{����)'�w�.��>���ͧ�����>�aʯ#�W�����s^��na�%���#�۔%
�oXZn{~ ��7��R��.���<�'�|[*�4垔�C�	k� �.F�BLY(7�Q!�,u� �e>m�p�'�*!�69	�|��LK'�.4o~��2q m��ssߢ����Հwo^�)1�@���1tH�{_:@P���̾�/�x`��T���c?z %#{�i����ò>�tf5`�{v��͓���!b#]�����[I$>���Aʩ�@�Pʐ��,f�Sv-�ϺI'⟩��ɒ�$l�R�,��5)��7����EFx�v�_	"L�^�5�	on����0�=%I)�?�?D��q��������Q��dd������ 0���i��	B��>ߊ�������6G���D���{�&��iO���!�\��̠����ca�ܖ�~�8�??fYѷ�;Io����?����W#���߽[�W�>H���^Ń6͓��c�Y�݋4��$�1 @��4�K�L8�@s�����<��E��\�e����C��i�7��˞6�&���~��X�<�n�5G>Vd���K�Ƙ�
�uVY�G�s���oq6x��\���>&	�ț�f.�x�LS�o�DL�7�m�ЭrD���р�@�
>�b�jUw��%������7���Ϳ~�ˏ.=:��E����_���X�?���k��������xb�NH밮Jv�K�Z��0�d���0��0��a\�f��+)"gC� ��ؖQ�.�#n�����G�9˹������\MXqN|�BM��Z�B�����#pb�N�?��-�_GH�Uҋr2�L�G%"\l�68��K[4ԼnO�VcNE����J� mF����.� 5��@3ے����lE1�l�_�YXl­<��8	5���~��y0@��	��f˳��g�tH�g�6x�v%h��/��tN�?bs����6o�<e�7Kd�P�Ψ�b�}�G��&�G�����'�1���1[>|���9x�0���^��/�́����#>����M��Ә����e�|t{��Of�0������c�Q�@Y.������q�#l`�or-�nͧO3T�q܅H'���˫�����9.�'�`�^L�����U���c�?v,�9�vN]�W\2y�4;l����w�pVӃ;@������Qw��D���#��6/W�=$^�L�»w�5�/�q�y�l�3f���o֛���Y�J���L޻u5��Mz�4~�_�j	�a 05a�I����������g@�����o��g��q	O� +3Ҳ���7�J}>�)�<�A	7�֬ЃFS�W�� �/�?�7e,|�F�M��n�x9!��u��ȁ�@�W�ް���:��Y�����l޿�y�`���k�xF�������p/��;��i��e��
<�&��oR[�Y>O]G�g��:�A��0����-Һ�f~�k;4w��4��+������K|���&}g��(�Z���}�Y�d��o�8J���+� E� 5#u�e����@�c�0�(e��]�!V%᠌��<hQ��0-�|���rF�6���Z���B�Տ�7�8�1�;Q|��&��C�`�.vփ̣`��g����V�)pP�~ʞ�'�^n��?��;�(x3�)x�}�a��M���,�kξ�y�a���wD��2@B
|:��I$���d��lKn��
�,��{�D:.�i����6�V�M�%l�/� �Ԡ� alй-���g:
z;���� /���R?	7���j�U.����6����(�_���$�Ә��V&�v*�i��>�ߙǫP�NY׏FC���5�(�N�I�']f��7b�'�W����yu��-\��J�«u��ޢ �p��������5G:���ޅ��5��7;;"c��{9���5!m��֙f;�Ca��.�us vd|����o����K
/�Eng8Gs�dxL�~�������o���K���!8����%����6�����!�_>�hs�3���:���^�z�yʉ��q����0�������H=������_���K��[x�	����W돇�zY�2���⡙�Ԋ��T�����啴�с(�����2ek[SV��/�W4�4�f@����C��zs��.��vD��z�8�0r3��P���^�=d�+���c>ςδ�8g��T�|kZϼ�$|d�}��DA�}r�Ðã��Y���Vg>��*�ٶ�~0���x������������=�Ə��r��k	mb�k(o���~BdbW�_���X���<�d���#o���1pM�w���T�S.�i~�"4��g����G�O���#�r+�&�ȝL�^�ߕ��"}�	��Ѩ�?�߆.7��9��l��=�ȘG���|���3^���}S�8F��mE�� ��>Q�m'y+�z���v��߿DQ���oN��N��<v�����y����pf�\�@�H��eyhv����򩇎}�����'u���gO6w��s�#��b���D]�#�'.�茋�#Q���WF\rĿ����d�!T��e2���r�af,o��N=�Ҿ���Sf�P��};v��q����ė�D��?���Lg�,�b���%�t�㏯7_}�d�g��~�HV.v�4�Ƙ��>P��PB�X����1�kV��d�p���O�6��>0�A25�ŭ�uҚ��!�b�I�Jl�%���gރiF.�t�3hhԄNԂ��7x����1�'�'�k7����}�6�r�� `����i������ze��S��o�x���Y���䄺Ƴ��n�ܡ�< ģI\r�3#�U^�*<��1��rYMq�	/8J|1�g�5&�0�{h<�˾��)��WB���k� o�����?xO�&Td� ��L�J0�&,
�v�&X��3�����̻��|����w�������"
_�џ���sX����6����nn����$��;>c��v��GO,��,�v���'��<�K���p�����?�1�t�9ia�R.��z/@��?9ρ�*���B��Y���<����ʸ�.�x�n��I���8�"�%=?��O���/�; 1�R�Z9"|��.�p���X��Z
�tK@�c��:7t�m^�p�A�wt�^�ڼ{�n��v&����,���63a\P���{���I�6_�^������[oQr�XF^lL)���y��Q�pʇ�ƒw�"�[Yo�M�M�~�>7zrj��_^�I�����x,g����5xF���&1��У#�~����*)� (�KtP$������Z��&?���P&:��%} ��Us�Z2���<OS[�D�gy�>�z����d�;f�hz���/}�gF��=V��O��ۋ�d]�]/#�q� }��S���y5M%����W�ʷ��mX˾e�f^��W��B�5��\C�A���@���  @ IDAT��3�=t[�۪�_�|�+��p}�M��n�� S���� �-z.�y5�e4����U2�4K1�V��P��%�pȳ�����hs�P��UN���tF˷�T�)Pa�@%MZ�<�y�M�
T�ѺgԼz�)�/6�˷�o��C��ˎn��G�u=����#N���톺3jL�Č��	�da���5��� Z�+;P��e��V ql��A�\�~��
1�(�@)�@VoБ)cfT2�� ����)\҈��	0���gv��P~�o��D�o�x���I�5���/�Z�
v��{�3���w8I��CҶ�.p���''2�r��´z߄Im���`�RraOE���4�P��5�dm��g(<!>�"���l�9�� �r�>	|�$�4|�+�v���T��z` �(x�֠r������AW?D��5�X�C�����10������e::������l����o����P�;f1���V�oE�|@�X`2�;{����>#�=g��e�@Bg�s��#f�<K��ǟl�9d�]�K�|}��Y�<�H˦[򗼃b1�@�n���ua^ ��:n�<ÛT-�y�4���O�쒣2eșlX���#8�����ٱ�Jݱ� �Y =�Y����x�YN�G6�1G��{���e'�u�O� x�FaV��zɛ��'RM;x���YJ�þ\X���W����I�A�{���V��4	�nq#l�h��e����*/�����:�\5J,��hLI�n��!�3z�Jd�˫ifK�.�.����X��O�C"�ű�e��V5F����v�j�G��w��H���P&�Ȩ�8	`:asO����h�.��]�n>�G��6О�E�' έ
���s�j���׼�#�`7��x��{�v�Չ��Q��0�jwX�;��>H�
��v&wd
i�u�s"g�@,���эƥ����2!��^���ұ��	/��z������N�ϫ�?��v6���GG�b��2��M�+�#���k���Ja\C�%.�MXo��Y��L��iLQ�*o�J�[��sڨs`#�)
2��%be���*>�����	ni82֠���S�a�������|��|����
�b�Y/��9,�����{���Q2��L�o�����֧ �F��͠��+�"п>��<V��f@�#�)��j�����r�	��M\�Q+خF�G@aC������m�֍-�Q7Z�>����^�]p��3�J~���BC5����nL�Gҹ@��s6 �9�&<,�Ԫޭ_ԽFp}&���&_�'!o���L�t����f8=?��h���v�A4d |ݔ]��@�(@�����5������|�@�Q���s�C>2+f�F�o�yb:׎zF׸�'``�Mh�#6x�:�-m�Ӵo���[g�sz~�h~� ������E^-7�Fq'��)3� C��]���Q�g�����0�|�Zc�>K�9�*�L+�A^�ǂ�@����	!�\�ZC��#FTss��oR}���9M9@��,��G�'��<����c�ɫ�uL�β�a���� �X����bsj�RQcL�s��\�����ׯx���;��;Y�Uv�g�
t�]v�Y�/�yS�;]!����\�(���r1�+<y�r܄��$������a`����Bƨ�]0�9�o��?�g�M0p���V,�i�Ev�M����"�[��[���Z_Z������#�D��{�/����^�!�h�_�Ľ&]}k`�4DDa�n�������3XzO���f���.��qrƗh�t�gs�Gh9������L:��7�6���硧�&���g��*� �O&��+d���g�l��x
kZu��@��/�Qn�q��ζ����3���%��cl�!1P�2�Lhh��%DЃ��%�b��(`S#�=
��}�m��_��)/���QZ(�$�}$��H ��NU^�	Tp�s�g���BC婀<�C:�����y�o9���'/���%���a��*>p���v������0����X^k�����l��°�@8NY�rK��I�D^a�`����:���L���a" a��3r����G��$~�Y��9��⹖ddeb�},-C�����߁`��ּ,�?�8���(�L��vTϒ!D��:� Ľv�T�o:�!
�D��G~�8���y�у�#*K3����y�9�-��m�h��3��3�򹖃�l��^FX�wJ�lpK�B؊�M�_�J;N��WK]0����ʡq<',��Ф��R��$'�Q~Ҥ�d���/�?�\|�#"� � �hR^��h,
�%93h���D�r�N"J���˒����<����A�BE�8�%����Wxߤ:Dg�px���M����r�Hϝ�!Mz(��o�^�}��i��`v�y�����\FQ�y̎�8�D�W%j�c���W)-r-P��a�)�<[����#��O�� �L<�V��B�?�˃YUƤsP���wV<�g6���H:�P����l~�^|`��Y6�5������;�Es�����u_��\�h�i��3&�y�%��>.�3|`�\i�����pg��a$^ Ir�L����+1����Yg�����P�cD��V��5�~�~!ƌ&��Vy����|��x\A����`Mh��nT��\6D3�Ĩ��e������`�z�8s�����m�gܕ�I�߼�4�7Ǽ@��I�g���d����x�f�{wx	�-T�E����Ŷ��I���Cbs0��^,�g�5��=t��m+�CԷ�)cm�`$�;0���:)�^߰�L��V���㋴Sb۠w�"�	K���M\��������.v4�@@sL�MeSY�*�!h�-Ô�4����idE���e�xvNE����"NB�g�8�ra)��)E$q2�܃Xɩ��(H�R3�~Ź_Ϙ���'���d����Z�%�c|9�����;�|���94|V�n����|J6�	/7$�,9�.���6n܊c<Ѵ�SB8<�[1��;���1�O S)M@��1�������|Z���=y�N'iWD�Y�$�=<	�[�I?A$�r1�q?�d"����`kh���F�}0
3�D3��1
���~��F�>�C�;�cFg�;|k�Y�t}Q<�S:�!��y���:�ڢ�W��M��$N�L�����r$>��N�vۤ胛���	�D�Oy��@�?K���T�
,��N_�޼��6���<`pst�^۵�X�N���,�UA�`���"fAR�Z_Ut�ȸ���t|C��J��l����F	
��2r }��r�� L�L�?ڷ��h����^�������yq��z�c�y�%%uG#�oV*�Ag��U�c\RO~��/�h?aE^#����8�@��0E5�ɜN|ҕ/�e̡�J1�HSTB���^�ѡ�2���K}	�>8���G��s���|'����KA2�����e]im;����/��\&C� r;�rS�f~�	� &�>��\�4�� �ǣ�uvٸ:e��g@�'��@@����3|ݏfY)(#�ff��CK���>� �,�2#�^	Z��Xi �20	�4�(o.u[�j2]��O�:��z�z=C5@��Nf�Hv]��'���y��9�Y������g��v����6�$�g��"!�uǺ�"�a��瀺}�2r��[<���p2�!S�4~�笱�G�ܖd��'���%}�L>����]n�,_�Y��.=2+lC���7�9S�����BOq���͘Q-L�	S6r��U�6���C�k�*�ʚ��8��%��cJ;���l͓��HV�� sWq҈����3��y�����c^c��{�^�`��5���l޼�3',Cbe_p�o��q��%{�.�r��1�vX~��0C�ó�9���+ڷ2yo*�����Y��[�F6��5~����o��!���Z���4<�X�0��"A4�$�fN�O��݊��26�a�������w���4
0w�!��5�[���k.���a|	�̢����	��U��!6&*���dm�.�uy��B?f����=F�v��^���z;��p�A��i�N�"���c5P���@n��+l�aV�SJ�;�	�?��K���ϣ!āOd���-7�-���$�����A��M+dD�y���9T� Ck��ێ��g;�IZ���/����[��}���ѣ�BE �.�dF�r(*�0�d'�MM٠��	`�yb�����)3ma�=�����Ͽ�b0Ҷ�-�ܓy�Z�*(u�ᐂŴ��]�M���4o"T������6���g�I���E;q7���j�]	�ܡ)]᥇��i�a�|:&.L�����-��ų{�ԝ�^k����8W.�?��϶��94�7���^���p�s�7ӭ�.����T�<���k����3Ӿ��s>n�8ˏ�;#v`;�<�F�kȝ0v ��� e$�̈́����m���z��$�Z�K���*�A�Du�ݒ]x�|��Ad�-tFR![y����UbfL��'�	�?ւ�)݀DL0�Ig�+��:`8�A��1���KA���&&פ���#����p�9y��D"~koL�xlf�/{��=�X>�;u�}זE��=ܝoBZ�.����퓙
��|�-��9�g��"��P��ݩ�5��A��M�Z�0y0�������q�����H3�nڛ�U�9�&<��Ӧy��t b��!���H+�i�}����5I�c��To�I��܀)��,V 
E�2���tb.��ld�%��3`vD%�[�6B�C�F5�ăSX91�F��װ��#���#Ø̪'�3v9��e	?O�Q���Lg|��{�^d���֪S�l�¶�.6�;v��i��:��G��臶�o`����[R�a��+p �Kc":]��z�ܟ$���6
�{��,I�� f����S.�M��/�-�����D�<q-
<��,���d�ְ�n�#,�1��$�b���F<�S@~&�'����`��"�BJP���Ɍ�H�C�&�r��E�*#d���̮^�ʾKg��0�j� <�௑e;�|���0UN�㦠�ζ�@H��<�w�.�S�	_��eAXd>��N�8���B�\%Ap�#8F"��rXf�TԦ��c����������_0�X���$:�8�:KӜ�HJ~��K�����G	C�7�~����3���ޮ�O�r�bo����$�B�<Ю�\�Q.��3<ؗ��N9bxEgq�؛o��<��?2����˪T�0�d� -sg%���&��)��*7|�a���;it�?�R��2'��!yқ��J��)u5X��1�Ɏ�g�h�)�ěd���[�N�:�C����q>�?:��܏q���.��jR�� �\9�<�KA����+O���,e��o}�+̬oɦݏ ɲ?��6Q��|�k��޸��0ϫ,�7q%��t�E��g��|i���G�	1��o���22�(
P�L��>�G��J�-��ߊW���l��M4�Va���T���,FK�x/��`_���k�|ڴ�K2����I��o��3�CW�����&pF�I���.��+w� �%>�	�\�Ja�5�>ǘ�[��(p�S.��ن��ٴ/�m���hj��E}�E�����F!��[,]ݹd��ps��������]��05���Kصz���gv+��F�3�&�(D7�j�Ȟ
#6$�Td��_�l�3�t֯�YC^0����������P�Ga��X�2>;gs߹Ɣ�Θ1*�(M�{ʮ%G>�D����GN�A��O�˂�!	_V��e�3��$�u
��ĸa���o^�k���C��|���q�U�"�<R�`%DŢޤ��Z�Yi��P�g��6�%���5�E���i�u�F�`�)n�����x��薴wKK5'�����΢�	q�~���;A���c�w���t�P�=����=����ٕ{�Q���Rp��S�c�AX�G��b���N#%3�U��uyF#n�p�o:�B��	Cd�R�Wf�ҳ���&kZ[�mm�KChe�7�G��i���v.�7�������?8m����?p��o~����Վ˅�����p�գ<X�����M�:�Q���ޏFsF�Kf�^|���=�6yUos�@�����_l��	��M}��̈:CDB���#�W�ֲ�w1n�3�.���_�?��y��ā�?d�.�]ԟ:f�2���4����F�	A��������@�,9���S�y�֝��i�څ���c��M��zk����*A|NΧM�c����k�d��9F�[V��{�\v��O�/?��JA��vR�o>,;pJ׺�>Eu�Y��s��La��]���L�j�%jq�*C�3.e����#ƭd�|s%��k����
ob�ǫ��Yv�b�������O�W�Oa�=uV��"�X�(�o���G�-�MD�7q�g�K�AW�ҧg�%�2\�h��d�t��FC̃3R���
��d��P�"�	{�/�-)�|r��RGINL��0���<�k]���~�9H�|~���i��5a�C��>��F�_^ �hO�S̨cs J�P*��֣�Ǽgy���s�����Ӈ�S����kަ�����W�6o��s���8-�(��P+Q3b�ԕ���g񚉬��W����!�@:qڑ�.U�t�͸����	^���b̑ޅc���ۨ�� ��$�X�\�d���e!�֧�̄�;#���U÷̹J;��hŝ�֊>q)�g@2��BǛ|%����4�7���Q6�
�4`���G�LT�Wej@p�(i��Jw�%�
�V��l���zO���G\n�!Ϊ�-R��<4|2A��3���jyNh���,�CJY(]�݁������l�M-M���|ڇuT������/�.�k����<ɯ5^�xyY�!ގ�M��������0��d6pН��a�w�
'3<�ʺ���o�O�x2-Χ�O���+;��Fr,=S��5���fj��3���/���sڞ�ruugVfe�6J$��y_�T���)���� \ �gG�E���Bw��p�8a��ȆvL�8D��>�̴>��.�ₗ�YH��8fI��%[v�m��:q�7D�R�����ͯ�X��i��C�wO�Q�gK��S����<6Je�v�D."�0�7�g��N����O��z��Y���?/>���b�[�g�Lg�ox�U�igd��i�Փ�XF�tnZ��d'��3�Z0���Yǧ����
�7�J�c�z짒��ڟ�e� �C�$3�S�� ��إ1��p%�{{��~�ҝ��ئ�y�F���v&P����b¯���M�r.�˗p���ﰥPE}��!�SJKK���Ux$�gmG8� �X����/PbG\�#u<v�܊���)4-�b2�}VPaG0:��+x�	 ��)W`gd�S��1���7�8b<���,�qG���IR��y��T��HB��=)�� �%�;Q��<z�ƹx���|����ʍne-H!�3u���C	6ϙA�'�)�Gid�N�I�	��UCN�x����W|���L�ޛ�/ڙ��{��)��fh�nhѠ!ub��z��fI�7�f���>%t0&�'���}�J�Eℬ��n�8�����C�DD!��B?'/�� �N%���#; ���K���sec3��g�9,CX� �h����*G�U��D)V|�v^�L�p���9ӓe{	Zg.i��N�w��F�.���l�9�y1�3]�:J��/�� J6�&���f���7`�����	Y(���k��-5��Z�����@՗+�Y��){�\Z�14��XB+7����&1���y�L�s�p��"{i��}0n恞�L���LL�9�3K�@]s���0�	mh��k~��[�ߐ�/<ץyp=���چ%�=y�D���������<+�6Ɍ���5<�	�ʡz)~m9`��8f=j�΀�15��Gu_�y�)��Q�؆�*�A�q�0��+��#a���z�yJș����yL�U~.vW�4,y��yC0��){��sxxɌ�3W���.~���k�fѿ��?.^~��4��-�����>f�z�32���5�@�������/Ρ��Popʘ���?����7|W�ǐG����m>mTˏ����i���#���8�o�q�7�7�������ݰ�6��ZV��O��EF�;:?����ʢ�2X���/�<�b�v@�@5�-2��B���y���-�zUTy4C�/��5r��x�U�6�]�s^��n�<��Z&8E 3����7J�A8���+���}��/�;�-=�Y�qJ����\�M&�����/��&�[�.�&��{n%��G�k��c��[��$3���=r����ԟ6�}!ጊeN���u�����g�2�kE�t~r� 4���2�Kt�O�0fdLz��e��(������ĉ���hgq�ц��;�c�83��"&��ۈ����n(p�^��bHz�"ԎS���1�-�P"m̲�Bx����h�(uҵW�Č�1�bIY�tk(߈�F�k Gl��Ҁ����.�rN���6~�!u��;����>ZL��ꭇ����7d�ǔ�hZ�Y����0�6�5 ~�D:�!ױ�p��8k��ѧi+".��c���M�.�ۉ�Q�)��'̕��@��%ڣ�-��T*��5�u|"��Iv3���$��/��� �!�,Fc���!�3�b,��V �
�z�7m v:�8Z�Gt�̗������t�q���!A��B�I�-����."�,ab��zE�|Wy��(?��7��N�*5�
]*��:;�4��id�0F���bJSJ�z���3��ӹh�!}�ͳ�B��,�őbfc�ȡP\ΣhA'M��H�{_�Q��Dl��@h��a崓��s�L-�߃NLP��9�}A��\܌E�[A�|�2��Yi���&M��F��1�獂���6 ,O���&]�)�Kf�jA&\���L%��N�gIw��gi�1%�+C���� {�и	ҫ,�(���{�JJ{�RL;G~/qX�����z9�^�Ns�7��{�z��Z2��<Ko�������Ѱ߆�g��G���'�!�~qN��ۆ�����C������V!��G�oV̊��W�݊"/N�����Ku䑚b�e�Z�����ǿ���'n���E�y��d�l}�Y�t<:����q,"�lWq��v��@��Ѣۆ}E�^8ٶY�]�M��T�O�)_V�``ж
�f��#��,V���I��t��Ga�2-�xmU�ղ����>����;�},n]8G�^������Y<���Ƽ�%�9���:V~��G�-@��<���6@Q��]�u���C�z��D��A�&�����LN0"���$�K)�ۨ�n�??8c���Cx#���HVH����&@��l� �8�h��枏T3W������}B�'8����/�Q_�۟�+}��L��k�f� �yLK:�����}���rK�#� `��.^���������13]�~���u
�a�(�]����x3�%o�1�r�gF����l�˚�f��ZA�� ^�͟��j���E}(K��Q��,K@lT,��8�����%��_���F���49`_�- Dy-�ډрM-oy�3#ў�����8L��ʕ�KlB
��
�+(�#F���Rlb�����Y>d��4�����ř���f!�e���T�bj���/��<"95wM ��T��C�Z(|0J��`��t��I�*iK�^5�KhҘ�����>(��+���ct!zM:�m��?�&�������<��y�	ݳ�5��qmLG��&)�p?�LE��0_a˫yt��������(�WJ8�XQ�T�b���	uԕ�����ݒO��O}�X�F��rK���?��٘�VȣK�i��Νz��9�"ξ�<�I?�G��k`�W������A��	�7��9K��2��m�h8��쌷l5p{�����u��_����p~�%q�6Y|�����ᗟ�lipΎ�>��E�=��Ɍ�W_���?��ٖW���֒����{�}�6�C_��#����]A��o���������b��AKp�^�H��7��~���K�N8�3F80����v`J���o?��O���������I��������m8��;۶���#�3�;�5"\S����:�/����Xߪ}!��iñQ�&g�V�A��y�(�Z������:���?ؖ��'0ĖN�͵�vN{��r<C�&hZlՎy费Q�U�A�V��k���6�)�݈-�O�<���\��KWس3 �����.��d�,p#g��M`�:��ڠ���g .��ͯ�㨘����y����^��)yo[3�ףe�Ųț���3<�9|x�}��(�0��2o�R����o˷�y��c��S�����^���q�/�A�v�?9b��}�c3�c?�5�`���U��g�^�N;i�)�8��)h�ʁC�k�R�٦pA(-��O��Dtn_�ma�N*PG0H�:��93+NYlq�T˷٫Ce�z����(?e�&>�����A%Sq��q�� _V��;֓�M��EyAK��o8@_:3N�Y3u�#�b���ct(�у�s>�tdf��#j�`ǒi?�O�3I����3ם�1�?�F	\D�����4��`���U6����	S0�MZ?|xXN�����fh�����p�8e�d,��W�&��̻d7�F�{�4��`�zb���a[�׸�U�4T�}�����u�����A"�6�0���Q8����/a�6�Ƚz5>�Ly��s?�pdJ��I���g�C������F����+>u`���ýQ:6�O;
>�O��P�+�9��Զ�,�Z8�Z26�ď�E}edc#0	!��>
r�#���Y�v�M}�:��%�8d(�fɲū��X�9�h}����D6 o�rM�D��������q�%3=�>d7rE��:D�7|ؘ��8{��
��ǡ�ݰ�%���V4FG�V��q�������/��g-&�<a���͇Œ�[��my����Y�u��uB�{���#8�C���Sd��1���_7~e��=��7�G�ǞO�|R�G��/�\��L���J��0��woxT�I����m(�U���Ro#'u)��9�Ge�`�J��l���n���Kx����)��ߨ=D��i��xp|L�ߍ�	mM�I`0�#4�:�}�y�gU���&��۶��Ƚ�eF�v��`�%P��B>G\�"�y�`l~�,�&�ϔ�S�S�%�,i׵�� ��lDZ��_�v�rr�r�{&x��A^��>�8΃_�իrOP��{L�En�OFЉQ� ��Y�G�	d� ��ܧq[�懂��,r�`�Pc���^{�#^��2 i�l�c��f�cN��Z��b�0{L�zá�]g&���L�N�vH��h���R�G�Y�4JG��Vɺj8�)�r�qΑ�(��-6�ݪ�8>}�j��#b"N
!0eZ�e��޼J���q�]D%�n}�fD��\p�42�_с��sf��v$�C� ���q���UEޟl]嘌��la0��Di|����-Rr�KK�&�z��a�8c�[L�L�x�l���CA�=��&˰� o4ri����ę�Nk6z��C�i�8_�k�#�(ؘ�M���a,d半�.����0���1���̐�c���)�xa��3�,`��a���
d#�D5��M8�>N.޵�h��H�󅬴��2C��^�#t�J=�6'���y7Cc���L�\���9����AJ_�&㔁�<�/��h�/���9�6�
�!������\ȷd}{�G~'t��`� ��	�0UpH���G\�B[�0N<P�
��{l�����Ip�g{�Q�]�`�ԍ��̺��|�ݷt��APX��y��������*X�rY*W#�qjg�:�ڒ�h� G8�:��0�$�T��l�l�a�s�bn�R<C�f�8uj�3��+�{����'��ݷ�oyx���N�z�3f̖̤�X��a���%� �ݵl��,&�v�y��-+68{�]�3/o`J�5o��Q�rq�L�W8{~j�/g,����Φī_A��el�2�~�lÌ:):�@c:]B�S������[㾈��x�eJ+�G���`��u��afd�6���1��Aa�}OPr����V��J{YEk�I�e�`�����1�gF8;��ɸ�DL��:m�ًl���_\Jwfd�S��]u�욵����u��U9okW�#;;_��<�J ���W�)� c��
��E.�Fh=W^՛4z7��n��|�>�L
���k\�B��u|�T\�_!$Gˊ��o�va�k#5`vhc�ƻ�1� �s����K���N��	_�P_�l$�ǯ]�in�*i����23&ƒ�K�T��4����ö�3m!��@BK��c���G�ԑ`�G
�
���6:�y�Zo��-��;:	VJ">K&R$Ȕ7G���u�+���+���=q��м��G����U��݆ź tM���V���m#6{0�dq��F��(��rq���b��mc"ma��<�L����٫��k`>�jI?��+:� � ~���"ou�,ſ�XD��N:�^�̷�t�ҁ�z�rZ@�;	���kA�p� smTr��
U&~&�����,���k^��5�le�\\Wt���i�|BG?Z4�"r�K���ِ��GB.N�����o�=��@oS+��8+�A�g(��Ƈ���:���3��C��/eK�ģ�d�;_�GL:�����SMŦ�Xޑ��c�m�뺓�zX9G.�g�\zz��Zx������B�mn68�9�V0���5���($�ؤqo��:����3�s�q�q�"$�V@�/�`3��??ѣ(D ��3q�Q�&�
�sA��-�<���I��6=���$�li��H���/������%1�l�$K���v,X�ể:�8^�A��5��6���O: ~oҷ�q�������ʂ�^l)�f�t�С��� ]��k��.ܳ���yu��w�7,�y�oI�Z���?����! }���m��Tn��cqLy:^�m��'��m�OF��#+��:<���̈���*'�$�Ag^�E�$���NT�HA�)�v���2��g�!��~�S���%yT=hh�"uF��Je�C�S���K;�2ipV����I�E ������?e;��7h-]j�s��En{eIC�2��0r��O�@�|�%�pO�җ~�����)6М�?�%����gI-�2��1�Ǳ�3��`�v.��|��3��8Z�pp��K�M:s�oS�/n8yB��6b (i�m�xm��o�k{$ťi�7�5'S֞DT�s§��GjY�r턈�D$^*C�xX�{��k�!.�	�:b�	 ��G������0��ŮA�v�aY!����-���R5IQ^L
]U���%����@A�+����������#)�� R�΍�DcdPEٹx�Y4 '�Ȣ�QI�o�cd���2FR����#I���)�Lc��4?;|$�}:Tx�&�S'ˢ���r��I���9T��)TA�Fg����}�1�`
C
���>'z0G
�]�r�: ך��on��I됹���oQ�y��bXc�X�����|Ls ^���F�,�����{Rƅ�9�yzi�=� 	���;+���X`u�z���c�?��7�����J�einZl�ї̎M�)1ؙ�Av��(+�=*��ړ&][Q�s�h����1o?������Fup�g݋q�ґYv�C~l$��bff�yz�f��(�C'),g>�� -���3�;K5�P�O%?�.h#ʃ�'�8�d��������~Y�:f�H�n��G7�C�	Y3S�����<��pF�8'p�����ݬ3��"�������w�cg� �:������L#�N9q�.�$��8?�qǢ}i;��8���t������j����V�n�b@G�^�@�+gW}=>ߠ�ޙ�Ά9��g�\��K
æM�F!0�9�R��� >����L�z#ho�j�#[Y��]pf��2�L%#�8����y-�sf��s���6��Ƭ)���rM$,q�;m�Y�E^?Ɲ��hw��5�:aa,K��Q�pX�������Y�l.Ni�Iɇ�#��#���)��}"���dʙ��?���!���u:SHd��s��"��'N�	�b�gLΦB{,3����Z>\�fe�qt�Bpĺf?��'}>���{ٿ���5�qvv�x������X�z��u}|�Xߎ��\<"&rѝv�^()�P:>u��(��V�K�tƧ���K'xZG&o��VF� ���z��sw��t��F� �)a�ɽEE�\�\�F(~��=^�O��R���"��4�G��L/4�D��7����?�3�,R������Wôs�������.���yў�I	 ��#K
�`a1r~3Q�b��y�7D�1�1��gύR�TD�(B1�7���J��ZY�c�I�8j"d$m:`�MN���y�)u��U�)q)\P%B3X���H�W�����p�}B��{�0>��g.��,��^	� �@���<rt��-_���_/oiԁ=Ca/�=��#�1�|�f��錗�;fT��;+y�j=�-�#u�9��JS��I%O�F�>�Ce�����!ס�����8a��,ׄ=0[,Q��ĩ�4��� �>�<�N3�=W�6&�|\kW���ށ���v$=��q��9��bv�\�90#�iE팅K	�)-TL-?��a��e�|��A�d ?���L����C���M�'sJ��P�"��i�#@i��｝x
�t$����g��4��\7$BX8[�MO1L�ou��{v��)k�R?KOlּd�#ppѱ���_�&T/~��G�N����ܩ���Գ�m��|l�Ù�u3�<�������Ĺ�B��sv!�E�=�fq� �bM֨:�E\�A�M�	��-g�7��`p�x�|��*g���8cf;��0��6���{Q�wF�r�jm�hW'��|x �Rf:E 2�6��MqA�����a��g��p�^y��1���=�YG tP�)d�y��+n��Z�Neu�e � �m������4�N,�#���MQ�����DM3��i+�ýrɅI	ZA�Q���-,a�I���	K���<nMNv �6���@Kv� S����%�Pe�%u�k��z}A������g�3�O8�;�~mz��-\�m�[��-[�>�����i0�,_��u�f"qI��W�#'PrC0�f��0@�k�YL��)kȏ�d��Y:�E[ӯ�e�:�H�o��+q���k�hJ:����8�����;fA��G�И~<Ԭ<b?�9�+}���^�-���p��sԓ�.(�q��4�FC����Q�� �%��2*�@ �#0��5���Sj�U&X���-l�H�iB��`DNx�V�pb��c��ͯ3����n<�Rq�$%N�i����x "0� ��QY)��R�{-?f���r�댵%�����ϋ���r?P��������6!��c���Q�-������DQm�K� ��]G@`S��x#��w�<40h�~������5��:c{�mS���z^aB��$���@Sn���a�lb,�-)�ɷ�p�8Z��9r-��*<�eRq6��śEN秃cKw����V6�#��g���ƌ=�xv^����Sq������J>�r���q��_��j��LF#m~�y��������y��U�̐�)�)�$(��Am�c�����4RҮ3�Aے�a�,��YWM�� ~ivv&�B��_�R��>e�s(�Ӱ�T�Y��^�� f/�L�eJ�2WN>K� ��ƴSʍ�A�c|�̊��5��A��t*j+�$�sf-���E�j�.���9�w���b���gCG�~X kڠ  *LIDAT�šÕ7(���탼Bm�]��e_n��_n��8q��|L�_����t�*_X�v�;C�c�@{r��ܫx]���ȃ���������m��R]�F�fO|�r�,��n8����E�<�T��Y�N�����>9�eZg�����o�\����[�U�'y�gy�5��/ι}�0ѧi���vI��Y?-G4jJ��?QФx)
���`�g�8k�)`.��#ho�Ѥ%Ñ��4d�-]�`�<� r��WxBfh8+��T���Ж}C��=-_�M�������{�1�-|��A�oJ����o�r}A}���]1 �I��:�\Ә�3/�%
xe�`8��"���;2�8wdA���|d$f�)W#-����?%@b�|s�zg��'<TH����=Y�I�l�&g	^�zax�Dnȝ<�~H�0����U�=m�;�ѾNh��=�����޼�#p�y�5P��Wa���5b�j�R�x-ى̵y�!ȼB�?g�#��`�V�� ��)�r$ �
_�r�i�(����16E͜��C� )���RR��D�O�rcNe2��Eh�5��BSg�\,�Ǎ�~]��]\yOG�f�o�������|����}^��\}G�z��DǽD�΢�\t���lBe`e�*��/�FH���+�x?d#H�y�Q�ʾ�l�If��ר�����M�u���ׇ����IcM�������`h�j�g�-2u:8�G��p\�H|L�GB��C:Uv���������*؋����l����O�:i�u��,EQ봸/ԓ3,Yl�5�1��Tp�T���<zɬ��R"��,���_��2�0�=��3mjXl�z��������a�k�"���I�ٺ�kd�}��kZ��6!�*{��H����V���8��@���7�9?yq�w���A"	�J��}b��N`=���z�.<�ulJ�7NWL<��K:!�M~`�/}	��3o��ɃT�<�Q�����y�H�I:��E;&)�Z,c������r�R��A��R��X��ppptT���Y9��S:m����t�����	ʧ^8�u��}��L��H���I^��N����_\��s�SҜi@���\��ϰ�: S��Dy7�A��*Y�@h�?�JS�uUI�Y�C`�grYg|a�q�K���2��x�N���@�Y�� �sP���m��?"��C����K+1�Mg�������b��bC�K�����x:�qdփ��M9�?�q%Z����	���33MȜ��E'`f�>:p���C����q���-�s�א��)"�;�&�~�l˲*e�T/�{ʋ�{Ԏh+h��b"��*���r��=v�Z1Q����\��)����5[�/]-*0�J��œ�7#Q�iD��]��zVike90N,A
��0�D8ШF���I+�a�=�W��A�eW�j#��kLkY)��B4�b�o~�K���4s$�ye�К���D�&��V(�� ���U�pGr6�+d��Z�+��OQ�ߟ��+u�xԵ%�Foɣ.���KF;g:`���FKeR1��4(���|{&���I��	MT�yo�k�gБoDpJIS�.��LJ�ا����ɮ�!��B�i��U>e��tu���A¦�o>m�$%g�\d8P�K��8S>&V�KXm?�>e��0�{�)A/�����t��e�:�3'��d�J�5����Y�����0�G�I�6���ˏ�����YN�e�4�q�hg���quN}�0k �Vf℗tbF����`��U��j�	�"W@8=��F�t��D���>m��M�Ȕ?��mV3�o�BFYn�;�����5'T�S�[?]�0m���3Cv\�x�3te�$K�C�틺�i�5�~;���9���2��ʠ��Oڥ�#yeM��5�Sv�#^�s�6��!���v�8;圗��� ��k��܉�8q��<��u���"��h�]��.�Θ����g�P�e����3�Fp�Xc�Bv�TZ��\({�c�����E'9m m��4-u'��i�J��M;�H;6���#��y�d�3���Sd��%n�I�ϙ�Z�vVC��m���U|��%�$@s�rc�Z�d��-s�;�7ȁ��׌�i��q���b{�#�v��\I߂D應���lǂ |�������.e���3d��p�(�M����<[?|7US��A����%D�Jƺ�}d���y��[��l��8y_��8M8��>�Kd�F�R��]�S�7���e�F��<�w���>hY�a�	9�P^��p��9Ƞ�vw�Ӻg�%'�~�X�3|�x���oZ�b�C&S���G-����(���u�u��~�.��%�(2�&�Dɤa��VI�z`zr@��&��\� ��X(�(��5��_���J�l��E!�:��4Mk����#�y,�+cs�u�9��D�3��o��t�'��r�^'�/���z��K�n^�c�ҡ�;o���o���X�x�
C\f�t�:B��M�ya���H�4z�SϥZ)y4���O�܀U�#�����<{���'>��%�4���mJKM��w�����kMMVg��py��Ǝ
�cTV~
�&��ʽ[��=���|{�����k`o��# d�@aA�X>�Il�n�#iӮQ����R�9�"��&s�^`��?�*x�!���k�3��'|d4̛+�Y��?����}�c�
�L}��5P��Bn���.��,����><����Kʤw`�,S�u�R r5�x��{��#օ�b!m<�H{A~�@�vC��s�y�y�,?D$D�f�B 	^�G;�dl-��s��6L��2At�䯞��zb�@��ë��b������BW�Sgi{)�@���ZZZm����2c�C�}���q&��G��|������ɟu���HG"�c@�K�/�),�6$Y���kC]��t��f���'B[Ҿ�NMy�]�����/�)Z2�@�@�M�&�%�<eN�3���r��}�t����Y
�@ ]���G2��S�������An�jɮn%pO2����ٵ����B��7�B�
^�<��v�d��}�%�Yv�V��tˁ�Cֈ��#�W<MY�-�����;	�̾z��l�W�K�&�4��2�R84˜�������3���̫!�~ ��2,����K)-"�tDrhˊl:o��ľ'UfS��^{�Q�svf� Bp�t(O����!�h��-OG2*�&a�m?�q��b���׷o^.�����fo��y#i��G4:[���G��oZ��>)1p����J�q�X�C����A�ЉN�3� �_m�i���V�BP�R��?�%kI5
?��يeIf��&���II�����%s�����~��8��y�'.�F���]���t����o��J���k�ƣ������X���Q!�����o˔Ύd�^�@�dY�9��
1��6p��֫v3�L���Ů�o5�R�a��.ex-���z8�#�'WVLi���>��Q��cc�c�����6��U2��t��_=����`����O?-~����O ��x���5x��� C	�[����c��S����wK�S�6γ���egcl��3��p�������0�ؔ��AXDq|b�_��|{��y�������8G8a���� ��1ΨtL�B:(���K$y���툵�:�Ú"q�K�$�iʫ8��NǬ�2�+�k�H�n��N=6���{���"��=�~X�N �-X�B����>)�gʳɑy˓~���Y�-0�`S��Fr�!�6`���ն���]ֱ)lH��P�R��8.+fQ}�*�O���ZzC<gu�����I�Bi�)����1Ηߵ���5m���؇�O3ays���h�1dy8}|���� �;���q���{���`q���|��G�w:dOl��M�~��ku�2 �Q:'�
f�nyM��f=s�����8��M�^������Z8b�|�C����2AQ}ki��)���;��78u�` g��۠;�5t@���nH'��'��<�7S�����Ƒ�cu��7�-y���
�y�AB8�>~|��|�~�fq����G��-a�p��P��؇�-P�]�6�EۚԦ��pR��'R�``5m�H���J-�i&R��6(���W��;$ތFZD������60�	���سr#�6��Ĭd�uh�A��zm�u�`i7���9��.���L��⎙�OT�P�����]�~\���4��ϱ-?|��0�r-�$1tvɕO8�P4HgXP
%Q��t�є�����A�"��5TKx/��_��li�F�L��⦁����t��N&nK�EMDK\<x�U�b�@%�a���U;y�&�?����-�<<�?�k��gY= ޸�`&��X����O<�:BY��M�M:�j?t|���D~$�W���{GC���d$|�1�>�6ʌ�?t��-�-����!tr��w���� ��yS�	ܫQ����z-���%��8��8mB38!b�׺epi����]čI�Q"k`�y�r�go�;Õ0;K�������??��o�/~���|��)�,Ч���NAˡ@ʉ]Zշ�L������1����2��`�د*��h@��Y���I;S�<�����֟ʭz�~#A��_��u�MGŊT��A9sD܂+dl��*fi��c��	��8J`6�3N��Ә�l�W����_��"��,�;c�F���%��ї��YL�YM���ǂ�]�^$цS6�}X;s�DG�C&�^��]��!YލX���J+gaC�"ˋ�<�9I���,ИY����G�h3s,�`] N9s�u^0����!�{�v�/�? س�Z;�a�qV>�KE�r�R8@ɬ�8�S��f-��O���A�ْ�x���C�J>��6#�,)oڡ��I�n����IG�����->~b^:2g�u�\G�G��X���l�W���yf@� �cf�t���at�4 ]�'��E]~t�8dzN��9�|�y:�q4J���6V#њ��d(�n�-�Z�t�2b6^Z�zD~�e;vd���KO�OA��C�;@G�%b[��iC�8��h�����Q<�?o��w�e:�s:�+:}�â�W�\���f�5}H߈�>|pd;���#��ip��q�]�jݲv�K,@�p�"N��6>lQ��d�:����|E��DZW��"q\#E`�Cґ���mS�O�������WG���#���dv�8e�m����휎�x�!mq�ɫNƑ
��w���ڥD����^��d �5_�~���o�^���Uަ��|�E=������B�r���ޝ��y�!���Û)<�+,�Ά#��
����o ���h�@��@��s��A�`\j���#i�����8����)�K9�\,/>��J/N��y��yxmh��{�f�d*v�.��5�-���}b���^���j{����,FD+*���˼A��6]Z�Q�X���y:����7�%�HA'IR��)��8��K�p�U��� QoO��#r$��?�9��,H��g^���,Sx��̈́��4�|��/z���?�b�T08M�
��@�=>�-�٘��,w��`���K�{F��a�/6e��l����t�x���o2� v�}�F����9wР��F��������9��F��1�_����kfXP����.j���)�hG�FYeSvF�C~�5u������C#�qNM�QS����w�3VY(S?�<�ڐic�C��93Oq��IÌuwzXz�(�}��j�3���U��6l�U���!��AŞ܊Ŏh�_;S�К��Fgo�c6:�r%�pN�ڂ�Ȇ��D��n�#�H05��"���%�Q�[�H��_v���D^���#�v�ά�fl�)WU�U��Jy��ox���9me3$ox���ݵB�C;�N��;o��=�S�0�ہٞk�:ʚ�m_v�3�����TҔ�) J�䵎<�6e�<un���4e�����\����ҋ�ϔȹ����gəez}�-^|C���p�6�g~�Y{S�ܴc�^<�Ð��fK��2����"�-W<iv�9��ٯ�\����.x�~P7v��O�
�]��+jB8�G1��?\��#�pvՎ�����R^���m�?���M���v��9+�7G��v|�l䧏}S���5�7�8�����Ҷ���g���6|w��x���>3�L�@���P>
��!�YO�$t@"�����5PT�d�AD���݌ۭ�3G��M6�2��X۟�{�ZG5�2��.ɹ�i�mJCA��C�m/��s[��x@7>W��n'��*_��kMAJ���S���C�,O֯�10ڂ����p^u����1�CΎ�p4�y����_�������8`���}�ݷ�Љ�a��c�z�|�'���6��Kc�3��Q`V��Ĥ��Hk��Q��D��(1���z�A�?�"�#A4�J6�R�_�y�B�5q�f-D�j����\��W#dd��T��v�GZʁJ�0^[��8���+�B7eZB1�F����a�+�q6��菆�]�Y�w�t�������ѓUD���%��ۯl�M�s���̢a�iXP��49;S�9q_��[�S^%Tnc��s<����`t��)�8e����K�N����!�8���X�]��7���ī�ᅿ4�T����F~7u�ଛ#�3�T(����f6�-�l]SQhx�QDR����8`��vΎ]�%��O4Z���)���H������]֩	�A�?��~@���.bԡ\�(�/i��>�� �g}��}��8���]^��.~�c՟��#G���3�0l_9Iw�{������F�"^�$�[|����s�d�1�*4�M�8��
��*Ӏ��$;���=�%��!+�w����'h�PVt%��H�	���a�)~p;��G���#����t�_�0����߆��]��~����KZ�8�ҁk��83��#�L��;�ヺ�ɝA�־{Ny�M��c�i�����T�K���7��z�tG�i���I�:)�e��d�-ĀTmm~n��5n�������83��r�.W	[�r�'Q;5�dfx\�O	��H���Q�
k��*���Ǌ��2�M�9"R��#S�"���N�Yi�>
��i?�o�8��ԡG�mg%u���
�����V̳��Ou鬄pjϴt|�7i�c��;�ș�m�v{� oV8���E�~zFGCGByE�r�eZ��|$�Z�k��~j�58�b��j�E	��>}۵6�n��GZ��c[�u�>�#����POEt�|��]L�T敻�|�-|�U[��٤��f)u@�bv�����I�N O�u�: =+^�Yv&T;qЩ�5�\A�pq$�ML}�#y�j� F��Jmٖ�\���˳�����A�|�O�}�K)�^�Q���Pf� Z6�>G����������D����R����gnO� �C���o�ÿ,���Z�x��|�'��_�˾ߕ=���!�^��>J87�����
���:x}y$��0L��Ӑq%0Q�,~�UvG8
O�5(�8�!-���
i4\�G�Aۘ��O�t���\�1()&?i���>��vh�m�T�ę'Ό��$l��ʋ�MErsHs�s�gC�T���g��O���hd���oq���b�$�-4:*�8_�}|���#`�a�3���� l���6��UC{�9tDү{�G���~�������i(��bC��r�F(��\�8:PXT
�K[F~\+˰av}�8*�Q��ͨ��a�y���!/m����=�(�-qH��{����p�x����-��B�Y8��A�a��8��8�7��}��I��Gw�ݤ�١�ʧ!S��**�O�훝8��V׊�c����eq����`������-�����\�N(��u�6}�!��x�C�Ҳې׹��*oEW3Mg��E��e+�ryd�'��.ξz�ˆ�7��v=�h;�h�:��E~�;[$L;���"ę 1�FS's���}eǽ����]��W!�En�؀�޴ÉO���x�nlh�{�k�>fs���������
�:��؀r��6lљ��y�'�vV%k�,k���Q�kμ�pVP>�ڤu�`7���9p���[���,E��De9�� O���b������as~���!4d�P��϶Ⱥ��6��9�,��r;��#{��ޯ��b���P��I^<�I�w `�v�BOf��Q(��$�ʑ�^u��{�(��忇ylw�l�3�
}�i�c&�R�(J�E����<}%=�g�;�����"/�8�,�ڕ4qJ�I�%��t�g˫�UV�L�l����dҨ�'?u��;zx��:�.�[�%��K۪-ESb��Y����G�v�y����o f���Gm�K��(�S���5����: ������N�
�v��'m�ɿ�2�OW���5�u�z�M�*II����K���<-ײ&]�Jq�z&M���>*;���a�Q�^\�#m�Wo�,���]��S�{���|����{���5/&�@hpl@�xXF�Yy\�i'��f���(���)տ�T*�7(4�ʂ��˼�F@[!K�Tf�KG���ťbUZx���ct �oi"?!N�ʶ �9�S���v�TpN;E�M��-��C<��)N�wƮO���Ye(������o����x�\�"�NUk�i*��Ɵ֟2lA����Q�AjE��+$���QǨ��^�v@Vi6��V�C_� (/a�T�;T���b�he�F#k9Vh��a3Hm�X+־\�7=mD����^҂��	�]�G�y���8`q���*-;��������0��FV��Υ#Uq�����]����^G�~T��aE��u�00P��Z+;hb�����}�@��v�,�_�9�1xx�C{�>�Ϛ�n?�c��t�i����Ӊ�#Ϩ{�_�:J��Hg�|�N�`��u���v�Lc�*8�2õ·M��.A0�����:@�s���u)�7Ζ8�-=�]j���|�K�E��aQ·�9�M:���`��V���E�����A^1��!��,d+�p.�8b����dv��	�p7qy�S
�uW�:=�eHl�2��~8�:��B�����I����R�tD�[r��:�!P#f�5�5dlG.T�wC�7y�>V�����Qӳt�e�a��&��K��cyҞ�V���[2�u��_��88_�}b�GNೝ Aω-��SS^�K�bNdQ�_k���J�N��XՁ6sB���%�I�����/�N���!^�ڷ�i_R�&m�w�Nj�LȔvK>�Gt*�@W�� m�^�D��M�T>����t2d\h���y4V�X'��=�9��x�|�_��A���`RQ�%�L��}I�C�C��:�FO��6�<�>�x�w�-^y���-xl�#���խ�Y_m�cg���^����A�~lGt|�8m/u�`Q_Ca�ׇ0q��Kʙ��
Xl�P2���<�t�G^����I�	��p�'�Jm#��6�E^�����1�����%�]:_�Ϲ�� C�N^�����y��[�M^����.���`$@�C�w��Ӓ�!4
�w�ʢq�Ph4�dR���@���Zy6��gp�UO#L	�ā��U�p�@�Q�Fn���X{B�K�2*�
�`K�H�xk���c�LzKW��b�-y��
���ؤ�x�'pQ$r�Z��P��r�l�LE�#��`X��<�v��F�-iCfCXK^K��_R�u�CZRI�t����7�=t���üY�,#va�K߆�H����j�6�s���~.�I�,�xq��yx�ڴi{nz�(Qّ��$+�VFe�;�V� %^=9��[���P.Έ�L�|�t�:;���U�8:iL�!�:Z�mx</�>>s��������ۯ�_���u��ǃ�+/˦� �	NHt�����A�,J�:��X�m��)�?����%rUf�Uf6��۴����UG��Ѧ��ȩN�K��HÉ�
g�į}+���KLU��334!]8�;��g̵�ktrǚ�#��2�6�5&�̐�wN�Ǩ�jݠ��;l��t��dk��x�Dm��t!����xK\�h��c�)�� o���xYA��Mj����hf�iۦv���K�Nz���g�u�q*�<r��5T�-(4m�?)�f�ʗ�߲�,���m<�Q��":xR�`���iێ]R�z;�-D�%��a�w��A�V�ڕrf�-�b#�{���.̗!���v�^'&q���ɯ�U�����7�q�n����P���"O�d�eV�v�7�3h<�}q�.���-X��+2D΂e&,�����C�S�L:q��c�̄h����#�I���98����o�S�qd2S먌�L�Wa�% ����*�5��{��~EH��T&>��c=R���J��� ��g��A
v��Ôwi8�Cڴ��������Vڸ�oȗ����_�l�k�+.A�Ҕ~�6%�!{e$_���/C���I���f��M�+�����:l��	��S��?�	i
�$    IEND�B`�PK   NM�X��i��  V�  /   images/c1791b9e-feee-4a68-99e7-b4273f4cd073.jpgT�\��0N��4H	H���H�� )�G� R�%� Gq��)q�!}���q��������]����ٝ�ٙ���~������&&��`ܯc��;�a`��cpa``<���$��FS��툁�������1��h!��F����/M����㵖��������sAޗ�e��qp���/��I<K�y)	�g/�Q�����^��X�X�ؘLX$��$���hٸ����"0��p0q1�=|����G�������y��� ��oL,lRF\~2&�2�䖞�x�'�R�6�X�|��k�m�P��u�7�֔¿S����#O��^٤�����XB��./bۤ�[��uQ��T4�k~�OM����ZTLIY��蝱����? �StLlܗ�̬�²�ʪ��Pk[{�������ѩٹ���%语�]����������_-�������_%pp���$XXh=���q�p�pp�1�6�&&e�y�/C���I@���AfKY
O�Z,�Eo��Y	���f}�Cn��2�����^
{�Z,�?z��QPD��o�W[���x�����)<�cԿz�����ZI��565��_o��4��Oō���<��Z�0�b���>z�O�	�R��SSSR�S���P��QҐSR1S=�f��bD�LL,�̔���`>z��W£Gd���4LϞPq2q�0�01Q�`�`d"gf�a`��yF����������������������������|eV\V ����o�]m���X&Ӭ\1��B���c�6�ї���1[F�}q��U4�L��x�FrrmF�*6��س���J�	Q^<��M����r���J�ٛ�G��8�q����r��,�:e4IS�Tn����ü&���j�^���=�~����o�P[���_�#��I����5u��8Qj�Ud�P��g{��I[%e��g`uw7%o3��^?�������~�{���f���*�0�`�5�#��MKm����rl�ϳlp݉m��vf��X�}�5�l����sbL�U���9���ƥ
r@���`^S|��.f���Z^Z��\��Ӭ����i� �L����U�K�s�Q�ֈ�� r�i�"��T���c�����89N>n�V����ܦ)�M0JgN}w!�R�s��i�`<5��T��IQ�$PS/e?�O�6���^s8#������3�����#��

Cgݞ���x�b�%
�N2��9Z����:l]�sw!�S���A:ǡ�%��W}�%P���5>��P4�:�듣�%Y(;���|N�Z!'�
��;Ijz��'JPPBs��_�P�����56F>�Y���(h�~��&�Y��W�'��j��]Pm�<z�z_��tz��)m̀3������9�\�U����v�L��H�H��?"��j�}���Z��1N�3X,�q��"���K�*9�ǕvjX'�����T*�_>wʺPKNdKL�3��$r���΅_�_�bSu�Ս�s��m쓞�o��$��%%�ު9eAK�x?i��	�q����2+AJ��@	�d%N0t1�?!�)d��	�����"턨��_O��9��fj�]���( �z�]��V3�F�N���|w�'�����l&�H�8Yv�N�Z|s%��c�B���@����v�q=ޟ߾n�����:.:q���&�#�����ٕ$J�X۬��FYl٩��|����A��7��g��j��,(J�J�U��%��Sz�Q�t��}�����Mm���m2�R-w���K�|��� �	*�
�+@*���^��� �.����[�8�V1d�B��z?����"�򸡢m��eݫ��!�������`�b��lޯΚ���+�A��]�����5�iw��K����ev�MNK�v�kiL^���ٚ5�� ����]�A�n����NB�A�v9��&����?빽Jp?<��e��si>�^�8u���)�K]7�2�
��K�L���.NDI��v��9���n��������ԥ�7^�\��l�f.'};!���c�[J�����n1�9/-
B:/I�2�au��}km��rh�}t���yD+b���r���jKo�PK����G��Al�k�F�Q1+`��ȍLl" V������B8�������K�ٜ�Wn���q�v��A͡��m�EuOXc���b�i �3�����-���‗�܄�����rҋ�"������牞��}�f���e*��R�佪�-� >�	�Ц�~�a.�ٶ���a�Lu8`k���j�9 D!���0��C���S�f��;��p�RM~:�d�Z�bǩ�l���e;������v���v����w�vϚ/i$�5o��h�}��bl~�5n��1�<�_��1�k��� �X�ğ\g_6�J:6�y?'}�����{���� �G����w�,�+�m�f֥ɡ��r�&x%��9V��i�,I���6a�NK(L���<�q�M�/�#�n~�����5�'���g�X	u|��uy��*���9����7����
o��7ۭR�	6��9�f߳���$Z�Q�|(0��R���F�6d���W�E��Ę*N��oJdVhwmq��ptQ��&�R���e͂�s].�^���yD��eO��V��'�5k�r�k|u 6 �1��HR	�2��
�4u��d�<Ŋ��u��|	p��S�1��w�69}��5�7~kx]��C����R\��ס(�.�*>܌��� &�E��P?c/_����+���QrV~U-խ���[�+x�ͻ�\5W��8s�Y���C�H*p�����J�t:�<֠RO�Bn3U:ӓm��D'��'�_��GA	�0tp���`����-��r����*!3q��p��'T���=�����:Y��,l�l�7��@Tm�M��iz5q(5�[QM�Bw���_1e��zB���;����	��P.'�ԗi�4�NYy�Q�
PPV)�/�1|���Wc��l��%�B����B��F��Xi�L��WY�h�˅�ʴt?��i@ ��@F�r>�.u֜���^�Cdwddj���F��|�����c��F-�ҭ���l�HRO*�ZQ��A�A.+�rm&��r�8���nv�ba5�R�>o���5� T*���I�Q�ʞ�]d�Z��TU�WP��1j+��ގ���4�����0���h��]u�%?�|�z��#�c����}����XB!����'��)���މ1�?�I������-)��T�y����Z�N:ڎX6T��[�3�V�
i��x�{��A/b�=�.
�`T(d����m>��t��c��+��4!���j�c��ښűp71A���M�/�)`���Q�U�����L,`%�|���_a��mv�M����"��j�󙈥6�r4w���+��� ���2ibV|�g�5[neU?;�a3�}zLܥ�Y�%�u���f8�˩�+O����M���.��2������Jo������kF�*�!`�-�Б�5UV��|MN��w�8����*e�h��ᴻ̀����e�C�n��`�t3������oV����r
�lt~2���N>
��O���᝚�Ĕ���U$��x=d��z9�-�ɲ�\��:΀��cZޯ���RI���a[\�]tr!��w������&�Xr�����I�+��d�d�Ba��@z�E�v�����'�9�����;��s.5�qX�<�p��&�T5L�2�{�Ѿ����_�Y�3��^��e��2w�b���~sQ��ڰJ���� Z�<�������Jy/Hoۑ k\�}~�g S�G�t�����(�����8�����y`�����,�-��z^���i@AU������t7wX>ג&Tb	Z�S�
[ʹt��?�V�%����2Y���kV�c2u�}鸝�'��޿P�ѹl���}���<�xC`�>�+�sA�Fa6$i���?WG�"K�S]$\<��Bn��d�6�:��P�,�v�u�W4rf�[�/�Y�+�������S,��=ܱ>���1�crgv�䳣��h��!�*C��w{�{%u�S,�%�td�4�9�8��29ԯ��t�+���@������n��2�&K�(��d#ss�|�@"V�3���,��(L�� �[l�2?�[ϥV.��~T\���v*ba ;��Z����ގj�0�px���ύ�V�"dY*i�i��I�T�w�5N�����)�%-�ɫ!d$0'���@Q��ɋG���<�B65�Zy�Z����F��^�^� �-0LݤU����,<?j��sL� �a�2�J0B꨿�:��&H~����WC!���.�de�ө���Ǜg�r{��Eu�dx;0_���z��b(!��(��C�[tkԈKgB&<��֍��f�����ÇOg���4�δHv��Q�
���kb_��(Hx6�J� ���EV����0�@����K��R���Q�#��zA��RS���<֯HV�A2����7w��W2^���Ӣ���uo�E(l�����ngk���&����$����&u"���ʐ�6����u���Z��<f�����h��N���<}	�G�_O����'�N4t�ϛ�cr+���+���˘Z5RE4�%� lq%)9%�s��5���Cu�.6ݜ/�Ȇ��+�ʕ��h�6k���-R�ŏi�΂��y	OӦ��N-�M�?`�P{�s��IݽKޕ>n�eg�
�L��	�&���Sl�?x�,�u^P�D2XS͖}��5�Jo�H��LN��')�*�8�8	�-2կFn��z���k%�?>����4궞�!�����	���5*�\�:g�	:���-�	����0EKn�êot�aڄ����mO?nҏ�#rF2����e^�f)�4^���j�}����i�]WLD�t�#T���i[�-y[�i�;]X�~��sg���r���ϫ�Q�b�x/V��_�&B1�lL)Мo�H�2J�.q����j3�ǪA�S��L�h]�u�pi��Ŋ)�?�>~���Yq��*�*+kZ�U6�7��˄	�,��(gR�43���	Gv3O����I�B�g��x�wX(����_mM���r��s�)eA����H��1lD��0�o@�*���bST,}�B�&�d���;��Q��GА.!�̴9f��i0Q3_?SW��Z�<E�vKE����B	��o�"3�ȅ�x=5nj1_Y��s�R��U�}��@Nr��W�[V��wS-��ZN�.an�ʼ��5�+��@w��T���B���E���κ~Z�H4uw?�g]8�>�������U�g�l���A����Am=�$#�#��L�u;��]�~�}�B+r6��$�5n�)��� _�A��j�FY��9ȼ7����x���W���%� �k��y�6u.�Bfg�Y�$�	O6��
=�⽾�	����o'�����u�����V�:�|�N�<2���Oɕ�_�Z"��~�/:��mUA�f5�X�S��	 2|�vJ����>6��)��qOB�ct&�U�ɤ=�㠫
�)�]��(����ٿ�V<� Һ��uڹ˯�\��>�&��5�>��*�;
���Z�]��YQ���u&�u:O���e� ]`��-��	3����}g297�����]�\E�k��;�nN:ζ�K�G�+�;)���6g��<]J�R��24M���l\GD�tf��"�ɝ57Lv7�;{}Y>�9`�cJ2%��[�}�qmac��%Z�_M���+@�2m��<'�"g�^2�B8F�ږh�`b�ݡ����;�����rF�"�mo�.�=g?�{���%;�跾��wk��`&����&V�u��Q�?����@�F��@�:1�����M�.��I�|p�R���D#�ș9�<'z\2.�l�K�����f1��糁��6��oC^KT���+3�� wQ����b��
�sq߽ǰ��`J�
�H�.�c4�"JE=y-���2.8�nS�k2�[��fҹ�l�0��^�%���ˏ6��o?���V*�vK*yC4-��[��0�R�L�М!ƛX�����+��<�h�/H-�ʟL��y�<��,�9[V��L��R��{�Fu����a`i�i��2��*x�y�Y"�K��7-mK�9f$���\�U�Ge�َ����H���aQo`f�jn��H�ـz-7Ov�[ZN`n�SHYzjg~%%�n~��|�Z��ݏ4�Y \���X�4t�o�3uet��:�)�Ieg�#��}J�ʳ9(�ho�o�x�>7��B�H��K}�~)
}��KC2zX2����Nà��d\(���g8��I����m �^�Q���gT�Z�o�m.�����$ Tt��������<��eu��i����$�,.䆃ˮ�$���3c*��Sd���$���A6����')��(�� �s���%Z����.�Y|���+�:��v���k�{��K^�:[�w���\���/����eo��%Y��9�DȔȓ�?�}x7�)���C����CY����w�^q���:��;DH$�����֋���?pҩ��q8u�'������l�4V���V�j����uR����;f��-�(��Ss�i�匷Ωf�ﮞ/�{*�l�� QW�׶=���^��@{���Cn����W���u�����_'5J���ǯ�F���E�߼)�Y>ʯ5墸�k�V���>8����8��l�rFO�2����F}��r}J���M�!rT�U$��j�ņ���� 
~Z�|�J��T�J�K��6�Ҧ��(����
Ņ��H{�5��-�\�lKL/���z�eHlN����+^�c�aN�P������X'B{��MFG�OU��;X��X72K�����I��b��|�:��7�N:�B"���)1�7��?�Ȼ3��7�ό��<�IS�4}c}?���$�)���(�;���ɵ��xn�)j���Ǩ��+��C4��j��F� ����=��+؉���9��RB ��]�t����mz�P뺋Iݤ[���2D��f)���ҡ��?Ǚ��p0�TA�l��ߔ���������FiEφ��Ɣ�E���ҩ��ũ�ް�����"�J�-�>	�?\7�1�*���B��
�6�H��>������[Ε��0NV(�+]<���龨F/r4��f�5���JB7�b�L��s���*_Q��Ś�I�ҟ���2�t����ݝ:��dN�PG!ݘ�����,�
'�8�K��!�У����@�7��e�CD���;x\�/�Zq<F�fs��g�Ŋ$���IH�[>�1Y��i����27��z�~���I�rR��Q�(GV�:1n�x��!h�M�2#��x�-��'�9�c��¹A}��=N��+Yq5�H�*H�[Ws����n��5��J��!?���p5,^a�w2=c"��B5Bq�]��� {P�@�3��c�e�p[%yW�w�5q���#�+dw���鯠A#� �[��ףͣ��AE1���1*�QMw%-���/|��Z�9�Ά>���+<B��)^s�/>W'(z�C��U��`��&��:��xL��p[���2m5V�/���Z=��<ۚx�,CU��fu�����!�.�"�M�LX8Ƹ9u��Rp��)V���/��*ޛ�e�#T�8t����pK�*B����9�"��U�dx����)�b6~�2[;���N`���ʂ����(l֯�Z�N�i��C��~��pt�08~Hv]sW�6�*8\1t�E�
���Q��S�3/�"ꭳ���M�tK�z���l��I��QBT����^!L!�r�7�*p�tJ�?w��z�+u}Q'�jӢ�W�>����%��K�bT���`_w�����Ч�{�%��μ*A-�V�Y�譨B[&M������DϚ~�k�d�#	>c6�N��ipru�gI��,*�3�j�,�a�)F�~������r�k�3��#Үŗ��,�J
l�!-�e�ӪC(>���~0�ʿ�5�o>��>1I����]�UovX;֫މ���T����M�
\G�&��߈�}9���>� �o���ݮuLԝ�ǫܶ_2_��T�>:�M��iK���u]Wt.���̙?���Z�s]�:=�=�Ev��- ��� 45���_��G��䇻[巗���t��Av��7\,�7�����1Ȳ S�>��O�*j�u!Qz��*9�c���C�%?p?�eֹ�b�B���ES��yv�y��pM{�q��#��n��/t2fuT����;�X�v�M'W���]!�yo�l���Ro�CP}K��o۠a4Y�~�_W��`���'�p�Ϻ7����KwU�4:a��Ty���-_����3t��:1'��H<�v��]|�;ױ|��d��s�A�U�+�P�vL�m������||x�����:~��&o�9C��>�^��W��'�Ǉ-ffj���Z�]�H�\�@�v�d�[����m��؆��h>W�;(׻YDH�,λᾝ�����Z��%N��V��n~���y9���T��>w�9r<�2t�El���yYѝw��O(Ԁv�Qf���2���z���1Tn,�XY�im�D�7��Ia"��iZ��e�ĕPG%t�)�sy�T��O|/��dҶZ��b���ڵ������v��¿3�V�V�����������J=�+'��:�����ƹz�<��.݀v=���ձf�Y���'���*^:��.��� ���xF���ڶ��{���k��Τ�����QҾ�׶R�k��_ZGM���oq��V�W��"�vNduߵ#C�0j�}%�ogj�-<��A�ZBO=��>�;�������9i����5�G����<Ȝ,�Q�q��z�h��Ѝ��n�5V�ҤEǮ��0�~�9o������ƩGH�[�0�5A�{	�Y�3A���C�3R����|��ڭ�q���ݖ�C��j�}�y�BGG'uԿ(�|�����֢]��W���)�E��7�)�pEP���h��=�ːm�ƛ=ÿ�@��*�j@��N�������=�E�n'ښ��ئ�s��:�Q7N}۲@��=2q����;i¿x��~sv6�����io�l_���F�׎��#�d��'��=���0�-�e�R�&�c��V�%�ɟ�Ȳ��p�����D���=`���*!3z�S�&GC?�u�������5 ]�/����{*���S����i�������qˌ�c㻛е��Г��%.ɄJ��4��0*n�1�'O?\��@D$&�A�G�w� ����S� ����N��1�
�N�7Q�f'�G��|�C�@������c]�S�.����6�F�	u�ճ�u��fg��gE���d��UMݪf��w��c��Ww����V$�j�w.�1%��w_��GW=/r=�^J���%]:�Y��^?�Qg��RƁ�2#�Z
�7�@�K�FXȺ�`CY�}��G뜴z��gT
��\�ߢ�A�'�C3�H�;쐥0q�{�|1��;<YG�Ҝ*	��2B��MC����M:^�v_�g���}�˞>�?׶��n�q��Dv���GY�~���FM5S�`*:��y"���*r��5��|�Y¤-v�e��m�$zo&�o�9��-���Y5�PN������6�*�����X��O[����A׉�@���n�!P@+�hm�b���&����K�)�Ǡ�0�]�W�NsAU�F�2�'Ik�x'����ߣC9�=F��!�f�����dke?������B��+��9a���'����?���RR>le,UW}@�0zs�pD���_�Z��|f�Q�}f�mThXv�]��w��0]x����u���2t��w�/I+_�v\�%�l�Q ��Nh�-�>�]H�	�<'��d'�Ŗ��h,��醔�:).9�&/ҼnU.�_]�ٌ5��"��p;Cq��]B�Za���? �C�	jh���A��M�zr"�|�HW ��UөTg����C�}�m�z(������1�|:���{�i^P�X�7��fN\����<��/$�]�&�<��q�O�K�����M�D��v[�P�>��� ��s ��ň�����$�W͊Ǵ_&n���$EǨOI����B͟�s�s3�D^��E�8gM:����4���޿}��`���E�y��p�Ī�����@�d�����j|������&�q$�Z��lnV��&p��qE0��˥����&~�1<��I�9�Fg[���y�)O'
�4p��uЏ^!뮊�~_曔�m�"Q)L	ӯ��O�Fò^t��I�?5^Pp+�|в�Q���Us͵pm���ziff��ϔ�}9>q���5�4�����V/����o#V�J�6�>��jEј�%�$��DT�9�Y���iD[���_NGS� ��*"y�E����dۑ�bd	�?
Ό�]Bߋ�����M���'�f}7V��L�(��D^�����]�#N�w�`�U>t�S3��P~vI�F��;{y�C��Φ])�;[P��/|0����`��ũԛ
�߻��}в�[5�ןB�)����Ǹs-��6ͬ�@5��|�B�^�v��<�cm5�l��. �z�"k���-���X�3���Oю�%.��8�g�N�.���q�����"N�����ZQ��Y]:�e� J�C^��d���Պ3U`��|]|�%{;@�-�K���4�J}��m+����Y��s�5�w�hv�&���]��/r��o���ggML���"���)����Ou��9X������YMvyʷ�Z?y�]2����I�~5��1U���K�tc���J�>k`klsa�?�����Ij�̷�{�M��/��W�z�OclP<�@��MTy�|${�q�̋�/a�Y@�5���߅��d�o�}t�h�zZ��r`"�?>�k<�8b�ȃ4v\+��T�6$#/#v��E�1ۍ��� ��T�	��+55u�eU���UT��īh��6<�ŀ�>�1��3"��g��bL�1*�.���֪y�45��Cn^/�ԭY��d:�̐X�e�8ùuSR8�G܎�)󯂾O~Z࿋\�ev\�B=MNz����C���ﬖ/X::���SY��:W�ErG��|}}m5��Gu?�p���Y٭�wDw��)�f?�w����|R����*m���&[�S��Z;yʓ�яb��O�H�2����_��]1�<<z"��ά/ؤmռ����E����2�F��&��iq[�Z>I��w��	W
���Zu�Z1���y�wuN~Ηe�����<�f,x���򭠝\�6��͇6����u��-�g	�$o�:���S��O��
&�'����u2=
�]\�+O�0JtZ��b�]��4�P r��J\!z���dO�[�\��P�2�$=�ߓ���bR&(6|�����\��[WM�0su�a��y��y�.[m�M4�:��#����à�ء�ќ�8�H��9(>�Q��;|�H��	�*���!��O���4�8�+j�<A�b�����{ݙD���71,$ʒ��}�ڎ�}J&�A�͞v7��b�	D�U�G�t)V�v�A2�k_��3_fsp�&�(��R?�c �1vI�x��&m�3D��J3�<����4>�7�W<;n���V�����)�rj��y������N�,�we��8S��0�^�
+�Us��7�pκ�s��6�+�/���P��Lf�[����׽=��)=�r��/_(vO��,�r���j�`�~��L8�I��k�%"G����g~	��@�����i�Hsk-	 �$P��O5����15+^���)�7�0i:� W�Vk�=��|R�=�z��uw�q�⡖�X��u��������Ј	)q���Cɨ�<��Y:�yܦ�=����C��Mz�A'��k*��t��eK��ߟ��`���%��n��}����ʃ6W�9io�9CC�������'MF�������S?�g�83(�j��D���i��܏�#�	.���l����]�;ap�cM�'�������/dd�獈��/w_EI���l_T�"��Hf4s��[�7q̿Y���������Cǘ�4����a����v�M���F<�1)���{��V�
��/Ɋ�h>������Q��M�k�zf�t]������j1�*�ǚB*Ʉ�g�jWeW9F�����@E|i8:PLɲڞ��Z�`t�P#Bוa<��x�H���
^&=��-[7�Bwd��[����1������Yd3r���*u:~��OȆr�E�!�9�Ci'lF��"ў=��(E^)h�&���DO<� �o���1~*�"��W#7\m]�M0�zx7���ڵS*[�2@<&k<�<�+�߻�1jmz�H�T�ʫ��F�|��h'���b\hJ^����(����]&%X��a�w�)��Iz��h����k��iY��������o���K�r�ݴ�{�~jg��n���rK~3s?N}ǆ�c�M,����a��҇��jQ@���Q;f%��/�e�}�)'r����]���=��i�ph��Б�I3j�:V5��%�	?i�}�?���)*W�N�Z�)}���������Iz��i�kh���ׇ����]��=v5T�:���3)U������Y.��?�0�M�b����W,o|8\�� ���a�cj�B5%h�������Ų�Z(j2�5�s���Mv�����@@>�d�Hm�(�� ��_�;��r�܆��Ș��|P�4*YQ�!�j(#�7M�61�4�e��pR���w�<Q��Um�Nf�C�O�3DIS*>�n|G��K������KG�Ⱥv�j)=<��]�1�q�^�) |����8��MqZ�y����"�w	�;�L�|���t<���	�m)��W�YZb�%�x}���aOs_[wZ&}f�ʫJ41���;��ʀ��YI�D�Zfzq���Z���:mD>�&}���eM0h�~�&�
�+(YV��7��w��Hs�H1Z�g�1�%��P�W)$1/	T1��	�Ql_���֭��}��.ӿ+c婧�([;���N�Α��uM�w�K���wy��Đ@��w���qPZ�E�ir{���Ba���}�J{�N���	�NA�阕���a��?��Ot��æK��[��OR��{��[��.�;�w�������?�cn?r^��<w��P��}7��d��I�P.�%����%(]v���4��u�!�*P4D�L��me�g�hWg��P�mf<��xŭ�~`�~DS��m�=Ҏ�������RA	W�d��yJYWUt�OBsc���n��ӿ������|7�i%�תgF�,���\�ea�OO�����p��d��T#�p6�䶚ۄbh�^|LK���B��y{���\kݧDt������#̴���W���'c�Y|Θ�K~�"�ś��y�$UI��w~��@�Xf}�JAj!�6�]xb����۵ f��'�/ږ���ew6���� ��|x�����5핎B��n���b������;7���=}�V^��s�`�kli�xa�,�~/D���A4����Ӻ�A�K/������p6>j!�#l���8�T���-aIk��'���� Gb��Fa�j㗯�V�4&�:a�P�6Ӟͨ����	?-��R��_��$΋�OhM���� b��Ԡr�y��W�;��p�a�C��pf7ش+U,NO�M���:��X@G�I�J��I)N�y����g����l��^�Ksgo�AjtЙ 1�6|j���8��ָ"���o�l?��B�Q��Y�\�t� >?ѷZ����+�j|�6�]��f��NGgs�	�n���+���li��9V�X̂�]���ƞYжL�ٱ܀��y�3�n:jض�S��+]
��PRI�E~�;@�uV6�!�9h Q	=jȎ�: �tpah���d��$���w��S�b��:~n�=1���B��!�ݼ ���6?�V%d�wXs�oT�%�l��ҋx�W����r�Jc�X�{5��B�a�
����+�(ȅ�������4��G�|�o|�{OWd�H>̐ڕL���e ��:,��i�ny�,{f�	@~5A]�l�^���ߢ�q�n��Q�#(��H���"�SL6�ǜ���%W<����ө �}��j�V��	�6�|v��4k��V�c�$���N�
�Kژk!�`��M�"O�I���OkO��7�ɋy�����r���j<M0(�{ɟNڮN�I[��5=�3Ф�Bl��ڊ��e�.�d^+n�%M
�-�8ۚ��%lnV�m�|Lj�M����J��	~~��WP.��{}`u�%�s�ݤߩt���,>�6D��&�{����᩟,}<v���S�4�O!�@s�j�M���S��k�viS�Ԃ�D�:v�� �{�;,�j1ʭӽ_ԻN�y���@�l��'���t������V�R��f�xvU�"����C��VeXg��P*����,�z�u�=�\�k��˰ڱ�5�%��ᇄk�K&ߵ"�Tѹ�5���}�´`��bhr��,Wx6���æ2�����@�f%<0����g
�~A�KZ�����u��MWF��E�����ˆ\L�ϙ�;���`i�?e�=�[Jh�����^neY��U�tz��>Ȉ 1������׸�KE~g���l>�Ԋ�Z���`+!��Z�9+�9[z�#P��!�����gG0���żKRE�Dl>~;�V0���z6���[����[�4Qy��Ta|�B���w<�5������\:,;�&{������?�߹'����]V��J�E��?u���@h��@ymOyiōnu[�DXH̂���l����A�]z^�w�]j.6�N]y'L���|���?G�����&����P�,�tv�������M@2�BF��_P�{s�|;[��/�-8�3�9b�B4V�J�����.�Uk�?��rIfR/Z����]� ��p4	tC7T��.�5��A+?w���`t�� ��.BT�݉���939��#5��N(D�
�PE�yp��Uɨ`��n�v�v~�	6�bG�Z{�9s�0#0�(<;r�]{��������[�P*�*���]�L�g�"���S^h��������G������,Sa�x�2[��YL�ь<��b�^m{�rp�6����8�Nͪ��m!��ƾ>��c�+t�jv%��N��c���PU��#}_���D�%�%)�a���
�caA`������� >]{!knt1o�z�z�F�e��	���*�"i���l���aCV2(�Y�O����#6�םԉN��σ�gR*aOK&Io������I3Iǡ?_	��3�Y��-�^�^��.R�������|�����+�[����1��|�y�~���tM.��a�G�{v�`>�:գK��hړԴ�i�:�'y1���I�L>ݼ�wW+�V��TqJ��k1�tPQ�І�E��T�[��t�!��C��	���6ǜ=�������Sr?��QbK���ܶs6VI�;9�8���t۴���PY�ه�[yz�R<�-���i�I��͊���Ǌ3���mC�b�ٖ��/�1b�[��6��������z�\��z��w��аB�Ļ����I��)G�>DLOU<"�uIr���.�Z2���n����G��A#x0��S���/U~� U�,�����$q*��]�^�ᯱ��F�}��?w��W4�Nx���{�˰�2�[�<�+�p���̥�� �2%p2BcZ�N���AkS��F#8�{�/��c�T*�k[�Uݻa��' 0��a�Q&���2����XG�*B������,��c7>��Y�aGۺ`��*�����Z������uY�f��Ɛw��l<���2��/_�<i��	}�X���`�#��_Ki�A�Sp6q*|&��Y��[�RյD7�3dh9d�4��(u���t���,����k�{ p�X��:�cP�`�Ȧb��إ ��Ʊp�A��h����>u!zzǊh����C��ʱ���i�P0�Vյ�P
Z��u�݁�Dh� ���a
ZS�_�*�������qA0�����fz�ZtR7����k�*4�5v,O�@I%ǆ4���@�~͐����-��kny��9~�t=��������̬`�K�k��kRp��k,n ���W�;�\�S�6RG2%����G����F�������m��N�7O?҄N�W})qI�=7��YJ��
a�w5
�V��g�e��gLOxR|���K������6)c����A��/2�5%��6�T^J:ޥ-ʥ`^�_d��̏���(����0�
��"�U��Gy��57���F6���"�4=�O4F��+���V�޵�2Wve�0R��:��ջ��)`�E4���;\�>��ۚ>��Kd�p*/5�����խ�j^�4���<�$#+�-��g�RԾ<{��B��?Aщ�Eh.�7�o�N�7�����q��4���8���C��g ���P��7�۫�P�J	]���A'�f���X��G�,����6���}�(B�l&ʚL
�p,��طO��l�����2	)d�ٳD�6ٲg�Ja�B�Xf�̙�������y���9�q�����}��}�3^3��N�Y�_�����ϐ�֪�,|��Fh¹Qz��x(<z�p�/�=�rc��?w��7��- ������Ĩ|�j=u�ʻ�G�1k[�^����>5�������㫞G5�x��`�_)�2�+�!����Ca�˼�_�pk�v���i�ڔ+f�K^	%h�Áh}�i�m5�_5�>�v���պ�__�z?q֒�/�>��"��8z�r�9���gp�W�n�z5�����輖�~䀂6�T����5��A���^�?�USzBn��� �����>0ҟ�5NMMc����@O�7�w�E�f����������\��c�f^��<���,�nl���J��8���	�����g��J�gR��w�i�'��dy[}7|$���.�\��$�����e!�'$���1���įr8r�i��	�1��U=���_m}mixf�o+����IU��s5�w6L�%r>���p^���I	k�Р��w��AI��?��bN71�Ɖe�S�����<þ�9��~zU{&�;t�ل w6�g?m�ˋx�0��(��&��æ��ϘF����5o>���W���z^��}��D��s��W�nNpޅ�������+B��QݩO����R�j^�!���p�g���Z<<pE��j1:!W'<pE�x18�A�'�]}��;��,� Q����X��\��լ�E-6�UE�^W���L�:&�,&������7"?売���Vz����� @?B��"���r lm�.P�s~�MR���Ճ��H_��� �6��mX�"9wW|5k+����������gK��FO4��¬+Z�R�X��'�T΅H�d�M3L�M
��,���!��\��e��Ҋ݅n�h��`^a��4��������9
��%vF�۴r�*X~M��.��g�wI��?-ö!�%y��%;Ą���	�`L��������ޠCڤOV��a��~��sNZ�٦����˦v~�z��t���$zH���$"��r%Z�D�Zկi����/އʮ(�j�o�}��IO�
��V�{��!���- u	�u�8?6�z��IN��.��B9xJq�녟8�
u�����y��2�WɃ����%�O�����}��_1�y��I���(�k}~a�E`��0ϟ^+{E�����#�����vA�)���r��ԑ �>P��/���o@�6Ţ&��!�D�b��Ɠ�k��y4�j�@dJ;��5�2�-ae��B_��˽$u*����8,��--o9��І7r�Y�����!S��6d��t�:�K6r,ph�ݝ�2����>t�A\�Hե�� �P�z�7�|#��c!,�K6e!��e#~����%�dkRx���Y��AE�̊�mxۤ�H)I�����/��*�?۠����x�~S-<�s��I�f����Ƙ�f[�*�M�#c���$�Dj�X��ه��~�{{9����k��
�l��'��m_��Ii3�V���̈�B=�@��M��F\#�"���(��F�!#)��#� ����u�`�ѨS�l6�O�Q�֙�2tÐ�K�����B�pI"��hGIgC����\iZ�ԇ��n��uj�Kn�ș��\��x.��'��?�Ӥ:&�� �Y�5�L�jpũ䠧���Uݙ4�z����M1�.m�:��ٽ��ֆbQ���s� �	�Tb{\��J�8��.�ik�gV]ȑ���-���v��/kiz�@{�pt��~�B��m%C����R�P�������s�a�m��"�P׾r-TӪ�1mbK?.`����X>e�w�yPo�S�;I�W������;֦U�d�w,0��4��9EֽM7��a[�����ob�z�����e�6�,�)�߼�������x��'�S�o��K$蝪�~6�p�-,�����D{�3o���%:��q���>�<�.P�%tl譌yn{����#��9�?ץ�~P�8�H#l�E�v�,�ۥ�h+GmY52����"	�,���/R�FѴ/�Im.���N�	j<P�9�!5���p�4n����_;���£�roA���76������u/����,N���r i�בí�|pa�Wn����[�\	g!b����3�1Գ�FN��$�OS`F>��j�[�u�%���"�HT������F	��E�`!��4B�vF����1��k5�k���3�a���7�	��u����r<Ӱ�@��~
B!�^a'5���8�[n���u����=�?P:aF��^b7�05f'۔�L�@Sv���sҴ/@%�?_�A�Yg!��ĉJl�8�Бi9 �ki��D*�1�N�c��ͽ���s`*qV�\�H���:_�Γ|�������!��M6�K'T����%�u��]�jV`�
Pvm�Rv��	:ɏѶ\��C�����m6��99��c5���<�&v�g������	i�x��ĺ�=䐫A/�z+�i�Ax�t�u��������<8IV�{��B�����(�w9:<?ӄ\m��Κy��Xͥ�v2K6�w0+�:�؏���f�O�O���0g���d!|ѾHCۖ������7�H�V*������E��Ѯ��Ή�#���\흡վ�֣b�G��蒝Z��3%�$�2�W�W�k��V���z�1~������݁�b!R�]��p�H�2J桂]�.i@��,�:~�����%��I��'X���%Őn3]��d�nU�N���pܒ�������ml�gE(^ЍWNd�X� �����mDJ��@O5FEƑI��.d�1~�o%)�P�QH��s`k7��3#�W~dYݧ����վ���`P�-YF����y0�����OЃ��	���Ȧ�,j�Y�4Li�V�$X��D)�o��4a~ה;��~����������siq����8`���(��ng�*4`d���"@F7G����\�eT���|����|�21+D��x{��T���������ч{~��#�:B�m�+��_~zJX��]���X���l3�⛁�W����d�ڶ�-u�{�+J����w*��?|�*{bT�m*2�m�/
��;�?��=D^�|�&��B;������I��[�T�I�����'i��ҴU�� ���@��H�|��$�r�hǷṀ�7��P.}b��x�C�Zo%׃K��c��:s�ޒ�Bڏ����D�G�!���ض(��tv���g@�|�-�M�%�i7
n��@V0����+�+�ڧ0��4g�Y7xn=@7���gPsL�_���m�n_�U��Sy�����,���
W���O^�ۥW��}��Ǉ���z�m�!�����о�i�Ge!�ȁ$Ζ��gAYq.W9w"�x��4��o�ס���G|�Gf�|\V�ئ�����EX�X:�����u6��Ky���ç�j���Jp(�8/��^c+��ҟ�� [����*�W-J;�}�r���!���9�ޭ]�׳�t�(�[�v��t�X�R��vgkh����J�W]����X�~\P kq�����@�A�Ud7K&��JT4��\ȥwn�S����2a��-#�M\	gzT%�Uա�,����ѷ���-<VC�rS���qd93i���&z|�(�:Cs"�rN�:��yHo�'�a�٪��%X�4/k;�~���8���ߥj+��)Ǽ��S��N����"[V_>7�du�h�
x����"��4Ӵyt�ͅ�ş�MD����J�/�e�CV�ѹ�*T��k`�Z�U����K�y��!EZ�X�V��%�1�ݧG=���3ѓ]����wx�lg����c#�L��5�b���*�N>����&�t�["�u����M����(��n357x�8�{���	bl�����DE"P��]�hm�sܜ�^\,�h�>%�� Y�2?4Jhh_^�e���Po4r>p�.~G�#tPm���=%ҿ����g"�l��<���_�<��Hx��	ݑi���f>�G+��;ڏ�	(���C�vژ�}
2�"�ME�ef�sJP�-���HT�DgC��"���F+Et|.�<n�]UH���=��������~	�>h���2Xz]L�Hl+14<Q�#]�u91��p��$�e!��� ���>����8r�!�)�-�`%o��]��yu+���Y�:W�?^��}��wW�Z�O����oP�1H�<�	d���f-�i�(ݟY��g�s��h��H��K����������$��s��^��k��0�4І�U��c���O�(�h�\~OL��*���)��NE�V��տ.�=(�t%lS������m�z��)s�dN�Jj����T��A(���O�F�a�8�֞����cfO���;0�X:��9����JߺDl����k�(g�U�bfi�^� :�xF�z%E�w>���x6���C�I�R�ɎhE�׏3<��VrŖ�Cq�8B	�0�rC$�#�X�̒mhY�#
n�x(�9��Ss�K�� ��1�D$�l�4����9�oۍV#c���j+	v B/�V�E��S�z��fuQ�����F=�?"r��Z�ݿ?=3�Q�3z�17��A���~��\w���@�@w>����ŷ^��ԡ�\�]5D�l�U�ξ��^��񋅽��ZN�UH����їN�Z}����T�F�-�zI����z]�C�F�ŧ�Ն�_]�Qa�&:�~CR3���I�A9ub�m�q�vHU���叢�������ƻڸº�7�\_wю�]��|���HK�]k�L.̲����C��cHob��+�[Z������5g�2��]:�'��w��4��w��j��i+�p�]����A�X�G�ֳ^5[����%)���Nr�L^ ���6�9$�FUdKl�҂��e'18���2�w<�LXz��[���Z���_���*�Z�2"6��T��� �r����҇j>郼(RG��3�H�oa��^�=!a�F}3���I�"D�*�2����L�Kv~Eh�����X4��E%z�G��W��q�i(��09�#02�`��r]�}�'w���b����G��r����-�G{�_Z��M	i�ץ����Ǔ��,u�!�5,�Ȧ^�g~�9я�z�7��_��JK�+~����'��;doȆe��y���s��l���{��r3NT�tJ�ʈ���Q� �h �f���A�k�#g �%���ɹF_�t �"ު4N\�t3<^�����x�IE͋-�@�+=W�8)�;�'����M��gz+�+�����C���1C�喌'"]<Y�?�i��[Z�����!9�m���c������	޷��5�Ul�`B�X�[���ՠVFCkd�5��z��Fq~r�y�V3F��|g�-4�k|܎�t�,y�Vaç�I���A=�흄�A컋�jV��H2\bv�'�e��cc�9����*-�* �� >��5z��f�&V)�x����b��E���U�c�@�Mjy���dl�p�D������F �d�-�j,�i!���o�:�/�bK)���C����W���hjB��B�����Y�]m�`�"�y>9��g��>���^��>�$�>���r!Q-k*�BWŁ1g���8g:bw���dXzBm�}w�ޤ�+����BlG�~ȼ����e|]����g��s�V�!���C��P�����A���f�R%���U>�҉TM/ӳ%S�kX��I�}H{ׄ�B�w�|�kio��6x��}�pP�pЍ?���1c��8� t)g�B�Q[����z��U�j���ړ�0��<�Б^)��
�귞��&��Y���n$"[� �W]�m���f蛖S=����\��F��!7#�-b���E��{��R%Ar�� +�g��C�5Q�jpb8�٪��1��IL`�0ߑ�;cL���W�UlV����Pj~���s,D�n��gm�5�.�����ڻ��ӽVb u"[a��<�l�0��/������e	��t�"m"��kE��<U��A6a���g��'��F���{U�d���r׼�"�~X�H�F���U��X��RTZ�l��ܲI�Y�d���V䶅�"~�}4���I�_ґ���+Z\�1���þY��@﫬�ܫ�أ�^���Z!]��\ +�ƸN�1m1	��@�l>�zvG��[�ɜBLM=���P��1��A�����*�w��D�7�V��U4�?�$�A�\��Y1������,�li��󝃚i1��.�e�cEL�z}���>�/���W"l{�~�.�����d�pZR�����EQ��B�v�C�'`X��v���.�1k|:�F���V����8߰-���YaS;�T"�2{
K�ۦ&��h�`��A�E#F��0Wo �eDb�Q�7p�P&	.���ղ,M�Q�Ș-NR&~x07�;�M�8���R���I���`1-3
p���B<��rbH�C|?�\/�9:U_x�sa Ý���*2#�B�3|[�
P��9LMj&zV�,i��20��f �%1dL�D��hč��$��ç����)���PI7��Q�׷�mᗠ魘U�O�����m�����&�?~iW�o^tL��K��eG�k!{(�7j���d�Ȱ靷#����2��98�'�ק1i����f�Y���g��a��&s6�=�R*��.~��2�������N�X\��2��k���%�b!J��� �͇��e��UB����I��T��ċo�Ƣ�2�pJ��IN�t���P�D^��#2X��DJ
k�
���!2�S�d`���ԉ-�M��Վ���5�ZF��"
kbb���r�ewL���q�>3�[�l��@��H?�9ݲI�� �FlN���Ka�X���D�������m�x0���0S��&���[,D���;,D��B��NQ�3�>K�����B����`ގ��=0�6o�Zo׻�[���N��VkQ��BP�w����_�
�·�����*=S~K�z������v�$�g!�	��_���׻�\����挆����S���WmfP�")��=X�^�ׯ�j��2u�Z��ׂ�1T"zx���C�p���%��]cʝ�_�a!B[�Q��{�K\"�t,��2X��8s��{lֶ��J�e!L>�,��mi�S���T��ܙk����U�6���=�y�/�������Y`���`kO�z�B���5Nv��!U
�|,�K=�vd]jc��/�~q��~%����{��7�d�}��8Y�"�������
�ٛZG%O�=dk�|���wo�ʠ��|���/�-�/�KVվu�1b�-�GSj���N�B�ۥ��ۊ���H�^~�	JD������ޭQo���ͭ��xu�:\a0jN�o�|3���i`28�1+��Y�v��I�_��m��Ԫ�D����R��w��I4M�$I�=�𯀽�,^ή6����P6b��;�J�[��G�� J��7�[�v�sn��kW�9����w���U����Z�e���J�񘀯B�X��|���ع��x�iK��1���5J�Ȯu��F���$w5������'��R/wG�om��7�������	�J�Ϻ#���H�assv	�	�ܫ�"��o����d�^k7�^��`Ό����ە�[e,��KH�y������w6�Rf�y��fT7�9.�����o�45�ꕨ�<P�r�����=�dӤ٠�`;��a5?���x2�f}I@����kw��6G�	u1��-h��X�g0N?�����3b��v�>`ĸ8g�5�;%�sV�%a\v�2��_�5�xV,�}KT�y�5�J	������]����q�� S��:H��\d��{�o�.�w(�",����S����
��Zb�kn,D�\5�@j�Fg�hPCI"�.�d+Bꉧ}d!&JY�l"�N|�:�������� oxb/8
{m:�����G�/>��{�~��*�NL��ĳ��y^�r�!Qf��������Wݶ���oZ�}���ʊ��s�塥5���1o��o�����
�-��VS>[=?��a����¥B����[ȏ��i���������O.&�?�ۯe�P�k��]��!�L�#����Q������+����u`�理A)Ŵ��e��|�sq�q�r�5�pE�(�{�U���H��?��[����Zzs_��:�O���_�u`�.v@F�~�
a$z������
вI�F���Y�"�:����
�6]�p����}�N妎��Ǘ*n)<�r��ׯ���f��xcx�j�|jNs"�����(�.��p�����2�yP�/V��;�)����y��p�[�����!s��s=�K7����c!&�����#��S���6ke������0+�g=ԡ��\���?�j��
Qz���&	lV��$�n�~U6HM0�##E�jߦe��iK��Ǘ>���@���9*�,�v<�1�O[�f�~T��(�?�ފ���I����.�E2�`B�$NU T�5q~D$[��~�g�
���}�酂vl��_lb�П�K�l�=�}:w�[�����Y�Y���N�95�b�&�r���/�P�l�rB��jA:L�+xa�w|~�B��*8G}�<)e�5GT�z�E�Ng�P�E+>��Y�Y��﹖��d��׶�2;�<C�]c�H�&`�ź7��z�G
Ks
\��HۜKIP&�O&
6sɘ�T��|���Y��Ճ�_^�9��l�ؗ���5�m]צ��ל�]��Ţ���h�+��ZB�W숕�����T��)�w628�������e�Ƒʆ�'��"���\���N��8�3br���C��s�e���s�s�9m~����j��zE��jv�$�h�P�X��;c��.K�M�dbD�R�S�SD�����1�!��N��:R�kə,Du��F<d�5>��;1
>�-_�Ă�^�>a!�'a�S_Ǔ�}8\_�f��W<�&1�N�@�K8��雞��Z���B8W삔��6S�'`6YBſ|��<�e�-0���[�6ɖ��e�h���O{�naZ��i�����$t� Fx�j�X��|#�n�67jw�~BN,M�J,(_}ֳ��"��m5O�@��d��&�Y��X*�O~0���S�^��Q������I����t��J���{
溣x	�	�:��6��|q�� ���@uz^�{b~\��<�O,D$�/�@S��U_��{�.1���4/kI��&�@J����-��[�b�,j�4�p�@�J��b�ٮ{�8%�:��Ǥ~���������
�F�"�|w_>X��w��� �;&-�ݐ�����B�#=h� ���1�0�0�;5������۾ڜ�B��9�fKR��V��Nd"���iMbf]	�a!�TQ�!@2\K�a��< 	 n��r���jzG`�)��Ռ�h��KC�Kd������(��- z,�l
ā�4 bǰ���髦 <�7 ��m��
�:���d/!{��1aw�׊֗e����G��i���O|�rS�]����qd��o�C��,`��
�C�&�1̅d#�A*|��������pp����s��{iY���k�_B��I	��,D�:|��28q�b������{�4�����s ���?,I~2�Aϑ��9��_���`���O_�J���B�	k��%x"#i�=e&,���`>Q�8��	����\��=H ��j�`ڔ�'�:Oo}e�@�1,��O	2R�e���-N�L���9��v��j���	*�D������	�C�K�[n�
��^z��<�N�?(x��"q�ΐ !�b	�{�����C{;Gh5��	�%�4pr�3�7���
0��J�RHÆ�do��Z���0�����w�`G
�@�$��c$�X�K���������.��gx�'��[�p �?������n(`4�~�N�W;K��0k؄�1p�2�x+��F����W#0�{����&{�Vm�9��G&�Ƽ�Z�����&��m_�T�x�ҝ-�;�WTX�Q��>��q�?������1>��x϶l%_���c~|d��N��>�=H%-��<M��Lڂ�#����zd(��i��>*��n{f��v�!xVQ0\�w9�8D#���Z\Ӏ}��5	��,hE��h�8a���N�����(RWz߅q����B�i
����>~5A��7ω��S����P`�y\��B�� )��C���/��B�;�<4*�s����x���f����<�@��jQ��x4��4�b��4�?����u�V*)5�g����Ht�a�vm�d�
�%`������ ��-���Y���-|[f�O�vɀˈ?(��@%G��t�B�ގZU�>�Bt[���d��ΕX$�C��=�]��|jz����m��^A��ռ��,t��T;��hĜ#�r/�cܔ�8��ͩXRPĕPX����P�%aP�>�q.87��n�|NH
	��-7�pmT�+2��w�':�0ܰ��[C����_�l���jv���%�/�����c(VZ���T��%H9���%��j�7{�f�餭��I�3A�m�x����Fx^�mV���@38!�Z��ns��$	����}l��h
E���k�W0�����.}��;e4�m!N-�&ǪWؼ?�������U�c����YD���c�IƱ�'}6n����S�F�m��h���c|���Xj�H̅[S7��s3���������2��e����jXd��4!
ޅ�������B6�������,���V��<�yӘb1y��T��h΃<LS�y�ϡ��޽~�!��}c�C7�=EWg��߃Kh͡KKЭ���ݯ��\l9�X,X�U ��O+�3�󆁿B��9Z������W$��]�
�	�2 Up7���j��-�M�-�ZS���0�ӈ�L8��oڅO�^s���r�$ے�K�u��]�~�z��hv��GA�W�zM�����_�_�A��,ΟJ��~a]��\wa��g���o��b*��_5ӌ�����o8�VȔ�����Lv���N��[|n6�1K�����������DS{
l���&X������3N�֙ⴋ��n0��*�i���S78�S�6�R�óL}<n��7�L^�����kz�TX.�2��A��2��Zw��yr��"�ve�>f��	s�!�:o��ެ��bjڊލ`L<`�����K�ͫ}0WMr�]�v��7����}mP&8��oP��P��`6+�\8֦�#�SvK�o�/(q�̭F6�wt������b_ D/���:`��ޘ�λm�Vơu"L�d��na?���>F�mT��?R~���1�pv�"�\_�ٮ^i��/�4%�x��s����M+8-Bap߇.\a�H�w���U0���L(��;�R�Nm+�so%r-
�,aB�dS���@a�Vɣ�ΊcG�����Fov���:l���5Y�j����#"Dv��X45zt��zr�������͸����.ZE�dhx;JGK�������)��77|�X�>cu��&}7]7R�I>a%G�bS��۱���I�sU*?E4�����ϣ��R.��9��*�d�M�_���Zs�i�8^~0��`��"I�3�fs���sݶQ먳l	x�w�*_NCm�*���v4�E���a6�}���� F�2���=����	�P�G����a�b�=��\
�����\����� �"3 Ԯ�.��u�M-[j� ��`3���T��#5��ް;���[K�wu)q-��;�L��yJ��zT�֒Ϭ�^Y�}Q��=󫞲�'?��77���А7zk呂�Z�y�K��w����A���K���]�YJ��`C5q[
��0;�� (6PK�J�����')�l~+�W�k�@��)�S�Z�v��-�0�N����Z�M�HG�e�����.���{�]�\�g��/�Qu�_�՞y���N<��D��SZ�W���O��!EE�G���K�N?�p��H�Qɂb�h)�jbY����;1���i)��д
��.��� ՛��K�t��K��[���M�{�-����ٕ�+����;���`�u�c����x*pB��\��aL�$c�adY��B� q�e!b���ع�0H���/��w������l�~�F麨�T JD**��J-�ry�8y'��'�g�D���PC�զE���*��6+�T#ݡQG")R���4VzG�<a�(�ѣ"��#%g�K��7����2keL�7o�z+Pi'Ϛ�x��ߤn���|̫��痞���0F~X����9P����M;Yt�ٰ�$}���y���j��R�.+��-8D�{NtO��5y5Y���2�ōt��F���ϓ����𖔕��i�4�[�n��V�K��B�j�V_�>�2|�����R����]���q]T��(�ֿo|=��r�+�۱pk�� ����c���o`AR���kiT��O��2�q�d'Lu��X��}��t�6$�2��'��L��i��68w�g��Ȟ�
�>�5��I��M�b8�����Z��0��w��N�I-R�:��Ȏ�D���V�v+���)ޥ��	�0�pMJ�l��R̼d�Q�*����6j3����Z�+ԛпc��GQ{�)�e}~x�:>�X��#�J� �޷q�2�}3
8�Q"�T���y�c���KȜo��<����;���l&�%1�m#��lĉЁ�bBu�����3�pd���)�-=�mV��3\�3��:��$/���d��$K9}�j���B߉o���o
"=3���^|��x?}�&�b�֭��=Ss��i�6��ܖ��%���S���+`S���dO��+�U�F!��?���P�
����C����2���.e��	� �e�k����+lbˤ��*���0�:QT��,'n��Э�2��s6Y�Ow/�](|}/�m/v<�l��@�gֶ�*�<֓H�e�SI����-�Gpa�鹥��c�=�(�u���{R#)���]{C��j��N�mo��/�u?x��b�'c�TG��ێ:��a����D���(��h�i��ի�bu���y��jיV�;`�'��'#a��=l�����
��A��6L�a����:�q��)�_��uіv�L�K�'���-�lt���<5��7A�f����~�cXx'�,��
B*�fv�x�#�;�^Z���%�z%	�P<"goF����Y�ж�hT�k��)�e%��Y����4Å��|=7I�)븣�!���s�<��.�(=�Ovjۀ�>5d�ߕt0������*ȡ�l�X8Lϲ|S�n���2��܆��j�&��H=a�q���i0mo�������V�3�\�
 t'�sL�xw���wM�C�~��q���"��sZ>�S�f1���rX�e��z0_�R�\BnX3"���Z�?�EL�Lsw!p&m�F�B�����ܭ�)]������C�Y\	\����O?&,+/I^�I� �^�;�h���l�e�,Tu���l�M����~aݘ�	f<L���>1�2]����yE�/��PI��ү��Լ<n������f�?�j���k��G��	�G�9�T�r:��ٙ��k�������U�`{��=�!A��q��G����e�X�q:��˛���i���"d���<���}�N �A���y�����+�?�3������HmU��|K�M����_H[.��~��4�q�ӎJg
iJ2�	a� CJX�h�}� �]���g/|층�JL��� cø����s�p<t��)����jU-�����)������!a�	���mR����ˮ���`��q[qE{��jM�)?[�ke1:|wq����w�[�I�w2�=V{8L�+s十�5{+t�ՕhG���cz�Qs�[��-xػ�������f!����5Z5^�|����-�'�4�h�~����g�t��|-_4j �ؿ���Oc놳�-:��7��x�k��������k�I�Ӿ�;J�aoʢJ���\Mf�^?ca�7�u�~�fʙe�'mҔ�{ލ��P��QAQEj���|��,�R�����������&�U�8	����\������}@/D�[�J	z���۰b�������x�\9�"�8���o�8��t9�<�\ݶ~�t�J��\�1&Yd�1ZS�a+]���K�L�ë�
ION=p@Ԏ�x�џ�c��C^^
J��C�/�8
tӈ���i
w�]�([�i��ֽ^y*��g����gR��@�J0=�k���V��f��h�!�i��e�9�>���&۝�O�'xa���w"J�)�]���Kn�(��6��>5�%!ۖ�d��~XکD����e�0��h��Gx�B0-��l��b���y�-u����d�|وw{�����s�t��=/�� O���w�n\�"Ơ�~+х��ڮ0s<�������MZ�N6�Y�p�]�
.���|��:�FLz�i
�-!�����˱Ww �B��:�Q��R˹5����ל�IF��?L�90�O_�8���{�����0e������ќb����H�	V�j�3�ŏ�%�l\u�i�Io��;��f�k[�,���$=��^ը-�q����<4��H�]&�dQS~�ٸu�Y�>��B��� \�/�Yv|�jߜ�/�Y@�\]�o�Uݯ@oC+�BR�]7e���`�C'l�$[�e���o�j;����b����GxF����Gڊv�*�u?b�[�v#ȽR��1��������6�-:R~;THSp
��V�^6q['X+�W��Nd���=�Bq�������]�/2G�
8��ݮ�2�b��I��u�Cz�G��<C��R��hϾs�Pff�R���R�Q�K���Z�@�Т�`�=�uv�ML�8�ZUz�t�$�q�Vkh��98 g����'����E��Y������$P� ��o��Y��S�?�<^�K+ˤ��Ò~�^u�.�*�?7/y��+��qO�ȭ��[���F
/,�"�.7_12/`ʥ���C�2��n�����1��Ǡ����s���12d��_�����p�� �t�un}��M��L�����b���ZW�鐣�j���߾BJ{��#���
66	�~ְ�#%@f)���sZ�~>��r�"�B�g]6b�o�L4#�^��{`kiAs%{E��w>N��P�~������/՞r�\�}���ko4g�|��%1��J���~�Q��y$SJE��t�־�1���L�|�K�b���g���}�B�FS����g���H����d +�g�㯶рi�5�I,����� �fjvߘ�Z��Ox���ʔ�]ee7��C
��rMl���Uz.T�*�/F'q����\�Z.j��i�l{�L_��3��-��N�Z�m���t�O�#�#��Y�g
B�~����y���@�C2!�X��8�A��h�}ꘛ������Z����+��g'�G��3��i1�|�����<�Q�v�j�v�`�s8j��S��8��S��.�R�0�0�&_�8U� �OLy����� 
Cѩy<V�F�P�D
�i����֬{v�D_O �e�r�q�Ţ�͢�
7�':7{ovq�N0M=`�*�m�e�e��w8埩2e���p��|�?�4���'A�/乶s�\J
�#tx?�sj6Fh��I�i�{u��Ԭ���u@伦����>�p�l�y�� N��gM��)8�ra��R�Q�U�P�����k�;�r�E,�*�[�Pp��$�$F��(��I`TH@>]�-#�ǟ��^>�nس.��긁$���: �!�� ��v(�"�_��y�+��O9��9���<]�2[��W�|m�B�����ZhO��0�I��j���j����&���Rv�����p�x�ӂ���4m���.�o���?�۩ �ns�[?��z��!�D����C�}:�,��c�u�/*ڂ��b%٫H����h��I��2��2�����D��"PQ*��Ʉ�1mv)Ǟy^�pob��҄\�� �z >���*�ƴut~��l61-
�|K�^��i�H
3��Aև�v`9�ϴf!AEp�Lx���X�`�vʒ��AP>��*y�@.EMlB�!��s���5��/�o3h�
M&as&�8ug�)4�g!�fX�7����W�C.�_2(����^	��)s�;���f�4ͺ,lGmBy����[�Ai@lV`*8ȹhۅ6x����L�.���[w؍��g:kp-#�~ ��A�b?�@�����\�6�UZ�ч��C3���N�Ö:�D����/P�54��lp���Oܯ1$'��U���;��Tڭ�O��R�f��9q3��hO�>fy�˱0��o��O)=��{4���[N��b�'�-�t���CW�n��� h�̎U�x�"B��YWJ"׾H),V�z�NQ��84���{sD����$~���٥	잭q`�����{Q���7ߊ�k�֤�6�X���uI��Ld��.�h�� $j����y���~�Ơzb�ʍs�%����N~��s'��F���t��jn�r+���2V/�=������g!b^�?�-L���d�wT�.�zQ �.�J��I��^�� %��{E�RD��;DD@A@zT D$@H��w�y��rr���gf�<��̐4��]#V;�����ȯ�q��"H����/��i��3K��jLF�ѻ���6���t�=\B\��z�ӳ|֗5s��0��싛R�ON��QA>wɣɹ��ʆ��%Ez�(@�������.���� �ȹ�-D))�۾�I�M��p�߲}r�e���FV�p�}�W�S>���IL96s�.�Q�%���j��F?o[{$E�պ%ܜc��U�����3�9qab��a�����\G�w�bm���(Q��ޥ,iK@:�P��ͭ�*��fl��&Ħ�^R<_������V�i/�F��f�q��^"��A��T��^����w������h�YY2���ݭDk-���Q��f����a�n�Ѵ��:d�R�;��w�!��̉։CP�;�ܳVʯ����MK.�$���xM�[@��?�v}�k���������K�[񿛾���OڛP>0����Dբ;u<��h��@��MLG��ٜ�z�����`g��c�S��M��B-�mh(��p ��==E:����NtZ9��t��K�1�ͤ\g�_g7:3�����{�x=��:9Ģ��`������I젅G,�=�CGǹ߫���|� ��y��p�����%J�I�����'���S�e/_kӺ?$���̝� �R5��4�x�yK�)�������'��6o��t����5�:۬r:ng����9���J�n��d�Xb��17�����h�i��}
6��f3��I&�k�~�S�t|!(�B��ߩ���b�gb���3g~��L1�"QQڸWL���2��ywT�?��a�b�'�[rK$�����8�2ӜY�6�����o��Tj�����=��eQ}�f
W��U�#"��V&�ABr]�LDA�㖢U7q��=Ί�l��D�?���S�h3�V��������8�r���跘^�h�6f[rjU����D��t�\��^yEtCm"��%�/0GB{�TP�Aڙ֎1�"e���C�o��7F��o1e� ��}��b>��Y��C��j���4Ð*�r�жڋ3��in��}��CMOmry�!��0ߴ���;L�}uuݛ��ù�:]��"��v��5E�Q�e$YVj% ^�`^t��Y�Z'�ʵ���S,ń�"?�d�X�p|?��.�2����2��v�MP��Nk���MЧ�������︞��_��˂��Q�����7Y� �9]��Q��^������<�����؇��s�ǩb�>5�3p̊�,�L���Z��>���R�϶�NA��|#�}lv�6��
yPJ ��
T0��3�O_x�;�;�LX��o�*[�t5wW��������+��*��?J�|�ƞ�� �V{5�c>�ڊ�@#�έ~/>Zp�S������c�����j�s'��?3��2h��z6}o�2�O��p7']N�{W��9]C	U����1h/���Q>��DA��r�{����O�x���p��@��ʛ����难���eHQ|2+�b��>�E ���`�0ӑ�aų�����0�~��a�χ��O{[�ʋ��FSv��>)3;��D���؅�N��O�[�_y�_�UMF��Hd3_h�C�i�LY#�jp.��G��I}0{`fl�W�+�'G㛳R�D�2�c>��j�6ke�����
/K�c�������{��m.ۻ.ul3��V��R�b?t����~������Տ�붏=?	�-��=;X�2���BLq:�:�t2��`Э�j���iZ�Jɋ�@�#m��0�:���?B���6`�آ2A�b���l����9�C�����|�h�>��}{�p;?��]�vd"�ݟ�l,��֫����>��W׃V^t=���ߘe+}�"nl��Y�qC?-��W�oA�����W��b�5u�,d�?���ñjd<8Bs�J�~�l��ۏl��y��<����Ӑ�_��� ą��m�d0srq��x_9��lEH��SZ���L��O���V�|����	�*�aA������K�?����+A3��������;w-�� �p���c\�4�wz`TW^�5����>I��6�������5uy:ޖ��_N_��_z;Puk�w=�~���}�~��S���CԆ_�\Ǿ��]
�a6��[�����k%K����bo���&��YyNcڵ./�/˙'�7����o����	�.�Y'��ٛr+ٰ���˨�T3%�!�C�A�yE��UgC���n)�ރ����ٯ{��H��l
�3;x"����s�������m���6*��˓W>9��P��iR.�����`�sW�ͭ������iG��qꝙ�y3v#Wm���f�1�D��:�{�������#	~:��]�y]�ζ�4�,��	"�;��_��җX#U�T�i}D�/1|.��.�0g�v����i1�~����;!�Uc�Z�#��+����!-"�[�Q�O�-<�������O�	����j��Ty)�bب6��m��	_f�l��S�T~����O�9�J587��eY�==���r���;P��-�>��2|��X���?�yw�K�.���;��%���*�_uS<�����]�/���+��Z���2��KkemL�]�`�s�~YVW��k�E��8�H�[[��Ҧ��a�C�V�^p�H��>�wPV(��AV7����%��NӊE�[�ڌ�;���,��'�m3{rf^�"o/G�&���bU�� �'�����|�bㇼ�F^9���SZL��ң%{��f@r�1����6D�	��b����e�p��*����#�^ĳSq�����V�{LL�[ߔ��=������w�xnѻ��dr'(�'�v��?�����>7M��`�
׽ �x�*��j>��o�N'f
�'���1�hR}vϨ� p� �O�� 2�U�K�4��Շ�<+Ee��p��STi*4�zפn&�c��/�1��,&�x�#�~y�V�%Z	�����+	U�ߴ��y�8���6����6y��~l�b�?@9?w����4��k�֍�l��1/���֠Q�����-t���x�����l.�'�B���h/��~׽�r����N4�>@�%�>y@�xz@�ݟ�M׮L�x���Y:6�ʻ��x���g^+ޛw:7��F��5#Jq�#�¾��?�����8�}��=1\(��͓���q��4/]ʥ��Rd�?{�h]k.	����DX���45�S�|�#�i?`Kt��f+w)	��}�L���{��^.��l?�JO��L���Y��� �����~��x{�J%�y�(sp�E��kW���|��E�4v��{��_��c��'�K'��i��jtZ?ޘ%eB��}	?L�L=��	���ɯ��Ʉg�J�t}Wqm�a���!�<w�C�4�C��O4RS̺�������G���ja��u���Lѻ͚4n��T�wY��oLw���P��Of�E�{q{��c�����N*k�tr!ùr���K )���6ϱ�r��*>7"��nj�C:�N�rRz0�3�l��zgP����;��qPl���{�9� �F
ǻqq	=�#)��ʅ[q���K)��E�h��������{�f�%�؞�)�q|�2����0_uZ,��KAx�WK�!���t�:�m��f̩&�t���֖�cʟ{�rz���|�Z�XZ3⑍�,�<�o�-Y�l3���hl^t��h��+��M���}��=��V�5�4#��	�:#_��y��;g'�A�+�w��;�U�u�����ő��;ǧ�ͣ���)f>A���Hw���0|���d�/��]�hsj��(�u�=�t�IM�R�HN�$s횔ђ(��y���n�5��h�~>l%l\�ֶ�MT��L�4d��7ze�țL9��%礩1�O�έW�턽�%��P*��lK'u��w}R�^��=�:��?��������S�M�����;Q��z�&�ӓ��'���:�0Bٹ�`ٹ�۷�͍{<��PZ����O}_��h�%8A�9Ga<U󯽽&lJ�½>rA�b�s��b���T�GKd�27'�e��e��h֌��}�0��Oš{�&=��Awc�J�s���x���MHފ��������Ƭ>B�̈}��)�e�;+i	��s^�~���������\�GU餜A�w���V>dA����%@5$��?���`�"n�e���� 84�.��4�Ո�X�-:��Z��ZJ/��vx�p�+�(�dЭ��'�j�h�����H�A���'1�X������	���^t8d�@]�d2,��3~��i�����Or��bП���F��$8|
���m�߸��>x��S�����"���XF �[(�.��f8 X:diwڿ?^?��o^��y�_)3ȴ\�� ��)"�>�rg�[���%Q{ޏ9�!�}����*�E�ڱ� :���a�%�� �>���¦�#��eO}	�f"��`'�k����Ob��Sk��F�]�U�E^1�e}k�~���o��4ɛN��O�?�+�Wy���/�8�brn�o)g �������*�:>�|@3��ɛ�ܽlRY�Dwy.vX"m�=��0BU�* -xjc�N��y^D���q-���l�ះ��J�i�~��'�᱀���wb���v�+�'˕�;6�{.�e��騱�b�D���M:�Ğ ��ƽ�mu2���E���k.?q�~�j�"3?��y�Ɗ ��(���8F�������Ӹ���P���ހ��.G�	h4N�"ԎÒA���H&`9����+�x�2�y?k����7�|�6�ɲ��B|���F�F䁆3� Tމ?a����\�A[�x����x1����Uܔ� NH���ȉ���b:�1���ja�򻨇7R�~�R�'C!��3�F��S��PR�$>D��<���MҴ�T�N6�#�m�C�����S�/ |��?��!����&������.����5�[ԫ�K����L!M��H9��/�=,L�nOǢ�qfa�����BUCJh7Nҗ)\~[lmR�6ݭ�+�jAY�[����;џ?�MZK7�A��2;Tϥ2����stKc�fu���p�:��+3)�h�qE��4�wT+��#:V��Rs��9'��%��'Z7'���b:f׊t?�/&ƽ�q<��x�X\^��G�K�6�t�����*b��'=�g�����δv��v�f������8z��� �@���l�R2���<�K��S�C���ӏ���o}ʤ�TQu�!)�]]Ezc��v����D�؏��e]��b������Ҫ8#���E�K�����[��+����:l�!�#ﱌ�g�(�:+��|�2��ٯ=�J��&ۈ������`��'c���AR�_K;�av'��*
���e��δ��s�d�>�����'���L���4���XN�uY�3 ���^|��ƴ��	���VY�u)�׼&9���hK�\0c6���y����<'uh�y��@��'g���g�Y<���7@�%U��~��hJ�@K���^�Gy�4'fN�6̓��g��#K�p^P�/��Y&���]&�sk�Ϯ�0�Ζ�u^�&a�@vAb0�iSyք������=FŬ���7C=w8j"�A��D��!��1�4b�;m�ib�a��$%�cef�]�����V_��"A���O��^��t�*��|���tB�,��C0��A���נּ�`�;\�[�2p)�Ϩ����[414�f-�5c��y �J��¿�R.L|�\4J^��M%6O5叅����@�3t�c��B��\���MlkH���e��p��0�$yǙ�����jE���S]�U>�T��s�E��A�ކ�����`H}�1oJ�n�=��>1|���X�>�.a�D[i@l�z�H E9�!xq;�XH}\A��[��� ��_7;�0��x�?�b���fI���8*R䔉ԟ}�_SJl±4e���_}���ox�� ����o�%�o%�5q�i�'���͜�0��i�m��>ʰ�uϽGs�R(�LB��������Qq�Z�,P&�rk�Bc�[�.�ń�����?�Y�p�91)�˝^!Is��"��)[����[�9��@  ���y-^9�4�U A�^� Jj!��b_H��Q�l��YP39���N�I�]����^g9)�.H��y.z�'Hwd�M%H῏	t��sE�#���X�T�/��ɗ��!�6�I���;�Y'���O������-�H^�`��2q٭d�!N� �B�v0��%`�pn�2�o���x(�����,>��i��av�Q�?P_+X����/�.L �gY�:�%Ո~0/��{��5�3'�"+��@&����;�����}�[���
��q�!uF�%�x�1�G���i��B�֒��>��V�߆,�?A�j/*�$T��(����l&1�5�Oy���E�P�H@-ʢ5�%4W'a���'��b�׏��~���$����8Z��S�G��J�G�FQ�O�UGY��i�@���Nk�ղ _f�����$e���k����r�; E'�x�6�+ʏ��O����:��&f�ꝗV\�P��6Ѓ�5S���N0$%5Z��7ғ�v���yEt��6�AC#1��C��w�U�BK߬0S�S�"վl!�1��$"v�Q/��=�I4���#��`Ze���ƭ�;�1<a�,���Dd�-3�t�h��R���¢� ڸ�C��6�Vo�F������.S�������g����f|��Y�##(*�J�1��pRo�=���m|��&4����M-E�@�h��v�y����O�R�fv���?[�r��9pҍ7�EWk����'�O��V��N�R�j���p��"eY�J��E$9�g�´���G|���F��j���-dg�d��R�Ԝ�ޮ��:4`���-��g�slGA��m�7X�\����Z���.5%� lN>K�<a@Cϣ8}�
����C:
�eHl*%$��A���x8q��Qi��t�����Zri�3}K��~�C%�S)��(77Τ*�=g|�ر�1*JP�CO^���
��if}�V%$�{��Ob�c�p�������?������u��������,�������7sͶ�.����SS�����"����;7?�����{>_L�{����"bO����

�ħ-a���$q��:8�I�?�!C�(�����B�0��FY�&�ݚb�{��F�d����ݔ��T�ؐ�������t�B��d��-(r���gR(ِ�V�S�E:��c�2�@�1^f���:Ǘ�B�T!��EK��qY�~$|$Y����ę�"����̇;��ݦd��?j/M����T|lK��{�Y����F �0����ʵ����] 2��o�9�)筸/��y�6��r�� Y���q峑����SZo���]f-�4��ǉ,��׏�R��;�6��s�$^��R�I���#V��q�!�x���"E�ac�>K>�k�C/3*��u��b*&KA仴=J50�f�?�h��b��P���M8��[qkL�k�6>��[�l��%�mа`.�'N�C�څo�:|��7�UfI:Bՙp<8�-P1������]����3������ðD1���}�۩��
]��������?\*�70�/4i���(T�d�)�`k���-J"�`�t/�{D|�<���!!�KZ�"�sqQ����9�̔�dy��x=��v��2��K�Z��a���9��3�Q�"�����$��XT)���~���V��ȭ��$�bp�7CG�K��A�+&�Z��{�gц�B���+�NG޽Y�U�q�l2k�͙���o�wPa��̐>�؞��SMԇ�[2K��v���CD�,"�R�o�آ�U�E���[l�<7X�D5��"a�?䩮a~{��a��'���Rǜ�"%��NO.W�O&�F������>b.�x�6�)��c�O��L��
�A�6���Ecw����.f�k�B"����lP���'� 	��oL�3�6�[�X�5�fs�
�'s��Pߎ�W�߳4x�Q��_ ��s����s!w��[h�4N���F|�A���%S�-8!���P��˔}��\V�nu��i_bժ2�Px}��Yy��p��C�		xQD�<�F��w�m���:Yr2�g�3�4\��Ѽ���֐�%����*}[	$*�B^�tj}����<�5�����)!��r^�CS�U��4�>���]���YM�F���Wy�����fߝ�,G��,���`�dk�e�����ڨ^Z܂��3R{�l`6�/D.��Aa��&	�l���-S������y�~�Z?tj~=28=�-|�9�Ʀ�Ѱ6��N�E Q�.t�>����˷�Ƶ�EX��Nb҇���ܲ��h��uڔ�l4���+iO�
�~G�n��E =ϯi5�m;�8v2�XWԐ}?�*�.�q��_,��	����1k�v�@�	�aiU�@�g5�#?d�_�H �%"�	� Y��Hhl�qՓW�'��x�g+�t��˔�?���)C�s��Ă�k��:��H���@&�!�����нm�@H�j'���hpTôw����B�I$�y�O?5�zD	�0���E�$O���ӗ��d�a�joJm�0�ko؛v,��&��b��6��$$���� Q�o���CA��6�S��,��=���ك��a�3P�$����Y�	���9��C�����p�=��}Gk��UI�1�&��QP��< �1=a���	�$@S&"ƀ|�Fد���k&�l�ɪ�oFn�3V��Qh�gE����-v��M����%�k�F�p��'r9������W[P�Ȃ	y9�Uio�.>�,��R��M�_��T�a	'�����I�����nՍl�.(@סz�Fh}w@@����0i^�bv�C�Ĝ�^f�q�=ϖ�Υ峋:
�f�Ql����Q�<����ݯ��ac֏_�YS���Z��Ghh�##'��/��_hq݆�(<�P766!��� Jń�����ؑ8�7�2��.d��m$	��g��A7x���{/�'q
- ���;�����Z���f�s��+�278�muA7�޽����Z�?����0��`�dX���|t�Æܺ��td`e����3�SF����3 j`͠ H��]���	��}&i�y|*KN�����N$�soI�ĭO:�r?po�j��� ~0E<�|?�|��@�%���O�N�΍�$:��ݰ��Q3
�����6�)r�5S��Uk"�ȭ����Q�}�PYm�	$�����Љ�8R��g�������'�~R��*�3L*Q_x(����K,|/�]jx�Ϭ�ɩ���Q��#�
�7"<��"	t>��T�s="��w<[
�����U@��%�۟Rl�Y���S� x��?���	4 2�_m��0��R1�w���ȉ7�����ځ�Z@�
�g�,��4e@#�-X3<Kޕ N
OJ ��[ ԧ�Q#B�
:�VҘ�Z��l���X��j�Β�C���r=a���Ͽ�k��Zk��H!s�_��� Zu�fF�a�8�<�؂�Ú\�P�;_4�{��;< QƗa<�2��+_G�\����!�kI�&�Xy�<���8a�k�t͝��gP(�>�^j�@[���@#A�?]m����2����������o��+F(� `���-W����q����������9�#3���;2$_RH�dX��KBH��£����*�T��9@����p���[z{=%� ��Ux���#۔�*d$ NFj)��u4�rȢ?�4;,"r�:���Lu8����}"���-ڀ�S�/ⵁ��빔.���ϧf�|���wj1�������02���s��iC7���ހ�h}�]j���6��u_�vE�Ȼ��l� j6OyA�$���Z}��:����h�����*{	������G�ϧ�� �hCh��0t��K�į/�>��V�k�w�j��a�-�ݼ.��i��vE���gv,�о��sR%}D�T��Q��_)�[c4�R�s��5�< �M<�`�aq����v��5^��B���K�hjX|�&tX��&h�b���\w҅�uo4��V���08�8� "G���!�n�m���z;1�-��ƀ�?6Cw˒��#%��J������S��Jҝ�����q��~8=���V�9��fŅ�^�t�*%O>O�d�����c��=ȓ���B�!��������;��آ1��7���@�{���{��wyq��{�������9��(Cw�}d]�H���N[� s�؁|�7`�
8��w�E1���5�߮ng��1���:�������f���qk��"�_�>{����T�U���|�k�w=�����4@���� L|��?:A�p=����pU��Fا/q{%��X�EK �w�O�h��(S���'ߐ/G�Н?y�mݦ��|������ۨ�3~�-���{�r���y�eHp��OlM�U���D���i���Z�b)��A
�x��.��N�Q�l
 �>����p�����[ǔ]�/��rsq|	�z���z"�[ �#���4�O>P���G�#x�U�}��c��u�� 4��v����sN�.����¢��E���f��@�@ȉ�����{Q.�f����2�޼ˆ�
6luC�^�V�qU�!���A�ƅ4U��Ԙ��4��$D�����ï\ F�)��gq؏g������l�ύpŻ���=�y���6.9�C�:�)�H��A�n�@��6N�K��u��0�94ɷ������^����uo@E��.M�NH���8y��i+M�sI�u���Cav?A�{���s0��rz�.����1
�k�ѻ�%X�~p�q�ߩ?�e	��u �B1%���ɾ`��Ƴ6�+W^��%H��i�}h���[e a��&�����}�T����~�\}揞���6k�a��DC�� 
�-6s��z{�Pӊ��|���H�c���}_���C�B
o�h�ۖ�z���z��)1+nx��^���F���[��f�	(�:�'9��@Bf���E�R:�J�6E�AM�3����(�z�
��Q�:���8kN��r�=!�P�m9�� ��f�����Ph��e0VN)��h}N�TQ?uT.��F�Nvf2�k��36t�-e��#����HJ�N�M`7v�/��myI8��FĆ�&%Vkυ�>�2�E�b!/r^�; gZ�=�W��'�M#���gU2�ϸ�nl77S0!���.��*Ц<k�|�y�WAd�+qN�G�:��P�@u�IV���d����ԟ���(2��=WƤ��]��f7����i1N8s�=���Y����ȃ��b��n��]����4z�M2�oZd1��H�/A��	M���b�K1?èGK��L�ŋ�������{��|��wH��*��l.hbJ�-s ���rC{�gOzrm�R���`�8�v��
gVBq�jɴ-��c�����]��������\8���#�����7���ٯ��Y�����=��p�@���4��I��]����*��˔�5�_O���mN����*��ND`��5�5rw\ɸ�0�w�6T>�V�M4(�Xn��a���8�]g����Cg��}a{Y�3�ts��1��V¶X�ySn4ő������@h��I	�ҜD����
�Ͽ=���ÿZ4X�����}��!�+3!�˄ ��_P���vÿC�A��#���R&��\���Y�@�:�� *kk���/	��7x>}��A2!c��LTʍ��u�hL�R$����"肁��4��X�����R�܎�P	A�)���=).ibV. ��%2T݈��Ό~�� Ǵ̞W�e��ٺ�«����E�'46!dF.�Ђ����b࿲��p5�_�E�?߲�?���r�=3�4��  �^gC�O�p����*�C�:��b~������Z�2�83���ӧ�6�vL�Ȃ�E\���F�f� �����&m����v�6Q��e?����[[}2Q�H�~�_���z\��=��	8����?�f�%�7]��r�Y��@�?P�6%�5��4_�(��@&�����s/���Lc���VG��av����t�/�Ȯ'b���m�8<x���'���>B���ٿt>�n��*�˗�}���H�3��1�91��?[��UK�у��I��L��htD�P�0�����ÀfyC�T#��G��9OY�������B�	���V9?��"KQ��d�c�������.�o �b#���0��o���.�b��d�/���!�5�r� �Q���jq����d���;k�53�!s0iၪ�}�L�g�R$���(��$�f�N2�w�c�X0ur���6���rp�yɬ<?���i�ba��) I^A��9���e���T�9ƹ9����ԩf;���A����Vl��E$K%���Wf��1�����-��N���9o�%��!��6M��H���>����Oha���e��x�<M��8/{�T���-@�/V:�: ֭����(��
�K����c�!+.d������`f��z��,B�ʖ�lW�*�r�5���x��L�3��͏���h��������X�T��o�V���A�olv�-|X� b~{��7?�a,6L���z<�1YԜ�Z<aB%wۚu%�vg�P�!��������6r��m�A���?ҐY���v�+Kwub�I�e&�hO��bLC�WB��c���^�>������`֑�7PRW=��~���F�&�����<�oD����>Ex4���u+~��MXH�O�Q�u�e:�r�����J+M��3M������Mi���Q�?��&�U�RC#\��X�)�}�zѥ��!ӯd�h�|	��k� L���ȴ��r����pδ=��U����+�pX��ʃn��q�R�)�D��Du1O_�F��}s.����1A3�=H����LO�,��J�_i�?c�/�O�3�\B��1H��)z�\ށ�hH᫖���L�cGC43\��v�V�z�e��4�sʰ|��Vts_3yJg[�����9����F+�:$��9��| �0Lj���T�w�(<�J9�U���B�lT5�hQ�Z>L�	ު 
�Ȍ�'���>¥ T`pM�7i���W�[0��xI�z��0(��n�L���a��=������ϳ�I/��T<{G����vЈ�׵BS�B�{
�*�H6Td���m-ל"apnKE~�w�'��y���zƙf�H��/��dءzAn��؇tD��.�u:m�X��Gk`|��,RZ��t�s��/D�8I��6o����S�I�"�l�a�i+rl�����|u�e�L������-u�6�8�7��g���2��
�O���f���SG��Ϧr�|Ps�.c�7E$�t:D�v���Jȫ���":����j�t%��J|��4A��V�|z������Q����ъĽ|
N�%%��>;t�Y*�K���"&���5���a�"4�1S�H�Q-D��#c���6������S����$P��3�LpZOj�Ht[��TQ�O�k}���x ��Qzl;��O��"��n�A�U��p�@�}B��
��O~e�ƗN�o�ɬ@��5O��d3ڿ���/�:t����UsO#z����l����u0r+�UTtl���<H�"=�������]��A��Y4Jn��T��7q��!���I�]	���ې���m����E"�{'����^�H�?ajP�zOaL_=���{/�,���F#�S��l��I��!�K�9������Hș�A'�hJ���.���$�x��"���n#��V1oXszt�h�ِ��/�J�*�ɱ����
�����%+�r�x��8���7��'}+�C��%�	ۭta���GQX�hH��;���{Օ�Qf!!�������?n~)4,~�/&��yޤ�դs�ZQ�48�SI�+S�+���pB���x��h�;�j���X=U��m�U�ٴ55y� Z=���)���d�.q@X.7e�Ol�`b:���d4RM��.�M�ԣ3���:�Y||���e�뎬������W��3�#7�шck���n>�*��g�;�}��Z��^���*���nɤ�gdiBI
��r��t�<���71ٵ��@`����(��P�B���q�u8E�f�"7\ .�@�u�a8�=ݏI�e�m�E�)�ޓ���y�5����n;���X�����
� '�/f��	�,}����?��y���F#�����P�^�;���6m�h�-v��(��3W
�j幉L�6����ClBO��5)���-� T^"We�Q�����N����_�@9n]����;A���� L:u�2���NCJ5v4 )oUޯ�Xf�3\~���`r�T��ν�jpr�?c�]R��$j�ֽR둔�(c^C�����k�q���YP�Ph�\n[kn!�Ӄ!
N�F=�Ą3&�(�s�����3�厜6��y�E��aZ">�L M^��KaJւU×ݞ+��σP3@^����J���K�Fu��E(v�C7��%r�X���`B����~�r�y��z�i]��xl9���.k�=�˼�f�ߠ��BL	b�*ݣiĭ�ǗŅQ�Q*GO����e>G��*�� ����Hg�-1G��1��d��rY<��}�h���>slW��'\T�b��զ�d��<��M�iȘ�����0*^V绐wLIS�E���r2Ğ>\�a#!gL�-C;�݄Q�ST޼�����X�,'>�ۦ�I7
����.|a�ͯm�E)�u��y��u�[E����N�������񷼁�G�Ċ��ZF�� �l�y)�uR�����w���j�d��ւ;�k31%��ݹ�@t�8܄$�� ���o�F)���w�sMD.c�ϣU��]��G��m'*:,$7��ڈB�
�i��Fn�ZT?�?�Owv��������$�R�c��ս��~cr����Ժp͖'�֤Q3qp#��z	�m�<:�tF�uп� �r<�f'���Г�1��g��}�Yn��	(��1p�ُ���J5D������+v&�zhid���%�/ZX=9�x��5&\;8�ӻ�4���?u;�x2�����ӫ�!���9�����M?hӘL�Ă�J�b|��o@)�CƆ�{���۠���\��l{\����A!��LIF�f]`�qF�Si8S��E2/���^�C� ��8S�<P�XUQtRsI*��?]���������f��9DN���K�Y?�_�Oi���6~�Ěi�Ԥ�<T}L�?����)O�d���&��հ���t�|�撆o��PC,���A�K14n��#fO�O�#�8�
���P��-��j�-�
֨'kZ$lO�d�$_�AE|�B�-�g�^�������[G���p��TƬŴ�<����3hgK~���K�&�p5Gj��`�$�O����2��+S���f�6'��[�ʄί�|�<� +M��@�F�9��z����셲�kwɅ���"��U�;!�pyA��q�1₢aA���]z ��7�V��&�t����
G�U`���o�O#��ї�~W�+��O�s��y�k#{4�Y�:0R�.���y���q��#��5����"�ќ"vĢ��P��nn�%�nD&�9Z'� Z�ỿl�ns�8��#�f�9m�n"���U��>qg��jb�M$�R��Pd�y�d�O���/��o�Ao��V`nk,;^��?���z2zx =�ƒ�j~�7�����t�fq�H��.�q�.�ot�����_?<B,����	��*�I����3gƂ���P�����3��������M[M�L�§? MB	�)&Ie��i�/�4�y��τ�YFy{Y��η0�@�M����Q�����W� �n�=�R������]4�'W�|C &�!a�׷���z��H�'֕ۦ��$x�g��ۘ�v�lj��\3��B�Wi+�ܙ}������؊� jk��>�񪣚Y'�u�;)�q�DA�ڼ]c>���J]e���>bb*%�⑤�Q�������P�9S�e}p�S���G�z�m7 G��H
�)���y����zS��Mq��i7��]�X �1j(@�E[���F���0�h+�°��FW�}a��0�0n�]Aˠ�n{���/�ˤ��c�H��nA���Wry���F��ϩ<>!'aCT����&�iewx�r�_����qi����=��[�W\�'@�T��Xn9���uk���I�F's���!�ﴍ�H���ŀ� �I�V|6�����������|��A���.���G�� ����]�����ѯ�<��i��� !���T.��؅	��?�*���0�&���D�_�4��,�� �w&1������ڐH���E�&~.YzHO�p@P0��b���)�u�<Ri�jxJ��I�e�n��R�mB�OW�YG����@<E��C����[-���	���틆�*4�(&�ɏ���x����0��r�@ψ���`q� ��$Y��䂼��ԅ'o�1Ń��^?v2�?4J|s���@ϖ��"^�}u9��60���@P8pj��u��#�>�#�8���K���H�����>K�2Z���D�\�Pd̹�hÍK�'���{ۇ~)�_k:P��� w������JP��U�X�Z� ��4���]?����VރcC���>~
�Z#P퀁����H��u�L���/�ĀJ'�d�7��SPP��i�~����_ꔏ�2pS꓊���HE��91�<��|�>�A6�b�e	RY""��qe
59�W.E���9'é*!�i�	���^ �(�}Tꠙ�2?ݜFy���QCk
�~f�i|�$���F(���a��\�}{���4BB��|�I��8>�C%��_�8�p��I�X1'#�"5�/
��Xq6kP`M���.����`�.O��$�u�R"���l�!���a����!|6CG��LFc����ݟ�b���'Ќ�J"�FB���Ov���_���{���?���V���,�?��}@��n�/��������+@�D�t'v#��bi_�?��榌ʱ
���*��}�>k�����Q�����Qs�Ś���94Pc3�V�@Q`�s� )��%E�I�'g�ʀ���K&��͋�$;�����b�d���H/ K�P?��O�3���$'8����Y�KøSHA��͒�"��� �)���1��ԋMg�Q~�c�S �GpANe#�6"W⑘�M���X���Ơ$YC�a��o�����W�;�� ��Q��`nt'���B���)I� ��A�D�j��$$�灋C�<5���+��>޺��� �}]�B�_�A}���F�/�{H����p�K��Bys6TC��<�S��� ���������g�� ��"@��`��O+`x)��+���)���~	�H���G�q1�B��X���`~�ͤ��)�6��Df�jX��<F{��[@I �(��� ���K�,��	���4BI��c�'�F�G�!�!�1'��*JCA��/л�V>�s��ؔ�D����|�nAӣ�1�� ��2,}�W�-�`_b���^�'��/@Ǒ?�<�� �T�(b����d���y�$҇�ƌI�Ѵ!���%I	�ȡ�� ���� �@@v]f�ɠ�����|M�3E�~5Fr-b��.>9��/y`�4g�L�W@I�n��b!
<���G"�戟�Y�!/�	�6�Ԅ�$���`��=��ȑ=4W�+ >'3Y8��X����~2b�;ˉ�m($���s����{mV�(�!g��1L���[B.��D������2�(�\��x���Lwx�lA�N��:҃qP�@g�,�6g�*GI��ݑ��O�� ���H8�?v�:K��"�d�k04� $�&(+"y�xF�C�$�EoUԇ ��i:t� �`x�xd#����� ���� w�>fn���u��2�DI� ����ne�0�f4��(z���W#�['$�hx�?}�� v8�ݟ'���.�=XO��W�TT=E��70�"����H� /V_���Z��Q���濱�+��P���T�I�\�Y�\S��?�Z���Wr3�?Հ�H9>?�5� ���3<���)o�T�Ր�;�1�ٗf,���?�#;��?t�u�
b���'G�wO�<�9��z�!�CH�A�?�v�\lG������ CA(�f���+<c��Y8��EG��H�����$���Q�����J�)?�JF�͉�{�	�P��c�?Ő�d�}4DބT��Qax>*t2�̈|	���%��و�s��e��#l�X�ЬmdY3��lI\��[���J�� �� �A�����c�={�܆W�7�A�O�D�pԔ�dL��ur2�^^N�E$̗���H�+\�A%�oL?���p%=�T`2��]%��/#�L2�9!�F�A� �nc��9=ŁwYc膊۽� Tnv���.�t䝙���� ��>鼶e[��L���>(�}��P��Z>z*�;�JZ#xF����/����ޏ�[��G�\�il^�`���r[�M?�� � �
9(7!t��4e$�Y���'���ϑ��+	�\��,Z�L�M��A?��ऋd<, f@�۝i�Ic�0����2����5Q�ر�q��6a��D%�ʖC�*u���eS��;<Í��YG��N������Pb���_�ZGJ(�pC���^)|��(�џV3��r0�I��@"c��k��xOyWm���U�wr�#��SI dsQ���T�|��_53aO�i�`��e���1�x+�c՝?��4��	�����DO͋a@AEf��"��?�NW��V�C������IP������*�~=��q)�H쳸e�JU�'��Z�(~)��Q��d�"a/U�i2�c�r�h�	����wuN|����� �5�C3}��Ψ�`d̘pL��V	�� �tG�byYy�l3`�R�+g!������ ��qv�t�2�J8_���Y�rOȩL���+H͝����ϫ�T\?{��I/ZE|����#'*q����D0G�B:�ؘJ�,��B�rV�W.�,��dY4WN�*�� t�R.�<��P�"x<���U�(?dЌ1�D*0�T��'��d��4�<XXF
�)�B�<�Y�?�U���/�6P�<A6RA�%9�e4�ls5؈����;QA!�g�e`�������|��Dh���e�'$Gӕ,�b���O�N,���� ����F�������7�ϋ):�0DeX"`�?�����P(e;ŝY$$���@��9���w���|mn�T� �?��E��Ir	-�1N\��I
s�G���E<* �ǒ@��e+B ���lT��?���� �"��Oz}����� ;�G�^��01��H ��j_�'��2Õ0D�6;�n���-?8Pf��%H8	����I1>��e��(S��f��L��a����xb'��'�bnGȌ��hI�F�=&��(PL	�i�^eUR~�_�*(�¼���f,���	�Tչ�c�,�"�Do���UN�Jy;hO+�� �?�G��4�~_6|�e���j�C㼴�G	� Uy��#��d];~b��4��E��ByA�� ���
$f�T��xR�8Yx��._����t�:P�8��kx.���j���8��y�+Ÿ ����P��^[��T.\�v*T�� �E���� ��]�dt6�S8|w�aϳ����%.¡�*�VQ����5v�/!�_	Zf�VTG/5�]��c�T e5�f]�X� �B��q>o��"��s��(�bJu�d�Yr�<E�_�NaB,'͌�:O&�,ę�t��({�����S��v��֪����� W�C�ETI$`�xy�!bL��X'�]	�I�v��<�r�|P\pA+.�I|T�A,�;z�=4�}mVTqϛ'�^����z�GP�C������\R���T���(6z��X�p�My>���ڂ�y~4I������(0
�y��h�D����Mj/�~\��"6y�<Vo�.p�4A6����(���;���ʠ������&���H����h���x1pRP�'������L(㥲�R��������g����X�a��),碡*#�� �� %�xFc�K��*Y��Z���-#%%�7����?�U���0�|Y�N�QE�������Pl��p���-R���^�'�d��M��+S� ,�F��������zap7���@����Q��u<V��?����B���*Ý`,��N�(�I�&$��*D�<����	0��!H�K=R:	.��u|72>h�\��z��F����U�L�9�X:"�#�x���g��+�����:���>�(I]�M�����?�@ @� �6*"�E��$׿�jŧȧ���� U����������c��(�'��O�f��� "~�JT�A&�]��
:9�ȱ�,x5�k�`)E���G.�CS��<s?=�ڰO��g�r_WHO�>f��(�ZBr���33�U��=���2s�(�)�y^.C���O��Z
1���GR��y�"OzW5���z��� ��:i^p5�W�jdnO��*`w�5����^��=Y�9࿫}���?�����V��Z�g.l���%� G�`�QGV+!%�±M%�A)>pҬ��z�Ǧf}Vso>Ov0�t��M�&��aB�� �E9�_�Vb�'�B.�,�9O�b� �� ���PK   NM�X5r��W
 zX
 /   images/cccdd3b5-475e-4e4b-8694-ce23b104edc1.png|�P\O����kp���ww]�.Y�Mp��� ���<�������[���N����_�Lw��9�Td1PIP  ����  2 ���p*:!^(.r��  �_(����3�'o-/�@�3A �� �?�_��_�g� �����?F �����Z��������b�Gܿ�< �	����)�)%/��i�;��w�0PU���������������#���������o������aN�����.�#������쯩�^�a/�ZOY�J��L������Z���J���ZPC�ݿ�?3���=<\�ٽ��ټ�ٜ�l�9�9�ع�X��`u�u�0�aur��G����[�ٺx�:;Q�57�p��y���5�<����ǒ�����s@��$�l���ak���K�L�?8῔	������m�x���D��������"���nRΎ���	˿��-��&���X����6��_M�uA�����_.�v���f�o������\����A���z�����Pu��sT����߼�����
�����&�*���&�(�Q�K ��"/-��u�a��F�����jq����u�ŗ��S����!!a�����ɂ���zi t�V�s.y���t+�h3��ㆺK ��s�ѻ�oぁ��`ď��y��z5�ggg�̱� ���8�oFSk�۴,�~������Uy�v��qNNO7NN0u*^m�{N�):�[!wS���y3�����?��	[t���)[���DH���I�ۣhB�R�[r���s�U�Q����C�܎��E�DbA7��|||WYs���kMg��>ʇr���3!��}��������,���R�s�K`��.���e��ht�����mV�Y��Эo`����}�����h�����޵��3� ����^O^{�Ɉ�L��g[�4�cݴ�@�Ss�]O~8����gYVv�g�j���*�f�Ɠ3o�����c���ƪ���?��1�}t��K�P.ˏ8=�ݕl1��ǻ�;�ڐ>`��]�.w�NX�-����6W�w�~�����'<�昻.�D,{�/W�*)L�.�2�������kw?��=�*�&�p��Z��mVR��`�J���{�$�!���A>�X�2�F�Ӧ�\b4k*� 7xҫm?O�q�� ��>�l�ʛY�'�_�z],��8LMB��!TgfR�q�%9OxF�%�C��Q�F�ݼ�,��T��0T5b(�@ޣ�����6|�<�k���yzt�"n+rBSPnN-f��8O_��8�/J�Q�5B��C�����U6������
"���l�+i�І�!���R�l5���5:!w��� 2h�a"��-#�(w�r�@@����/)z] ��5hГ�c����o���ۤ���a�ۜ�T�Q;a.�P�ll���RJ��4�ق���틩�C�լ������h��N�+��ϛ�[<߮�ŉ 4��w��"�p<�8�~�E�/� ��q��6D�G�9"̠��N	3���7��&��	/c1$��	A��_�*��N�*EgA���^�H�=�oи��Q�!O�B���C�;<^ 
/x�$�����X{�!�=�8�郙���Ӕ�U�,A���ǛS�$ִ�Y�i��+au����v��JM�2;��z�\LT��3N�W�먏�i�FUs�Qz��"`~x�.B��py��*k�1d��_D<{'\@���Xr^{FoiA�H�ӟu�!�i"Z��Wḋ��ӥ�t;jG�|ɁԨ���a~?�\(��D���gw��jy�(�{�Q� ���G�יE��������8�կq%8v,��h��ף������^���@�/���Ƒ~�~���o@s5�PT~PX�؇��V[��`H8���SP��3�6�Sl��_��T]z��*�ց&ޓ�����
��ҺS 0�j?y4z�-B4����eI�q��MK|I U���Ⱥ��"�%�Y:��p,f���2�˔L"��d�~8�y����Kv�{7@(�ū�>;��������U��'��\��q ��My'��nT�D�i����b��^"�*3�� :G�T��k7�\�ČU(�:u=�!���Y�<�c���z�V<8څ\�2W�(���:J�mOpe����9�Yb��I$�d S?ù}�C�c� 	FV����6%%"�F��Y��'�����!/�r_��Ю~����[��:g�9#��R�%6w&��5����h@r�ySM=��Ʃ�LWl��6X��2��^��l2��(��f>N���z����|.2IU�N1r������;����r�s������q��I!ka.�d�kV*��0^�����W�v�.��!�u7OO������	����,d
�)A��i4�����Zњ����u�^vD?�Vʂ�_h��fb��#�8�8j��c(G�<>K���:Ӵ�Y��'�)�'-^G�X����%�6 /�	�{!�+3�$�:/S!83�
���M��:/c�$=I�j*xmgns/�ڍ�ܵg�;�d*�>��r���A���.���$��zM��tT�R�Пؚ�������:&��ϋ�C�O�]s�O[p(��U�H�B?�ߩA��ω�뾵�C�GS4�v�|\��t�W+�6g�J3�>p�g��B,�r�Z����B�Ƅ= �����{T���%�2cL T T�iC$ ��|���Q���8�C�$E:�����)C��r���������]��� ��������tr���o�(�%�|NgGt��e���90a�ׯL1��dD�9�t�_�>Y�5'ܷ��`�Hi���՟߳w>J�ՃJ���bX+�眉�\��YM���4^�Zj��R>�(������4��_7�6��7,�Y�W����t��Dl�����'���r�G��$�w��2݇A�v��7\�v]��P7`�tMc�׃.Ԗ_���yd�T����:�}���?�֪�x/���ǟn|��Ce5;rUt蚫�n�5ٛRu��W���d<�JP^�^�Vh\±��/:8i��:�t(�lpj�-~l�aa��N䟸TEw���5���dZ�|��i8�q���[ҭ6*$`qf��1cv:�Tg}�=��;P�="��0-�,7�u��3��{D&`挸�\3�-�^k�Bܓ(�ξ�W��p�Fr�	�WWn���H�P�'��f_w��|�^�ԫ<}�ť�l����Ou���XG#\/�kU��%�V|ġ�ub��T�>���9u/f�,;�R��ℳ�|�l��VI3s	�l&dT��'���յ�0�8-�I�=��D�k�[Vz��M�3�]IOu,��|���2"ç����]�}���S9i�D��p��#�!��H`�����AU�n�9�V�^-r7�hF���v��[Oj+����������X���+o�Л�"�Y�0���T�����@@��I9��Qe�?���5`��[�"��J��3^3
j��]s�]'AhB�x�C�
g�4�|�®)Y^��tH4�
 ],���M"$�B7"4��r�wid���1�T����v0�
zt÷��䐡o;�Iz�P����e���ԛ�CZ�F���� � ��^����5���C�����T�:J����g��H��� ��頧�W��ѾZ��Ş�ޅ)�a#����1�1li�7)���d]��{�(771�O{/�Di��@�5�^���O����}�h�*mN�Û�?��N��lM'��ג��#7�LL>B�?ki�I|�f(��5�Viؙ�][�h�.�BI��h����'�tu��F��vH����G�pQ�:	�X �����cp&�en��͙'f	�_��z�<~��;^�,�٪I����c�zM`_�~U��L5>�7C��Yj���u�6��M�++�me�;��t䋬�D��6�6"�$J�V{\l��	�~�0y��/�����g��.�1E���)
	$i�kJ���x��P��?�K�#�G k|	�B=%��	kXXP<W�5.���E�iuuՒ~h��XE��}�$����7R�� eL�7�8Ӊ j����w����f����T��1����2���x1��x��Y��/(}�E����K] ų�T�c��W���1�0M�8\+Hs���a��m��C��G���'�$j�+�;�.F���D��b����cP�ұ���������.�.�V?�+�EZR�|"�J��/�uѨ���ʍcKX2az���8L�U�/r��]׏��1���Ox�Sۨf��Cl
�w�a-��!:�kH�1�l�ˡn��sq���Q�[[�)�k�߿�[Q�(:d6��{;�)�Z��}�Ԝ���Y%��-7���J7vY�u�:l��Z��t�ޣ����Nf���6��� =�n�GkIFH�m�}���qd%ަ���g��:�;����<��G�[�ɻ�����hfe�(�U���r1�q2�+mi}n����߲��!��:LBD.ۂ!�L�̾+�n<��,Fc�����M*�0�(e����ʪdOl����{�Wz[�ޞ�?[s��Y�5�P3��oj�ҵ�j��X���w���_�ë�����?~��s�x0|�Ԅ�M���P,�Zr~ɘ����b�E�j�O^��{��cQ)k��8	n�g��!N��E�����I����ֶ#�B�I'���;-{27ɭ����pЗ��ao�B�'�p�ؾ�e����v�v��)\MbFs��&��U8:z��b遦K^��%�Y�ڜ6��_����C����h1���u���x&��� ah�����D9�^#/�">і�a��>��+�^^���Ѯ;pnBhh��A��Kw�Z�
�#:L�{a�r����TH6��QN=�E����Y���x.��b�eLT�X|ʃ3�͵��޴Fh)i^@�}o߁rὢ���>5����qwh���n�7=�z8�2�'W�qO�wH 5����+`i�Λ��9wfS�8���E�ډ%a,Qf�)������]�T���;���7�I/������K�d�Fs�{�������e#�	]R.� �R<���w��Ԟ��]E���po�p�ͽ�����	!v�'�D埖^Q�x�8��dÝ�VM��g g�L����L�`���O7͌br_2��Ų�=�V�C��z� �����h��p=�Ƃ}�C�D�h��P�� L�z���zF�JDR�Uyݖ�b��:|CM��q���W���O���^m�KR�At�s����0���򍯋@a�&x`�
_>��j������ ����)�wgUm�xEu|\j���z�r�LN�����O�� �kr�O�^�L�	ΈS���R�Ɵ_�޿S�{�V��	�ŰC��ܧ �r�dd@7�c�(fW3{=:��P$Zk�v�t�m�zΙ�]K�h����oo �̥�����;Ř��_W��Ωj��G��>�<��v/�乮�z�����a<
��E$����9-0@�yMoK�'�6'0U=�v	�D3����p:�7����պ���G
�1��9�<
��p�'�{���s�>,:�6���NM���j�%w��!�����ȧu���9���1��{��#9�_�������,��f��^�a���j;�vY��)��2�,�����K�;�2ϧ�ٕk#{�0d��dQe.�@�ho�6:�����;sE�TUʩ�Ǒi_�`��c��#Vb=�@a3H=v��<M9�yn���7����\A�TUImX�f6딴L¾�VH�D���iN�h�b�;���+�w��>�AS�$o��[�_���r���̑��� ���v[><v
9�K=�1��~2�(�~w*�W�����(6���TO;� F��Z�ۣ���W/�+�n�E��L 0�]W~<-Yy�A{_��;m���Se������E���W4�W�EB���P5����z#��,�]�Rk��֯���d*�� �!C:�!����\3�����C-�藥��eC��ި��ù�>D��%�&<B��%k���;��?�z�0���JƘ��,�E̴4q��~�æ{X0�/+燐�:���̰�4!�Av�A�1�?�H2�cx�M��^�w�vlT�6U�b,�=��+ܖ��wD[&��&Ѡ9%6���Gom)p��+�ߪ��R*A�K���,�[9y���ӱ���3S˟������� ��f�Ft����{���Cb1b�e����3u�I�v"�s"�����n�b���of֮~�l�K�rz�e���RAv�c�r���ƣ�	h��T22������+F	�#�C���
����*^7(հ���/�4d����Y�s����M5\�+/��&��"�}�~�D�/YH?��FGP'�0�t��ت`$��om�!:�^�Hr���쪉���=�SVZP��P�����jv���N�yv1v����N4kn+<����?;��:l���K,����3(��]#������T_���t�|�|�2PW��y~݀����^�������I^�hR%��6��o�4 ����&R1,о@����n-d���Rk/��2͝���+��M��.����r�$e�Y�z�V���Fw�/.�x81�@n<��Oz�M�H�̓�B����=5X�Cj��1���&�o �"xS�`��Ի���'�+��h��n��O��JM7S���U�<��&A{��t4�jܺ9u��ĽS]��XZ�s9�tq
M��)y�rm��k��f�6
��?9�QRR�;�,���y���s�����rx��Q2|&���K��A�nD���è��'�4�E?Kr6������f�O�z��}���!�:��ދ�Y��)�O�Jt��ch���E���{��������v�U���K2˂���<G{��
\�$�Sfbz��ʹO���.;��[)��8�?a�l�ݶ�C��$����B���c�.|axftF}���'����b��k��tݑӔ1h�9S�r��'��" s�����)E�~<W�Vd������7�引���U�i#*�t$�k|�vx�\5]�ǲ��٥��Q�GIN�.��g_弱��B� �1�"�,iDq?���g񋫔��ͭ��n�]8���\�w���P����G��ǌ�x(�\�y܅K�v��R(���:j�K>sd8YD8����$?���;��P2��<�YW�z�R�=��eF�MD\��[pZ�������m�3׫�q��fe�Ɗ忾�x��W#j� ���_�������'K��ޅ)�z�w��i��/� R�xk����_;��`՛s�@�~j���$������L4�;c�[���z���S-�k�	����'��e�oЌ�=�t�1Ar�}%V��禓���%7�P�)�ߵ[�tQ�GQ��04zk���V�;W��l�=���W n�G`��9�3�	��UYZ�y�0��)"8)*�ȭ��@ߪ�HX�ӄ��G!I*R%�,�NVdR�TJ�}���Sp��ntډ���)�J͒�֣}>�_�j�eg|Y����l��.�g�4��ь�2���k��+q'��6&���K?�6�=F~��D�ĳ���>txuijq��Y#|2i@7c�/�^mA�����}�x�#���a�U3z(��W��ETm�+/ҷ�l$�r�s��x�z~��h;�F?i|� �k���W*K����:}�۝?��o���V~�2�G�D�	�7S+fR��.�<L�0�_����Y%�j�}�h7x�~ж��:���d��4x�o2q����<�#�
֙"�p�?�3l�Zc���3����\dF�D_q�W���\	y�T��s�b�lC������M�8$3S
�E�ҷ�= �.jN�&��秲A?~q�%�`5;�Z�lr��������u��`R��#^��
� sv1חn�P\�d��XM���������%��W��5���9����ۖ�+շe�����-h6�Ns{��u
�'�˳1=�~V27���A��$P��ES�+�E��瘅X����%���A���\2��!�����|����y_�iy;���c��ӭ�qd�#5x���U�v���J ��Z�'���;mY:���A+B�JQ��(��&A�X���m�S)��V�D�ˍl0oe�q��]Ns%Z��\R8b�˼�:�@��*�'D����$�巑���M�� ���ӗ�5��\4]����w9�������xo�jk'�s����Y���nCD��e���D�a�JY���"�Q�aN,k�%�1����կ�"���@j�35�mU��f/xߊ�"/^a ��6��g����u��hW�B�p@1R}�w7���G�^�_j{�O
h�i��j�o�7л�7�"�2�@]3��u�.S�#[zj�;�wխ��uq���Y��K2�ڭW��hBf8���`��큐m|�l�c�k)O�O�d�ŅB��Kh�p�֞"D6���w@n��@6���L��y{��]�_���w�?�����Ϊ�*����jտ��e�B���.]�y�����:8�M/���C!����YaU�|#ߝLY����� ������=8o��0:�����;���2?3�Z�`@Q����X����N;���N|̷�^��!­ue��7˛:S�t����T�l�xQ���\�G2R����L�^o��{]4������Ht�:��Z���vB��R*��F�5q�.���ɽ�a���um���#�%X�������]s�w��m�Rݻ,2�r����6�b��y�1݅�xr�$`�M�9�&�48���,�~=�}hkK�h��x> �l釉9���~�
͖�)Z+����l]��zml�2R�d�>�k*3-"?_K�������X�f���0c<���t��.���?����Z^@l<'��y�<V���u]xn��H�l7ae�,�:���H,��o�E�З#��,128�xy�'�Yqi*���:�3�^�Z���m����*���ÞX��@¥(i�ꯖu�]%�����>It��'�*`X�ޒ��\��)L9fK%UW�������d�"�y|$�f�kie��f�by�7�j�kN�q�����G	s�w�a��'��5�1�F/^I�H{�_�Z�7�a�xݩ�c�9h|4��@b�� �g��,��[�V��De�螶4�r���c������etL���9�*g��"�?� ���u�L��΃���-(�OΈ)�%?2KQE��	%`�cP�����"�]��¼�;-+��I�yQSz��fT�%̎���m���}x��b��%,^���HR�K��T۔�Uo��Gܖ����l5�O��_��E���]
�0ԣʹLNVvsu�;
r��MRu"�)��"Q�Uo;l�ײ��\��U�!CL��}�s��8Է��x�I|E��͐"�c�I�YI=V��wB2I�Ôba��h��C�@#���y$a��q
�S���5�� ��z0U�cOe�P�!�+jؼ�p�)V3�?�4�i݋A�h�����'�J��T���$��?}a�I�\���ج#&��?��&G�uڗ�R����O�q�Ix9�Q�&6)Ö�D�K-��� .p]��rw�SϬe��]�� �^�^]'�K>��s>�#��bGoƻ$v�[�_L����I�E��ǄXa��{D�]����S/v��B�C��i��X���m���^�&,Xj�kK��>0�+,��%��6�>�,�`���(���	=�|�^�����K�$lB!��xc�=Y��y�Zw//�B��P'�^��)n�5� ���H��:�,��g�Xs�ș��B�A�o��[���p\����������$V1N]���O�rԊj5>lc9��]�'m��p��Sl#�-�I 9Vc������dqa�Z䦐6QFc��3G��;˃5���������X����R3a��T����/�ՙ�a���n� ^-E}d�Ud#4"�(��<$�E܆��J%C#��"���#K��Ş�K��W�7�n�R\W8Ə��*Ek.�>��h.^�H�Bg{��>�t�9���� q�AoI��ړ�'�g���(1:Ğ�:o�:����U�[Fw7:�jG���2~�Lk���RS���-)8������������	�g��w?��x@Æ��]fɖ��N�Ԍ�����f�	վ[�Ś����Cv���~ﵩ%�U�TU=2�|$��[��a>&�H_;��Nuq,Py�W����t����X����z������ů�B����~���G���̒C�)�쥲l���Yq�������`E	h�������6�cy�jjd��GL������rGX�ƫ�u�MQ�)�>������|� ?Q(s����3"D䉄�F"c/V�� I�ZUe��QS}���Ӻ!LR$�W��q�ҳZ�K��Յ��IbޝC��������^�G<���l3��1%?~,�(��<Rr1����N-��I!���K�������*�_�W5�o���.o���T�里��_���V�&%���f��g�9�O�{�e��^�B{���d�gUꏳ���	����E:�A5���2���v&ߒ�P��Y�k���6���4�5U>��F�~��e�I�Z#!Z���ͻ�L���?:n��b�&j�	�!��ن߄�6W��2���`�8R�,1�`"����X��IY	���Z�K�?TeB��0V�E���V,�K�;ݍ?��4�%U�r�Z�i�E��:��۵�uY@|��aA�^��%)I��Pn�)
�~9�i]`��X��/�
j�59�-�h���O�	���=�iU؍�TǦ5���a��� z>p������ñ�3����MwR�(ի�]��(� Y
���MmN,91�'w.�q�\�_����I!�0�"'R�mI��r�4�4j ����2c���)mQ�s�*�
m�݋@'-���*�nts(*g����-���'EbM=�����Yl�G�+�2�9��v�w�nl��oF���9m�.!��M��y�f��\K^<F���P$��JWߦ�%tX�=5�ح���f!�8t�9��N�r���d�;F��>n���{��10'�0	$W?�M�(������xo��()(aѩ5y�;��*�﹖+-C�j~��x�4�?]r����/^-�%;���Nt�����3i�9����_���c������jQ;��û���C}�1��ވC�͕w�FӾ�[C��gY8�O4��6�/�d�ݎ#[��A1S�����۴T2ט��T���ݴֵp�oTM5����9��0F]��)��bi贈C�=���gt{��F�9Ṋ�����V���n�~�1�Ђ���b!����\@j�}���|t����Z�9i� ��a���Ǉ�\[�"���:=�!�z����Z��K�����@f�)�o�f���>"�w�y��I.<I-���p?)w�'�wP㾭)W*M���+��������WQDL����C���t��4q��
/�D��E-�0�ʅ2)J~��1�i6=�$�{-��9)�ЛD|����#���qN`xnt��۱�c��B��H���>\`4:s1m�x������q,�_�U�֪�.����1�wZp�{�"DF�*r�k�����Y�1�dwx�����͌a���]S��7���/A�g���U?X��̛��"�cC� j��\�,.���F�~�>��X�?~1��o��u$j��λY,W�<��)�G�Z��L�D]o�C���n/ǘ�B��
?�V=�Hy2�.4�Y)Sw��L�ٻ�ߚԄl�9�孏Z�l�H`�E۰�����J��M���7�i�1n�o�F�n���ﭔ�׼AC�F�
��
<�9�40r$:fO�-�&���xߎl���=��Y�q�qM��S�Kz0,�K�I_maɂ9}�����p�I/2���Y�y>m�\���Ɛ���əG�Bf���Y�F��WO	,�s.�cۆA9{����)���?���G���/�T��b(�"�Xry��?��#�u@(�e���/��,!��hر9�͈wI�&��@���`�'���垈�G��u�z�3��U1�귆?�j%7��5\�u�m�]O �v4�IErKf5{N���b')7�Ӽ��;� w���(��%�,D�4sq�=�]���~�Z�)�����X�����C�o>,��>,��ڝ���
��u���I�j�Ga762���R�S�}��l��������|��[_�74MXG-F�ܱg*MC���>	�^�d�������(�bc���[Gl2��^" �v�E����S�q�%B����nޢY@�|�z��y��$���~b�->[�
V�����d(�!7��񛖼���v���]]���<x�'�i���5k�Z�F��,ʅrm1z����0L�J߶Z<D�2��3�/�쬮���Ez�]��blU���!���xdF����O{�ȝ��Ik�ϝR�v�<��:':>���}��e�u��ւF;8�nm�P�M�v�߽��b�3���L>��)��I�Kj���B�o�s���ː��p*�2$���ɲ�?1$l��<X�;X�x3�&m�-��ޯq�,��/��,�-8.>:|O+�"�>�%9:5c^��X��c�p<��W��gp��J�������}��렓�<�W�2l΂�V��1�_Th���o��C�zɾ*ݕK{��i�R�	_����ln�65��V7Ü�vិa�����Ȏ�(���[�Q��,�Y/��W����Y7�]�<���,�ͽ[n�����6�b]sYG�w�r=K˹��|xQ��9�0or~����m�D�e/����-L
��ZD�Ǐ�<~ب������!j?����9Z���32�I\۬|s��^k6�E*�^q�$
�
m���5�i˴�FbW~��/�`�ֲ�
��~�R�B���(�!W���
�$߮�J���:�	�)hz,����n�vȺ=�}�'*(`��c]f3����B���ys���� ��80oN�[���B�}X �xA/�b�3O�-Y�7Y�,��:��\�|ۖ/K��׽w�����(�.c�g�S0�\m|���{��ϊ�^�Z�
.E������Y�w=$�`���#8��$�:��";��h���������q� �O�(�����B٠Tl�AhY�ý$"6���x�%�4�_Z(N�\��:�Zҩ��%��U�d=n!�e�E��������/W3�F����ѷBﶘ`s�z�����]d��u};d	&������y_��ۨb�0�[�d�it$����R�1s��)A���Ǵ2�F��F�Ead3���bj�2�-���=��\(�y�ɤ�P�ϥ�Pjn����=?(�t'f�¸s(��se���<�h_Y=bs�S�8� ��ѫ|�mp�C�:��=
��0N�&���\#8�!<�z ���r��+���ΡNo*�����5�ޛ�Y6�ߪ���!�z+��;��+'{� ��7L5IJ��]��'���QH�;�*mi�Qf惡,�%G��s$xɌFu�������A�ڀ�|�����OoD�ͮ�e1ی�ԥ_�\��~�P"�������H�z�!�7ծ��X�A����Rn?b��Nmvz|�q�o4<��G��2�H�7�y���gX�u��[+��<%L�ŹvuH?��WMTӂ|Qk����e�U5M)�~�<�ϒ�BHc��)`�����B�D�l]��@.���Q)1�u�lw#aI�vo��-n���R�+�{�J��4|�|l��$�<)3�uӚ��B�5��	c�j�� ��u�%�Q�]�zy��G��W�=_X�S��ե����Vd��.�iI)N���/%n˲"5��c�Ʈ��/M�-�_\|���A�V����A)~��.�7��Z5��IE���p뷷���۟�z6����a�TswP2�]����EpE�+�;�/�8;݀��e�ɦ���Ξ��������V��>���KRrǙ
r鹁GE�
G�[*�|;���2hAbc�d���*i��g�0�9\����iM�\���7bY*�J�¶av$_����N���_���C�ե >���D�ɱiQ�BS�i�#%L����^A������ᑐ!YC�>^���&]#�|g�X5c����#���F�<%^n\/6�er��y��ٷ!7CB� 3U�$\.��\Rpv�y��E�l�ؑ�цc�B��a�Al��-Ҭ6�F��r��iY�[14]o�m`jxK߆�ݑ �x�*_
65������O�Hwۉ�qތ�c�䭾m�+m�K�X�o��,69�"�L]�6��u���4����ˮ�KE�.h=W	���4��@<r�fL߀q���(��_�ġ���q��Q�2t�"����},΍�[�p���J�kD]�b�/F�i����`�)��
��@�r�x��֥	��[�h�O�C�E7Q���;5a�:����� g,+���W��N�8�`��x��^��-B�L�����r. �;����)M��ч�Io(�n(Ӊ��:�su�P��J@{��3� ���&<��n�Q���u$��[�.6����䨏@_�4������U?�}�l��
�$ժ��e�yXo6�'<8�%6+cr�X�o�vk֪�Q\)�u�ɐ�m�Q����c�Iy{�Iܛ6��+�Zݳ�	S䨎֎��3ow�13^<�2�oh�O���d~�\e|�[4���I$�Z�rI��lv�_~]�,�B�d;5�<�����|*o���'�d�!�" ��,��~nSy�]a��ϫg&�dU1�+�����JY��p����h��� />�~kL��a��P;=�@2,��޴�+S��(�o��,L�y9���u3Ε���Su�zI�d�j.��}��4�Q&6�m����,4zy��<y�*ł�q�W��\�X�� �,�
��w�բ���p�MdWI�ʬ�)��?B�md�����?��D�)��ۂ�ͷW�2�h�P�63�$u���ۨ0~+��.�����	�k&��D�#�@)r��Χm|^6���E�E҃Ly�-�T��'��i��G��Ȧ�� }$ r�e�����0u�����R܎��2�S�3[�L�3�eȩ%Ŏd瑗E�洟��:���im��ˤ9��6�'u��.i:���	1WuDMQ�wJ<R�#l�D��෢�i[�� ]Q��ռ��vɅE��bGuࡵ5,;7�/��A�H-/����w�H�wǪg�b�����N�!�
?�0��w��ݯnY'�&�"t��G��dG�{���ɥgWRM���C���P�$��9F�Bj��]͙�[���@���*�p��s��.�$���#b�_K�`3���:Kf �`����>`��6}.
6�c�c�!��Q��z�1�m�X�'4�?�g��������0�N�ߞ��_�:Kl�������?��qUU�b�D�z*{���с*[q�wo�B��/(�&�[���������W��B���P�'`"��~�9���kB�QL��:p斶7�V�s�q��}y�O�pj��{�o�QKS2)�� ��FjMKI�P�$�r���6�V�O�ko��_��֓�Y��A���+��0�ԥ\&�
���~s�Yb�#&ȿ/\����|���Ŗ
w��+R� ��²�G|���]
e6�,
<�F�d��Z�F��2��9��"�?�������4l.J�đ�\���g�|��֎
X�J8գ���^���"Up�x�W�Ri�4��]z��[@
���G߱N�=f����C Kn�<���g�O��/W �x�ۧy��k{�+����{DL���'�F����� ޷e]s]LA�.ȷ��&U�g�:X�����nrץ�����k�U�{����w�e΅���6��p��Zi�갗����z����^dG�0' d�5�H��0�gg��E����=��=�Y�=�)�RpU�;G]�ş�}לlt�)e�HP%��V���G4V��,c�0�X��ew����������0mh �d��4�/��0C��Q�<t�)�n��ʊS�(��|�����7��CDh8��nI6�r��>���ݺ H	�u�����U������:[��ӄ�w����TF�K��t���&�BuNMN������Jؒ�Bt0���ceM�멗d��]E	J�A#Ro?o7a�uO��~�6W05$�м��pu���ج�Fo>������6G�3p�߶�f�����\�t�㲲�+2�+�%�f����h{�b0W^���"��N�a�o�'�6��{��%yX(}�8q�AO��-�LP�:r�ʥ�2RA� "@ݿ��'�6H�a�����'x��~�������wo�����ͫ �؆LA4�6k�c t�'5`C+�ޕ�45�T�mWpw�@+��?ï�} �3|��% �GX�1S�(��a�Ni�ݗڂ�m,r�Ƶj�+UG��`6�	xYc~��JK�4��ڳq�S ���0P�2d�j��,�/���y��+(��"�wZcd��tzg�:^N���$��	�Ջ�W�����i5���{xx|"[��z#*a�����GP�!���ic�~���|�Oz=!�Q�bHu�a\�8�*C��h(�]�|	�泏%����Z����X�5-�ijء �|�\�J�,M�xj���+��(��0T�m���7T1��h���kX<=�2�ܵjj��/e��0��g��JX�5�L�͓��2G.]�46W)�Hr�rӑ}i�m+9`�5m� ����J3d~d�|�����HH���봛���%���u�]+�T֚��HRaz�*N�^; ���- ko%��ܞܑ�F�圣a>ڊͶ�s���i�� Ƕ�<���}����	�����^�m�c�B�`�٘ƚz;٪:���v~�
޿G��~��=���>}�
_���	0[m�����x���9�"�45���S�B��3�D��& ����Ûߜ��^�c�XvǄ��t2H�)m�� ��f�x�.4��m�Q�< t�I�%��*-�z�7�2�|k;�����W�0�W1-M����p��5���{��?�1�~�������?X%��V�M�����>�=L�BrR��P�?��!�c��0�\[��k	��Q3�{c`���P|���2Wez%�[c��%���a*�4G-�����p�>_�C�nA��U���~��\���z�BH��nm<jm�y����rq����v-�0�zqW�����܄�v�ԛ:��݃ހ0g�ȉΙ�U��H���f��P�ΐ�i���⣼�uL�j�3��
�$�A ��m�"ceʗ�!�g��y/���>�������E�����A�ZD�:��c��Z*qg�p����"��j���2�_C�z
@����w��������3� lI�%�����L&�G������Z@U���=|��~��7����_~�� ؗ�p�
�C�v
�pŀ��g������b�I�5h�nG�HZ�M���`/_]Y�]��7���I�N� }"��؉K5$���T�!76g���
2�w�g����9�A�G������o��w�6r4n��n;.M�P� ~���R}&abk��g�
��5{xM��T�@�84�3�N�1�/�՗�PkL�! �d��~�ҋ���O���-�?E����0�d=k�Ŕ�^.n�z��nO��IK�Y����UB+`{%q���NA�i;a�x��$��u#�i^�tфfKZf��q|�ν0L-8Q�yY�f@��k��w�..��u�,�&y�y�PY�cd��Z�6Y��{���N�w�7��Iow�3��-�<�lHo��2T�WA�S/
�y/��J!�n�i�w�4�ī8_;�3�� ��O��}���\���G��W�3�z��젙aS%���6�M�vw�ک���x
~z\�]׿��/�ga�> ���'_O� �P���� 0D�sh3_�Ԑ�0P��㨱�I�<���$�:!��Cv5Q��ӧtm1�kF+g c}^��R#{6�n�3��"åg��mn=�����-�V"+;t�����{��Ћ�3�c�ܳ��VTA�����/���~��̑M >�����������_���R2U`�y��	B��؆�m��A'������,�oĶXdtԾ��W�˰��;Cj�oj6ES@����g�aF���k�o_�����>�N�Ԯ�i�T7W�?ލ���9W�^�nH�.�[�������x��fM��@��g�F.rv|��0���9	��g ����g��:Q���Z�gA/��+�=N�I}�&��� �� ���T%����MG`�~J��$�N���|Ҿ���#�!'~㘱J;�3m䀉y��S�ʋ{e�T�|9�"��D�����8��d.���^�A<�SbO��h��݄f[h�I���_`���`������k����khॆJ%t�j'd�cB�ww�d���_����Ͽ�/�~�란�y�쬛-n�Ŏ��6םz v�~l��I�+ѥ.��@d̘���j��C��g-���d�ؕ��j��V\���x�`E�>�?���w�s�۬gi�tU��ά�(Km�� �>ch�p>���V�&߭�ݛ<�v�;&�����#�����;���#�^]�r>���ف��i��+K=�l��\�H���4lŹ��m�Ԡ:Ǜl�1LS¾j���s1��>�cJ~��W{f��֦c?��0Q&�o��J;:{�r�G?���aj9*(;SI'
`��ӂ2G5�@AB�[��bo�"kK�.zvK�����^�z�
�֊�Xw��6e���Xr��ڰ*j� M���hq�ݑ�{ɳ��RY��W�"FR�U�1���h��H��f &9S}>�/�V�ju�xb�7|Vm�\���_`�LV�Kj��ަ�a�����̞�AT��]V�r`���#�L�:�c�\���H�	&q��R�Ė"�ڊG��H�l��H8 `�������/�X�o��+��o_�:I�F�,b)S�Y��c�#�������ߓ�ן� ���	������S ^�+�=�
t��m�.�����X��D���<�m��[�]Θ�46@F���㢺�)5��X�\���4d�o��E�Ҍ{39B�#	��"V�������9j#-s2^��*����t �N�Q$zڙ����ވF�\�<���!��A&�ƥ��� �q���n {��kh^����Z-<>>+vs}��X��r�A��56 áB��B��?}L�ؽ��T�߱�/�.�/�ynpuh�䫦2<6L����x�� {>�T�a'����5v�$3Gjf�����͌��jС*9�r�n�y�OO�zz�q�~>���#�S"�`ǻ��4@���PF̗�^$�P��؊� S9]�� !KՅq��HO� ��_���b�SoX�Śb cu�/q}�2Xk��.��d`��SiÁ~v	�|�OBK�|��S��zJ����nL>�� .�۞�<6�dj%u�D�ET�X�y#.@� �A&u���\����<`�5����߃|����������ܼ��-��* ��vbd�>����+��/h��~}�>1V��n�x\Cka�h�v�3G���n����	^[F�Ml@ѣz��w� 0{�%`��`7����5�IZ7l��س̚�t�D���{�"0�%��$t���+����������]u� L�;���Ewd��-�X����&�p}uV��qu�_om{Az�6:��H�Ǟtl���P\z/.�*P�0��:�:��0E�t�4�T�C�ƀL�9��1-b�T 0\��C�MaO��R�k���N^�{�'���U���a@� 	��pF��#�⹴I�|O*�0O�Wz�G�y�!��ս\^+�G�m�ڶ�7�p�(�C�B?�D�`��7�����7���v��o�,P���mzB
U�9��Ԭx�$�U�L.����,��܍Pjk6vO�XAmdLټRf�W��>��� �X��7�]ew�Sw�oc'��a�\*����~[H���AS���U �O����Oo�b��_����B�n������	===��/_�ݻw���A������l�xL�w����{���^ςڱ�u��m�#�yc�G-� �Rxu[����L��۬M�:�X�L��O�8f�r5ab�,�y��T�7�,��QՈ3N�R8�mC��~�=�a�G��ղiY�& �:�@W�xT����r;6,Tǭt�x���ȉ&���� �qW�H�E��/�.��z2���u]e��(���NNg	T��s���/K�B��ae�q���[�G&0O�*��`KY��z_t�of�Ź��UY����N���ck����2�����³�6, �n�G
�c�-*Q:!!�������+<v�m���_P����/����C���F�h����x��	�@�r��e��0���R����3*T3NX�ι��>Ԇ+�G�LI��(��!���< =����Y�Sl�b9Z�w]�O�C+ZENQW��w���䈦��U &�����(��]�VӰ;�F�X���p��A�|�ќU�3D�k2���[��Y���
����N�Y�o���|V	�T��0��_�ޑ���޽�w�?�����5<mZ����̍.�v�Ac�+\OD�<a2��$��+���
@Y,��dc��et�cj�c��J�D��e�����'�7t�NK�2���ܣ~R����<��=$���'�7':�r�u�51O ��6_�������~���Y`^c5@�{��i`D�)А9M6\T�W<j���p}u	�9Of��h����]�G��Ȍ)�Ƶ]ێ"�,�ɱ$t��y����>�3SX���9M��ä��[��(��o
[�*þ6��8���	yPF@�/sm�m�EnY���X���!��ph���@U�
�ɹv��Y�W���fml�'����ϖ!�' ]�{�e��X0�����®..���/�~�W�^ӎʧ�kx���ٻO��~��c �;�d�AA������?sH�@��|���=���9�}�N�4?7ʂ9Yt3�5�����|7V����?���I��j����
�>�"�,X�M�Q�8g�sѸZ_bk�6�H+�Dc�*0��0��]��ĝ��E��7N�5J���6y���3r��L�f���;a����~2�����N���\�,L���YW�F�_|}����~��=|���l�6��й���ΠYp�BT�[<��� �����B���#��r"�h���^��3Kj8]-���9�̙gufd��DPf�X.5�L���_@�s�D�S:�E2�v�wF\y���OY���tf�4>F`��tw�z�磀�e[dĴ��6��m�z��<Y/u0�ŕ�.$�&.G�G֧�����OM��:���z�����|ɅH�t���v&y��QF_��t����
�R�b�'K�7g�J6����^��)��P���uf����e���V�Wj�g�NKK1Fy��v~�ͬ��se_�{'���6~F~��6����&bw�5��2>�*�ɖ�iD1��o��P{/A�����������-\��\`����.�r9���+x��K�1��� L_�˯�?������l�[H��;Q?z�
Nw�"K�<"�I��d{.�l��E����l��~�6I.ʁټ�cut.������̨������adGGNm1�w�8���F�H�&1zM�i�8���+X�e����5_b٩mo����%xtq�en�D�\�P�UB��f&�[3�6t����� �cZ\��KN��d"nFۮVth�/��' 6{�
���L~�M�8^����:XE�����������#�!2��!�3�r��;)�ƒ����M��$��pAX���L@ �=O�]��}'1�5�@��`&����f٢�#,��@G�m�N��h+ub�����'���v��)�u0H��H���,uu=:���f��'�AYC��I�TS��
w��*i�����V��@m�B�A�`(G�X�z��ŋ��۟���+x��Op{u	w_��fu�f����i,2��}�8���1��TW}�����a�t��D���P�c��8�@̔|=sjPQ�<$�}T�ә�;�R��sf'Vg�քM&y���<�+dAJ����@�
��������>l���{(��d�����a�ˌ�'9�6�;Y�6l\�~�B~�8���s9�ps�^��y���t6�jղCV������|Y@Ъ�4�-Q�Ҵ/�Z-:qA��2u���*%�g3��o/�͛����=��[��Œ}v�6�HH�䵀|;R�9̲p_N6V.��Qumʘ5ed��)y���>˽&�ԋ���v%'�Y���D�0>H$�]���O4z�����C��u�ۀp��o�>ëW/���k�q����yv�U��[p������}�_��q�a����4����V�9#R;��	ڌ��r$k<m/@�{����v��t�c�)�~MW�fJ�0S&%>��՝ ��k:r���KY���e �a�p���>C ��A�x���8�tm|��׸p�mف)n�%w�ĳ�wY�ķ}����.t
�����P'='[� ����<�6aJ��߆��`>f����� n�����EG/cg�#��y/^�^������-���/���]�h/�抽X8xw{�w���'o�o�8�<<�����a
/��\���U���((��� ���_i�FT�L
���{��Ta��)��1B�֩T~c��}�~,p�����!�o���i
�u��K��/I ;s��bY�����:�[��h�EU�]$��!g��{���_�1ݫ~MI�kYP��&Kd��/`�N~����1f�S��p��Yo��q��v��5j<����2���h�����/�~u��\��A �Eu��\<飑S��1H�U$)�L��4VA b�� ̉�O�@Σ䇪{eZ<�\p,��'�?�`� ƺX���-��ܶ4/c�H�E�H��;Ӧ^n��/E����8�]�HSD�	�v׵�&G��z�3���]��_{$�w���^�Iq�7�&�ȱ��y�<ɜ|}�ə���$�ض�?Fb��ǯ�:�?��Ǹ��r��]��z�>��ۻ�~!�C �m�l\��ݎ�y6�E��X��
�S��7�:JG&���&����r �!����јk�XR��u�	eS���K�Ʉb��<\U  Y� [4�x�
�l��:T������D0�\�zBԃ�u�{�i1k0a V#M�>Y�I �T�0Z�|4��1 �j[����|�YQ����w���w��ݖ��ʃ�RGm�x���p�}}{	��[���: �?�Ώ�2�&m7OD�?=��׊������h��g4��'���kW�J)�O��C_���a?��}L��`_~��W_�S�4�l�N��	%��|�G'��;�H�.�O��>�.�2����	%�5�~O�h,�Pf�C^�QO���pk(��[�t,���b�6:s?�L �B�VB���=Ђ�b1�:��<:<\,.��2�g?�&�pO��/�	�$�����UՋQ��>��	���N�%�Z.�)`څI5O�h���0'� ��n��x���\p`Fщh�n`qy�AA�fb�v�ލK �u�z�%�]��t!�6ί7���\i}�X�ZE�J��P���ű�8�<M'p
|�K�fԶۙ��:��L���w�wd����/�gl;w��@�RQ-���x�Z��'öWx`�����_�}�O_�~�^����h� A���4/�T�D��1�{m��st׊��\�gi7�U[��L I;��:���h��ڸ�!�L��ҁ#�sd������������3���
uxV?�y/_����a��`u� x6<2>Kl�5�����Vd�.�Z�t-�1n�UƌU�h\ �l؂��AXxe��n�d�>N �G_��r�]�3R�b�6���U��62��uQ�jǟ������������P0\u^�U#������ܡ��\CZ�wg�^����I�o �BVl�@LKϦZ#0��5�|f��Y�4�ʰ �LӷL�|�T*�1��tj�*���9�(��7�۫{��4�ֿ�.K��?=>;����T�/��������Ӱ�	�I���Ga((i�@tފ,�2��������K���?�]�r�2 �9���%�ݟ���������	Pi��y5̟;:~���Ͼ5��L�F�D�	|{6D�i'%�����&7�pu�$����>��~���Q<��W�p�^���z�;X�9�?��7���nv���Y@���	,����w�U��uZn���"`$g3[�<R��K����H]����fxϘN59ao^v�&���xɖ�KY�5� O�����&T�0�].���|�c�7��x���� OFv� �����g���1_O�zܸ ��3-������R+KQcD	٪12���8�L���}F+���?.����@.�a���z��F}@";�$�GF��:��;��o�Y�W���#�Ce_]\���u��� ��s0�w��{��03^������Hgk@ю#Q�F�2��A��E@��0��|=�Wd���"��0�..f���C�A�$j�xĘ� ���^�T��qG��޼�?�����?���Đ�\�<��R�s�"�=�d����:��l��/U��6u��>6�
q)бA����>�k��+Y�S��l\% ����7:,��`}�<<������I
��Sɧ����Y��]�i� �+v��H�U�5�02���!�fB�.���Im�F���m6t
.�_����[X���_��.�� �3�S�x������j)+��կ&*�S4�/��z�88& �������<<>����>Ѷ�,ȯ��]�c(�e�6�4�81�wE~)���\�����.�ZzN��n�����H[E0Բ��6m�SR�=hS�
S�U�	(,�Ue��X��F��������a�r�y ֛��&��}͡?�Ǉǀf� S����׻{���+|�|�:ʜ�촨&C7�с�̤��]`C8�$#�X�N�O�I\�d�q��OP��ںT�H��2`���i'����qsVE����0I�
�l�v���lp5���}k�����va����-o_��Y =O��+��_���� ����h�$��_���*L��7@���C|WαM����|��ϰy|�HX�����7W�����1 B�����<a��8T�nB��d��������-����5���-��`�ܙ��d���	p��8`m㔩��N\X��>���ݑxd�|�C�8x��5�"	��i���)·R���c�������=�ԡ���!雨;{�޷<��?���K��3#i���X����"��Jp`���_=��\�6G8o�B�A�=>�ӂn�\�0�Ϛ�(���~)�a��-��!�A����sSXX������+r����F�s��W�K@3�,�rE�m���t����ku.2Uw�+�Q�,�2��4��ٱ��/Bޗ2W��ڠc�5� /������F��Xź�9�e�f;�fF�\|a�vmz��x1����H�8������?�*��D���cS�m\�����(����:�|�r��P0��=��y'��nM�]h��_���}� �5�//��b�s�%�u��t�rGtٚ�p��}R������B�);�c�u�]���H��"`���A� ����FA�IC �_�ʓI�(D=�+`�h衠�g%O��Ϳ^���4'(�u��i6���������2��j 1�[�"���b�J�ˎ/R�e�x�`���~�F ˝�=��<|��߿�O��u~@���� �E�,npE�6�ìC��Z+T>&�#x^Z��ؾ��n�%����~��_�%�|qC�j6�Mz����࠶�� ���QuNh�-{�W�A+2�?�gq��c�/��/*(T Vw'�vZ�c*��
��a�	%��c�l8�J���ZZ���1vo(V��ڳ/oC�_q}���m�	=R~l\iR��H^��ް��<�u�vn'�8�t�����d�c:�cȤ9� �b>�bP&��}���#�?�m��S�!�J-_N��l��r0q棧��:\�e`"�U��]�l�ء�%���V��&('�~%0��D��,�tAm�*�����Jv�ِgR���1@NkA2��e�W�֋���3G��	?��u��b "S�z��nb�V7jt�|�u;���1Ǔ0�;�|0���;��܅rl����'��z	�7/Cԗٜ:���������h{j�d[d-�@�P��Y嵘�J:B9�e���(&{�6�t�����4����M�Ҏ{3���_!*m�2�Ýl{��:UD��i�/���'r��� �F��"ӄ �t��X��!�Y��� d�!���\]�,��&ܲ�Y-�J��2�1׺�4}FgZ��{k��+|�� �>�joon�A��-�7� 
�!�Mhǝx��ҩq��F�hЏ6_��o�s�����W����':�qN_�8�Q��r!������"vZ���Huƪꔭ 0�ܡ�:,��'	��|<� �o�u\���S���E��j�mھvO�䥼������g���!�|����t΀=�~ӿ��g�����`å����鳹�œC�����LHZ0��kޡ�����>j��Wt��a���	�6��4�����׌K`ٴ��;gsqW4�1EO��Κ�H�bp���<��x�{b`
	x�ؖ��pFm.v��������1dȄ�N~�,�޼�*_��h�[���iW!�Qv��T׵�'ؠ�x�BƇ��LT�,�
��g�����%Z�F�2��~X��J�'?�Mʧʤs`�.b{�9��m a;2�A;�Y�" �ZC�̺�{_>{�Y�y��4�������ghZs>�.d���vA@� t������U��1|�'�-2���s� $�]"Q���,� �)����F�=�ޥ#�e�b X�*�XB�J厐|��<5��]qL8�zh�<�ԙ��\���g[���2���j�ػ6:>e�#{cNe5+A��ȼ��f�s�D%����G{z|"@�~z�N�\\���&�h�9�/�r���i�U �k�SAn-�_�ۿ8A����������o���4!aGG ���V�;��a�bh��e� ̊ڳ-"N�zX.v�rR>9�8y���së>���pJF�0�Fij������PJ��>������	� kC�35t����'�o�}�a���\���Ǹv�v=�G�ߐx�?�7�w�BD[��}��4����4jg�ʤݎ�f���V+O���Y��$j��U��a��3$i�Z���i��j �-��9mO/s�Ϟ�B���;�̑�$U�)l���	�;�f���lݒ,@��*44��y�
�no�uR���DR��LvQ$��ܥn��Q�K2ݳLb�6t��n�W�m�������.D-�\�b\����ݱ:3aN�8�f�8�#Ɲx7�~DSEp(�&� C���9Ո��^����D��7�-�`�~�w�C���qhV�����|���O�C=���f���74�:�+z��5��'*`�0��SH����P�À�=�@@�`%�Hm�?�J�ƝԶz5FcIa-�A؈��9�E}6�b��v�T��y��"W #F�N@�'��w�.)�T�����?<_
�,>?[B�%����gfd��c��40餩��F�ual��^m ����F��#�� �%P4#���/ޱq����G��Q5go�<$�/ܘzFZK�] �!��?���?�@;D�{� о�/4RM+^>�۝����`TL��s���9����m8�;B�S;�j�(|����W>�Z�{zR�������:�>0P2e���٨�Pkf���)��@L` �K����♹�'�g���H�N�c�t�e- ��鹻��-��ɏ��9	˄���-ϩ���o�����Wbh^�xA �����V�tr�L�Z{:70��ZQ�4�e�X?g���+��\qF\���7*�}�cW<o�A�g'��5�Bp����(F?e�{����^��#\ݼ ^
M�Щ(ʭ�֓�H2����HKͰ�����?2]� �|m�@PPXX�o٭�������3s�0^|�޼�8y˰hB�@v�2HF@��+�~4�/:�4F��c����܇��>� �+�A.����"\r1`&tH�*V��6�ΆT���<���{�y4 [��G��Ƶ���+X����;�X�(?�0�xf��HC�Î�-�CNW���mjT^J8qN��A�o���*��U����%��]@C�w:�>�+��e���^(���⑳Rt� ł]l ������@�"�th��/<���#S�d_���exa^������gV5����S���.�l �v#X;����wG2-�ݱQc�ZT�zsB�J'E0�>q^�z�_�`���Mrӡ@�����K'Z=rʹt*=�Զ��$[/�gٸ�����Ah�F��ҥT�PQ��cs����>a���Xz�Ʈ��[_�䷏Q��c-�ӪBs5�T�s({�q��~�r�k#ة[K��� ��!T��bF��Ϳ��93w��\��sI�F��Q� L���Y��8���,�w�F�%v�#�BS��cr2�6�LP�5��h�L��B�t����j�(GAJX�!���Qn7�V��]Y����^�"��w\��5��5� �;�wS��bަR��L��ML�HZ2��$?Pݸ��kѠ٤�����'�4>���k.��FG��'��|���$�W������K��)0�sx�,��\.ft�&�Ɍ�gG����ē��x�^�]�}�(��kwkxz| =�n`� % �e� ��"h�(�B���p:��N�1>dZ� �8l�gu(�G
 �Z$�,��J:uT �l���ֈ��	` ��'|�L@�ex��3���x�h����*,�4��\B���1B��Ry愒�p��5�޼dZZ;h����;��QNO+x�h+:y�^<�{�+�AFq�#�ڛ���f��"�yyuV2[x�}���n`{�H�g7�t~Ն<�o��ky����VO3>f��� W��no �� �ʌ���bɫGd�f<��A>�z�����j ��#�<b�����>	�Q�ݜWR�"x��1Pn�ק۬�)�����s�LC��M��S幌f5�Ư��<$-�V���Θu�72�|���?y��ӣ�vm��״�zb��ls�6�K�-��3�:&� �d&�@2�&�����5싳{���z~Wf�MFtbO��m�n��61���}B�4"[�j��ޠ���E�T��Ǭm�l�������Ǟ�[��(Q�E�Er-��z���';/rZ�"u���-�>��stt>O^��"�Ş��b��>�;0�k@|~	TmS�K������6��a{>m��ѩ4-�#��&.(/3:#�%��i�}	��^#���7�Y�wɒ
��g�=�$G�l1s !SWU�Q;�w�����o��<��Y���%R���k�݁@�̬��;*3#���p�~��ZS�Y���T'H�M^��X�\�
�/c��)HZ��IEVGB�����������V+�ǂ��J��ťt�U+�E���*���*)���(�Q����̀�?Xic���0eq2� L�
}��e��~�:�y�4nd�[�,��i��M�D[.���K�v$�q�k��SLf�<uD��ʧ�~S��e($��US�^ � �
+�����<�f��Ю-׫Z�j^�b�gP¿b=J;�S�!\�8��nK�#�OsN��fS��i[��2��p��=�k�5]7��X�W�"��{�ݤ]��ZF�����v��ʐ��5����{���S�p�ܣ�l��O�~ߍw������������AӉ��r�:����۹��I2-F�įd���b#\�z�DƒP�\nN܇����\ww6���h�NX�-/��l#�ò�t��e�:�[[���ԓ�q�.��2&i��'��0�[�*��)�� H�Ǳ��ھ�dB�c�r�M�jIasL����}�O�Z��8T";�To����+�x!�?�Ѓ��������%�*v�N��ɹ�L���$QUvO�бLT��?�[+ �m�L�ܛ ��o+v��.Ƣ�z�ُ;U*X/܍\E�H`� ���F�߄��@�b��)�Li�q�%qE>���ֶ9����lF{O��g�0�\f�7ף�� �&��^��9eiP��� ��{�u��5��n����0�PH�l0~��j,^I��nW�q*��E���L�:�[�}Z��=�e�j�q�6R|���y\�3>�i"�uƀ9�����^�k��j_1M�������z�؍ 	"a����M���F�u���Mh��{p�8�R�fĮ�/|�)e6Z�J�oٌ8V�o߾��"ĂA����O��p˃��k	������Ug���6�f�l��-�3�f5���i}��m�k��w
��[?~�9n�_r;�`�}`�Ê���{�Ex;��� gn�3�?ĮH⯝9A���Ȣ۹��F)���hd�Z�j�ūe��z~�������d��D�*�/؝F[k8٨ό�c	�qZ���ה.�1Ko �v V����x�O�UaInI��?�Y^]h��߰Z;C��L����R�kG�.43GYu���ɑ��]ڈ��K�
u-�j�wN.>�ǟtM'%]̧tqyA7ח�~L�
�E���ؕ�G՚ׇȪ��j��sq��=@R���`��$��G��Lk��(U����aJ�1�"�'���ƵG���ܬJ��@��#�p�:�m!�l�Ѳ��.����f��l޴�ct��0f#�tgd��gʴ���5-)�S �)ł�K�UpR�U�Z��V��pP�=�� ����tK�``G:�k
�խd����a���.ŷ�l_��V�Tv}N0]�hv��~��MB�'�%&�?*x�`E�*���Y��I�V��{&G1x�\�u� �=�8ǔ�i>~�:�����\@1z$�H4 ���Y1+bX�γ�U� �L&����fo�?�D�\������ppy��oz�v(F��~�����0E9�9d�1=�/�e��������{/���>�簃ǎ{lK�Q�}��q���r�Ϲw�5𾁋CF��kv��.S�ƕZ8��� �BC#"�Ni�1��,
%fqD`�`,��/&\jm����Xl��m396�Z��17]��4c�|���?���/�i�X2:$OK����U1sN��RH�jT�lO�]����F{d?�j�/��,�fͱ�P���p ^���UC���`�/f\�U[�x��M� ���X���˜��^�L�+��W�d��	|�H�O"`	�Ir�VI+
g�
���p4����k?>��.�S�=�`	'Ъ����m�l���z�F�f=��h�~F��r��Cƴh"�ϚbJ�z�s3����׸zT����i-~)��c��+Ѳ�S;�5�����_]�����Z�2P�����.OiPe�`���֩��Z���\�i���5Z�N�f��܄֞�SU��d�Z�fD+�Z��C׉H`��!��.{ �˗��W{v�z.6+�O�f�Ť�f��b~yI#�SV�v#�z����0Р5����Sd��+���s6��l�Xt��ȏ?�,��l�Z}p�1j��.8�}�p>öļ��xV�	Lӡc� 襌M��q�c�u��%�=�����;�X��Tiʔ��1���Ϊ��pM9��Mm��#YJ>�WfXU>�� K[�V���g^B*0���%�F�"'�\T�	ΌQK���͇�Ļ򱪊AۨF�c�Z�[�u6�ַ��e�z}c��0�[�Yo�?����h'����+j<�C���}��9x���BR��mu�!uaRS������:�mp��� c����V����ӑ���9�{sM_}��� �fv;r�=d��`��Vr�`�q��e@�@v"6|��*�&�����

�(���ֹ_�|#�DŌf�����~��c�Q����6ٍ
'�E����.)U�3m6���"�o#� ^,�ߪ�&6�^�F�*��\p�:~r��F^r_�Ȫ0c�l���S�@OY2 qj[-� ��ͦ�L�M��n%8r���2y�ep6N(�b�g��Ht�2� @�Z�PP,�����Lz�"�Vq?����l�$;����6��y(]�\��u�Z�ӕ�	�6���[�{�9U�W�0�
G�+n���KV�Ǹ�}�|q��ZD۾kZ<�YA�|�{�6Y�x��EPZ�l����EA�}�c�>���Wj�ks;������6 r*�q�|����`��uN{���9�s�x}n��{��0�6�ӹ�����fG�7�����3��*��݊���~-�e�؟}���F�9
���ߎ�K�M�bܵ��gm��5�;#	�繨��h�K��l �ƃ���s�5DW7���ǖX�z�)�d��]�A��[�~��x�dio9g�!����b�3��jP�X�,V������|_f9�ݲ@%�޼^dI��S��-W�d*��݆��Z�j����ftw=�7���Ż7��W_���5�C�8e�y�vK�J���*�{��k5>͠F&�'_�t)ml��b��̞��K�P� �4��.m�#AU�1M�]zyLꈮ.oXt�`ƺ��OJ�e�X��_l���E���H�+�d���-+:8|�h(t�,[������T�Bi%w���@��Ɍ�-���!�<nV"�a���D�JuK�:=�a���#� P��w>}����Gz|\��Ӓ��XmiɊ��d* `>wͭ9�Ȝ��m�p�	E�8�	��qf�H��֤r�)��l"hlye�O�����Ґ�i�,M�=*6e�.>�(��<�4����� �;���[�	�����?�m�H��Լd�G]5�����|�DWml��R�7�i�l��Ui,Z� z��E|��=�7��ꞵ�Ky��q!�E����=�����^��!�Ω۹���}�C��A�>�Ծ���\7�P����T۩m�w�S����=���FF�MJ ����K:Fv�����]7羶��1�1k]���P�l;�0+6�i�>��MX�y����j�Y��~rAh�r6�2{_���a~z��~.�ͻ���4 ��?����)�cQ��+�(��M!3�mk��6�h�+Xhmo��Mﹳ�@�{^ߏez����8>�V�w� 	�y�њ�X&�w(�1�mR{ϒA�����<7J-ǖ٭��%JĚSM�� � ��E������￦o�zK7�s������+����'��K~Ul�����&����F���8z�,`�E����CÞ0/�����yѦ�	�ͱ�##�H5?K~!�m:��/��:�:`�}���M�f�@� �,W k�{9���7���W���-�0P��͆kj©�-��X�L	/�����6%��t�[����"UP1�(H܎� ��d��ެ�j�
�1:a�U �>]��' ��'�xO�?|���%=�6�\K���i)������ٿf-�����O1�s��ZӬ*��U�-�2)>CZ��\�i�S��R�i(H������!�kb�,59?��A]�&��+�e����^`A� ���c�=v38ŉ�(122/K6��3b��E!'Xh�>��3<��S4�������D���sc��mǾ�\�a��>���`�wI�S�S����צ�>A�N��apOi�K�}m��Rd���n���]@u$�ǐ������u���׽��8��	���,<��*��8]�9�E� Tўp��M�`K>R����U��Ĵ�G�(R]����>�lb����p�6�e�0E�,{[��	��t�ۃlVFL�Ү^�u�N��Fw��"��Y�ϗܔ��X����*8�qS53�`�Fx�'�����7o�_�} �<`�Y�Gu�F���m��q���S&L=0��Ţ}�U҉��B0x!�2��2��X�s٪���gOψ$ I��H�	膔���5���;?��&\��-�H�ߐ�g,� l���9�������t��+��oظ^\A|l%� �)_,*.x�:L�g��T�$�Wn�F]
S��
�-�G5�%���e�Q���8��;��I���"Po���Jٰ���'z���V��p� �Zs��(]!�q�T"d���7�;�q@X�@��PS��#�!�,S|����)���Y�櫗���c$0��X2&* �yI����uQ�e�(�3Ɖ���p휙�T	����ዣ�ꀩO�ד��� � ���������BW2�@�ִ^�8VL ��x�]�Pi"�嶴�����ݎ�! {h�c���ɿ�R���v�ع+�Z�@X�c�N�[����J�~z���9�t�����;@]�<t��6}�M܊�͍.N�9�4@�IK��c�?ǓQ�2�0aH�ȏ�g��8��#U�6"�	�a��<�_��� ����h	U�"�$�ޠ<P\�-vq��������"z�қ	L��=��ŽO�/?d���fF�� �L-��J�&Cu0`-�	��a@X+�_�������%���_ӿ��+��7_����dC�Ⱥ/�X{`f����c���D���r(&wTL��yc�e9�ܐ.�}�!���I�A	�S��x/Y�R/�dO]U��%��6�8�e�|I��WtU�9.m�7��B�؁C�J�Я�s�_4� ��� �ް�)��" ����I!���a �}�~)�#ʳ��Y�$	�7M��DҁtX��gV�K\b��=%@�KTwT;9��e0��y8����ꊞ+� ����>�| #��EP�$`����!]w[q�.��W9_�� �_ZZ�â=��SrR6�0W@WH�NO��=є}���S��.�<�ic&o��� (N\qm�f�zd=���]���t`�pz����6�lVK��&��'��_k;�.$.Md�h�ӕ�m��c�O���� ����?����@�����>wv�vl;�����7t�S��g3��̟�s���t����������ͭi�Z��*wa�>�����r:Y
�%�.cX���Eb�ew[�-A��8��>г�ϳ�?b�d t�no(��i��F~��2��������ݎ�49J�$�QÑ��Dߝ_�^�e@__����}����������^�h.hF&dB�$�R0մ6���IX�I�2�I� 0������y!��T5H�f�\�3Q�C<_��� 0�~���@��Y9.��q��πpz�����G�rDf�+�8V�-Îwo�bv
Z'o�n�6�=�̹X'j�U�¦|r	h� �xw���qh�d�I�!b��Si��b��#�6N�%yaT�6,���>�Ϧ���r/�EW"�ф�*�woD����#��|O�~�}��O��~A妥�vM�f�n֋�%�%�W���ƓBEj��6�c�',�����=g��xKl��U���;[���� JH�&}�����,9Ĥ+�V��14u֨P/�f>��I }�Ln�B)a��c&�1\�x�. ��>k�f!Z
x���@'��'nΝ��Z��x�kr�ˀ�z��m(����9��{�������ې���J�*�O������K��s��$�;d+L9���4F�̹fN}LzB2�8ˎ���F5#��*�b>cW��F��S���l��)�6�ǥ�*Ջ�vR�%̗%egRj�밆�mW����g%�!��f����Z��[�K��^��xůi6��S�U�Cu ����Ajb6��ջ;�_��ҿ��Kz{;��ޭ��\��{<-6����1�lZQҨɥ�6E2d��E @����C�1�]_]Ry=b�t�:gnI#X"��ox�gY&������3��Q�)N��_����X����..�\�D�'���|Y�U�L�������ߢ��x��M����*���R
"����Cٌ�2��&��4ө䕡L� �*S��UA!�X*��4Rr�և��Zp��tJ� ����L9BL�
��"�=���n���<Ng��������އ�ܬ��+��|5sb�L���kSs��i��P� ��o���ϧ�O��A$:�L�H;{*��V4�j�����y��9v�_}6I�/�UA�#���XZlW_�9��$�Q�}�̅6·)�0��BV��=Y��^d�
�~�v�X�U�s�ldg�a�,6��!е�{.�����)�:�.�4ܷ/�/G�ܲ/9������~�5�}G�m��}r�/�y�����q����T&#�3`d+O#�7��lW����^T�!`O���)���Y7*q!L}�IE�$��e�ot���L,�`�J�.0��/�����Ҽ,�{_:3Wg�oo)X�����q�j�����՚U�QZ�#��^b�|sK���������~��[��z�UoWr�R!��-=-7\E��u)8��R�&9�/�풸�Zޓ,X$�m.X[N>�%2��A�\h�;B2"����Ӛ�"Urrd����iW�)�ۯ�����B�;�<�0�"µ-�D�>�SCj����=}�t�.Y���$�d4�
Tf�,�ѷ�斱SLI�--���Ix�@ v9Z����n�3M��K�AA��00@-"&I~�9 ���S��������& ��~��[������?��_�*�,��b�����K�*�����7�Ǭ� ��+[�ѡ-[��{*�C�v�!��´���U���,�(H��I]H��]�y�r��B�}^�O��{�{@��!�:�J@%�cS^�\q�`� 8�%6y i��8�y�\@l���~����c��s_,סv���I�P�c}V�s��:�\�ٶ�_��$K��/�3r�&�='�C��i�/L~��>��i%�DN�X6����Ə+h�+i����eXk]?ظBB&RhI��E֊�0QV�R_.��5 ��bO/�Ol�>�k���c�i���l�|-N�">�ˋf� ��uXnB��B)T����������&�����0N T��f�O�K������Y 3��*Ka � )g�= �b�˅��E�Xh<�%���a/�o�<a���"��V����x�r��2�� � 2���rD���- �Mg,E1��8ِݎ�Q�ߤ	L� ��[ֽ� V��hd�l[a�t��g�ՂSQ9M�lp9-���u��bЩ>	��ڪ���.i�]��"�.�5)+-Je�(����_�	�����K�X/EY�hX]\]���Vd���K��M�=��_���`�9gn }A�EZY�%��}�F�8컃��|e>[�d#|��K *CB����[�L�ug;ġfq���E�@� �jG�4�΄n'�ཤ�f"�x��Nm}Ǔ �#0�N�v����@�/�1	�;���8�R��\wߩ�����{�����ږCl���x�_�����v�{ͭ����A7n�蕞[o�e��u2+�%w���<5x��2%����K1��*�g5��Ѧ���=�٨�L9���`>�*�;���R�������.��9��Po{��9�e3�ţ�����*��_��7\�51d�OU!�,���-�+.;�Z�\L��ww�����~�o��r�Ux��1�G�i�J!px� 2����;��~���J!�1R�/�-��:� �u b��Gzx�H[�v��<T5b,�NK,n�3�x�C��E�L�u�EP\B�;J!���ꊮ�oX|��+��B.�j���+ ���W�ʿ���(k��VDV�YB-7 Tl%�$G�:i� Ud�ӭgV���ւ���$Ķ@���#a0MHݜ@�b67䂃����Cm.d=>-�f��Pz>4� p~PPv	�X�u���P6b����w���0=�ƒ��ɇ#r�ǅ��M�)��@e���,8>PC�}�OFg�J�s���$3a�(�o�˟�N`���Y,�ܷ"R�����K�FA�V�d�.//%��de�����Y��o�A��:��_>������c��}n�����)�\���<w���fO�>w{^����!����K��%wc0�V{\ƨ����:Y�e�����ea(B���[\��ok�ހ��0sf�$`�H��ene~����!dň\��:2��� 7U4�{f���`i��>������o�웻�R�~���b�t�8�,|HZ$�HY%⚎[���^�xR��|��o�����kz�����[)D� ���j+�~���d��\n��L���R�$��� �f�0���Z.��ӧ�����݂sT�	�	�b�Jfl=3h`5���Iv|�=O�s!�� �[�3 ��~>�~.���S��2T���1�Tb¬D�Bs�)�77����A"`�V��P�\ nV��YY^:#G�Z�qPȀ�ZE (I)5�z�
`A4	Jo��q^^^�;4֚D�D�t� �F�������Y�S� �Y혗��+}��v��?��RTޝfp�����-ԫ�qp�s��GZw��`Z���;�������=`�傴"&�M{��a}�:�+{l�Ϭ�b�bv���Q���T��]A|�I���p����tDUuX�oLo�=����5��\{Ζ/�9��:f���̾��}.��2K�2V������jK����A�� �A�%ۆ��> �K��s�����un��rs
�J���w��i��3�9��(��ܔ��Ъ�)'��*�ss�1e��k�"ݵ2bxO܏RFH�W�qξK�|�̇EA�h5��u���+�&<�4�{ݱ��ba�1Oݏ#��)�C�._駋�u\T � 3���� t�����w|}C�7W��Xo$�,�[]�* �1��� �*6a�Y%*R�h��"B��{���J����|z
�\Q�kZo���A�9�J�z��iA�`�
�c��^HTO�R"i4�Ѯ��	�S�>b��o�"C�2tJ�鵬洢8#�&��m gk�b�<A�:f�8H�6�n�Rg��:�������J&$��3������M����/����n�$�ŞGcU�o"m����V��h���˙,xP����i���(..r���������������O����,Y5�mU�Ѩ��J�(�W��\|	�;���X��u�Cw��
R�E'��������y1�;����l l�
ؚFj�����M�.}��UⰒ,�N�r�Q��Ve��s��6��X��*s��kl���Ţ���s�������k<��wj[��c���������|�{s�����P[�+V�8�f柟z�c�kg,8G���b���{�*�ّ��_��+��$[��:��AtZX��x/x/
��!@��v���8;�D�gAp�1Ȑ�(U�B��X��I�p�R��|�1�_#�)�d��耴v\b�3u��t��2���ʤ�~���)x�oL�lkh|���k�'
iڲ�������o~����p�$Ak� 
׎ �7�,�0��
�9�R���z[�+0m�1��R���$�nn�]���zAO�t��gZ ��|R�������͵�lNJ��(܎SӚ��OB��4B����>q�:�,���j±����%�c
�RkpL�zq��(>�J-Hd".
�jFe����5���]Z�����4�L�/�m\,���O�dW7t{���~ ��-ko8-o$ߗ�5IS}y��L'�?<p ^�)��zF��3�V�u=w�ٔ~uq��˷��aE�7��B'ͤ��'�@�D��zS�0��߀����e}a;P~ߍ$2�{�m����l�TL��2Lt��N��X��Ƀ�x���eJ�������-b�W<���Wt]j]qv+�ˤj�/�n}�˶<��z�>�<��>�� ����Hǘ�}�;w;��&?���k��߇|����s��}����kǩ ��I�u>[�Ʃ.{�b�}Upϳ��0� �OZ0���,_ٞ*+$��f{"�8S�up|!N^���*@2�e�h����(w�U +,���'�
�=E�F����M�}�қ{p��B���|b�WDb< E�a#A�H>��qI7W3��z����zD�CD��`G���,G���#�Q�p U������-�Y�|`MQ蛎J܅;�a�%:]�c�UsJ���$����w�r�5����9U����D�SE�
���@��ns�[��?*4�V)� ���3�Lo"
��8�*6��)��9���r�%��֧:]�֜���1E^ 
b��[d �t�&��+�_^�ݛ/���;�!(�-��"k ��&�K|�By���;r�0���YJƬD�Yo?}�V�x[�|}I���z ���;z
����r��
�%��U �-9�����v�ي�>���+��Œ킯���I��]� �V�w������b�<��BT�#�f�s�[��ɩ�%�(u�h�5[V��@T��X�hk��e+;V6nT������1r��I�s��yJ��?��������۩,S���u��YNn�K�9�)�mϽ�;1|�}�l>|�q�ejl���[���9e�39�b8� y�Z�%��ؓ���0���[�O0�m���� 1�(��Gx��r��*l!���TlVa2��&s/l0��.v[��1��*+����������N�bެ��V�����h����)��eı���[�y74R�f0��Ք����zΙ�����>�#\�B�F�L�1tR���)It`��$ỲX~�-��j~qɉ��#-�?��6����wM�a�"�K��I�u�1�K�M��9�1	i�c�i�ߘd�Г���B�w}+sc�N�u??8�S�	c���m����}P�� @E^�ܪ~
-:]�`� o:e����]�!��& �9#c�t�t$O 
���U,�NA�=?�L� *���ʦ���
��BF�¯~ ���~�3}|��		x0���1pX�� �N�͈���6�<1i��q��}���CģdOS<f"�\�JϪ�E�_\!)��]���� /OY�>��	:��c0�YFeoPF�VzK�9Hui��^gK���z.Sp(��P�U�_;%p�%�ƾ�\��F�6�[w(��i��w����c�۷1N��Clԡ�=�����#���8� WJ=��o��3p������I^���RK�U?���d?|�B(�f��w.�8�Zm:.�Y��5E	�k߰�>/J�mA�΃lKҺ�2w�!N��Ӓ��=��$2>h�Q�q\$c��<d|Ca6��A���sj6�U{�׻��,��Dc�D���	G.���Մ�.u�j4�8����ӰsaR>�	 � ���K���*��N ��� jU ` jJh��DL��g^��~հ܂ -6�5�D����ʩ���?4Q�hX�:::�g ���'C��(�n>,����ʤ��;�{�����(��A��\h����18�i;l�ȯ��LAn��87+Z>=�C4�r�/+c�$e@ۯ C�������~���.U���rE�vÃ͕E|P[���@Vl��R��+��}���G����1e>朘�rr�e�ɡJ�8� ���5��H��wWѲۘo�n�RD�1"3h-�vg��ee�ʪ�{f(9H��	��ǡ��؟�Ix�v�Yzm�ol�?�M�ڮ��<�)��P|Y��}l_lX�=�'��������ܶ6Ӹj˾�cch����]���`�6y�x��|�����cfj[er9�=Y��_��`� ô�BU�������HbRQ���w�PdgA唐���	a+� lPу�#u�5�f Lc�+QH��1-m�(L�w�Գ�7 ڕ!�e�)�W���FI0�O����W�+���ÎZQL�C*��业ӗ_|A�޽�� �.�&�P"�D%���ֈ�����/�}���'�x(@�k���*��K��Z!�H��Zg��6�� � _�j�(:q�|޶�l��e���n^�Ǽ�U�
�P��.3f7Fw5�M�!Y�I�?nRE%l��y�u3�ځ�dp�[Г
g\߽�
�@�QG#�_�Fc����]���Q�L��Z;ę��w.I���P�HRi���C���,�w\�j��zLR�]���5+���Tf���VV�g��������@���f���eY@ݡ�v?ۺ�IЎߑ�h���^�(�7z[��rd�$f)#��xg+�6]��Z�d���/��hU�%``��t�z�O���^o��Ow"��{�����4����M���K1�7��!�U�=�7�����S��)۹�����l� ����s�|���>q٘�b����ڹ(�m�aA�����\,��(u�P��AP:ߊQ�B�\��8_j�q�Sԍ" 0A oR�۳e�X�z�`�M~����hl^�N�4���i��<�K6:sף~��\g9��u���<e8 ��3!$zgR��Z)D(�t-�{��/,��n ���NT
��{*ś���f8=�+ң���h;�+U�<����"ܴ1gn�J���������c�
��Jv�����u��K�^�e
���=T.z�"N����*�j԰^��z�7ś:p+9�xK�R�o[��K-X��S�#�9Eg�sN|�2�g���rǛ��� ��Y����t�m��#���;ԐQ���rFon.��bJ��X�l�jؕ	64�A����z��K?:p���f'O�>��E��G1l�(����� v�l"���Z얳�����o�I������.U`0���p�V?���z�F�)Nm�z\�IT��%�>��ǭ�$>c�� }�V*��d~��8�H��yNp��s��^�j��c�j���b��?1^�m�/�sE�6[u�e�����k���h���:�?����:���kZj�0�"�y����H�$U�����f�bk��8$��;j�������_�hb>�H��"F�6����y�5����g%�H<��5pc4r̨a.��z��}��3���n@���Y�Ri'	}�ό���߆�|�h�|Y_G������ahm�	��E�p�>h����@���Y<ýws}Gw7oh6-�{�X:����\�K�#[�ǒMva�5:�4���M�vJ�a *)��َ��ա]ۭ�;��m5欈��@�<r�Hka���^ܔO$���Z\9Keή��K�A�q�?ʆ��#�u�+��B�e~t��	/.��&�v: �]�e�4M]	 8��t�\dW�W����0�h��v1�Q\��� *'����a������zZ?�U�,j=�p�0�ژ������;}d̝m�X��@��F~�2D��e\~}����B��C�d�dKH�s�d�pb�wI�N_��S��*��)Q��&�]m��e,�9�{(��_ bؽm��ct_�����f�۷�O���v�����_�~�dߍ�8��<c{��(|.�8��9�.���qM��lh$;��N`�NQ�|���:���3��@X���z�����i��O�q�w���V�#�n��e�5���2��Z����@�.��]O&����q_n$��~������	�/�npYJmeԐ,�\XW��S�v�epڶ(T=U�Iϫ�&�K��s����{ �k=�G��)�o׭�ϵ�v���|ܒź�)�� �4M�*��˫�`+�lgS-�<V�4�^�1�%;���X�'M�Y�����gD���VX7��G�X"�P,*)X�~����!��cѽ{�>�w*ڳ��x�gh��x�J�`�,
;�bW4�80�ǁmcf�|Qt��l,D�-�i�M#���i������QX�6�uZ��Bv#���n�Y4q`�햼j�ᧀ�R�88C�`����]��0L�5+���]��P�(U�b�H��Lp8ɵ\������H@��;|�BXF,^�����R�q� i�z�U"�J�����Ma��^y���^�V*��V�\��$i�j��{I��y�P:��]_�}����a��}�9���\WU�h��9<�����{�qOu9m�2v� ̡}Ni�9m>��r��[��в��}����1�����n5MU�x����JkG�&�`l���wB����
xi�	g�O��مZb���k ��l` j��RVₜ��]^Л�;�kݮ��\sl-����Н�=��#/� R�xߕ]��������Y�Y�R�ܤPz��9��Ŏ"��k����l��90?zlz�Ѯ�
�z'ө��݇���.���VF
�1�0�ֱY�Ι�U�R�;��0��ݺ�T�?�]�$~�?N��:
A��+sDi7���S�~�"�����pE�� 2C����#.4��ū�2�Љ`�sE��&X�� �n U?}I�|I<S�~��B*fMj�w���z]9�՟��1��2"�GZ
<�B@x�{��l����{�u�:;�4�ע�ը��d��.��ǧD��	f+l�n�+��V�D�������B��ā�����uv=���k�O;C�+���ܦ���R�h���\�B7�1v��oC������ש�Ɩ�;���4 @=��覠$g�0׈���$����PYx��s��Q'��H�I �H`�+�=�^pɺ��=�ІY�`;F��O�@Թ(/��V��Φ�N����b�H]�%�l9�?@�Bt.߽����\z��Xwf7�"�,d,����g����<&b ρ8� �Ɠ1_������x��ocޥ�w�̈�w������`3�XQ���%*����_��|�����Oσ`�,�~��O��[wjݣR�-��2�I}�h/�?���ݑ#Շr��� 6G�����d�[�!gb�A�[��= `��7�MC~����ή8o���a%B�(��)H2���z�흾�A���XE��V��6�sv\|�H�R/�.I�ql�ڼMnp-J�"����x��2y�Ϯͥ�b����Y���X@��k�slqB�����/��p�� ��)�����������6����s:�s�Ͻ���<σ��m'5󒊩b�B�QÕOZ����J�3]�r4�UV�I�* ����gf4����]]^�����H�[�)�h	ܯ9 ��%��d(�����7�w����3�ˉ���|�QAg2�.�FDN1`9Y)vg��0A��� U�8ϳ��1�.7�̲�6,�!	u$�é�$�_������ W�t��xc#���)�vɞ83�>���-ԫN�4�ʁff��B��[j���20��b?$������3�T�gn`�xx�;喇��8���$0^|��Q}z�x�24�2�t�(RG��삛�����͘��py"�|�l_��&��{g�9�/���G��f�������R)��t�|^�ت���x�'��nO�kM ��O�q�}��u�cTzz,�����)�O+Ɉ���ǠƋ����x��KZp���06,��"]���"[���m�x�����/��~���ޯs�j�s��k�q������Z������v�L����`���f,�ُ�}�驵����	`>Na��he&2�h˼#]P��Tq��Dj�M/h�چ�0BVd ��A9���:|W[�S&%@W�_��^��F�#��$�H#y]�J�"q9��b<z���H��h���ͽ���f��E���a�P�qP��o�۫+�ԭ�P��ߘI��Pҋ聿}��<�=�1�d����vh6/8YhY�2�g�yJ	k9�������mOؾ���cf�	�vc���X-�2~E��Wi�4�FK'�e�N+�m�F��+���)6faV�U������q� $cK�H�lYm�+"+�ޏ����\XO��'��zud$lrr:H�9�wR.����x8�e;0�T+�h
V~F�&d�\���[>�D b<�{�l*e8Ux6�G7�� �[2^}���gn�����X�Nd����S���¶��[���n�#��v<��� ��Z�����{n�\��;�,�nyft2�V;�)��G�m�P��#�^Xv��^��?�8WI��W�ˎU�{QbWm�Ǽ֠�޶�9�Bm]b���
�Mf�
��/�ox��q�ڶ���f�M˓<*��P��r��]����-���β]�/ �T��|�Q��u-��5�j� YX�~�����R���P���t����2�+����V� �"'�kv(�$XL]�����;K��N٪A��s��I�Ä�*�F��]�wq�x�fH9WG7�qw�dG��}ꍠ����%�w�(`x4O5Y(N�:~�{�dS��f��LM�Ym(��~g�귽� �<9���w�Ee%�=T;K��-��ű�4:�飊�� �jK��3�w�{`�V���ɤ�+��s�0���,�{?P=�Z_�j8�-��q����3��9_�\ʄ�o���G����;o��ǟ+K1?�)�z�}���������ˮ��~�y˫�!p�2C�_p�y^Ӭ����e��@gYu�7��� �Ҏlq)��j#���z�\�eƠ�jIl���A_.�u@j�M��cMka�:��l���2_��B�UD[��^���R��&�{'�T��B&%���v��\��.�Dd?Zu�� �dDv�V�=�~��r �ww�;n��Iz���L�*�h'�r-^mx������d���i�QC#�j��v���k� AO ��-�5��R�@�8���7�~X��]g<�.;6N,A����Ԟ@]�v���`�',��y;G�[��_�#��?+ș^Z�a��B	��x<kgz��Ev}��(������$��li�Z��@�#TE,��o�8!����f��Y?�R��Y#�.j��I�ș��v�����w�.F�;�/9�?���d߱1Z}��X�W?��v����#m���f�����:�7��,���m�ǅ���ީ�<=�16�C�Ak`��X[Q�'���b4�9R�v�����Ym
�O��V�}]@��jj�#���Ge��`�P�c����>��LO$V6!85\��0���ނ9��}���v�9�4s�%x�=��n�W�ӹ�'��_���Ok/s�D�bRsN�0ְ��^���R�tj��֬P�Q=KN2� ��'�>R��gQԱ�^4�TO�� �񲚿�Z�=�'\G ���RL��l��y����x�f�#�_f̴I��_g�n�J���AK��S'�J�H6X�����wo�w�T�8A�tT#o��Y�w���#�jz�"J꼗�����:�+^Y��s҃��\/� �keV�K����i��$k7[�8�x�o)�Ѱ�N�,ź���wلg�O���|ـ=��܏�ktmCY��a}.�?�1P5��c��a�r0r*���Yw�]���'��������|�s���q�R&5���{�����'y�˂����ii1𵆾��6z]�Ҽ"�L�9�B��QV�Z$���|M���bTe2�';g�Þ�$un9��B����2.2����
�e��p�`�A�����W��-��B�(z23f�����vw���PH��T-㽅x$ٺ�K5i^�A�޼ |�!��J��k��d�b��{�E|�g"���}���S���	�2 #����0�l��V�_X��K�w��V�&}�����������M;"{	���l���4�d#d����i(2�R��yE�Y3.�=d���kZ��Z��i�a�6M~�	I5������n�dhW�+I�kg�)QAy٤���P=���\|�}|F1G�Z��gS�j���ِuTï�@����Q���
�bYʤS�o�OtI�D㓴E'�#g}~��w�.���>7������v^��ϴ����b ����i�T��aЗo���y?��S��<���EX8��P�و2�V���5x,���J%)��q�T��5�N��o4�L� q(��7<{J�\έ?׍&y5�$s9Y�"N�ch�q  �:!^S��Co���XǷ��>�(��^_�:�Ϻ�ơ�/	��<�/�^ R�R}E�m@�g��vP82���7��e 5�����cW�Dlt�ɉ���[����rm�S``�8�Od��ԷD�Bc�H�1�qq��OA%{�X��c�]��k�'�H	��'΢P19�i�+eD�J��P{���$������Z��ʧc��y||����M�d"�A��j���|��|�(5��d�߷	���Ӆ%6.vL�+�6�@JC9���}f&�d�1��l�{��I����V�\���&����i6L7��2�+6߹ǿ��Cf���`����mǘ���c�;�V���s ޹��sc�'��m=�1���y�u�� @俶,���m��q-k�~�������7�J�o7.+4A𼅮��F>�3�b:�>N��x�B �qc@p�kS���0ϗ
�����FIfټ�JԕT;�s�gAY�'�2N�7	�V��H�KQ��9خ�Zm�i�>8��>.�S���S����ĦD�4�T�q�V���F��#Y��E�����
Ϣ>f�@Y��
K�ˀy6�"��-6>�Lk�g♅ۈΥO�L@m��K]荴٫����)k��(���V�[#�]ОO�_�0�� J.m3�Ad*Ŏ�����`'����ϵ���9�ՙ�� !�2Ǚ+>}������)��:݉_���ץ�Ůp�Cc�޳���8p�����r8�;�5�%yZyR�|�~�ܕ��T�Xu�ժ�2![��ׇ��E�&g(qЪ�k��������r��^�aՉ��Ę��&�K��2�ū"0>���{(��m���9���9��v�}��s���s��9y��Ŀ����N��q��l��;��m)��9�,�H�y��fK㲊$A{�l^��oZ~5Z7Ҏ��hU"�j �6b-���[T;�kXl2Vg�% ��#J��Q�$4�^+\�E�
�Q�&G���o#��Xf�:�@���W���� ���1~EAb\�s�z� ��c��ΰ��d2f}5NrӲ�|g�m��*|�`�Z���H��E,��%�y���GHNȖ����ڮ�a���$�b�f$#�P;lX�^2>K���TF���1pm��U�pϊ3~7[�tvϠ�SD� L��7f��F �(j���0�i�:�e���W���(�R����l6�}�D Ƶ�J)�$?KN)j:�l��x��H+�Ԏ�@��~dM�A�.�@^$��o�j%��N���f������tĖӊ�s�B�-ǃ�B��dQ�x�+���������R����6>��U�q=���$CqĀ�{��~�i�_ӅxjLӡ6�}*st*������9[�o�@�������^t����?GtAv��o���������r*q��"���v<V�	�e�I���3c�6֨�d)L��
�%�
�� |J�R<��A,Z
eQ�/�>z|Y,���X�����D1�ʦ�Bm��Tʕ8�/��Kݙ��3��~z��l�F*G�S���	5�7�U U�A�	��i4���'�D{�x�(L^�TX��DϞS�hw�����3Vr��$Q
�_��\�X���gA;���:�f�T��Ci]\�,�H���9xu�g��|�x) c_iM&�������] bl���g@ح�8��*5�v��M���.|�v �N3�Д�!����h�|HC$.\�S}��Fc�Q|�`�&
���v��[��#S�V�E�~� .π$]�h҃��}[�v��c^>�����պJ��0�Y�4�1[M�@� ���ۍ�/�
��r���|9��m%�1�m;�����>��N3/������3�`�ª������|�9M�6t�>�3ǎq��R���㿄ɲ����ɝ��3�e����Y��l�b��F@@6qomEV�S\��|�PRդ4`��ރ��z���A�0$rN0jV�����b���R�{��p�p��Ȇ��Je2�[��߭	!e$�6G�>k�%x2&v��|ϳ{/S�G��&I�dg�vn��sfiL����[��:�$��dˏ��H�Kh�	��Aol<-��H�P����I,�Nt�P�_�#H�^�h�\�6�0��){���F+���\�����J ��ԃ�}u[ݪ�@I�R��7q��N1T��	~`����O)^���{Oo�k�d�C��1(��iqe58�9%�ϝv �1�h��/'��>�v�P7�&<���O���==<.�����C����Ͷ� �Lb7���F�d1L���,�M������C�Yr��h�Q���ky�QtV�w�v[wFf�YX��+������𪴂���v�Z`n�J@W'�RFMn��6 �$>b����S1���e��9�ٱx�}��s��^�{	�x~_���9�����=�vj�ع��\�y��Ǿ��*���>�NF�����b|4M�P�V9��<�
&))�,W)̘I�X�+��لc�d.l5VH�-<z��6
�m����,J����6&c�Qm�kK̡�6�f������)�5|3��UؤrDV>.��>�b6 �a@���+M�8���p��� f��R�B�3h�Z�;�(�1���@YM8��c�|���%>e���t�F�����.Y�]�& ��z�6�����L��b��ɥ�C�`�j����$֊�ָ3��.�	�Ui"0�T��2V�ݹ�����p-mX+��.�k-ٵ���_�����8K/����������������5�R��`� �n�&X ^���0}��D?���>�?p����� ::�����1�
H Vљd�WH-�	)� �)K#����#ˈ�VS�]�{�e �+�!��	:U��aB��-�k*bو��_��<�Q�t?4-cAS 0�D�C9�I_/�a	�"щ��:mܲ��w�qݕ���q)�]c��<������<7����1�t�r�c�>w�RdD\��sw٘�L�S��s�}@e_��q���9'����w���ڹ�"�ݵȾ��13џ�<�N|�L���d2a���2L(i1� dH�*	��nuOB������3e xb��Vps���#�[9�B� �9�e%��n���<�{��Я�yN��l4����1�r*�+���l�n��z>K���~���Bg���Je���;�e����iMKzZlh��C"�`L��H�xڲ^n�����޼���5�K[ �x�A|���|y�t�6�{�\�Z.�����
�P��ضɶ�����u\1�� ^4�ִ�/�+f�F�)���pb��E)@^�W7�~^e�{�U�A���7>�2�������jj4}=�����׌��d�ؠ��D\�����r�e�H������T���k[�
� ����ρ�������;~�?.i1BvF@���+�Ta�
4��O�)��%Er��tP�5��2�M�`_�]�~/o\�DPf���u~�ɨ��;��y+&+}\�գM���?�e7����k lV?�w�����j���i������>�(`]P>�Æ�%ũ�s@ܱv���}��%.�S�qh�CqR����`��9g�S�g�����5b���Yn6Ř&Jl||��5�<�>af�3�Y�5��&�v;�W�#/�B��#s7�}�vL^r|�֕dCL
dQ+�)s'z�v2?��k��z�.5Kי��C�J�_�Z�G:�'k|9��9)o�e��6^���x��N�MjMԣp�B
�����q�v������n���< ������,!�k�\S�Z2#&l4��j2�rPe9�E?g�}IJ�P %�-��,�Z.�xz�s�J!@YZl��|1�Ԇ�!$㦭ų�%qI�QC;��LB��r��`GnӋ���K�.���$�����0�A�*������J\��~ ,�%�z�}�[�x��X������V
�*��q�;I�� #��7���Y���3�af+�B�z�00?~z����?���'Z��b��p��:1a�Ϋ�FW����1�3��@���@��ƢJ,��B�@�nW�@TA-R�լN��+���<C�	�X֏��T�F��z[�>�Z8)3D��F�6��nD�|i�a,�����y*���Tt�1��#
����N[B���fz��U��L�ˍ��!W��W��k:��[?�?wݟ{�}��3z���9N�s��0l�w��������j�إ�ҹ8��Fe83;�z��i/~b�Y����7�����F�����L>��r�r5��5���O�ÂkLA��͙��#�� �Vr�5�h�U�FTq�z��+����l�(x z�RJ��w�]�CZ�}*�E$��g�����	{]���IE۶��~�@��9��k���^�5J4y���b㚼W�����~�[h��4�����[��~CE c|� �`��^Y�׫��D��iA������G���� ������=e�]r��$����߰�E%B�ƓMg,N&���ys��I�"h��m\>��1�ƹ d�+�ǆA�*µ�u���Qr�@*'+# �;��+��E��ͷ���=�)�a1�V�\A���6�vDg�
/2I��bE?����������T0J�|��͋o�0:��(1T.�Y�k^���iBh�@����
�Yf3Fr,������9{PlN�7]��l�cc��l}��]m갊؄~Z��͖&a_^���/�,~7"��l~A���'8���3��,��W��I2�-�;v�k ����t���h�@�A�w_�t��9%^��9�ېa����L�/�����\����k�7?߱�x�%;�k�/_��|N���o��z�����mf�lb3��w��ٲyP���༸�`�/>t���+��y�-�ԍ�R)	#Z	���I[6�Z<���u�5҅�S�' Q�U��}:64�y��>$�Pfi�`��8QQT9���kU�2�H��؍���������<\)nN'���Ъ�?>�ŏ������	��>���wCfc���;mVl?8���`WƓG*�	'Dpqt�7 +1�[y��-��rA�'~T��XI���#��V�����mܵQ7���UD��T���Q�?�j��8���c�2�>V"�92���T�%��
!���p� �*�|���N޴XO&EAI��(J2�_��9 ?���7���4+�z���*�
L�HC��Ѵ���X�7�+d;���@}��_o6�Ï����~��O��:�=��y8���h:�* \��Z�7>��肰��ڀ&�m��,a���A��k<u���E|��qD����ZpUH��{��|���$��H)ˮ��)�>U�j�׎�J"4m��9)��oo��v^�T%P x������^o8��c� eHg�u5�I(nʾ�
�2��g�t
��{-;���ϰ�3�/\��l}Û��싫z�;��/�s]�/��>���Z�?�NN��KغXG�}��m��Zc��VH\�%�(���a�0�#�
���]K�a>�|z��7�����:�_`b�� x���mkq��y� ѳ@d��@Y���x0��z�ȳcI�Ί f
�������?�W�������'��t6��7o����f��4+�>�p�~��˴,H�lM�#�J��_x�!o"�R^�e9M����S �?qg|��[��ODK�)�zdƉ��L���2	��s���O�.��b�(dP3�L���
|����]��`���p�Fe�+�r#�?F-bq=Zn_F9Pb 4ƍǊ@05���7Zt۲+Y�-�:D�����;�_\������B�>�r��')��P�Da���X/�툠{fo4��*�GfC{N�8Y�{���UA�x�ih2�`m)vu�0>Z�����u�"�O�q���̥)V��[}ߴ;W���|O���o��ex�B�Lt W�P�����B��dz���t�^�-�r�(j[���G���Q�������֧D6g� 0*��czy�6s���WjWtC8����V���?����.&oi>��>X)><-�C�L&-MWkc,�J*7��x���dT2)X��<cK-ƭ��,]{�Wgc�����r3�v�ס�~j0���O�������$p�
ǳ��㞚�q�۳}��} _[C9L���=����/gk��Dd����ґ2�-	�҂O��$�۳��-��� �����P�Q2�ZzX<��Â�l�)yD|֗��?�Y�F�]���.�@��[h�.|��"����w@��l��
 `d�3��@�7Wa^�oh��mYC�;�:r�Eg�����ј:h4���������������~�3�5�EWU�4�&b�݊�1�@�$��D���kM�Z��.1]k*��o�U��53^��� tT��8��A�*?�n�U��(��V?Ҩ�VCp��蘪���C�Z
�O�S3�*6�����d*��� ���W[8�: lb�k�`@��z�����%�:U�?�s���_5hH���^�������/����3���W��]X�2Н
��"e���'k�0�%(�	������'�����_к���'.��ڞ��t@��4��� 񹋓C$��$�h\"I���*����Р�g�T�H�lp�P��TC�ivD|hI�����$7e��V�򰑂TI<xZ����~�7W��o�
 �*<�+.|��cv�Ng4	�Tk�����1������2͂l#�O��:�K��C]��+���G��Y���6���9����g�������%��N}�yO?�fֶVe�����l�Ϧa��,�'�)+�ր�]\^��5��Z���.������~���O߆E)B4x�ںL9@�T�_#h� ˮ8����;\�GqR0=E���}�2���b���,Ev��sZ ¡5��4��(h�߭_Q�U�Y�')}�ڌ��"��M�h�P�����U�Y�
Ћ(����	�����>q���?�Ѧq�O�?�/��a��Hi�s;F,�& ��f3�13�Y\d$`��a��]���hr9��Vd�#����$�a1�V�P+���`^t�{��! a$�+�9���'%��c��d�Ւ�҉�����-�/%pͨ8C�<����l?�>���j��Z(%S�Z܏��3�*M_DA g����2���s�NC�Z=1H�Â̅I0��@��l.�X0Q�W��y��zI��2���������*J],���ϟ����/��o����J�����Z]���&��1H����Pۙ���;����D�Q�4N��ie4����M�+��iJ14n$j���5�V�5V2_�g���[]pz;���� -�*`�׷���yuy��$-�!����~�f3a/��(cҀｬ�t>ِ
���f�y��*�w�����V�qFɶ!cr(��`�_r�۶��\��%L�k�6sDi�;�=�b��m�2^���S���!��T&3?�_��<-B_��>��{+3`�`ꅖ!�I�a��J�9҇�uD ��5#LG�8,)D����+���~��O`�|�4D�G�L���`�� "�+� ���b �Ɉ*o��	���)H�`��jf��Ӱ���9}���!��NX.H�7R��p%�5M��b�� 
 �e������?��o?*�qG�Wc�� ��t)Sh�5G-��ɣ��6��@\�&�ƙ��ͫ�M���e�>qD����R�Nf���`u=�d�|P
b�G+6�T���ӂ���̈Mf��ˊ��U5����h=��gr�?��O�dI��E���EV!�ސ]��x�u�B��p�uX(h�A6A�`0�g����ۿ><�D9��`�onni�< �7
-����2;g/���Kԏa����A'�W[�������������< � ��)߃F�3
#jB2ͬ4�W&-�]Ҕ�3�忘�yNb�bH�&g	a`�{�Y �-��Ŕo4&�d��By�����+�Ѯw��z�6+�wc�%���0���?=<�߾������+��ݛD�@.+���2�����j�n[h��,�ZG�	�	P�2��0�����?	��Wާ���nt:�Q6V�����l٣q`��c�܀���|��0�s6|0��8��m�oy��*�j�X-�	O�a��   �[��V<��6	�V\z�4O���~��G�k������62̏���,�*t�v�
 �<��2���
%V���n�8���)b��ZMY�\�xUG����c� ���1S�J��$Y�pEJ7f�mf+�̛��GR��)	��*#Ē=F��EC_<�����HO�`��\������Y&��qV�QSG.��+ψ��H$���l�|6ѱ��=jT߭�$1J׉6��8a����A��m|���b����ȅ�Ո��e��`&������z|X�����[�����ے��� ^쬗\{b��u�tppl�j%�v:gq;�D!D��*l��4�z���[		S��̘&&�+�k������R�ɂ���<N�jY�΋����ZD�P�ܷt9��V`"3�����?����o��g���?і 5�L�YhӔ\ c�A6�/�}��M�plY�m�@-��|�Υ;M+����*��0p\C�fK�po���|��..��b���(��u�WH����:Pb��J�e͋Q�om�bR$�<q�8*K�X�7�ӇO���}n�u Ȑ�@� �zj���&��yL�;�x�G���&�?��W?�/����+ oǹqR[���='K�5�O��u���2���!��s�H�&�>{��1V���>�X�ک[?��u�"�o�~;�s�=RiݜǰL>�N�����`�R��m}�m����s�v�۷��J�-�#����cX��@����C0�53+пRr(..��Eg��ޖ��Δ�ߟ���6��1e�C�R�U�[Q�"Y��q _�f\\��ް�(&{e=�Sİz�{��c���삩��9���]�f1�='+H�G���ǅ����0dl�����1Zz�uBťɽ�����7����x@�s9��q�i�wƢ��0n@Q�,
�<s���M�1��@��i}"���S�Vq���������@쁕S�~�7�ZpY��ꉙ0߳���xB��A� �`5�����_k�C�ՒC�у9Ǫ��Jk+"�	�����B�.�8�t�>��O�Qj�Y0�H�`�(��1�쒌�.��Fg P|�D�ނ������?��ǟ����Ӧ	�, �`U�w~M��%�Q�87�צ�r<6��I"����tG�$����R|�㰒������MJ�7��==Ї�~��Ygd�o��;z{wMח4��i�AJL �nж���eZ=��N{��*U�~�T��W���Ϣ�U��3uMAa��?�g�������K�gPA~B���_`5+�썞f��Ҋ�v3�D��Qy���low���\<Pn`e�6\�c��i��j������sݠ�f�忿������^O���~��${��7� �(���A��ֹ:[�-v-�p�f@��vMU4�Ŵ=��l�FP3/�!؉����)�-�k��x���o|}@�
�/N{��j��G���h���.8����1�� p/��h�*��ǧG�� �L���'��q,x������͕�Ѱ/�8ć�8Ūz���)��R�,#�".W`�&�8�,9�ކFl�k�=��J��ҟ��sh���xO�|uK��/��-H�vZ,���(�0�Z�9cm�Gޱ��BU��!Q2�9�J��e��
���o��'�ش�1�edc�R��n�O�j��Aűz ��̨�gg-���&�6W��-�~`���o8Pl�:N|��Y�/�nG�^�ڬV�=NT��
�'�� 1��P���ZW��B��	_.W�X8��H�	3�s[�t(�PPJ7P�9�Z;�]����} [?����3 /�_���1�ꑀ/���~O�`�B���¸���Ȉ�ne��O�r�6Ź"e8�n��(���j�+��̀!�t��D�22]�pƨO�
سZ��{/�o{Or�)vC�����D �$n���k������wё9��IF仪��VK���,�X�������bqgF#����̈ ��cf���`䫪5�������;�������	������ll��G��ͱ�9�,�qd�c���q#���%GT�l���z\�'�{!Hx��\�_�<�����i~ɨ��x��{i[^e�#�v�s��U@Z`JV}W�27�09�D%W���^���辡�����ǸgUi�AܴR$/(�-�??L��3H������������������y7�����˯�X�HP23܇�#�� Vh;�0}*�T���q����4�,Ҧ��'����П	 ����@W�+�
2�u�� ;�X飢,Q����o=hm_��Hk3�%���$����� `RO@��Q!獘�>�ğ��#���n�&�\lk�#�^ Pۭ��~�s�b�h.���M_,��(����՛ΡʁX�cF)`*`VFTǆ�IW.��gl䀠?{��sI�]R�2=߃D��Z/�RX	>����+v�%=C�l�{�ZAY�/�C:s�.�6���5�ч��P|YR��F����� +����$�N���h�xE:\�KQ'���I�ҍV�b���VX0<,������ǟҿ�۟ӟ���	�}�4��i�t��k�>�a�� �eڞ_��������Zf�|��^`k),�⃚�͸�%�f��ۭ<[��.��u\ηHP{��yw��ޜk���C�z�F2 #��� q`&9YhB�& ��\�/�G_ �?��Q��������������L���?�߿�1�����#�}�p� ��Е�tr�S,7�V�-l����-X��?�:�`�ͨ<��K!�\G����/uh��_i�����^���D?t�<l9�I�R2sL�L�3���k`��od�! >+7�@n�O���y .WW���b�SkI�܉d������|}���Ⱦ�X�,ǃZF�$R
/�O�-��-�M}�X<�Qʈr�䆼Եʼ�G�.�/���p�M��ݷߦ�+��ms~&�"}�gi�U��!s�#gJ�d��+X�'�,QY0��H�RsZ�}�HA�_�}�SVdχ�}:�J�noӷo����ޤ￹I�N�n;������3u��,�bu�т��F���|�� C����@�@(�e&Y
%��0g&�_ʨ�+�	(LG��=T�5"�~�壀LV�т�����A�.b����h
�����������EY/�(="����=�vf{%'���`�4.�ՙ�ф�B�):ѐ*Q����,8��k��n��.=L@��`{��_�. �?&��׿H��Ņ$qH�Ś�Q��;���+i��%�:4G�6o(�d�7Nײ��桟)���*K
mĬ�Γ�x^L��:R����P�.6�B#M�M��y��K��L�*u���v�ӡ�qP�՞}�p+���0n��������b�$��#eE��)m������������<��n,�|d�4�\M��/�S �k��_��@�f��\ﵦ�g��G:u�5�)K����̬����ёO�����5|���3���?{Q`�*[�H�ִ7J�����
B�$C6�ͦۨ������58S���Ǐ �u�:�0����*��f�-�XURx��W��k+�ldwmD�eI 
y��A���T�w���� 
�D�Or�+�WRJ$AnOq��o|@�1k$+�\�Q�қ���?���e�v��<���^�/{�Y"�"?!m%�R#�RC�.���.���>��E�~�͕ ��{7�.�hQu�#|ҥ��E�nPQ7
�N)xge0�w���P	& 3�#��hd�Y�h�,�� ?�9��� ����F�\��~��=j�����+���h����s����(��f#]�=u6Mҡ=��k��^63q�G�B��!��a`eYR�$x�X����M6d;M1��FB:�/��K,�I?M��_~I��?�����&����������	,���{��9�]�E�Zd�=��{D�=�ձP�3��(>o�w��TX��pZ9-[4Ŵ	8$�_�e[,�pm��3�4�F����F���X�$�WH������q���m��m���%�������	`e"�Z���F ��6�������#}��1��_�2-���ݛkIЋ� �m�iD\����/cY���W��
f/j��l��� a|�k�ݾ�_�c��K��2"_z��>�Sf��ޫ��_�o����8o�s�)���󩶜j�S��x�c�ґ~�;�M�d]����~��,���"�Ĭ��� �{�}���ӵ% 2�LPww�\@�`�ˁ�=�"����wA_���*-c.[է�Q�#���*��槛Ij�,'4�Z`��v�r���Z״����*�gڣ��6rm�D��/���@6�k�͐m}V�|�%i�f��e L�6Y�V;Q��ʺU8�DjV�l{;r�~����8��M#4}�A�������"��&]�)RA%��@��������"�6�LR����1�*,�%����ɣ7u(�N��c�<l��o-%H&si.:��W�[��0*tfj�����4�?"���R`�~���t�M:?Т��
n����9��kj�[�;�h X�����j�,i��﹘Fsr�(7�G���X/�M�^?V ��L���&���BѦ�@~��IY��C�&���v�b�)��8]<�Ge�N�V�w�HܧN�+;�T7�.�_^���M�LaRIN�N�c�gm7-�>cB��26������0�Р6r�7Xoa8��̐m��5H�"�sfT�~A�������n���ד�vZ@��k���	�|���Mp�1�	�n��G�)�����Uad[g�)����A�3���zn��]#����6z��=��+T��w�>/���W�Q*{Gm,�t7�����/ϣ�$�S�V�� [|Ǚ����x�����{�����0S �;.�S�������g}�ً�_����+r��Mq׵=[E��	w�4��n�#o�7	�۰�<L���PdŠ��}O䓕��Z��a.̓1A��^��<�0�49Rq����v F��'Žt (�d+.�$� *�?���H6��t8��� K�� ``�z�|q��:F�-֟��-�,mzș%{�痠	~�(�=z�H��l��r3��swwc��<$����F�WJ��]aޱ��v�q���2"ٲ,��%��/�F�a"�f6�XC�1 &��d1��V��X�Zq���w��6���N�W �-ঌ�H�\F��R��p�i��R���z�i����WI�����T� ���P�آ`���6�σ%�'�[� ���v��dqj��Y{{��Bvv�]{��e2!�c7����Ն���"e䫚��a�	1i�����is������NQ�g�!��u��J6mK����,]��V��y��|;m(�oR{q��|�>?@��s�f3��2: $Q\��)D�d��%��lL�Q��h�i4�H�ŉ�%��5�A�אԞ�HG��S��4�[ltS���\��o��5"�l�h'5��:H��xM���3��5L\�_pD!�:%�����O��CO�m��~�����a䏰E��-�ss��`O�0n�|��̳s�;���������ζ/ۧe�����̞W:/�����V���z�Q/;�:�_V`Uϝ�M�A۷��󌩣b����8��Y[Ȭi���<O�����-�{]��z��;��J�:˓�)Sz1i�̈�5ȇ��!rp�f��`"�L�=p��� dP&�@��c�����}��Y�
C��WB�T��X�!L��p/���$�����������K����������AX⯾_��6�"A�^��8�lW�����rfgN���  W�NQ�o�܀Z�]F����>k��o�싶hZ2�q��y���η�������	���}5����<��{��)�@K<�:�3����\R2M������$׺�Kͪ0ͽ���N.�̭�T���P������٭��0 ���4�B��߉��@z�a�2���p�YhViEc-��,.qm��C����zq��E�,���E���C��cRn�z&�Ҥ�H���d�WN�o�P5��mz=���09|�K�L���w@��d��"�_�j��6�3����,=L ��n/Z��@�R�c�0�X�p�(C,��n/Z([�P�i4Y�>e�$��b�$w��Z�S�����L��0�O�����tq���k���o���K FӚ�Ј���{�~_Γ/9�O������瀔�E��bb���@繾@��z��sL���9�$(Ku�U�&��ٵ���e�*Y�\l�
\k��:ٶ���׋��o-�sЕN���#\�*�֝�{��elʀEѸr9��E���5��I�0��47*j�$�j�����C��a:H?4�\��nϲg3���A��/���n�A&ɼMX�P������-95��$���D�_O
�"��l������^�NL�Ţ�P��`���CR�4k���?���l���í1 �r?Z��Ӷ@ƛ��������s��9�k�lh��G]��pyd�}+J��,Sa9��� -;S���w!H�6����m��{���Fj��$P�媻���L0V?h�:�,�O�s�NR$��]�kzF��~k��H`D�b�:�:Y8��zkI����*h�4��!��@�R'!�luВ�7��7Һ�X<���AɨJp�&ǩS���N3�Z�)w/l�(K�8��K�Y���.��:p����|kEQ��PIM皽����;�ϦQg���w���j�מk��+$|�h��K1Ck_@��Tc�h��9ZԎӸIY��"s���$Pv�xzV$�E�����o��ƒ 6U���7��!���&��1j첰d)��裔
� �?�x����k�D���}�k��c ��c\�}�v��8��x
T�j�\yH&\_v������#+�+p�:4q=�(���ET|*C]���,��<`���$�H�$��(�I�9����i���~���ij��je?�yL��� �<Yt�O����H�F�p�R�*�j��Ո��xy�Mk`&�ps}�~������r�;Ϳ��H����������V#�!�pE�@ߒu���̾_�Uf?	H�XA���s�n�X���%�M|Mr
�F����e�ehZ0S�/N����9qD{B`C��@om:�Mzm�o�yUe}�-XcQ��~�=�RQ���}*51K�j���A� 8$�H��#��DJX l�{t����\Ce���k0�e�N^Y'"[o�WC���tm+���k(��>g���:MV�kT��ʳ�s��n��
��, l#��G�^�:��l����h�Oh~a��	��a��19����Q����V�P���^��H�|#�]K�ר�K6P�{j#V��6�b}<r�1~ �`�_*nZ�ӈ�a����"Cy�w߼Kח��S�����ue|�V;q�<��4<#��kг���3��Թp_�u��R���6�}u��;��6�	�������x��9�?�٩�>�{l�w1���W�o����-��pzZ���]EL܇"CD6%-ޏ�Yzϝdr�ިם}c�o�ع	��qٿ��<>�%���R6���S����*���;}��u�wװ�(0g��}�2$�<��<)���J�~Φ�_Y���P +���F}VͣeQ���o���)W�g^%�z`�n�һ�7��|+���r7�]��t��AL�c!�WSv�R;N�%��9��Sl�{�ᘬ�
@vV�imoG����(&G2VM�	����9��lu�Qs�ֹRjf|՗�w�%f`L�Becg���߼�HK1 ZN���K�k�
 H��"�Z!�D��|��n(��KHh��pқ�.���3�/��9LSp��T�^p�Z�z0�V�A�ٮ8�ոc�	�V�`�,{�l��Ż-n82Q�Zs��6x4�40�K4��ZAh˂��hLحECh����9���i������X[RL�P��ԋ������fP`��/�P�SM�vє*����X��QC�(�"
�8lD�\ ����z�o��ćŪӮ5_-y����6����|{}�~��w�_��O�|ۥ�����l�<6��q�Lc�(�_H��B��`��ƚq�ױ��5GI��=y�i���آEޮ:Bd��ms��g����zKi٩�{�������ض%(�m�kPC!5�k������/Q�}�D��-Oϫ��RP�{���XQ���8�q�V|_����S�s�~�:��NG���AY���6A�pפ��w�)�~��R�\$���=�ut�W�6G�d�β��f,�@�.5�k ؐT�R[dc�PR����tuy&���d���Gw.9:w5���(�k�?�*)	\F0hp=+($����ͩ2`t\�l7�� @�"g���l�d�߫�E�5)�9���<���9[���6�"{:G��;^O�P�$��wZ�����&��v�@�m3������ܙ�p~d��qO_��k7���U�G�}�����i0{�>(��.�#��;�+[�,���Y�շ��К��ug(&S��&����^��H�&�-��H'�47jq���E��¨�0���� �,���  ��IDAT�+ l9��u�m�6T���j�.9'b ���i�İ����l��
��(6��(S��F �+Z���j^���j�YX��KO2h���N�����?�A��}�MU;\�N����mZ�M[���/_�3�Jm��k����y��W���ߝ��4����̑�iֆٙ+߯@�X?|>�/TO�/��ǋ�^������G�Y{^*'��ڮ%ċ�g�� eks��?�s�gf)���x�f��U���`�t�i��a{M��K�vZ���C��y#�.~��n'� {���$�iU�.	��2�ŠZ)u���*U(O�{�������&ݼ�Io�\M{�:�jh
��)
��/jZ�7�35_Jr�p��#�+���-/'�{�M��-��ю	`���<{.�!��"��ݻ�n��x�7Ռyv_��2f+�?����{���!0Z]I?���.�X�d���qkV��C4 �=��wC��v��J��o$g���;��A3��$��~m�E��ma3ר`���
фp���iҲQ�8�M��e��PЦ��_ \(O�v��JAY��.D��ˇ(��$[5��[��-^��O��*���Jwz�1]X�ЛϜjU���q��Lہ ��`//D��^O�$Y_cQ�E#	�Fz����U�o��(�"�I��i������;o�麾�No޼Ѹ��F͈��Z�F�k��b�cݔ~=�5׻R�������&f�!�7��@�uN}>��� ]2�W���6��x |h���'�k1�����ؿ��k�Z*Q�m������\z�PڹM�8�/6�L�O/)�����1�j��|����ZJ��)q��*|��$��1�i�	�6�f}���8Hj&i�
vU��:@��v���ۛ���	|�sT��O��k�������0B9���4��ӝi��X�I ��尒�d��9��F,R�w��� �{ �C��6�0�0κ.B�4��q����CRB�R�u,�j+?Qc��U&�`���@;��k�
����d�������vW��V,����I�B�'�P�J�IȢ��4�ʕ�XsĪfP$XV�Yt �j�L��ꘋ��!�!��s^X����2|0����EcW[�Sg�)ir2Y#7`iF���G^-Y�ls�=��9�=�d3�����&^�Dw�1�k����O.a���%�H-*�i_��%���<�hm,��S�Wf�����7OB���Q 5D��ϵ�UQ�L��rgW������c�CJ)�n��tR���
2��%���P��~${od)u��ɭc����S�����%��k1O�uXwp�l�-�wy��h�kV���}�;��x��>������y�����3~���|}=�.\Í�,y���TA߮���S��1[T"��#�!"{+J%�jJ�����RaMn�`~(m��dc��4u��/�ȍ��̍L���R{-N�Y�f)	DY�
"H�p>}��j?} L�F���J��׬�i��9c�0�t�2f����kʣ}�
�t5�d�T����lXr���*K�rbT�xt��Ρ���y
�[�1{�i�s�g�F����.���k$ˣ�2p��3I�ىp"�&@��q#Y�7 ^e���:��ޫY�ojd	��o�nL),�,�b��%�H��}�(��_0O�԰�J"Oc��]��XؖB��͚���0s_�ޑt�t�[j��9��M��(�cẼ��3���L�+�ٰd�W�Ш�R��fpֵ�%�R|%�ғE$�T�S}�+��@I[�x�$ l���h^����r��M����N����e(f�ծ��0����s�r|�αЍd0K�k�(��o?���_�P?W�;��6F'��K̡QX�k�o��y�A��_�{y<�_��a�V�'�']��$�W���x߬�Q}Κz�if�4_�=�:��J9�W,�*���SsZZpU��n�2����C��E����X�=�#ɍ
�����L�b�QY$�G�6K2뛛�tu})�ر6mDV��v��w��<�����.��	��fjwVI/����k�~�C��j�3��?����|A�0'��V�v���L�I�Լ�y�O5�ɏ��\��3.`"�	y���,'�Ͳ���2��{e��/5��x��7:��񹾄P)L[4�Оre�ʤ�4�e+�TJi�#�V#�S�IǏ�L��Z�5��?�S$���rvG}"l�_�1憝VBg�H��Ո#c��܁{.��qt/k��L�,Xm�����Ĉ�"9�a����W)�q�G�,��ڦb���15�0���?|e&�k�!ĵ�붖�+���s>צ\��g���5ZNb�(j��̓���qt�D7�i���\c0��������_�f��#y,`���:,K�Y�@*��-�C���n̏	���9�'��:u���]�����U^��ꫯ����S ���LD��t޴�%�%�Z~����$(��Y�~��ۏ����s�Zm�t��)�cؓzOZ]�m���
.��ۺ�H|�U��O `s?Q����Wvs�Y�چ2����n'��V�R�>�.�)��=W3 tR8�3
���iZ�d�R͝ŀ��r 6�� � ��:͇����R �sX�7�-�i�G E�Y��%����+�k�j�Ɉ~r��5�*y�w�� a�fSJ�K�\T+fb�d�w]������5��]L��[��ɷ�A�\��\(0!��A���ҍiLl�0�	�G�tY	3Y����'����& �\�4@dEY����f�9[1v`���"IF#�Tg��=j>�qo�ǳ;��Q�zq�B�k�3F��T\&�Y���lnP
XR���6b��p���i�J}�z_���
"��*��`�f{Lt1��Oî���1�H?m\ R��N�M� ���I_c����z�}-�}�x&��g_L����O\䏙�^c�z�=��Gʿ���l�ژ|MS�Sר���R�����S��OW�O�)�3/���L[�$�:�2߇~�K�>j���������t�p/����Ӟ5�w�[�s��E	�D0591r�Z��U�#��9I�0"PhQ���&tE���ϟ���>]�o&9�O�6�{{�~�ݻ��oH��Y��t�>~����������Ǵw�/����ӈowe��Y]�U���͈��%���7�4�533����o�LX̌�>�g���r�O�����jv��TY��GAY}���S�Q�;:�%x�IUI��L�gG�
��1O�O����*���p�V���6�[U��Q[���*o�d�B���a�Wm�iȔU�͊�kOU4;?n0u�W��_��2+�"2
AU���QJ�U��J�%D�D�#�d�|��}�g�Z[��� �"�R�I�%�T��xc�Z�#���!�0�ѐ*�4SZ߆�VKi�P zR�Ѧm0-�`K�ku��"8��ΰ�r�}�������y����S�ʪ����0��VP�7/�-˶����Qf��z�G���)_l�{V+^v���T�������<Z*i���G=k�9���9�嘮&F�%vÕv�^y��rZB��!=[��e�ZI�� ��a_��ނ���"u�T�$��p�Ւr期Jݏ���BL�<J���s�iw��u���7�݈Br.��I�m����|?糋���n��O��g$b}�I̎%m���1���9+e8��Z����l���p{���������Tgq9�f��r��~�����G������9~�թ���Nt�%��b%�j���e���:Ϸ=�~�y>�8�7�ֲ�E{ T��Eѵ�8SK�����Ɂ�d�/��-�i]�r�:* �M�-"�V�6�d5U�p�ڏъ%
&GRf�8օ�r�犫c�gڽ#n�i��-���������>C�¹t�KS�� f�K
������,lH]�Vυ��hm��,�I��1i��^�4"Qu��������4�v���q��������,�x��Y��.�ɕ?09]���|�5^ˢ�0/K�9��=��⛅�y>ߟ����~@���><Qa����Y�
`O�a~��g�$�o�f#^- �����x<6گ	�xr=����/[�U�f����,i�Xȧ�wF���d�L�~����t9�D�+5W�����m���h1����L��]��m������>ߨ�F��[���=���`���I�U~�|���������~ק����7�Ӊ{�
,�#%�����s�|U�m�sO�����ج+�>6Lnn��Y�x��؆����g�1��>~5��W%p��A@:>x3ѐ�Q��-����O��'1u���X�ј1˝��d!��k��ۢf�h�A_����	�7�g����,����(���G�4s^ ��R�P��|)�X|p��IC�Ξ��b�l��*���� �4N�}^·J�½�[�dG�.�0�Oy��pj��� I�Z��J���Պ3)�x$�+Պ���a�_aج2��'���v`^���m8��O ��#j�!���0���UZ�m�R�4n�i��
G9�����H�|���	A�\���� �x��_?��O��������r����k����q����)��S��s�W���3?r^:q��}m�����x�Z[�N+e����*�~(d�%�"��J_W�w���
p�0��ڨ�W#	�G�+9���F�݄GF(0C�:���l9����)����w@E������!}��O?}�8��H=q#@���UU
�F�X��"5!s"��s�ZI�����
MiيVg��{�kɶ*�o�Z��z�����r����=5�\
 6�^Ы��%-tɕ)8C҈��.�	�5k�Үi��X��D������FĲ����l妟 A��a��E]��4�f9�ŕ�˵��ɴ�c��[6Kp\����ԂQ��Bq���(܄�L�26��9mˎs�"'O��@E~��%엁�рp�T][M��M�6h�
����4[�}����]���jo�cf���
�������pk&}%#Vʙ�Wþ7S[�S���t@
]*|,��h�����Ի. �����/9b{N1[%>G�y��O9s�f���G���K�ȯ�w�܃�W��ט��`f�:���ʩ���̤K�������uʼ��|��T�R����5e���aX�+d�����i]��T�5���MU����2�� ��H�{�����P�f*�,�g�et\��>Z�ݦ��W�/��y�]�ߐl�T�V0,̀��tw�$���S)���j�FY�G�7�Gz#�a����P�h٢�u�^��2r�h����r������^�)Gø��p/�R-*���q������1�Q9�,��\̛D)X�R�@<x�a��v^�X�i!�P)|�����D-&�-��o-��ﻃ5�����v|��rNj(��]AD�̆�Κ��i���K]24͙�l̂F�]��|�GQC03 5�ƣ�E'u��) �C�c�/I]ō�W��(>��-H������$��\c����5�.�@��� =��R�N�G��ãº��o��Ȉ.����K���?/��[���4��I\���t���qa,o��{56I��J�S�Lw�m[?榆z>�S�kͩ����,���f*���$�~��k�W�O'��z-��10���c�`ٮ�8�����A��0��鋃l��(ο}|�h�_��o��N�E2w���n���yH���:�2q0�	�����xuC��3c�x}襩k�a![]��N���]l��&24�A2����R���g��<F�@�L�z���Ŏt@��^��՟,LMK�M��a�ʫ~�ij���|X�����fB��;:���*(b��|�^�)G��l��Ɓ���qqB�MPH�PQ�<�|'o[T��=�Pm[�С*K"��:�*6��@8����������r�J�� ���es���U�7ͨ���p���+آQ.�K�$����+��ab��t����
Z�m�v�"��!�VT{IV5�G6꼕��Z�Z�Q`�z]`��<X�0M�ޗ����Ic�8�r�l�6�F��Q��KQ7=� ApC�%Q��!@�1����S�_v���ՙC�5>5�r��D9��-y���R��k�󫤙�Q�r�:o����������D��x�>�Q=U �[� �?K�V�zE�?�f��n��*H�����)����kר�,[��k0�g�.��C�2�F]�ט� �ҼHL2av��6�n�����(�r�f{XN��O��1s6T��{�Bp������3�#|���5�M��	�#�U͹��`�@"e��a�P�H{k`�.Dil1�0�(2��T|��yr�E�4xb�,�@������ݢ�_�"��9�7@��T�'Wg#�,���l��O�ɬ�½�����$m��e��=�����GM
���[Ax�8��q�7⊸]-�\���R����q��/'_�cΧ.�'�H�u��W���{dQ&����^9�D���5�Smt�3H�G��GTFp�Á�O@�N��`����@���	D���&�o:e�q���M��N��Q�3c9a���VjS��T�K���ZG�L}&. ��M�iS1-e�<_{7=
3�J.o5L��t��;�)�<�zg ^R�?���֖d~��*�M�p^�6��lv��ww�i7E���6Z�C�0��.,u��Dפ��'5s_a_���.��4�i��7Š�M�3�x�X��jY�>/�fVA����<��M��0w�Ǿ���9�۔�P��������Y��0h����Z�q����5֘/3	L���x�瞅�Ё������b��;��J�]����P�`��R�"yԯ&w���i`��u�#�o~:=���\��?E��dso�k����Q`�ť��8�Ƣ��}�HME�x0ߪ���vq}~na9W��S �)�>&y /5iy�YЛ�4�l3$�	&lg�/���Nl`"{)��H7�D�&�.�{�;k?4����x.��
����qhMb 7P·��k�\�Qx�<�&�>G�q'�'��~r�h� �֪.��B�|x~ta+ x�&Zo~F�>G{����z)j�6[���< 4�k��A� �CY[��
��U�����8�Jd4L�9shrm�v��f�T������PAg��%�bw�8�:L��̎��,���s�9��./��(�6�XbS���aJ�|靴,��-!�:��]�]�ϧu�K��%��Ç�_~I?|�N���b����"�z=<3r���N~��T&<�c�k�Ǧ�/9ƣb�������Hs���%�Vk��<yɕ�# &2$Ο>}�:u��B�����f�'X0|w��F��'����ymeEC����Me" � ���i���>���'�9l�8^j
]2n����N��L�<L���H)�����X�(b��o���q`�p �>�g2���n>���P�����'�Ɯ��Ƨ+*F��d���ߎ�z�%���#���  �Feױ'e��v�#�/��ɤ�����=���Ӿz%��r�3|�k�$
�D ��C�'S��k�,�~�UU�Wz�ʑ�Q�ɀ\ͧ�T�������N��!��d���YP�}�/�6+�rL!k5MQc�AV�j���|}�W�7L�Cy];$�\%w�����|�����s�+@6<Cv�5�_4�����-D4��8�I
,KԮk��-���ɆI�)� eV�]��w��*�J����M��������9\7 �DM"��!�K�O����k�p�e�/ލ9���s��~j���݋L�)uD���������a� ��2>ZRc#̗ܶU��A�Ӄ�R���&H�V�	h�q�J%Oe]IlX ��+$�&	����?���o��Ȋ`*X	�#���;��%���:'|	.-{�#���$6�W]�o�"�q���{�?�.0��?v�k��^jj���Y$c�� \ paޅ�����猀s�xZ�>T��<��������U,��7ZL�����{eT0F(!sw�n'�Ť��>�c�Ϝ�#��6>�:�R�v�Yc��4�=�U`�gy��k�;c<_y�#�Ahd�������o�_�����}��"ne����gȾv�2G��u�H0�b�B��%$� L�fٷC�5�@� �����4&Px^�{���
�L�VEܬ3�4��=���,�sL{G�+�2,�Y����>ޘ�ENV4���`�D��m�J�"�<19Vޜ�+ah��q���ݧ�u�>�z�9`�dh%kNU��ҍح�e�օ�P,&�z�釸Fk��8tf���2Xj���ces��Q�Ń����Y�9�*M7� �R�|~7κ7�y����K$l�=�4~�)�f���V��K�|�^�� ��?���(yhl������m�:=�#h�l�T�wfT�E'zIY�HI���4ˍ)W�^6�Q7 �4�v��6�ܜk5cq�c8Y&>�lT�Ĥ����p'�<��k[��*����<�D���:_ԗ��Xa��Tޛ��<�}ٲ*���Jc��2[������{̻����V��I>�i#|�+0'�+�C��l�ccH��p|��5�FD�9��>����5f��,�֋���{��9���Q����1Q�E�N�L��d\0��0`Ⱦ���2�����}��(/s}�%��.Eq��3͇lfF�/��c�T%��f��Il�q�2q�g�������9ѧ�f�<Ӗ_�R����>Tb�*�V3���G�qn��)8�ɘ�CI�>}���(B�?���ͭ�>����'o|�(��Jɢs-Ɲ�5�h���$�{ s���`�&�JcX��Ӣ_�4�i�rHn�פ�O{*����`�M�����R+�pkjߣ�8>��fmh�9T�ů�c:����I�c�<H-y��Q���,~#x���8j����1
0�v�n�k���|�(\&�sS#�^���O�����E;&�\;�A���8y8!�g_2B����򬓳u�M�9��<���!Y�O������zô� ���.��Q�YX�/"�F����d��d>3����g>_xI�r����H��-��i� � �M����?��c��yif/����P��Ṽ<��4N��L��]�8ѧ�="�������ߌ���Y=����5'��n��k%�Ǚ/�O�&����M����x1�6I�%�G9����*F�������AW��ٶW��	�}�����9��*ԏ�i@u��k������ɤ�������-_�(�� �k���L�e��X2J�(L��� �b�!5��>�٠O6a��͋��Н鸿��ɪ��/j����_x�#(��D����jv��kC�wp�x��:�E�L'�dl�I#��#�sM��l�0�.�(S*UA	Gw�*�#[�L������`.12�� ����>�l�i[��fz�n���{�b����3�u�c�e�}m�3��Y�j�� ��*i���,']v����?��V���&<���~�a�`1&'����ܰ��2
��a?n$K0Bm�Q:3gʬ�:%����d��İ��V��r�C���1�vR*�C�SnVI�\� `G�������F��pQ8pd��Y�!���+:۫��^���z��@k�$�0�A;��l:sl��5��(��̎���=ߦ�s��f�����-zc�
K���<:v]����A��Wg��vv��t�O�I=�A7��]q�s���h���n�_zd��dsb:����,��L�`MX-���j���8��D���\]]ɘ�gN*OL�0���K���ؤ�.��M���ܤ�����F�#Q@���m��V��D!=����1�׸X'��<7s������}`	�^��=�攂�z��8������Ĭ�$�L��Oc�1�u�� (�!l��3����ե�����'j����5��pL�̆/<b��$���Q��/_��!/ ��(�\��Q)Y^��O����T1�*K-Yy=+�W�4O}egES��	�㊿"FR*�C�d.>�Y���g�w&7�U&2��I��m���O}����g ��aH����Y����*>�&�<)g�1.
�y_�R���O���\��'��T̣|����>5����� �?�\��|\����	ּ�˨.C�R��Yگ.Ȳ<���4Y����R�#!r��k���I�����B.��
�*[��+[9�;�E�X�p�f��)�Z���8�~�<a���6:���`�YZ岕�Һ���3$�Z\k �Y".1hEhk�����p4LB��!p�T�i��~��Vɨo��0[�f�R���A~�9�S#��.��C
��}h���j�b��0u��6���xl�
�5'��I�O��F�������y�l��.9�����㠵�Z;m��7��[�d���n?~L�'@5��޽}+�G�8i����f�>X�� 20a0O�9=��T�|�O�����%�rb�^��5�U?<��b�������+���en�-�PQ���"�ݨ���Z�xT��%A������xOҳL�80[����͛tq~!e�����~S�YS*����:�틏��*��7�ڇ��\��h 	�3p� �x�V�V�}(e� ,�~��g��o&���LV9�CaM�)o|��3sN��/:��<,)0Hi<��ƌ�0���lu������<�T�j�q��{��&�&�-J;(�)�z�� ��.+6bL���M�����r�Ii^n�Rc�%E�ί�dkgM��T	��^�r}�E��
�;75d&G�W�bE2�d�DLN$x��Ʊ�냬 М8*�q*�����(⻣����t)�Kp��B162ǡZm�?�ڐ-�x�́�HΞɲ ��8}�S�Dec.D�n� *N���F���G��V⇙�%UŴp��V��}/�W�%i	�r�nUȔZe+��o�Ń 	�C��}M�X���h,j���g}���^m!�:�sI�=�_��P�X�x��������w������)���s�t{+_�-�4 �T�dP�Z�霿��o2`K~����Sti�b`�pq
@0�%�T����J1����$�_!��f�瀰�����z�6������b�YD#�#�	���רa������E�FƓѐ`� �����d������?����	�{D%| ��-�2H��*p��Ϗ�߼������ac��E�4#E ��QOM%9�īl���X ��?_L.-L����JG�7��2��@� ��VjB#���5��hF��m�g(�!�fb�Ǭ^���4R�A���1dKiB�� $qO�7�ڕ�o�!:J��o*���I�K�5u>'�k�ڗ����R,�Uߛ�]��q��4����Y�hU��s�^g͍2:F����%>��@?~dN�Ǘ�le� Ϭ�A�|����ƍ�g��"��Šau�j9<ؔ��PG?W4]{�����N�	�M�l�����`o���ߣ�0�1kKE���R"`��sg2��Py��:�_�_�/�V�e��8�X"���v�M�y-��Z�.؍�0�����؋�~�^�	�(���-{��%�M%�[�&��^h�V.���y�76��qQ���M�D��덉�}_�٧_r��E�c�`��i�
r����Y�ߞi>jj��ɼ_���7�䳦��B�%I���R�t�՛7�j�)��6��-�k�d�8�����y�˂���`��wn!��̆�_0(e����z-x��,4A�֔"aر�YD&ȍ�x{Q��P=}��7�痳��l ��a��
���Sd����w�C�߇B�-ua�v6�����Zc4�� Ȏ��7�@S<��QX�6�C�\4��H�yt�?#){*ƥ��� c�.�U�f
V�6ʙ��ĆbC���B��\�
i��5��Ϭ��`
���yX�=:��D2B�JQ��(�Y%Kiԋ���;䷂�K��!���A�B}
&x��n��Ĭ}��F�{qR�Fَ]�AX�˕�Y�?[��d��5"@y���'F�Û\,j9T��V�fK���K$�v�P+
%`S�^F������ n�	|��~n Đ|�7���l<;d�A�B?m��R(���ov�����k�A���G��8��oi'����D���ll(���&7��Ge(��#fv���F�|.���N|�$
N�	l�.7����n��O峋3٤�!��(˃U;ZT�{Q{1;�іj�n|��F���%�����ZRðmb��
� ff��Ӛ�'hdEk�=���e�bC�\�`�R,�v�TG_�1�S��׬�E��P�2a*�/�%*^����Yt#̑d�訏k *�CP�}�6}��w� צO��	��w�sG�G�Rя��\��?��ӗ����ϩ,{Td���'^|�Y�O���kJn;�/�s��`��Hl@�?� �D|��W����qø�s��2�{a?o��8xߘI.	����`���h�FN_� >�-O��W��c6���\��"�g�e�`���hL���>�������� �0J�K0�CI�[����ŉ ��^D7'KI1#*L���d�j�T�3����=y`�{Of�U�i#L\��y�([[�U��b�j�ZAez��䞻b_���^SftL1]`9�#e��f�9|epp�M�LP<}A����1��9����~7T�����V�:Go��(9�Z�M�X2�� D��|r]·� A..�� �	U� ll�M��Y7N?{	C��&�;���9k�������5��{��|bU����W����
&�w�#���~ٶR�{��O�tb�1M8�-��7����4 .��`�M��s�{{ݐ�rB��z�+�PkZ�f;��O�h,��,�v�@u��H�hf�@Y0�m��67j��ڄ�c�h,��s��d��n�s�u;y݃�sA�Cs`d���	=^kM���V-�~A����ƪ�&	~`6�W藵7���U�iqg�%��o|]^\N��&}�ͷ"�%@�ۈ�*`fhl�uɲ��mӺ�]
���+*�H��R㉟��+�'��죔TV�<��j���g��:�%�{�a���/�GG�� ��	\C����t�(b����{���w�[��& tЁ_-��d>1	����4[���Qu}=�U��뿏��8�ŀ.6�g*>й-��d��$��FO/7l�gS���bTd�%F86��y@��+&��*�8�O�(���1:fX�-Y�R>~1K��k
 sR+�ԟ,�4ˇ����V���h���h��q5i0��d@u�	�f�{���@ԭ*�j���ރ���|tV_�&��N)�_��z4bȝ�R����}�+��?\�X�k
1���?��V�G��HHI&�-���퍼r�"�܄<q�O3�,� @��Q��,90q5�%�oc�޽v�%y����������N�o�:AJZ_
�8��qS�W�@?h���h?���߃�"�0v�! �R�1�a�P	Ӡi�ݱ��]���X��x�@�rp�o/����fz4g]S�L���t ��t���&�޲�,*����F�}�=�;h1�^M ��ZB��Rs��ً��?~�K��I[����O�~u��|TXa�H���Q��ާO�u7�L@`���Ls��-|	���n��O�=�D�!~
��b�"k#I�T.l�1$xva$�< (���I#�W��ME")H��ñ���/�;Sf��5�Y��_��CH5��
3_����i
�F���t��mZD�	������K�D�s9�����e)(���5�߼�q.6�\M Z�C���f3�K������ag�Z�������~�EHj;���Zfr�\ߩ�3~ǧ:���?��\�(=c�0�	M�r`�K?5Y��A!�\X`�.�=L��:���\`��S�_��2� )9����~n:�,m��k �Q��r�z��(�g�~�{ʴ�zF{:�'yr�0��T�ZM�^,� esCI*��~����gL"�0GJ:<.����
��m�#�L}[T���jGV6��'5����1 g*ã�H� !��tJ�lR=+���¬�$��b���P�y����gF3&��P��� k�!m��J�T�������>� �yu�G�  �-���n��%Y�)�P��&M�Wޥ���y#�!�̎���	��`��̊:��B�%��7��+��ᏹ�M¾���
�
�%���_9I��r̡�\t���k��_V�f�-��i=qW�/���՘��` N���0��HE�� ��-RUle�e8�8^[v|0ge�r���яm���HW��)��RBc�A���o�޸cye�2s΂%Q209��:{V���k��ͳb>W���0�����Q��^��55��ց�hQrRbʘ��X1l�I4uM�(�34-������2�M���ozC�<uG���)32�s�|�qH~��'��+]�=�f�}7����A%�~�ùM�H"��	��6S1�P&6�,���AX��sI��-rqy�|���e�>��_�JD|��>L�o��Y������cH,��K9� �FK}�ά~��E��D� �����4�~��O=�|ڍ0`��c����qa[$P	�p��V� �JMk
�$���#��y���`݀[��ľ�$:�$\֍N�t)�O��0�tPQV���hLQ(� s�5Zު�~��h3�b��-�>?dI��|��t 3'��y����qcʬo�� _
`�l���HL��Fd��_���:��C���933A��ShCS�M�D�+]�K3�s4�!�A� �Xu-�]G�00���?��Z�|�y�d��-��n���)[8�]y�K=2r��?OB�va{�� �Љ1q\��f�5���9y	��3O[�FE���Q� @��q��5M5m� C�߼��(�k���KڣQ)�T�e_����P�R'r��u���2�t�Iss��ōe�W�Z���)`Ek�5?n-)jr���p�Wv�9�s�V_�j@��(�|2�3b#��I�px ��w���`��Ogg�e�}��Ӱ��l�I�R}7j^��E�~���GЖ�$�>g9���8d�H�d�\��C01��EK�$;��}gz�! ރ<H��{$m}mY���ߋА3��}L��@;vH8��P��28Dᆍ|& =�h�$x�<�#��ɳ�%}c߹c���8��=	��<���Х���#:��Z�A��fw�=q4g}Nx��`JN���\h9��+H�w�:}G����:�Ѫ��s��wwۣ_o�����9�50)�6߆469�{F1a��Hr+nj����5���t������K�K��a��{�ƀR��s�ilZ�����2%
v�ϑ���4N�  ��&�]��j�C{#�r:N }s& `3���J�� %R7
�j	:�U���y\����5�@+���8h�|�>�gg��0�M��܁�ce�:M����siYМU��Z��Fu� Ke?!�������̥G����ɗ{/e�!�є�S�BA����b�_I��6 �b����u#�D\J+�P)�נA��n��9���I�R`�h�$�$�DL'�a��I�ޤ����4g鰟�õ�yn�	Ly�����#�_�y��:�Ͱ�M������,3Q���T�Q 6��-�� ��>^KC�sz�&���t{�O��j�G�Ȋb΀l�G��:���n� c�bn�����'�o/@1���2�7MeJ0!r�L��2f�d��E�5�+��4����B�Ӵф�̌�sb7�H���*�e��-u�3��2<���
�EP�	8g�9��{x�R�Y|����Ϻ��R�r7&��4΄�>���a0܏���ڍ�Q�:�F]4�E@+���&�҃�.Mй @�KwwȠ��tyy!cx~q�Y���.WV9<zb�˫�]���:��x	j֙�c��炡�y��=��x�y�35�i=��:�DF@��Hf� ``D�����!�e|�>nk�O^o����P	V�i�sx�(w�f��������MoY �� ����x�/���h<�.��.l��ɶ(�4ti7ZV{W���
f��0W_���n��v�G�IZl���pX R�) �X�̗�/}a�֯ c�$`i�� Q
�k-��9��W�"=T!��L�M�ԉXh��"�`	����?;��l�p�y���+�X4J3��Z/@i���d���L�E�L-��[��b�aP&uh��|P���=�|0����^��̰^W}�:��Ae�~�ur�>lx�m8���X��x�Y1���`�w� Q<�n\R4@��!���XIc�:<D��R;!�M�J���~o��on�o~�m���V�0��qe���敌��ƈ��@~��O�[Q�� T�v�Qi?�P[rd��f.���.,c�J����e|gM��	#a��/�.}$6�������{����{��_~N�O;A�
 5��`p�,It�M ж`��dU&Y*�fB���l#�P�t�� \
rkm��no�U�,.I�ڊe�Z��|��"�wz��]4��hw+��J�P���8I6Y���P�*����^M��&��f�ͻ7�:;�dQ�\�y��]ۆ�g9e���S���7G�(i* �&�a�J�74-#J���W.U!D�I�i���}�DX�Ndǲ��ъ?�oN֝�0� ������Ï?���j Sl.��0��sA�\E){�~����W�R/���IS��}�AY��s���0W��D��k-��dѠ ��e)W��z�;)0����o�)��N��#�|T�$����m��W�e�ڽJ�K��dP���/rJ� ۄ�MVY��Xm���jK��vM4�Ygj;�����$��`���IԽ2��)�XY��dH1omR�`#�9����}�"<�WM�x��Jd�^0�4S�e����O����O�ߧ�ۏR�?��5�h����Y�\��)�T�˾&j�	ֻl�4S�$���_�! :��ڳ���U�u+�.�Ӟ�L2K����� ߆���Ԉ !��-l�R��`Q�⣬�Ŧg���{sbn���8�X�1���I��h��{�@KR�5�:�}|���xՂlk���8�}��pvΡtW� N��쾈t�{
�/�uڷ��A�"���Q�7bvVE��&��ö�|@��@�������W���.�}�fB����ք`!j���dq��*�"�u����|�53��$ayI,9\EҶ��i�Pk�eC}�č�f��Ƈ2 k�L�ٞ7��Fg�$�B���m/��i�������{Hno�_J����g��:��l7@�Zg�&��\P�0;+/d���] #�|=��yw�ڎm�:���x� B���|���>g�v6��9q������"�^#�����z�g�`yyإ��\�dp$�n�e��q�k��w��7���8��gIA��� �������v�xs���ij��9�$~<�.,TL��b�Fվ����"�)�&�g�H_0�ߏ��)D>N���O�0����I?����Iy:K��F��:#�{���{��zd����\�e΀���z�ͪ>l%�y=�x����u�h�V��>D�͓�?:�h , �b��V#�'N^[�~�'�iƈQ��^�P�'��1�M�n���L-ҁ���ng��:�s�2g�m���^��S���]�j�LX��h�%����
a�h�KS���C�/w����!-]�f�-R:M?v����<��_��I�HJ�i?��~�T>���l�L�����Q+�11��� Ӂ�ͭ&YRs��k��d\�~���%<�\��/�����I�g�D�������~@�$ۃ+�xh�����Y�.'�t&e&���i���+-����N�;<���¦]��[�0A�9 Oq�0��� oL���r�Y�����ޫ?>+�g��,X.%����,�7��:�����#���F
&��E�~��U���o�7o��ٶI��iP;�2Hx`�6|Ydd�j Xԟ���Fˋ"etF�3��p@�J8�9J��{��,�:�n
�����Bg�&�����xf���B`�Z�^JMVp����6�K�F��F0hl)�Բ��`t�T(
�$���[�+K g�_�/c��{К_�݁I��:(���hG-/�E��S_�<ͭ%�ٞ4��/��iQ?�b��5%�>RT [��$B�3#Ŋy��8�F4��7o�a��ﾗ�#�Ћ��=|`Z�6ȕ��{�F��q9n�q��G� $����~uʴ�s%
Θ�"�	�/��Y���<"PG`q�����T�sM|��/�z�Pj��Ⳕ�����k,|��_)��:hbݱ�eE�I�1�A���ج�Έ�戣��#2^/����g?Q&s���ON���,ǔ��a����s�c$��ۊ��9JMP�'T?��m�Ʃ ���s���r�aM3X#&�?_s�>�ң(�	)Ά�t4�1�v��K�B��R"L��Ca�w�#)����^n�y��EQ� zo{����ɴ)�U+Cp�2��Q�Z�-��%�f��_�$(�����ݴ��M?w���i�֜ng���\���}�����ɰHh��ր��1g_%0�ę�1��k�_��Hf�D�wZ>�rX���h�Q݇�ʥ�j	��Ӏ1qUٶ��KJ��ҷoߤ�o�K������s1�BH#1���7 a{M�ԫr��|�gק�Y��$�wߴMz�9�Q����%��"�OK�:�Y땠 �s۾.p�nt){~q%����Or/�(�� qtRk���O@l3�0A./PR57�@�{�╬��j��9D�HZ�TC�[��¨�������=�+>S��22)$Ӭi9BiV]֤��@�Ҧh�,��J�^U�C��b�j~��:��a� � ,���&����d��a~8X���|�L��@w�թs6��riH�%L�D����f�澍��cEM*��~ة�R����Pm���ڌvb#���&}�识z`���eZֻkZ���̼
3癘Uk��b;�h���g�D��_��7�HF,������\U:˪	����͚�io
0l���͐�t�0S����p4�e��``�$:�[�?��� �ˡ��0�>���50g$Ǐi���hީ1�@�1�`����u���c�}n{f�K�z����(VQ�l ��S�$�c.< `1�1���_p��t���5����٥��h��[Q�$}x{iKpr�Su慨D��z*�2SR� ��k�L��A���B�B"�q�K��t���Ϩ�A�5��xtS�ȳ<Z:$��d����U���ʞߨ)�c
�� �[Fd�����p{A��8.XI�j1`ʙƲ�Ӊ�Ϋ?*!�~-Lu�M�Z��D����U�����U�4KJ�͇�kl[uE����yzw�M���ߤ��� �M��N2y�Ģrlvn9�:��u'�!�.�~$��M�U�Q�HM߅[ϻ�o��=@��[	�콃������X� ���qV�2^�I.�]���7�=@��� N�0�V�:��Y\gR����!������5
=Ű�d�F�A��Zk% �����qq'8���t�m��1K\�j)2	��s���0a�����'mV欨m_盱{��K�6�,ml��Kp��vg�L+4(k%���E;S�a�M�VB�1M�u�q���&�\���jE�k"?-K��ǃ�D�	�8�!��\�r�����{�A��߉vF[�Q�60w�NT��〆vf7i�_�'�M����O�|��l�+�S(�s�N���q��YHaB�X�yM�/8f��X�Ϣjm�d���F�G&�YЋ�J�[�$o!�IML�E��'[+C�9a�22���&����t@;���/����&�2ov"�q���mt,���������>�y'嫺�1|����Y�3¤�1�5�E���h�����_,�*�Q�l��'�	 �P3Ԧ{���0��d��+�:���M�Z�����r����BK��Lؚ�{l�=�bl����6�:�@�+�t��	��Z] ��ࣩ��ٺ�b/z��m���6��?�n;݋7>&Q��������k�ǲ!�2�@�ΘH
�ZeyؽMg��p�)4R�C����>�k�r�4��� ,�"�1I%OH*a�h�c�h���,���x(߃�s��k�'Z<X��$�Ia#�� m��M�usަ�~�6����?��7;OW� m���#������������,��K��t$�,��	Z����,�</�sq��p �WWjVԽP}5X�7f:����:Z)�9~=�{D|�n�y��>}��K�����g�.��ٴ���1b$YF���e���r�J� E6 Un�G���?3/
yif���>Q�JU_bL)9H_1�8*+& ���6�1��߉�B���T�f��	?`_O�x7m���2@��68b��&lỬ�H��l�T#c���Xvr��9�RALhՃ�vp�X�mc��A���2��%ճ9�H�F|����&���65;
��*Z6�|��30;X�h��	�3Yڑ�`�7^:*�J��D���,����l.(�Vߤ�����M�q﹞0>�@������3y>��fF'���	��4lᬋ������q Gc����=�k���l����K��g�T�M#?g]�g��s|��Q�k��f
���`�4%�pg�Oj�C���Y���?1M��jt�6ވ���p+ƍ�q�o=Ō畳�C����F(Vd�(D�ڝ�Es��e��T���wǻ-�Rw���ܫ�L��ф�[��#d����� ȳvqq�AO���k(���^��a?��T<J:吶�Eq|o4M�A��������e�o�7>VNb)8?��Z��3j�` ��fz�� TF)�`� ���V��}ͧ42�`�2���7j���۳��Ј��l�s._xm���
��<��w�&���I��O?���杀6�.�Ϧ� ��d+�v��PΧ��_9'K�cN�fF�l=۪��0�);f��&oYj�����Z��(�ߝe)(����X�Ju�R�$�����������z(	�/:���g~x�X4<4�,9b�eP�E]����0,�	e]95"Ґ5����]����hf�Q#���A`O�"� =��.Q�
�\�m�(څ�,�TLf����G�D�5��f��[0jSX�`��$��%��2b�;��V�a���Ll���5O5�T!̎d`�~́�%{�I�Tc�	���h��k�����fG�O$Q"�{Q,{+�=�,6��o�G�j2;L��ajrCcc�꿷Ze���7��f�W3@hlC�?Z�&T~M���Pu�Ɨ�]fr���&,��ݠOP��/�cg��{c����@�m0 �R�����J>�	�b���?}�����jر˫K�|�pH���_I}�����C�����֠���̣�5~�cFa���L(��&{�K�|4�.�a��NsT���T�>�Z��	X�H�����
�>�y�1�Z�eO����5�0l���������c�E_�Y���5 �s�x��m���|o������ll��E�^eM+��]h+�������rf���>�Im���Z�@N+��QV�`��׊j�D�c;)>��G�A9�V�A#��N���A�L�b\�뛷Ӛ�������)1�<xVL�v�D����Z�g�๒�weU,ˢ��L~!�`n	����A���<7|����C����?�6��?���]��^���U4>���5�J4�� 	�+��I*P��ȏ�j�f31g�(x�f��PD3$�X�0%dϐ�-����W���0%i�:��D$+��6�����u�7ߤ���uZ�L�ܧ�	���S���pC�Dm2�留*�fI��:�\
N,���MI�O��6̪�D��v��	5�NԲ�/"5%�7	2Y<��U5r��kk7�gRxe�5%��5 n T#{�����K�t�c��-�y�<�W�XK5q0���0�6��ښi(7�����uF�ƾ���6<�����g�/rR)�T�͠��I"���l�����)4�E����fT�F�N�!�Z������c��+�:<��D��n����wuM�����3`�PMｷtx�7oߊ\k� b2SKZ�H�\�^���o�*Ɠ@�`�h�������u퀏��~r,	u�!��^�>�3�\��9�6���k���z��7��A��v�����_�a�@c|4/�ĨI���V�L��� �{�<*�ht10���dn$����?��G��-F�1�>�9f:�[��c_����.��u�����u���l��&�n� �	='�I��q�P�q'���%�x�$	�H
c��RL�L�n0�)�q?��o$Z\rAM�{�ij���L����N�f(ao�~�./�dm�W��~/ѫ�'��b�{��^���c��2�j���ۨ�UwS�ՍHq�h� \dָY"�/��%@�M83���1����'�M��H�$15w���pU]Sս;K�#����)�����UP8���h���f��
�G��Jd~�)*�*��<;��y,��|������t�	��!���u�	r�dn��7&6�Y�6��~Y�S1`��S|�����ބ��by�~d����^���P�vL.���E���X�Ro���F!�����D��U�bV�k(o0�o�T
��pY ~���X��@���^%RE��f�K�z1L1�
 T��>����5 ��ao��(NN��E� k�F�'��K�Q#ݯ�u��h��P��=3GC��T�Ѯ�C#KY(P�CU�<�3_X(�֖�/H��"���uѷ�B;c�4�d��u���P_�cV�;[+k���Rc�7�m+�.�����J
���yU���Q�g�px��m@�Q�~�#�2�얯�~\Nsǟ�E�Tl�bO��}�!R[$<~��9����o宴�;LV+���#�������9tvv �j|A��3���f2�e��|9C}��<��!����Zc ���;�_�^��,>{P�@5�mY�pmd���Ct���h��M�>�ޗƏ�z������Y,�3J`x���Q�sЎh�ׯߔ�_a��^\@Y�J�N�{���Zf68 �Á�h��h�`��Ϫݧ��,���W/��50Yuʒ����b��z{\�u�:s�u�.�Ϣ�Ҙ�����݆_�H�vl8NX�G3z�Hd����T�����A*�U ��F޽}��k�Cl��������1|I�$łmY{����nW����~Q�~��i�g�����԰RS��3\o�}(}��2�Qf�5�H�%��u1�;��2K1#��m׽�̔]«�3��w�8�d�a�F���RV�}5�s{K��L0�'yxy.��÷��) �<</�;ܪb��C֪��źb-�A<��2��0Q��c��.���k�+VrQ���\���\.m��A߮t�x��A�̜B�"�L�V�v<��0�G_h{�\T��r��퍼y���W��QW��2מ41�E�p�?�]uy%/^|���ƪ�l�q����vt�%2��dLV�������H&�fH��c���c#գ�;�ry��g�u���f����X-���f���XT�
�������+��"�{��Nc���t��J�S;�
e���j桘�rX{��-l�ZԘ/�T`�<���S�YwO�ȚiAoCӰ�͙/�n�VOY+�MzS]���͠��'J!�a�c���n�>�iO3=����C%��Vc��N�Y�}�v���0��7�WA�w�N\��Z��Y�}g�����ke��:�1� ��K(ړʶ�`�-�1!�Y}P_��j�k�Ν����yS ����\K��Q`Tn�t�d�GY�Oky�d����3�����k����׼_��{�:T� s�믯K�X�ύ��Çt={�d/��W�7ǊD��݁���]ɘ3�-猲[e��嗲Yэ �{�� g�/��N�gS�v�7���v�����*s0=�s7�����	�s����'��4�ug���qM2ςf�g���0����-�\�|�ѽS�B��1S�H�W��w�^
�3��Q�.�w����i}Gğ9�,�#y�g�P���ꝗk�y�V�\��Ѷ�:�[�n��/J( �cB�;���WI�=���Z����yck��&�u.	�n@����S2Q��2�/�Ow[�::Q�ɵ�"�M����W��1��0b�]��c�`cg�M�
�?yV�g��P����:�S���d2�oB��z*�ӵ���ܼO�fe�n6�N�]=z�D�>&W��ȦLRП(y�؃�@+m��ֲ`]d)���\�'A� OZ�VLkg��fWbJ��˨�� ؠs� |ds,���HPI���:'O��6�LNP����}�ƥʁ�����ݨr��/�M��֚�Z_����4���9��w+fRe�6d9�eօ�* �~.*�A�뭩p�A���T�1f*Yߥ��Ɖm���Y��7-3e���0~��Ю���{��\��92,���:��� �9G&b�O��ǉ��Z>.t�_�G6��7����O
�����?+ #�X0��[ $�?GM��O����kΊ�n�"ɼ�W�9{�����k����&/_�Rׇz�G���w+�2q���{R��F�ZQS�_7�c��/e�>�Xt�)��[�ڗ�g2�����>��vg�.@��3�`� �~���}@��12)k9/�>�
.*��%��4>��B��Np(e  ��}]���� bl��
w�,b�
\&�ZX��1 ʹ�/ZV�_�0VJ���f��g	>��͔{��@`]"D��*������Ũ��^�krL�}������-���r�m��egT�3�ڷ�3�z�ao���S}�NA4~3��7 ��&��Y�`���S)��T4Z,�x�:�~�	&��;e�H<�o���6�����tu��O���<���w����[Y��=�X��1Hsx��]9�M�S}�A�M�����s]�!������5������`����a/,cC�DA�V�9Wƒ^-�\J.��vu`�6�����4��N���5��y���G���L��CP0�o��"ճ� ��"���#yP&(�9�ܨu���+��%�����Vu�9����Aa=�}s�.!�:�;R�{jh��
!`�Ga��@�%2���ج4�J�Xّ�R2�0��>ƔTX�S9[��ו�`��,���^���0�JZ��iv���"f�3��M�E����L��ԙ˚`���D�H( 3u��'k2��%л���V�����s�A ��Bf2*��B��7�j �y�kn\0Aa��@���LBc��n���#yƟ�LHa��砬T�c�b��� ��l�84&lb���e��P@���ңGe^���R�^�4c��`�,S�A�H x���`b�#����O?�����B:�@� ���o"}#���K�1v�>��t�{_���1w�Ǯ�[G,kr�u�v��d��(��j �z�� �V�K�"|V�����^��l\ ,��`c�|�C0�Z��\a&�b�߼�F�={�c
﹀p�N��i]��7*nZ�=/ْ�vm� �������d�����37b��]e�V��`=$��k�x�S����e��׽}��XV14�v���8 [���s  �5��5{R<C��=@7���i
�����]�`��Fs��b��]Y>_�s�A�O�>�	v{��ɣKy�`��3U����u�
D���&2S�&Q��U7|. ��Y�؋�/5������Q9'�Eh�����J���޺=0�sL���C�N���F�@L�U9&b��a��,T� y�Od<n�XJ� �W���u~����U­>��:TO��d_m��׷L���e\6�3-�<Ġ�m�f�����jSنV]51�M�栵��ep���k� ��e�m\��gI���	�3Af� &�A���\覅E��j�Y#���$IRS�9`UZ!Y�H�w(�9����~$��"؞,��z����z�|)c���;����:5�W6h<^n����
rOV�Ճ�k���qc�|�>��j���j6z^�AA�������kT�V�]����}����*M���J¦��T��I�K1�#�<I�Y+���Ҍ/���ln8�m���;�>%S,�+����!*:��g��l�{cY&X�����qt!�T� M��|�]i c?��������WW�
�VM� ���:X��w���҄����[���?�T	6~ee
0��|���f��ŉ�������P��s��f�����6�T���1l����Ę-۳�p?�6A�WW?k?`������w0N4��,��������Ϙgg*_@��p�eM{��z����[XD�~�ٸ�N�~5���ӿٮ�����?�p߄Ĝ��T�콅�t���d�Z��Y�K��kR;t��s�I+oWfg���a
[gL��+��}��Y�Fb�Q���T��BM�I]t��]0�J�b��ҿ$OE�WM��.o#��/w�y;�����Y�I���G	���@➨se_z0_���O+{�݇2n��5/�t���5)��+�݆ͅ|��o��򑂗���jh�ק�<=+�� ��.�Ո�+k��N�		���  ��2S��v�����"�-�4i��Ë�Qp~ .��:;+k|y-���`s�};<���P��VKDw;0���M�pڹ�mj)���t�[���%a����,Se��G�jL��}s�?[X	`��,�(3���eӥ�)��у��u�v;���B�\g����z��B�{B/s�
�;�TҴP"V�0�
���IW��� ��.��8x��*5ͭ 
�%tAO���#���ƃYM��`⏽Ŋ9p�1`_ itL�U���3Y���q���չU��|�lR��Ήt8�1��b#pye\Z�_���5�p����|q��|���3��'w�����穮�|�R�m��&��_X��z�<K���9����`�
p�@n��O�^W��Ȓ�Y��0 > 7~?D��Çz-M�(���xmR ��n� s^ؙ��پ �gɵ�I���/]a�r���1���a$!H]����{_�}���6�_��-۵����M�����:��U�
��	��&�ڕ�s�����X^�P|�K�x�Y�x�xF[���� n)D���~��/�X(7��uf���|�f8%�`���#�?��k��Q�5��U����2^)��LmEv*�������euui�:k��T�+��az���t�呉k�Z4�)��\Iu��� ��^Oy��\��M-�D�[5�1�P��Ie(�>~$O=(�6���"^>Ю�u~}j���������*�!Vg��R���}K�����{��[�g�{���me>�I�/�5�=�7t�?u�2K�OH�5�.5��B0�qtA��z��7pv�7����Mhsm-JP36�������h3}��f5q��y��r�ƪU��:'�;Q>�(wy�P�ְ�
$�Q�_�F_����� �w
.6+��V̔���<�0�L<h�m95����b����8�U�5w��w쪼�� \k8�Ί[O��8x�y����/_�Ɋ!͒�m��9Fz;���-\ݾ3�����/ҳp{r�U7���`v�и�f�i]H�
�1V�aS�+�U�ag��Yl��A*��8����T 6M���m�b�b��%�K�K�kV�B��%{�I՚as�nh�	�@[0P/^��F\� 赩���|�|��5�l��ǽo�����H��C7ucH �@���~��^������Rgߝ�\�m���0W���ɀ%C���4���s�'ٴ��~���u���C|�R1�����];.F����z��	<<�>��Bԇ{`���:��
��1���,���u��G뒌x	��i�0Z�wu�S�:�̝���{�iA߈�5�s�`+Ѡ}�+�خek�F?�`���^��7��Bڠ�g��z��#"k������N�k���J�u�:����ғ�LvB�2�1@������-� �P@�y�
F���r���e��a{�@����g��,�Db�I�Zq@�;�k��[��
=�>�eￔ�j�jr�>O�E�	���i��b��|@�G1X��}�x���t���@�b�f%�陽X=�
��&$�m
�,��Z+�Va̑���"��MAv��)��C�B��dt��Y�?0�-�o��g٨ڔ�`0�H�/!Ht�wv	��e*�ҰH�E�� �L��Uـ����U�{ǒ-P��L>I�J���di��t�4�;&^�(ĄVO�ڶ�s�}����kr���,R���V��L-���E�4��<Q��+mi���j&v)J�P#�PݎS6�(���k�3n�R��8�~G�	��
����@�Kθ��օ�83���LvM�W0� ����$N�Ū����|͵BBW/�c����}�x�Ԗ1.���uc�7���fe����mm6G͜� ���_s��9��9���_���}�j�Qw_]X���+U೼W���|?+��eƐ�c�c�q�3Z�X��g>~N��쵯� p߹��Im�.6\Ct�I0�������8�*�x��ok�z�����Ŀ��܅��Y�p=�AõO���~5�D�֩�'n�:���}}��ڴ��9�,9x����xLX
)�Gw26~0�+��� ;��.��)�K�!v����ʊ��}0^��W�kS�]�̞�ǰ��~�8�������,V�/-��#���+�f���{���2'WL��ȗln��*�Lf���}��+��,��s_��e?;�����Z V���+9�(f�cL�~�Z1n簇��փ|�g�S�_�/Vv�<yi��4�\�T�g��g7 (����W�w�:6'��S7��Al��?����Ҡ��F��/�*��Y��W�?X'��|���h@�wP#�nǻ���n��rL�A<z"���Y�v�U�	�j�.�*]0&8�*����^]��?S��.d�u�  (����s
F�b�b�Rkc�Jd��@�s�/�$�ꪬ���nnUwm��ف�ŋmL�Zu��s�5�/�7�J��S���x1X[���:lo��-�F�� ����`-AƋyP*ۆ��cBY�2�wK��`��gt�}-:�4qv��\��0o{>Տs*��_~T�N�8ܽ�g�k�I�zr��HKW���i��^�Ļ Dn����I�6S�wlp!�* �� `��6`��ݔ|(����v�CZ7te5@-V�7���0ՕP�~�aGV��}r��{-P[��ٿ�ǧ����1iK0���=�e�~� ����:	��"e��"S���<�u���*�Ivye�?sy�h]'R`za+/�.2˔n۹��6����ڡ�(���4�<JN�����.(�Tt����cxسXU >B�rgMi<�����9&�.��,����e~n��n"������xt��J%�!��Lh���1��Z,�h<�{�����=�R&ge��~8�>��-����5�&���I�]�#lN����O,?���Ա<Qzie]�Z�;��#��zl,i��[�#{p�uU~.��\%��1��\#O3R��	\.��E���t���kM���z��q1P8o@��Ɓ��k��	u�p{���!���ݩ��I$�E�LJ+ YP��'���x�O��>[���A��C� ��C�b>���T�]���8�h���P0@\���� \�	����R#S��&�k�p�����1��
� ��֣�^�Y-���-m&b��\3��3�o#Z\E'����A�h������u�5}���R��b�zS:���84E�'�5����mJ?�)Mm��CA:�NY��_�-�4���@}�C	a<օ4yܯgv�� ٯ�p��cSA	�<5�}Lf�1W1�4u�z�����/�u�h��?�&�S��;�����3$�H�o4�Yz�X\�A��ɓx�{,���d,��Yg]��8\$8 ���o8>��/l�|tGm6븧<�f6U�O�Ԃ�%H�W��X�S�Y��T��h�T@�),�}.ה���̜�������|����@�ދ�O�;�w��e롪�?$�nK���!~�I$~��4-c��9f�٩�j�N�n�zsPƾ�S����1��� #Ӳ�M��7f�Ln&�y�uU �B�e�xbzqƐQ�»3Z�2]a�ks ��֮�T���#�w��MX���\fU�×մOmoo k�{��m�9y6?��Y�d�����\���<p|�MI����S�WU�W �yQ��2�K`�:*#8�g�˛��\gEj�vҾX��4�q?���z� �z]�5�B��+I��N�3hR��WJyr�����Ff��0 ~�ي��5������j�%g�����gZvb���fklWz�~���ܨb�2_�<e������l��޽I0�0�xe�� `(~;"LE�E�ݪ˦���<e,[@)�@�	��8����e����lU���ب��^3cQm�� ���x�{k�PХZnA��^��xν�+��5�+e	�S�P|���]T�DSj������VMGA�>�K�
�
�*m�����`!{J�Yrl��k�,��U���HB�L��:_�ڡ������)��{�U|��;cQ�˲-`��r��������-��Ŷ�M�.��n�tVv�-��5�qA8"��Ɔ�6��2�Z������#v_�v�����ƀ3@�r�ܵ����{�\/��ގ[��p������������k���g�б2����;�p���Zz�3��y�aX��F�ﯭy9ZҊ�R���U�0����Cl��2�u-NZy��8�o8˭�_�z2.�aD�X]H��;`�wN�xE <�Qa[�)����0x�n�ߟL�z�bO#�,�3�=kϓ�F�D{?���#��P�<�\�_� Ҭq2_�|E�U��!g�V��ˬ�܆���lX�~8�ߩߨ�]P�$"�b����D�Se�4)���r�Ww���3��}O��;"��E۝�f���)��fP���x�n� 1��_�F�dQ{#�i�J�L���pF�.�����ss"�h?>�ą�l�q��:�ep�{01��P����
�����W�P'%)�Ś�>�H�ƕǃ���X��ִHgB2����9]o�XGe�'s?QQ�e��4�z.�ʉ?U&j�7�k���Q���3����nَ3�.���I}���>E�vUw�] FV���l�Of�
�����n86�|������+X���`�*��2g�F|���p9|�-}.�b`����rͦM4|�̠Hr�Ս��1s���FT6%+�l���5��*�J�	�������H�ˋg�r�#԰0�&�Vl>4gZ2}K7�om�K���?�9z�����5OŻ���$��1쯳2����)�R���pט�����=��8�Nbc��M�� $��֝��v���ձ �Q�v��~�#y��G�'^�3����J[[<Q���X{W���M��^���P!�dƹ�Ø��97��!���,��[)�$!@.�<�:�m�:�Cua	�F��z89Q7��z����^�������0�ߊ|=�$��C�������lk�l1Wi�~��F]y�FY�d�-C�����R�a3�2��PTx��)����]ki����>� 9�C]�V� �_ ;P��S6�7�(����tbE�u���7�wf��5@�y&ki$
l�ab��`�aS:�\V����R���+�$��T�>ՕDtbn�d��G�?�n��'�Y����8�Y}���?K��-cÁ��d�'��6�({�|yl�h~pg�t�Zu5�����*�Q��Z+��X*}�xtSG`6 ��|���(SXe @��� �%y�1��T��$���[��2z�e4��������2��Ef;��Պ*�ʃ��r�[~���%�5��ظ�V�r`���IK�"����-���1%�h�*�Ȍ-��4��,Cw)j���gvLĘ4=}��_�������
ܫ&�Gg��6��C�w�-�`^���Y�:@�`�j��w6N3w~�`��o���8� a	Ėל�N�Y׺����F1JXu�c�]\
����u#[_�`������h��Ǒ˖xA�΁�լ\u�4P6��-7,<�ߍ�%��3��;�2b���k��5�ɟ�U���s����u���ZZK%U��X{<���������,ufo�D-*�����Y�\7��y0b�^���;���Ў\�Z�Y08���h�a"��y�a"��5әZW��f�s��2j�u0׿�+r��C3�;{��K��RͰ!]&U�;@��� �!�3��OqO9��14$σG�u���)������S��M��e~)SG\��j\&���c۽j���냤j)�,��~���m/� �����z�Z{����`w�Q�� ]�x/-���A�>�&4�a ��0�,�=;�)����N��	B��'{`+S��vѴ���@C2bn�x���1�b��x]/M^C�$R6�?�v�*����Igf�ƙA����a9���{1p���"�YL�u��Dj��ݨٙ��h�b<o�
�6��{�U�Y7g�W�٩.k_uA��6�Eyѡ��g2]�b�����cC���P�'�4lD^�9G6�&�]T�ޅ�fcCe���S���|#^������̴rP���.�x�f��!��O4Nf�aÀ��?�/�Rv���?�[���9�3Ki�ֵ���kN������)�>;-��K�.]g�v	�pP\�f3�`��l�'��a�k�Z�6������ۮ�ε������h�l��ޘrg9�Ԯ 3-�ͩx/7"�������T�(ͼs��r�}�O���4�\³��i�%U����\�%Re��k��Z����e��	�������}vѦ4ީ�N餦��J� ���^�l�+��Ծ�f�8����Z���a�Ś|\t~O�d�x�Rb�Rg�����z)�ҟ���m�ſ�$j���{b�k~q��uw*!���9��!��IVت�h��IZius�:#��T�!=�|�ҧ�y�j���($�� :9:?:��,^��XZ��Vk��4[��0t~/�d:�N������A]my���bÏ����w�Ж���e ��u�j�l9�����%-z]D�,CMY�r��D��� �&U1Yqd�]�����l���`ޙ\�vgnGޏ
��[ԙ,,N�p��, ��k��Må>�V	�Jl`���72��d�eX<����Ă1�U!�v��m�#��/0�w�����ͺ]$<��.Н���U�Ni��yR�LZ��:J��j�R3�� ��%0@/�A �9�����Ϭ>(Y�\e
�额��c\��j+wP��\� ��P�:�[���>�~�}�a�s�u�w�܋��w'��ߍ����o���h������md��w{���3���șC8<��u	�n�9<��ץIp�v���c�6q���3�v>, y+���0���~�ѹm���
k�*͡I=Lp�����}{����2����j<:L\��ˡ������Y{��d1o�X������ފ�#�|�@,���+�Aۍ&�]vJMR�Xa�j�eM%�9��f��g�4�g�1��+��Ɏ�y &.�L�kF,����z�H��}�0��)�*T��6#<ni=W��B@�<Ôٛ�T�P�{�f�Z����=�o|`ک�(��qO߸8rnp�:�kZ)�"�u����T5���h�W�c]�Bhέ��WА�>�[-�z��p�Ec�H��O,#�]K�ōu|��Zټ%{�W#;��2J{a~�n�	�3�2|6��'�[���"�Z[�y�2� �i{sg�Fc+�(i4X���c��k�-^̙���3t�k]��Ւ�L�_��\6��NV��]�1)sâ�L~l����	�t=.�����Z��6X�Y{Ff����,%�@�i6D��Ϗ�|苵���,��⻼�m�)�N�Hsc84b��T�g�P�����E�.T񵾚-��H�nJ\��g֥ڶ�mk7���e��v�7u�?9�z{���y�ǎ��>�����-v�ǥG V��f�q�84�V�n�h��٫�jv�)pC��	k^k��M�uW���)�k���'m�z�ύ1�����<Ⱦj��[]yzT�����ű���R��3`���~���:O�ʊ��&�h#����:�T���OY�N3��O문���[`d�G�Np����tV��W�L�u-pc�{55�mh���pԀ����a�1U���m3�jls�ٞ���,�����X�F��KF0��U�T:6���~���XT��|/���ώ?�����M���T����;���) ��Y7Tb���.�Ё����˷��� _pS�`���D���f��o���Z�QZgSPhLF�ז[oj�h0���̳�K5Ѡ�"XU��:��H���s�r�		���o�[ha���IZg�w�E��JMTW7|~o�{c��5!M�ubY"���.dHM��2�	��XQ�(k�fօ�S]�(},�c`��F�"��~{|��@q���۝..�/�َ8��7�I�3q]�[�� Z}:V�S6��9��n���^D<�-�
���!{ω��4s�cqX�)7�s�瀲�P��qŅ	�nX�<S2+�-v��68�(����0sg��;����&�����ιab<���Y	���3���3ִ�g�3�ÿ�) ��wgn1��|���-��>&nyx|U�ژ7��d.��n�(�� 2�����L���W� �q������w@�	R2�n�����_k(�j�,��ʞ���T���	
#�E:��lL�ϧ���5��8A��˦m�,Ȗ#L�W�������g�&��j@�,����a���qs��Z��u���6#�c1�tN6%�N����n}~�t����>�@�pV&\��{��Z/�no������AW�ō�$A���1b.����٘:�q��?�nR�cS�T�T������C�^m�|���o�R�;�% c�|��"%ۃWʂ��k��)Z�䎇�0)"u��頫�';���G���Kpr���V9^ S�)�d��6`:�� �lJ��P�ųU���ნ`��>��v.������2!�4�F�����:��~)�h'G`
���	0��`��[e�r�����M�i�앁=��z�[f���u [1o�����X"�:k����َ��jnW��XMH��~���lqj
���KX�̲v�]��-�}Mw_NaƩ�,��ړ�i��$�����Y+����y�B�o��֛�]l7�����Z�6�֍4��X6M�@9;`>f.g�\mu~qޤ���e��1b \m���7C$v1�+�
v�%�E��Λ;�
P/AZ�f����?y�]����^�{	�!��q�s��6�����j�mSF�cӯn�>\�+�ޡ[z`I(�
�;�H�c��>�Ċ}��3����0q0`�z�l���AeW�u�Y�:7g��Y��E�W��(�y��%a���.��l�3,�����$�˻��#�[����9ڙW������Ï�'p�&��c�涉���\���[Y<ZM�a;rm�9�]���\k�@Ju��^�SY�t�{�Ht<�.���yQ��X�SW%Bzȫ0TI�vHZAҨb+�>Wvy~�58�Y��&8,��L�Z�I������D��I� �m��Y�o��������.���FiY j=!�ǜ-�h��9ܠ ����*�[�n��B�u2���o���OT��Mg�c6V{��q�.������b�+ǿ|���=�(����/-�����u���ӥ�5�7��#b�w����E�.�Z�q~���7
�a cv[ �^c����9U�>�l�~U����\�e��Hu��2�OǢ�(u#̰�Z�X���"�LaNA�"�nQ<��LsSD7�?޴�w����}���85'�etL��tn�^�^�,O������lj`��%K����?(�;c�5�&
����7��\��m���{�͛��
��y��q9�#�-��+�-w�?m�?� dA��:G�����:�h�����;�c�N���������)����Y𼹔�f��@�EqC�V���l����2	�]rW�_1B�e�"���B=K���$�Ԑg �}8����5�>�Z�БCs���k㼾ylX^�F��k{e����-ݯ]�J�k1ٝ�����Y �>�l���&��AR������ײ��~�F޼/�������v�1hU�&�Y�IP��-�0)b<9��F@����\��B7�����O5Uy~Bx�͍��P�� n3���L:�f��XP9Y�$��l�#^��B�����2�6��8fo�´��1`)ͼ�:��"�ꟗ��|�/�;u2�q����^i3}�4Y��H�=�k��;}�4{�ar�:�ypkdTw8�&�=cS�ţ�zW VY�e�뼹O�
Ζ]ch9�#u����.�K����0�&3���΄(�q�`�,�V�E�XMcf��5@�>Cg�k��rI.,��bMI�õWF���ؠ�\cj� H����bc2�� ��\�i�ā����;��x��d�?]�&�lS�hm�2���� BX��MՒ᯳f��i5g��R���9��Z�({��l�,�<e���&6ɗ/_jB]�-e�6�'O��`y��=��.,c</�HZ�����f����zw:~�g�
���y��c���6���^y,%0.�N�����c��M�?8��[�O����kv�]�T�ْqkٲ��_��sON��ꋕ��9���{eR4�OĊl�Y��p�;�q��bS�9��v}�A�3����9*�1#���&�O�]/s�k���d����g߼}����ؤL/�sQ@�~<�ԓ,`�ѣ��@kO�C��r�To���i����s]S4{B�x�=���nS���0=�rd;���g�����ُHh�`V�b�+g�V���,�bUP�0�]�h�S���lb�3gc��?��VޢڗZP���kZ�������9���h�J�u��Ie��0����Fϻ�����'5cդ��o(���4�P.��G��	��<�%�'���(���sF��oǢ67lW�����_y����wi��-Y6`����A�E�������A��� /q9��[��x|w3爵���Y��V��x@Q��X1��AL2Qxw�ܒH�j|>�{��,�M-���Mҥ��l�fu��ߜ�p0�.2XkeS���a��`�o
�Vn����b^��`\O��$�]�a&*^�!o��Zh��2�8�x�L��N��`Th��j��Yr�~�x�G��~�Z}����(�@�M��yҬ/��ل�3���?ʯ����
�w_�������q��H�ک�M�~�u2g���;'�u�G��ǀ׃�q���r���}��i��>{�L���[��(��J�`a�FLf1pu���p��.�ܸ����+�_�Z��c>N��u��j,�1=
}���//�y�,,|���9c�Ԅ��c]��i�\�߬ɺW�͘�;�����ܬ�.	 �ӆ����=�@�_��1��;X�	Έ1����s�o��_˸yR^@��$b�z�����Ys�kNlߞbX���
�ؤ4�(c��>�zP��w0�(�<�:�(��������Ok+Z�&3��u���'��>�sy�19;��~60���XNj�� �x�5�*pG�ǁ�T��b�s�PR�n�=���{g�}��9D�S$��}� v+k��ط��؇&f�Oj��u�hxL������ݏs�94<��O4 �
���t��κ$Ꭾ�G�4��@,[��ν��XG��<�/n���e���r:�4�x�?�A����Q�~:x��|}j��>X�w���	�l�Y0<��5fW����ٶ��7X����.6xݨS:jI�EY�+�Y�٫��n��rD�,��V&���X3Ѿ��+[�	�3W��u�6�ƹ�uh�w�Q��k#��tb`���$����f�z�Ru�4�����e�l��h�h*�b�������^��W��ǟ~�������>�&ֺ2��z����좴Mr�3�ؼDB<S��Uيi��j�z9'�#l�0]�o��`��A�o�Q��J˹�Z���q�q��n�r������q��}�8h�w
.�׽�P������9��O?�,��?��_�H��� �J7eM���M�3 cVj��1��m��K��8�M��D�a�hƠg�ec�B �k��FdVu�Z����L)X��ke����{e�4�zM��ǿ�V�bn��k��v,�rm/�=2~Y��|NG��h�S�h���Y<�+�u��D,n�)�;r����S�����q?���پѧ�&��I� �3�c"cO��Q571e��!Y	4�gBQ担[H;�*���hkiƶ���!g�j,�+�kq�r{s����7a�`D�9�����t��9�j��5`�C�x����k4X,�-���n�0ϓ6�M��b_��|��=ӧ!�j�4 ܞ��|F���tqp?n�٤��a�N���}� O�V�r��m������{Q~���׌�q��7«��e  fڧꎈ,L����5�S�x�4YMJ�D$L:[PP�p��� 25h~U�Q ���P�	��S�ng��^��tkݻv�׭Cs����6IP�:/Ȏ F�����
�{W6!�j�Ň }ַ�����5;���|<�7��I��a�,~�ş�/(��`�Q-.���/�ʿ���-����(�z���2�E<��z#�
 ��.�z��ʋ��� �{0b����q�LW��4�e^��Ҋ�81�t��^]�q�a[]�϶����E�%ܙ������!؛-X�����#�>�e��|ܮ��c	�����ڱ)$��;p�5��3�?�ǟ������?�8Ѡ�ɅR7p	�������&m��!krCb�
v��)U'�H�<�р���U�����_���F�� ��t�z� ���?�/�Oe��������^���0����`��h,%*>���?npd7�m��d3�p��#�3F)4�<Dcb��M��Le�D��CV�J�ΣW�0�F�����ݴ�yEk8�-���c�g�xda
��Lם'9Ѐ� �n����@k��Bg�a�il-��!j��\�V���'Jy��p =q.�'p�!�}�N��&cb�����I�����(Ӟ�Z��t|5�F۩]���+����4{��}w�۸�ja6������4tU_��蒦����Y6b��U��|������q�Я%N$u�������������Jj��߰6�/��n���C�Ԋ��c�r��V�������xJ���7ަ^�?i��l�>ũ�4m�R��rvyj����c�s��X�hc��Q��.DT������E�x]�EY�QC��q�����۝\l��.v^����re?(R�)�^u�������c�36d��J׋�b�p�0 b���F���O�����/��"Ƈ��k�)YEɐ��/��"���:H���ђ��ް8�ZQKh�M�3��J���&q���z����n�gϞ*3�/�����;Y��25}�dc�q7�t�/�.���>���:��;��~����w�wTȨؚ�x��bv�m˦�������o򺌛��u1Gg�;�A�둷�c~
�=/�� ��ϔ9��d�Vط�[�Z���o�Xo"�0P�~R�
�#�{F2	�s����B��kӺ�y��Yw����5��]�]�}u�2���� v�9�K.�@�n�
Z`p��]m�u�,'+?Ĺ�ڐu�W����q���������)�@�{�Ѥ�H5��^?�LAKhKpFN&����l�Ρ~�6#L��
n���0�ִnfX����U�.�rr�?����7����5�fB�I+ؘ$�fA�;���:�d�8|M����O9��f�H��cb;��B	"���8@[N��L�)^������^�Iy�����m'ir��u�I�z����	�7�'\tq��k�k��rZק�6�d]�aUim�5�w�A��][%V�?ʱB����:��v%P0;j=6�6�� �4��-)n�}ǎ�E����)Y�}N^4��ky���e�Z�i %,ta�2KL}yy��+�}P��`{����d�%�:_�gQ�uGa�[d�����i�	��@��T�7,O���n`�������|x;���Z�=y�� p�+^��OM��.�[C4����$�q� 6V����_dqbG)d��^V�J7���w�n���M~y�k�䶪��4��=����6Ǧv�g檌~TW��\�Y�]ͧ������2�e�9�an���S��]����ȶ�aTN���7����ט��WZ��� �J���NZ5�׬M���ԾH�e�^��MG;���������P9�צ�=�r��;\�8�z���>� [�������W�p}C�>�XW�>�O���L*	c0��8�e�௹G�_���׶�1��X�s#�����$6��V���k t���?�߿�q2�Y�r���{1\����!��g,�!���o��oS��L�������-_?��s���g�W��W}��zUֽ�����J�X�C1���q�'�t�?�ud�2E#�»�VZ�'���T�'i�)����1l�n�nλ���{E�e�V��ޔ ��hQ�f�|����jRρ��=E�CV&��Gyo?1����g�3d����NA',�UiGT��ݵ�z�A���e�Bx��fȫ���ƿ�������j˕�� =E��T��m�=��Db� �kve�߿{S���\^�=pM�a=ib��Ī�ʀjU��ݐ�:�g�������MM�&�*@�z��h�1`�c��_�m)��J-R���yf����?�u�OuNl� `����;p�|��ɏ�f	��j^~�onvǩ�W��3ˏ e��5����8���������S|Ӵ�Zb�������n-�H����â��q=����e��>�A'"&'Y~Y� ^���b՟G��oood[,@lΡ�m��h
 vFU~�T��P|�%�R.�@L´�G�.L�o J�(>p�H�TkhJ�O�ڏ-��k62�R�{B�f/���˗�
�zU�d�������nv��|xr�d����`ngtk5:̭D�T�����31�g6D��]�R�=�Υ@��I#��d(��H��DL\�=����˳[ٔES��&��k0�F�%�ԀfY�_.��j��y;�����(L�;LO,@B7�����T
a�^��X��k'*11�k���M F�ag1�}_�Q�9�9�������zƒ�[�0m��u
C�4C���� ��Ÿ���֝Ʒ��o�( �J.�/5�l$Z&O�Ɍ�u&Ƕ�&��KPY����u޵��|�N��/�D̮�	0d,��
�b#�(���wM����9�G~VAaY77�Ju(wqJ����&X�:�=�w�Y��+�,�s��XЉ��!=�	eb�g�P�\���+��Jt��d�6E�)� S�OA��P����>ȯo�I���*B���)�Lݤ�L��~w�PWjߙ@�Y���;t�|�����	%
�ȧ����
����*�=�6(��Y��XPO�]e/,{b��a͵ԭ$�Eb�����?o���U����Iw�iD܀���������*����E�	�� ��x�~e&�
��-$o[{*?�l�6kOn�?�3�8���B�3U���f����={�ӐⱈJ�+[���{k�������Go��s�~���
�:�7��6�Cyu���8-��RL��Xݐ���6��	�ZN�/1�w������� ���0��V��'[$��j���q�nM��:����;�����A�����۷o�}�ԭ�K0�5&05`���06��ț�{Zz���Բ?��̥AK*7O�E����%�������$x&<;2����1���e��f�G2�<;�-]�K�澮�'�ݮQ�]��Ygr"|q����ⵯ9IɀN�;���_�c��q"ܘ#3���8�
��� �awݙ�?���TW�yV�p;�o�s�x5lX�F������y2�H\3�k͢��lk��A~��'9?��/��O0��W��y-����z{���{�#VϪ����L(�����9�1�j
x��L��W����́-����RV�[ n���<F����L�\eͨ)�!
}���2��}�vA���\̐�������,i
.Q���j.�b��4�@L��yf���Ԯ����Y������m�R-'�Y�+H�L�`i��ʯ�ޖ�*d��@��pa�E{��;��T��ݭ��C.t(�ꀶ�e�*������Hcv��Je))q�k� �Պ�{��wF8X|���y₁�2.4i/3��_WÖӐ�|g��\�rbweA}\�1dGp&�uȜҋ��M�%4�1/t�T)� ~n"3�%6�I���|s�I�L�Լ꯸��ɉ�~/t�D�_cSZe~f�Uf�K�XU�ѣż)�3�ul��?�\�R,���"ă���.���)1#G]�L�@��+�# ��$,�{Fbo�bk9[3^Le*�%(kv��ָ�����υ!ن���eJfm�=o������O8��/D�l�b��R�4�MwQ�\lsM�x��\�&P/˴x�ǎ5����.��{<Rn�����
m�W�<g�=����:�<��;`���{�q�^�����jDH;o~{n�3�?������qp�lv�S�w@W81�����={&��ql�oK[���
�@�p(��g$[�b���5J�.Z����� ��	Su%Z���h�s�����6YS+�ӵf8���q X/��C���Z�k݇q63H��k��G�w�M77�Xe2��q��5�AD���J�;��e��PJ����F\�(h0���ט�Z�FOR�7fM�鶸���ke�ih�^i�в�&��bȊɜ`/�,�_fV|<���ce�*�Q�ѩ�7��Fv� 5���L���3�����ܝ2Jh���"e_y��F^�� ����&�z�t\{��^�u4Z r��ps����\:$ٵ��v{|����0�6��@<t٧n�a������V���-r�,8(�OS��d���]f%���}����s p�/3�-t¬$=~�x���~��X�0��gȨ1W�Q����~%|"s{���לd�:��K���?����kL!��q3N���;( ��g�n�u�>i�	���Y�q2���=G�h���nnc�`_,��N/���܊���O��(o���g=GꃩNX��{pY��rW,�ҩ���[��\��젰f�9U,f��|Xn�)_�~��n&�e�j�m�L�ѩ�׫W��s%q/����m���A4��}F�AZB�c�3�, �T�f�깣�{��lc��i^������xg��Z��"J�k��| ��Os<����l|K���ZͤO��??��9���|��~�3(��.�K��k�(��w0��5���:3���&㼱�Y���-�We3�Ή��������<c�>u�71�:�����[g�5����A�����ھ
<�wt�d���G��ъS^r������U�E��G��<�|�Ϣi���2;�*� ��[���7y�⛙�?4��ϟ�����E�Mͦݷ&�#���}g�s�3��Av$X�KY��+���2dJC�ƒ�t#�v,N����\U���!�Wb�Gu�)�a�]�m-0Y�c4Ǧ�>M�Q�H�6�BQ7x�m�E��V�ge'lCh�VU�������wW�i�7w���S>X����=w&�ÌP�c��Һ<۶<���/eU@���i,��:ז��=#�W8p���5[�=[y"���n˺�V�uq~N��L�q���lRx��E����V&�+�����^������J�Q����+��u��c��5-�I�*�����j����U��l��-F4vp�q�ݠ��3h)y�`���`�n����XA���gQ��p|�-�A�����|tʃ�j�3ic�����ڗ� �k�h��k�T{���Q�o�£k�G���Hq���x�T꘎ޛ0�i����l���B�oo���\�pj6����4$d5Z�c2�/�M���b�B�B�/;���,$�}�z�� m���ۊc7�U�T��s�d��1^��ZV����ߛ�8#���3���|J�xr��?�F[�Eg�d�ۻFBa~�s���]'䧵��S��C���S����.^��{��4믏�7�*��l�6�ǽm�:4�ԇ6�a�ծ�-�[��)��K�R���{�DI]�s6A�؜M]�}O�����1P�X�X�nz&l|(��4T�o��[������`�u����W �Ճ��ￓ���*l�����&<xx%�����_^�*o?��Ͷ��^K�L$��f��2S!4 -`eE�ziL�sݨ�iRU�j�bi�Z�5��xʝWfɪ@�+��I�Z`6ΰ�gj����:�������܎���Ì���P�%���6���ǟ�����x�H�$���a��U"�c��7Z=D�ט�5l�Ȃx�Y���]��Bi���4>{���5?�9OG�xb��@%s�{�Kc�2]� `�A"rڕs�P����4��濞 �a�8��x�Ն= ڱ��Ju�q��6�;}�m�ԓҡS,�Z� �0v���-�y��l�˕erW`G���V2����uAIl�Q�#����t� ̩�vW��Ǝ��%$>��٬Rc54��G�!� ��@��}�]x{�8!C�X`�>ܰ����9��lOw۰Y�������@/X�m�������@��2E3Xֺ���uaNdyt��)�+�n%�*�[��ܯ������hFdu�j�v��}q֡9�a�:bѱ�X �[K�#\%�q��}�ȅ�\�u��,K������4j��p�t7�̍����@J�{i�����D�}s�}ґO��G:��r�s�u���5(]l3�e���H��)��k2�X����s��e�IɌNϮ��'7�[rus��q<s6c�x� 2����y�e��\Ǹg���|i���n^�����ӹ���:��HPoN�6��>T S�m���o��v)/^<��~y)��O����� �;Q�V��x�̕�w�' u����� �aB��I݅ʚN��A2����`T�s j�Ig�0:�0��Ѡ�3k2��gԸ>sGj]L+*�IB�I�������չ��m5܌1Wx�����qn�K���?�E����� v!�$2�n��M渴���������;y���\^=* �t��S3.#x�L:(�-�����Z��=��/<����$�W�5q6��Z��SZRX�y�ve��i8��m�Dm�X�R�R6<�tH���6���o�1՟��k��j�_����ذ�� O͞�o��|��|�&���I�U�����EL���fY���P�ȁe�$S��%��s�-��&�fюE:7W�������Et�b��_�_N��;~�SLLA�if͚���U�����!�Ej�j�ZG41�T��k�|m�|��j椺�:���X��E��-�����1E�����ޘU������vG,�-���qf�f���S����i7�vc�{s�C����7��s\+����hA�8s��ud僥���x�܃e災� 䚬3_���ɗ��;;���1V-�w���*K�ޒQ<�{�[YF�-Y�%��_���F�!R��IMuw%A�3`n�E��1�+K���:���f�˳y�*k���fJ� ��I˰��'ҬSȸ�ì��>#�6{wf�~�1��b\N�� ���᚝�����؝�&�����&�@�P�rq�Vuw���%����\[�0^��Q��
�4�/��+���)Y�^�Ϯ/{�����<����9�������xgIL�a� ,!���t�R��X�f�za�����p'+��j�0�H7�S��^��/�^���Y��y�`S��drD�'C7-�����o����
^&��a�ֺǩgȐ�jHh_-۵ոdx2�no�`?:+�d��,�x��T �f� ?�q�+���S= ����مf�zazaֲF��讖׉y�����p�	�zNt9�;R}RSD�[��c�@����+y+g�qϯF���Hkq!�g���5���������e���f�����\���6�)s��>_���dN�A�A9x�����!��lI*��r�����ә����&5+=�4E�3=��.G������ż�/��|wwS��ڔ����+��z��:q�nX�l�VqO{�\�5k��'a`��H��WY��B���mai�*������Mh�������EQ���,�����"���6���g�k�Z ��fЦ��s��sч� Q�5���^|�U����̯��)G�t>۲4��^��i�^2`K v߽�|���Ɖ&�f�����_�e���Y��P������>f��5kK���Z���KY�K53�e���Ml�kEf	�������R���_�,�r��H_4{�Z���k�h$Ea��H�GZP8) Ҁ�1��n����@��&�QCl��;f6Ȕc}{py.?|��#ă��pm �I����;K����3f�o���1�vRF���b�X��fXە@'��J�Z��JeDC"t۴��JT0&�;��hLXg1��1���נ�\p����ȶ�M�Sͬ��]��#�J�������]����{Y�]��Kq�I�^��Qvw
�x_~|p��
�V����Z]�n0����͵��o�dT�7W��e���!��D����4�)�l}�&�Q?�Zx��T�ݭ��7�F�Tί�w�6Vs(�r9*��V������1�^SV�rE��r���#�K�����S���V�U�N���Mi��jc*�5nb>3����3q����D���%S#LP��@�0f.bΈٽf�F��y�K�����n'��.A�rS�@4- ]2x9�vT�H$U��i��H0�1's"���*��Y���Tip�,w��9S��S4�/�E���+y��J���c� S�n� ���F�%��۹��E���'��pT���\�~�M[JS�+��.�`%�X�~^���|s�8���a'*���I\'>+����Í �o�]��6�S�_͆� ���/�o*��ʳ���.3X�m�Ά��D���>0�a����w ��a}.5����$�T��Uz�c�
-��c�݋����O�g��<��-�}�}J��2^
�l����#=ݾ��G]�����{V��L��^ЀP�'�
S�fƺ�������ɔ�{�c�ǵ��#����z�|SֶGT���Wo��~��$����_F��x�L&���΋��Iu�^"��ہeq ��C�!+3�"��]�u8p��������~ػ�9����9�N�������L��]T4��P��WW���n�����s'��<P0tu�+�W^k���V�q��?ww]@Ν|x70� �S�����Iդ2�O���F�@��y� n�����Fw��A��f��/�k�,�rHdQ�'2�r�"��희n����FCy�����X����Z���u8��� ���0a��g�M`���|Æ�ŭ���>d�A�N@��uv~�@?~�V�o�R��ȱ�P0*@���B��������y�
�yftf��s����Jn�+�P�"��Eyy�Jp �,3�Z�͋��jyX`�][���v3]Z�:S����������Y�Z���M#le�&�5���kn݋2������O�+��Bٰ�����%�󵾠�;*�酫�-80ik�h��v��:G}v�f��1<��)n˕���q @���sK�W�)6�|-㾖�_��I���X�e2W�k�N}͂tP8Z��9��ߴN�O�hs��{�����1�3�N��#hg֩�h�;z�i��LL�;�Uŉdø����`q��F�ٻ�u�@a`ucĵ��c��ƒ���Hn�vc�rn�6���;�-�wr�/��&=%�%,�~���8nޗ^� �l�Ȋ�o$�0K�}��t��ݪ���+#N�b�������NY�����Do�� v��9Y��({����r!{� �q��d�k���k"C7�˸Q43]��������,U�;�uk�h�aġ.�Zc�����;��!6�\L7{����'����h.��EO5�/��F�d��\����W�Ϭ�{��%�@���|�* ��(~���low��=��ԥ�W�$���:�vO���u<�O�<~$>�+�J>����g��d���f4��C=/�~8G�Y��f�1��:�(;nм�7o_k,���5��6�
HF�ӊ����ᱪ/c�j��P�e��T��=���mz��f�0�Q&՘�'�E|�q���<����twsS�إ�Qg����ks���5�T�[ƥ�_���EM�� iM'�	2v�xt��]8�R��S����&�zX�О�I�f,�ؐ���tz��k�F� l���LR�Y��MN�U�jݳ[��j�y=Ic ����rV#Y����Oe�<���Z޾����4����Q��IU�K�^�8{�Յ�K�9�m7���\�wN�s��?��k�u4}/�����ڲ^n(J��ʑ�i�Y��Շ<I|/[���25V��୏\�}>|a�~��Ɂ�|%�}��4NN�k�pr?��o�[^��@\=w��ԲBs���}L�kЀ�1�㫛�x��z�P��^����P�L��:�����E����0�`~7+x�-�q�F8j��>l�F�}#��?���ǲ�r����k��,bw9�M�@ri/��0��F$O��ը�P�gp�
c�����o���a�W�_ˇk��qM5iFû��WǲE�"M���@q���J:�\����hF��:�7�[|N�|i�B��yn,<b ���\@T�Zc&3"���g��TV(���){�#�9���T���[y�v+��/�_��W�J���/�?Y�6Z�]h�x;�YF�'ȁl�K��;
���������5�a����ۺ<���!/3j%������e�<�J��g %�����qO� `�y>��
�z{�
��M�!S�d��L�H�`i�����4��i��}������a�I}S��*����Yf ��퍼~�����Ս,أG���ӧ�������NLE� ߩ;�@�4>	�J�`]��a=�����Id���ڐ�N>�F��BW��8�2��]���r�e��AR����js��$�@���:5�(��`���tl�����3�V�ֲ���B�W�8jm�$h�� 6���A�����D`Fdo1�Ĳ8}�W����#���n��A,6�/:�l�~��0^sWc ��v#�M�eI��>aUγ�B�KǛm�
�j)!o/�l<�0'_��<~��J��f��!`�lP*�{qa�����.6�ʬ5��>L���� ̦NZ�S���k����#.w8��������WZ�)'���,&� �� �����|�pKX��>n]�)yܗ���V�%���	E�X��7�۬E��������
݅{���m�_ggT+�f��r;����;@��ր
��L�2�5k����e�p-@�/��B��c�j:�U������G�w�Ғ<�Λ� ��@�\�#�UΏX��v��0�X��de~h�=A!���M�C��Ί��c"X�8��۽�n��MoN��j��dL�߻F��-�:�ćN���r��§Cw!�ۃ��?~.@�Nk���V��ۧ���$�X3��*m��������f�3Fu��C6j���UxXz�SB�Z	#�k�
�z<�c�������ƈ_3;E��K�� � �c/�q]�O"���������Ъ����%�݂��.A4�����Ϡ 1@��p(�3b�0U�d�R5F���2�h�`cڱH�������K7�.������k�������;T�y����\��,�h�,S��P*x�#@����8��|K��c6[GâL]k7S3��{�[�M����k:�8�?�]���dV����-���o�j����=�:�'�.��9+����Z3OԷ^�Ϭ��;�fXj���-�I��i�_��{�����1�~hj����ז���Z0\v�d���G�:�F���rN���^Z�>�1i�v��.ZM���M�:�`���: ��b=�X�Qn�"���{�>k���y���}�N)��̌-�@�1/�h�o�2`�}�����S��E�I���?��'&���/&"��G��ɏ:mL��k�cԢ���|�]�M=��c��u����b�H�:O_������z��NqoL���πx�~`�[uUu��{�aOɃ��M��s�F���ˋ3�}V@���\&�LTZRƫ�d�rLpH���h�rC	;�h�-��x�d(}�Γ�Āsc5���	b�2��J�r��0ۗ(S!�txֶΔ��K��y�R1H�3I��u�-�~s[�F~W@�O����y�P.��]��Fg��*���a|�9�q���|����F��W�ѹ�������p�ՠi�r�͌����lb㼴a�u['sÚ����>�$	�xn����S7&����Z�-2�����y��1��A3�~*��S}&�#]�d�)ƺ0y�v��2F9X#��,G�S(�>�M������1c��w���k���M�=Ǧ���^�e�Ym�nd�w�
�s:�&�wP�CLrd<����|�9��ģ���N�E��iT�~�v�>^E�(��_xU��T$�U�fe�����
g���;]k3��^S��ҡl�+y�������<;y��\x/�߽��
��x�a�ζ�����`9��&^�h���>�h;�m�d@�b]��GVo_Y(��g�-��8���������1�cd���h�(�@`!�o�(��Q�6;��H�kcI������:;�X�<����ysnƻ����{���J��#�	�:'���@���(eϨ
�k0VT���N�[ք�������cşi�;�4i6���ə��藦�ڠ��Rg��{��h{�-Y��J��#2K���sp���w��ka�8C�hud�~��6���:����TVdf��6-0�q�Z�Ę���ު�8���1[~78��/<N�*%���c�F���Ж@s�0�;�p��0��Њ�I�bh��LB��4���	�/_<��n���\��LUo{{v����φh$��1��$D��9t}v!�7�?��u��]�A���>�H�X����06D�)V|/d�!��(^@�(;&�7�
����,}��u?X�뎮��~Cx7-���o��l��o��Voz��-����������M<�*�Uʇ��2y�Ɋ�,e�R��&�l���:d! <Q1��2�?�0֌\˖� �F}Q�{ %$ʙLE��d�{����w77�^���]N�4�ݼ v���ߌ��>!ca�ٍ�1��N�5����bŬ'��Ы)�7{�j4r�pT�olFm]��=ۜ��x� �Tpehe�ެDp۾y.�4����6���<4a�	�~6/qJH����\�\��<ͽ(Y ���FR�=R+u��_}1K-�k��dN �G``y}*��b/�l�)���;U�ŪFĞ��_~N�� ���R��L�}�8��^U�!��[8���Ǟ�r�a�6�����a���ň���s��* y���Bx�Æt� ª�R�!.%��,h^@^��*8���"5�� t� sz�Y10�|��Zް��!�_Kb"v�����@|�\�P�a���_z����ծŊ[�뙴�bEW8 (N����-��^��n��%@Vf����W�(H$m�BTP�H$�o6�70�ˤ�ܟ4��)�̙�;�۸ʣO�yɏ�*�rU���^ ���=����Js3j���C���u�h�P}yAW��t{��B3��^�|��'J$�W�|����
)�:XJA����{��&k���̡�r �l���F����}p�a� �ڬ���a�UJ��1��>���9���;����|�1�G����(� �r�@�[}�{�p����^�/����۪`Lzh��i�X�0�#b���Q�TT�cO�6v/��`����X��(�3��k��[����E���Ю��yn>������޼���+�'qL�}�m8�����3q^0���((�}���I�V���)��Q�sk�@*@�T�#5���fUA���Z�`���\����yZ��>Y�9� 񘊷��J,<�\S� _������$wsa��\'#%��X��!��˹u�$�E��/����?��l�q���P�镢�,��;�J�4	!��Щ���W�<��>G_~�)}��]��ɼ2����a�H�tqq%c/䟆��^��7�/������U��2�p8����@��ɫ�̋@fX�{�㈜-�M��_׺MqRi"��~4���a�Px��j����NJu@qՅb�U����C����;�Y$KD��ի���'�����`ȸ�N-�yN	ζXOyO)�_2�X�O����1���=��	`��Z�3��O>��no����^sy�s���'�CuC$�0�S�q�舯9!��
�щN��!����Y�M�R����B�;H>�*Y5��u4w��W�yM���f
�dLu�*a4Ʀ5�_���b��	b��Ψ�'o�̯� �<�hd��*�Z���&L７yi�VOƀegQ�"�?�لB�Ǜ��Mٸ^���uĹYFN �电��U\���n�]���5�j�_�ni�J��<d��B�Yà2��S�$�K���y'���j0J4)�a�ȠVQ.M�"���g��;N����,���;z���>��}��s����O_��l��8����q�v���n�"j��i@nZ����
��A>Eyʨ*Xd�����<��k2������qC���^��r�{
jGI�G��68r�ە�aA�J���
�!5L�υ"d
����ԼeI�:S=H<�+$�����*^Ƭ��AK��� 0��RE��I����Q��@K۶���3�����H��ŐrZ� lF��a,xMV��Sx�Tl�s����MQ���%�����c �JV��yXϮ/�zA/�_�#�S8T%+�� �W@]�j�	���g,�e���ظϧ��Ͽ����������w4�>B�kK�R��A���6N�c��{�� �j�o%�<H�yJ�Y��nn���!�'�σ~�Uy�8�=9�~�)�|�B���c�p�������Tf�*	\���=/�qO��F��WAXﺎ{}���$�K���-�Un]���k������JΟ!tg�gJ�Ai��o:o{�{-��0�z.�5M�Kj���k�����h���1�8�k2�]�k_�WM��	W��sTK��O��O/
V�ZE����|���^��|������y]�C�(׼�J��A3:Oz9��r�pT� ��U�s���:�h3�A��ӜC�W��J�����u0O� 26�n�<8�/Sk>���@�s���϶��7�&�|�&�*D��D-�Z%n߸��߼��o?Лw����U{��z�L�l��B�_0 �WN�PXk	�r����&�Z�E� �hk�A��{�Ș-�|���O� ����4����~�wts�2Z.� �߽y��NBF�݃�4�]�x��~���Ӂ�W��~�\���އхQ��`L#��Z݃��L���������D�B���M#Ӂ�bA�r� IeF�����G���3 Z�e��`��2�u(2�t����-�ͬ���P;~�" �k�A(?+��~�]x�������*B�̩ƍU_�xFϟ_J����B'"T�8����������5Q*�י�$�(a�0sC��}�����:����o7Z"�U𳱷�����͗��t� LvKQ+��Wfc��k��]��K{�U�j}�(*f�	�P{jte�>}���o�\$_
�^�?��?�?��?H�s �̖'2�5\VoZ���}�>2���^��	�S�|o��:qO�$���ޑP!}p�ëW��y���~K?��Z��xN���߫U��T95D���&���#y�v]N�9�=�$g�+*)�|�y�'�C��X�{��K�O��:�@֊�8�\x�2��{�]��œ���q�����Z~m�.u��]f]H��*��Şi�3΃�\0��E@��l��U�b�Ѥ�A��/�����s��S�t=dOϨ$�KK�:W#Yզ٪��{�ϷF����y^��i��E0����֐&
�%�C˴qް�2�ǹ�R�^�p�m��?DUx̍�(�Q&�i�'a/8h�$�}���NX�z8���{�p���_~�����.�G)���n�H3ҊFXg���e��K[éW�F���@��s�D;��Q�c�������h3��w8��u�~�K2gN3 �?<HK������ƀ��(��W�]��_b�1P��6�ݑ�T�B������� P�>��k��ox?�m@��j��/��&j��Q1t��8�'؊/q��`��gF�(=2 c�x�J�[4��M_]瞘X��@��z�Y�M��&�SP@��i�+(?����m��ۈ�1^>���/�%�=T͏�0��2��A��� 4ϵr��x��J�Jy�>�(��l�M���M!� :Hz����1x ��U�q��R�EH�mW�Rݻ4A�O�Ϟ�i�Q_ ��ԠХ
���G��^�eOק�~F���o�����_j����bG����� ��J�!��<������Ŧj��[���R��G�Đ��	U�&os#n�~������%�4�	`%��}�
���N�U{��<�W�T�E�����`� ��9~9Hji�S����7�M�}��[ȑm���7�/�-ɥr���ze��Q�Rd%�lF�' U������ū��u��#��UL���������3cgp�k����[�j;�! �T�qJ�ѨDYUK�iV� l����?#W�Y��t3`����-�YG%g��%g#9����ʚ�j�'tu2`����ż�I�[�$	G��#-:�4�C34ճ�Md�R�8�� .���  �ӒX>� )Z�Z	"7<tv_	��ָ7�s� ���⸤�RP�@��5���Ò�vg�7���pg4l:(+a�`6ʂ9c��� ��9�©�mS��*s�~����6W�ϭ̥�w�VpL��$%}G��pZQ 0�O1%��&��g_�N+�40UV���M=9�`�����0�{�M֭�/v��VJ�˰�A�/PJ�1ZȎ$�l8Z(�|��)�qK֥y N��c�<?>Cٻ���G�s�"�|y6J�য়<� ��6)Ը�b7q��ä���z�¢0PfL�n-�l�#��@8{��X+������J��H�y�L���L�)����濻�6���0{M1 c7.[᧲Ji������	�g��j�~����O�W�>/��nWWW,���D��g��׿�/��B���@�+�u�i�`k�h67V���B��Ǡ*���-Ч��c^��̞��^k���)���!���!����^�����N�	�x�[G��`�?	����x-�A��'<�,�ʤd������Sn�5�Z�mW�j:{�a��m>��������sZ��9�d�������˫�����|�~x�9h���I���ݞ>����o�w���V��yUJd�šI'��Oi�/*�S.�σ�k�Vos�$])�pq��Cѓ��)x�&S97�����4HD:����ːs3$��Q!�� c*_���g `����V9=�[T�󱈗k ��Z���#�(�V�a�g����s�=�=	������|c��$ߣ=W�5�C���\��ԃ�5�����ӳV#q׎��ܶA��̈��|����Dٱ�o���'cfwf��M�(�E�վN����B�rI]�}pl�,C+��@�M%U����,����(��&6C9�
;e#��l��~F��I���Sn8�*I!W�����~,L��e��E����&���kzBLj�%<��s,��ڢ�Ž����'_���`�Ū;�~��J(�oNN�g��ų+���D����vg*޿������}��skGKA��ު�.�3���k��p��������`x%T��K��ڍCC
����5 ��֡/(>��;Kn���r	?��og#U��I�Wϱ0���s1P��˯x��1���.aGX�k �ILH�5����g��G��b6Nw
 ��h��~�ۂ��D&#�Խ���HU�<v�?���d���o�v��
V�~����xto��X���p#�"�s��>fk��m��� �X4�����Ǹ!�j5��8y�8Ο+EL
'�8�ބ����[h�}�g ��`�����8ɜp����ͣ	�S�b��6�)[�b��<ӣ�,�D�%#h���]C�K�N�A��Z֊5>����z8Vp��A /PϹҽO��#�g4����\N(�:۽�sQ���Ƌ�����@�-X�9C�#F�3�?';�������Njdp+:�;�8"���hƤ�KK�D�W�܍(*�!�(���4\�/�g�W�TUV�J��<�p�~��;c�� `��'�p!��qQ�4�Z�*�A�����O��ʠ뜆�%mΞ�������L��V��KX����R�	ax��T<��O���B\�,H�䥥���Sĝ*]P`
��`�}-t3��N�O�#�Aތ�[a�*�U�Q��Ę<a�{�Е F�9�ѱY*'6,�&�'N�}B���D�6���@q^l���������Й��p�邉Xϵ���o���޼}C�|�g	e���������}�"����T�^^��Kڝ��eXoy��������6��{�/��JϡUf�V���@�^*�A>���A�>-�����Hڄ��z�a���(�3��ʟ=R̰�7�1
�9�j�3	�]__�O�жF2.���U�����AL�81֧�)���\��T�������5x:�	3���5��N��Vq9U�^+"?�����ݕ�zFY��pC�߿��`��ڝ��97�_T��sR8�߳��{n�,ǪB���K��//�]l(�{x�-�%�cv� �bm��A���b;��+X��J�����~>?<� �q㜆����sΞp��>��oNH[��? h5�
x�ԙaCm�����(FZ��+"�tqh��)~�^�� �&��T	�1]fa�2	�f���|�eZ�1 �k��2.GK%1.B�J� �c�{���� ���fe*��sEn�C��3�Qp�����g�ϣ�MV�6���P!leM[g��I_�jI�M+�������֒���SE��][$�S*�s�������S ��_�5�r�g.
�d{��S�W�Y|���abB^9��i)ƾ�y���G�(ab�&��GA��A9r"\����^�����
G�$� 
 �ӂ5~���9�9�h[�=`��'�Ea�d
$>�ئG���JI!���Dv���lה�ɍZ���߇�u�*���@?�tK�o����n&B�؜$A��YI�Ɋ�J+Y�2b��uA;P�(�ZZ�����>�Z�K~�G�;*f�p���%����d��o�z���؅݅���}����������W��si�
�!�$ȫ�i,Ċ:�2�������*���Ri�`Ƞ��Z�8,�ǜѦYh�(�Q<�$��?���Rr�>�V\ϸ��6�UХd� _�pm��.����K�ZT��s�)�-��0��
vS�ݚ/�!��G@��8A{|��k���ս_8�GT@s�#��@8��={�߽{+�j�f0(������q�[���^
;��D���o��9��M����A�������d�!�^�%�{�k�A�S��Eֺt'@��y�p�d3`����k�`�F�v�����.��O�%o��A1�5@���D�3iG4Y�|F�*ya[��C:��H<"�(d2Ϗޫ��bt�U�CJ��vy��J$��
Fv t�]*@��ɳ�c��	6ɸX�H��,囿݋߰�[���=���[���g���e���a��Q�k�}>)�94m7�8�+D�s�ÝF���*R������#m��Y� �M�x����ߗ�M�>�m�qR70T�+�����VHA$��hy�cD�ћ�r<v�7����w?��;��}��I3-��S�PT�o1Ņ�Ő�qR%��JM���fɀ��l�`r�੒sۄU�l2���J����HLm�p�Kp�Ѫ>ɶ?;u� v��.��h$�6�i��뱗 H���!
���s��G��.BO��R9u/�7Wx媕GׅgQ�Au�V��9ʦ���J����;z�ʅ���ne���'����Zr�������篤[=~��fc��7��3�r��U�2Sr٫�ao��C�9A�ɱR�����+�bX���m�I%ǃ������x�_�W���yY\����2����"D�C����
��
B]�do��Du�*�����z��X\ٸ�cZR�O��S@�t2��1e�C������� �"���X��#w�|�z�«զiٳPA��BMG���/�͇[�����?|O����_��c��<���lNk�B�1��Pl&!�s�~QQո������|�wf���.�,�f��`J�>�?u9����Ez�ם���-Z�p)�T�U�8��Y�����hZ�?��fҊbai���t��͙T�1�fl�B�1�l�y_�f)?I�F�yZYƊ�m>H[ū��1������G"_��ߒ�6%�dk�Ĩ�nxf�ll?;5p��v��)��%�<o��?�֑3�d��C���YĤ	>��S�4t�0�vb����

)Y��	~"�nu
�P��)��VJ�I��=�Wr4�{&����F�fyM��) Ca�8��+�F:��sbkf�(�h?}�
lY͍@��R�Ęc [�~��ڐ���%�>P��:��EVK�� ���&���zl�Tk߱��⨣����/qɂ�U�ö�P����O���M�џ����ba������� -���[������K��|�ʺK�5`|D*��#Wyi����q{��o_ӛ7?�r`R����t�� ���+��w_�?���?��zv}���+�F̚&����i;�/Jc:��;Y�#�>���l� (�/��
�m�V|W���3N����G�SB�#���_��!L� ^k!s*���딧g	hs��|cy-���$�P�~~j��^W��g�c>ߏ>��@Xzߓ;6�Ҽ^i�a46:��Q�O-�^�3��� <Y�c/�*��춃����t�����{�u�k��}ʤt?��3����K�nz�������10.�I�� j����h��̺�k_a:�g/�<���޾yK����J��o�& �����h���y���7�LƐ)�2����k�p���Z\�'@����<{���EF���f�Q#�F�K�ٓ���6
$��,'�F�R���1�����-�E��B�Ej����cަ���6���:�?8X���Vq��Fhn�rx���$����Z�z�)<Cz���l&�淟���\`���{c����{��*Gx�t�=���\["�[����sܦ�z�S�(}o�A��F��T/����g#��f����᠀�O Ւ�2���Tx@����	�	��(�E@i����G���TuΩ/C3�{�?���x��c�}h�`��Mp5f2�qG�g�حp����i,���������e�/B��T�I�O�)�����E��A�3���qI4�v۳B����MW0���z��������7?ЎC+�ط�\�޾/����+����ě�?~�?���V+���7��n��x����)7:c�s��;Y� OZ��]	�7��k����#��^A�}��'�����G��%���3q�w5W'.����K^y-e@���58A�l���ầ<`k�������<ZO}���ɏ}�;��g�5dU�2���7��S�Ns��a��,zU�-��%��U�O��o: ��o��
K~������O��~��'?��e�x��S��H8.{O��;��A�%$'9j�=k��i��x-����С#�c��Y��`�������>V��Q�����~9���<n�A`�ۂW�
���PM1�dp4��KU�꫒y�s*
z��ig�)+�����߲��¡���p�]��>�H�]���uU�P����<�uPH؈��H��d0�*�"5�yR~Q��b:{�E ŝ����� i)�(9Z�����ߜ�?������5ĕ̈́}Қ��������w1�z��牣#G���3�y�( T�'�?�f����&���%/���B��������~_��7S�tws 新mH�v�k�t1��V���QeУ��HKv��~������xүZ����Qbg�DjvJ�v�Һel�Wc�Ee�S��e����W�� `��V��#�<	L>�ǔ<�'�( I<e����/���
e���ao�����Y�`j��t ����qG���������K�R� �������J^W�.��@�t?J��=�l{�s��jʛ��x5Q�oTk1�~���k���O����������mg�����޸��i�""(���(��=�{V�v��z�,�'��4�����=^�0�z��%<X���TK$)��wI�\��0^�x��B��W_�u�;��0�/�bG��r�K}���ȟ?��P��0��Rt\jo��\�����Q=�/Ι������ͷ߈�Q;��DB��{�y؋a����M��7����zl�F�@���A�\#�3i�L�%ט�]��Pm�f:�,��Y��ە W�)H���9���ޤ�&2Wss�joA����  r6`�2�K0V�80�+b�af0�+�B�2��X���Jx��8��+������7�/�{ �ꄸ�z�23��)Z�3X(r�0x#`���N?�	�D�0��A�=W�l�Ҭ̖�??��ü��A���ѧ��a�Ņf��Hp'Jzn%�ܷc|!�4������K"��/)� �1Ư��|=�?��}ɹ��[��8�l�6Q�
���>[k"��f^���/y�2WJ����_�,�����f�o��O^��q��yZ���%G�۩ty�=y�������������M��W��)�÷l���#�_�x�� ڥ,��~�)��Vfl�ٕ���x���d��RI�hH����s#�=�*(2������T?��l������-�'�źjI��W�ɾ���́;��ڹb���ɻ�"'N����- X	o�S!�_����K_���O-饧-���~d�V���#��`�m-�نp���D���k��D/���s�OW��ׯ߈熓�o,ɟ��c>Q�6�m���)#^��ʻ�=��˟�B
+�ј�@��+��n(�p�ҩH�\�3���[`>|�or��W\�͹y�f���_�8R�h0�K��8��ܫ���3�;�D����Tn��F�g�/E��8�H�SZ�|~�� f%T��s�ɔu3����7�fr� !�I�YaB�!/
+D#�����1ĺFU.�R�S�r�#	9���&`ĺ)^�Z@�P`���Ѹ6%_{�!��f�<U F��Z	�QK�.�!�{FIw�R^�L҇��kk�(�6nuS�>+ض2���l _�<�&^!��׶/,܏3��n�ƙ������LEq�|?���7����;����b�B+˷�� ������=���d&b�#>�) `��g.v!߫�� h@��a($�j���-*��40G%Νu^x/'#\��WŗA�F��
��S0���iP�����f��E"䴄�+�X \\TeO��s�!����&�V�%���i���$�s8෿����v[��RG���_�*���&�rLcE�y�.iN��'9U���Ek(T�82  �=������!'A�pwKS#����p�l�rͣ�:�5�
� .IЕX�-���x�{��+u�ﯟ'���'*?�)���|U&�h�i`�������_N=��֬�J�UI >� b�pO���o���'�n�4t���	e��rJ��<y� �"?99�1N&T�C�U�]��gtJs��^��CVs(!�.��t��^0dhUt)�VL4&	K;�)��h�B�<L���
PhwX�2��I����`�R=�G���5g��G�%}�9F�hfCI�FsіV`�����4���\'�o8L�������Ϸ�N��W!����������b�T��=��5�4�y���U�2s�S�UJs��r-"���	��V�s����3�!�"�6�V׏m�N�L���_���$��Tǋ~�FXz�M|g��ݞs�����Hx�bq��M���jij	Fϯ���'�C�\[JhkX��-欵�$�E^�8Z���eދ��!���})󳸀�5C�p��������}�j(�f:-��n_ x��6F��ȑW ,�	�dE���S��o��}pw����:pxF�W�'�c�p��X��E�m��n94B�:�s�[�������	�+���2�]����T���c��s'�%J�5���?�!�ɾM�#���*~�b����~�������#�#���ų<������YVW�Ņ��~Zc�G��G��H���v�����7�>���(h^N���y��%�
W�6��{ZQ��i^�䧎au�@��0�dtD����3�ꫯ��~�sι�8��B#�h(�%)(���l����`�����"}�\ə�U�5:�����Q�Nc?$��Wr��nE�K�����oݫ�H5�r�i>�%�%%k�_wH������Kօ�?i�fN7�ƾ��̖�L'�$Tu���3�G�S��[����w#���eT�" ��0����D㾢���D�3qNv� 9Ն2���ʐ	��b`�f�$g_�Ř�c��W�sq����ʲk��~�۲x�����)�n�����<ijls��f�s|'�?ht@��\��E �$o幒���;���*�N�$a�l�vS _6�d?��+�!�0pE�� ��#�6���N�V��H���$ ������8��b�:�7�z��p0��2&��c����:��ŻN�|����EN��b���ŕ�`�MI�l�5��Md��.W.k�v ����`^��ZW5%,�Мp�4�9����av�s���݃�dc3�Z}��a���ī-~,��p���%ݲ��T�U�?�O�2�a���!�O�R�Z����9_��ƭ����#SPHB��G��|n��q�i���$�E��q.<8f�䵗��c� =<��	Sx Wwtb:Kz�|��R��m��rh�g&M���!T���D\��M�-"5ؖ�?����`P�@����-漘�=���K�C�M+��\s����֞A�,�>����~&gc?(=�q�)���O�����<+ǥ�4=�/\�����>%�=3'�W��y�܀{�9ƔDL���ȸ	����e;���Y�� E�pLm�PEZ��wDU�����'��{�:@�ļ8�ftO���z�*��.d?�oŹ�q���XdIV�V1�<���/�L���c�/�@��r��&�%&{�I	��,`8Sx����Ț	���>F����m��ҷ�⿎m��vm���ޔ3��j��A���<wBR�`bz����'�����J0'���\K��T�����N(Kz�̾.�SC��qh1�����B�e��ԏE<�.�͛E���2)R.�9���%u��i�f��ܿ�P!Lhw3�@rEV#N��M��ToJ�	�<��I�N���E�F @����4�I
BYɒ'Π�=*+�j�ؒ��i�u�f]�qU�V�G��.����ܗns�1�%�����(&i+�:�yj�IHz�?Z)ޓypz�;�8�r��~)��%hē�Jm��@�J��bPE���m�=�w�  ��IDAT�/fq�`�&Q�4S/Y���� [�7p���HK�ܿ�_-�2�*�u���Yh?zAa��b!�Ņ�3�y<�0@ͣ�ԓ��a�y�}��f<m����t�8�lv��<GG�tj�5���C����� ��V�V��H���e,���h�3��WW��ó��5a�bc���ۆ�f���/����
���&��Z5�X��j��b��5+¦��qZ�'��>��]x��#y��#s�m�k�C�¸���o�Fǭ���`S��F�>�5x���P�5�U��������qVORQ1��")wO�P�aUʺ��k�ж��٨b��w�F�Dn�׃��7
�8x���֋�Lwȡ�A"�t�lTsG i4�є!mvn��4oN�����wN��K7Y�%�k��c��)�z�>s������?^V�;s0Nd�\1Y���

�����Ǆ���o�+:��e|2S���	h����U�K�#T���DW���w �@�j5�M���ȗA���L����Xh�0������kh}�s�������~��$U෎�Y��$�����%e{%/
��t�5���x ��4K�`[���Ul����D�KK�)-���3��7�l+���� �I�����`�����c���"m��ذm�5xT�G3y���j�Bk� ��&W@����&�uj������G���<D�E
7X�X;b�/��*�yv0�𲆥�HhB-f�*���z�-�A��IX�Ǐm��<�G�J����S����k �T,x�kX��1�<�)�N�\�[�Zs�$�2o��^��,G/hM�<Cn�2w+<���I
r1F�	(�|��E>g>C��������}A
����w�~{.� ��W?�)82OEq��K��ilD'4��#,�m��%�\)��������X�d���(.�+nU�4�������w��A�`[=�gGr�AU������R�,�N M��� �u=K�L�]q�9�B!sq=�ywƺP08� �����u^�}����8���H�����Dc6�6n��X82CUϏr��q�&?�L�C�s�9Ɯʺ�]z�K�J����L#c�����̋�(΃��Q����!�|��*��0��y�*E��YR��}J^�I���j�Օ2k�V��u�jS���J��t�(͗
	?��tS7��K���F�E/�f���dt��A[霟��7��;GpY)�=�Ż�j�Yd�O���N�2����.'=�4���h�˒�t� -�´o��5�0DE���O�d<��9,!�R����˸�u�.���_���޼���[�|��F�E�C00�b��(Nʯ�R�+����Em�C�haԻ[��Tt">��{(F>�����N �mFcヵ���4U��X���*s��M�җ͕�`������/�~�#:4賠3D�P'<�Rr�8�P�� 0�����"W'���[�k��4���z� 0�dE�w*�h��Uf���ٸ; 7�Ӆ�ϟ	y�$�^�z���.K!*R��I��ZS*�4ԣs���A�����i�ǅ��Z��S�2�Y�s�z�q`όQPQ`���gN=�н�+���_+�V��"7�� ����	!;���&Ş%N	�א;W,"�����?S+�b�T� =�X����a~ի��X�Kˮ��!Tj�QdT3�1U�d���5c㌻�G�� �WB�f��tUI��س[����쇹��.���M���<�os"��0�����y�T��o6�Er}/�Z�y�N5��v�~��Ѝ������-3#!q�\��97���5�Q�i˵��'dh������˟��|��U��X_LU5���r�7Ν�<=���ժ'���`fWD�+P�Y�Ӂ��9�����#����1h�g+ި�*��NBB���8X�ɲ�!m7����ϝ/%��x���AAW��C��d���Ô��Ά7�e ��%l�Ǔ�+@i��r1�b[4_�E�J!(�e�����J���e%�#𴤏�4�`з�[�X[�o���
`c.~f�>�� ���%&$�O�v0b_x:`sx���'��6�~�,����b#�����\T�!�8�hK�$7,�V��)n�-���;�zH`�Ew&���tQ�N�T`x�,n�c�}�<��ͩe�V�K13���	Q<g6F�Z����9l<�b��9۷�A#`$9?R�#�w�P���b�����!q�p^߇%M��&��fiά�����vaT�$3q��&R��Qr*��0��2y����fs�tLav#�T�&-'�ǈ,$c7+�(,
���?5�����L������h�J����Ώ6Z��B&rx2�J�F��¼�!��F�������} ��SR�*�I�K�E�K�ָ-���"�Es{6Fd�k���{�K>!����呴Ë%�o�8-.�6t�����|x+-���o��_~JWϥ��y����"f$|�^�Q����� l�#�3��ECe*n6@|l����q%�y9�_i\T7pW���S�c�)@ج�	�tcE��%$������>c�(����: �M�O(\ճOt\��Q���')ɵh�{bחX���+VΎ��6�:{ �":s�%�<�g��޴�&I����ч�����i��˗/���K3'ڻ;A��2Revd�d!:��}��ڲ�G���9%x�B-[�x���c�_j���_p�,�]�@�=�0��5��hӐ�~��[� �l�o\��p{���xB�G�O�}6&#����g;;N�vF�a�VO���OU�8��[p�L|�"��RQƳ6l� ŧ:X�-B;���V��ٹX��]�p>��QWw%�˿�%,�j�ǰ��9zsυq�	G��x��@�	��<.��r��+�jZ��MЋ�||m��-]��0s���[Fn֪'�'pF^Q�3݆Y����EEb�ߦ�̅U�B+�N`�P!�d��X�iΖр��ϴ8/@*U~���� ��X�5܇���]�d2�jՐI������,�'@��ax�g3��:��s'}d�s�p~.JW-։$���XjP�sCU�BZ����W��Ps�7�'M�߸g/b<�1����Rϴ�O�����5�:��n�I2u#tg�q!��j������dl�~�{��ha�d�����q�L�</�����i�����r�AX�&����w����þ���+���W��_��~���Au<���Gί-�(��/�_x�5S�Ƀ=�D��tA��A%���� b'^�#��L�KN��wj{�ɕ�VZIqJ�Єۍsȥ+Ar!���8�ԓ*撬�Ƽ�E3���S<a���$o=��`�g��PB��cT��Y�1�0���*��JF�OQ^����� �����ڷ{z�pG7�����A�g���.������� �o�yϔe�IiyM))����e�<G``���$P>�Trz����-��ɍ�)]���T�le���L�=]�ϱi�J��B��Jݠ�]&J|�����{�����3�W;����W�w�C��\7�� y/GM��V[_L.�W�b�ظ�=�՜Y����������s�8&dV��x �!0x�!�8U(`�W0wyI�iL��   ���Ѫ�๭���,�9#i|�� T��C�xW��=Ք�A
(�h� T��t^� �A�g�Њ!U��[-#or��m���l
�C�����/xB�8j�c�YA���
mR�L�ne�u
��p�I�s.�ѣ�=��	E���-�˥e����z��nR�w�u�ī,[�}�:!���z���'��4�v������hۨ�a��C�� 5bL�^>���R��u S<�	l��n��(0�Ii����=��%�Q#�J;��xq��3���t��@wo���?h�݃�TzvyI��@��q��f��{M�ꪆ���h�'<_�Y �����������ǜ�o��`����M,�o���C#��k�)����l(FV�Hk�d���N>"�[~��p�B`�dBXv���6�<�XVřv���;��"1��=�BXY5AJaG�
V�$�Zʮ�Ͷ���l����St�����n�����J_\_�5�>�z�O�����ݞ�����v���جn��K��\�%����T%����b�,�@����)�^�K+<OPs+D�ĝ��5t�=�I�f�W}��"|߿c��[������I������4�������/?�j˖��k��^#G��k���C$�*���A���b�����A��>c�M�,����Ԅ1^� ��F�Ph-=�r�๠�jP��;K�c��>

��Kq��T+AP��@1�y���n%B���E�vN�&�G{����߻����.Y�x�ve�	a���rc�D%�nn�J@��)��s�;`F+(IЮ��d��r~v��1����(�
���7�����=cq<�i��9�!<h�����F�Y��N��vN-��^��ϥՂ����sr�u\��o�vH*7�ۧ���6" k9�xxJ<i�64�kٗ��_?�����Y9�R���TR�"|g��6���9���݀��rդ�t������&�wn��@
�Ր�F�qN�+���(3���`@+Ә<�+9OX?���B��!��<���Q��3��͞��+���m�<&	G�A�H�^�y���n�Yv~\\li~P�2"1���K]���@�@�SD1Z�,V�z����G�����ad���� �?W�2�:�p}��ڌL�T�l�Vu`��������RR�ְx���u�VpY��z��R^#�����S�F%���l�7��i��K��i�ހim^Y4Kן��9��F�:;����B��$;�4�Q�����B+%���j7�sc� ,+�B+@�唼˜��<?�RZ(h6����Gsd���]��2a&�� �s��{l�h�B"pg��{A�=��~��W ����Dw ��+nm��o�GI`�7�'�O>�}�R�����HV�@'K[�2FnW�!$�T	�'	�B��xv��6#?:n�]��Ŝ=���Q����2H4ݛGk�sNW���\8+�1"O�'��R�	ɺE��C��Bŝ��&�2&K@��]r룆��'��`{�����
0�(��Ņv-6F�9ʵ9GV��9�K7ܤ����jI����X�>���}�"�$�J!����V^V!}<6_3��`��r-�0��f��Jc=QR����`� �a��H�9�G� ��
�}��D���������O��m�2�5�O��e����~��L�7���.�Vh��t�k�%IY��R�N���<�c9�Ш򼚶-{'� �̋(t�� ��q��k%N��U�LI~��Yߏ�T�������a'�j#�J���F�p���}_{)���d YvN��%:�{��3�P1��D�F�Vyq��w5��7=}��W�g��Cl�ŞA=�F��;e/rz	�"+�� ޹
���d��e"��ꤠ|�7�PT����4�.�[<�b}A	`#-��0x�|8
@�9�09���;���R~0�Dl����k6}���'�>�ˋK��p+m���k:���[F�~��Κ�Y�^���Ñ�ީUίZ'+#��eq�c��$�O ���s�\��71�=���=\�bG���Ɠ��
>�d��fBr��' �h��;n���[J����+�X~���t����x`�����*-��&�*�i�"P��̸�Q�9�ps#��e�"e�G#b�[��CJ)�_�%���:ߎ��4�Ζ?UlӇ�ɝO�������%�Y��������ݽx����~gU<�@��$�m��ynSX�_�	��oZ����k�w)��{�
@f�#���f�=>��`�0�6�fy��A���CK�cB���.IFW�ǂ�EyܒgzeT���3����vcU���&+�j�������{����1�f4��[����JU��G���^�ܙ��+o��C�Lv�4icp������󪉷��m��![��,	p_�������s��]�|��7��?(�0],�`�X�n��|���X�{��"���6GT�h6s(&��Zݐ�����Jx
# h�J"������wO���C/�p�����z��(���!��N�����dr�� ���<K/���Ie*�3�:K� ��2i�q~��M�9�����^f�Z(&�0_��B�D�Qț��~��Ic\|-����V9��	I�!%���-S�vܲkvA�>�D�(���瑏l��l*ӷ��7@|2�����J�/�4v\)sT�!��b��e�j*�M�� �&���ZO�X<&sb,� �h��#��[|ู�ߏ�Ƴ��P�-wJs�6��XQ��'S���D���X�r̨(U������ �q;n����`̈́��$�7n��F?N'W$
�$w��&Ù��@�`��ޘ�HccK�'��rB���2I��ϖ-
-���%+�P4'�_����t%8m~����!�� F<�=4WE�w0�s��=P<�����2�պ�\�q�|�10 ��� ��	6k�D�.@3���b��z�c��"(��G�T�m@H�`[]s��4kWc���p��N�!5Y��{<��g����Wh�O�o���ތ�r�E��\������%��'�#Ƶ���a����J;C��O��8�B�4@)�q�|+&j}����D����"F�ƀ6������jm�RG��z��~'7�z�qx���������;����P*ˈ�¡��,ͅ��0��I�$�� ��2�B(�,�K�v49�A2h�u����,�3�s�M��y3��^��V��t~uM��$�?5]��>�Wϟ��Gz��JWt4�3;x�� �!�k��B�	������8��G�s�:}�Asͯ2ޠ�M���!�_}mU�$f<�|7���-PgYN�d��@>�D�������j �i�x{����������v�;��o߾���]���+�s!`��㸺� �&�>J[��K�/�����|dE�C��ܑ B+���y�pH�_�4T�%k`�����H�w���R�ٚfP�yN�r�~��ƭ�$j��`����|+���|#��^Jmjy�ə��m�ґƻ]��s��͝( �);Z~Wk^_]	���������a�����H����M�GI�wPN`����S�V?�ʴɒ�Gy6n���x��]\�˵���Vo�-���zm���݅��V �U�{Q����s�|��y�q��Z�1��hk��w}l�q�},��+��<�H�}b ^gkPBD������͋�c�-L�&;�#��DJ8�׷�J�o�yU�i�{�^����^r�лP���t;3/�:��iEJpJR�˞Q^I0&����K���c̀�ז���G� *�&����d��E����u�D���oN|~��g^c�z\x����ş�-$� S����X �x����̲�dw���އM<O��e����IK-�g���3;O��k��r���ǜ������A��J5 "�������M����g~��'��.4�#om
0g[���=mʾZ�W!��8�L΀��&j`�[� ����+øe���!���:��Q��=��V�0Q8���l^?IC+��}�辯�����W�ҋO>��ե�N���Ⱥ5� Xe�:*xU�6���V
(�Z���'�{@��xE��G�C�z\�C5�\�K�_�o��HA�`��,[��fQ�	�e�m�)�,6/�,ð�C
�c,�b��ă�X�#�հ8���4PEq������3!{���Aԁ�?<�]^��EIu�z���'zǡ�����
���~WuNu���T=��G(�\j����sǤ�"+a�����\�����-�p�����#� j�-9v]���`�=L�=��:�=(�ꗪ	ļx�;����ŵ(��/��B��x^���M�s$��L���0`�q+��A�g��kaO[�Z����?9�	�Z}�I��h�\��~1Wη4g��>K��pSB�q<+�o��V������̠yv�E�%oi����%���E��(7�w���[�*��?��>��S��Ot��D
��w����rUUh�͹7[�ܖ�eVb��q	 6Z VE�wRCD`�Wʊ9�M]?<��so ���bu�����(z�RP�"�A����{t�E6SxT��������J��d���v�5\�4���'S!��;��"�<"y^r*���9-���р��{�8ٜ��I}�᾿'7��h��U^���<��M�rB[!YXǼ,��s��+�AI9��˷�$��E��J���V{Z��;�޲[�'U�u.������tܨ����x������������޼~��|o��H7�ݙ�	4<��qN3�@/��H�єr� ���"��m������$�=�58hI~/�����o8o��Aք���_��Q��c V4�m����/h�6N��1��:�zF�~̞=�L�֦T*�y#/��y\Яd��ȸH����Ci)uO��B�t`��-�WY��,���gqfZ����!���XF�b�%�[Q�7X���jV"*
�@Ia"��	�$�j�h�������?���[��yG�9�=���e �ۢȥ��Q��h����4_������������� rE���X��)���Q{d2��*-��A9~�R���p�a`�x�%�=�@���I�΃F!�Oܒ*�����\��g�4�~���
���H[Ql��'����-5Q�Q<����p�y����f�l6 ��?�g����K����(E��	��&��3�o��ܛ�b�^r�vN+��O�Y燽#I������G֧�,���faF:
�EPK .�f�K���a/��'�����c�=;��3 ��g�{�3RɃsQV���� ��-9Q�ؽ�p�n�O�e���mԯ�5������B���A7L��|���b"��9���P�l��s��q2/�U����i:8h��&����{R�8��^K,�����)9z�{�ڄV2

��V�u�hv�� �Vƛ��O;X����ZW�f �C\�|�-}�A{b8��s4e��/�˺�&�"o�,��o�-t4g��g���t��yQ T�e���l]<Ms�Jn�>y-M�V�)��fl�{P/���9�{�s�;��3 ��l/����}` �Ix[�^Y����+L~��x�3���퍬�R7:��� I����^��6"�y��b�@�+�T��=8X���}c��m{���~��SŻ4�&#��E�&�k�]{/C�����uK � ���2huJygkJ��Z��E�VS1Z+�ڡ��d0"�_v5��B��%]_\���IJ��/���Mؓz����[@�G���
��E�{�d\�Q��-2\��]I����>�)�֙9���/e�Ⳇc�;G�<
]�Qн<H����s��/�:�)��G�mZ���/`$�RC�L��C�2'����}����@^�P�L���->S�e����4M��d$J�(���1I%d�]yl�0�B�QN�m�3b���_&!dݙ�5��}��B�}��΁��"?!wgwe��Ox�j��n�L�#��q+��x���!$��W4T���i����2�Y��Ɗ ě*k��"56�B|Nno��+C�}���IְV]YЬ����Y����z7搇zn�ڀ��� D )�(T�5/�&��0je ��(����\F�}TCF�}���w����~����&��
�X�0 ���|Wv���,��Ãϝ�D�s(J�EQ�^��0h�x}��  N`~��-�I~�z��]��A��\=>��� �UAy��7[�$1i%�ø�	�g�Y����9��hU����rA)����ab=�),xx,�y-G[C��C��E#xɓ3 ���K��:�U��arm����<^l@��/����?��=7 ��:"�Qx�yN��Z�M�OlZ�a�Jr��s�y5��|�ى�z-�" Xg��iU���!����F�Cm�����A�V�$��K���HN�!��7!(U 6���FU�;�뺟-w���xg�9�}ќ1>������{�uU	y�8������N���m��U�`���ɫ�����@�� �/���P(�6Π `Z ��q5K]��vص��e]�������|=j*Ͼ0���/�n.%R ��FAԫ���\��Ç�O��9��+[��r��~�K�3�9�e5|���G���Ԏ⟁��
X��aI,G����a�_�|���Iւ	s9��9���*���W5�-9�,^��� �ң��{����h
�������ޚ-���h�k5�
,�K���C�
d9�Lyl�{��2 ;H�(b'˕3�o=y �9��d.�=��˗�b�y�z�򮅕���{�jXI��;n!]��; WKkD���2bէ����u'!V�l�
[��V���"�d6��K���V>r/,��"�7�����./��Q�6!�VBXG��%�B`����'�8 4%�BF{�MS��6� �竉!��܉``�V ��K�c��ҫk�4�RAq�k$��;<�L@i��)��EX5*¾{0z��{��B�r
r4D�a�����|����ˋQ��޽}���k�᧟�I>G5~#V�hg3�L���� @�d����xҲ4��g�Rx������;Z(P=8A�BC([����4�`z��>���ځ�H�}�d}����8\��s����d���6��+�{ 4'�#�W8G�a��kh	��4�š:�u����%�˼(�䅶�i�G����i���� ��=N�7���d`�O��o����P����ժ�z������B.��WG�qp�)'Y�E�e��j��d�;�g�e+�P��+����z�F# �mS�;�����:��}�x�bP4�s�Ӧ�S�܆�
�imD+�-:jd�,���ֹ,��E�H�	�\̋�'�ɸ��, �|_����4{�$��� Y���m�� �-�fK��r;1�,?o>ZԄ�Q"*�'B�����O�x*����-��g1!+��e੼��Fo�����8��g����sH��i�&b-�̀�1q�9�f��-�{&w�; _Y���29͟`ap�Paĸ��sp��"4  ~@i�-`�gm���K&��'�T̫���HY� �rA7A�R%	�Q�8�E�s�86-x2A���/���e��"�\�Hq����s��Z���R;�gS���s�s�gK*�ThO;Y�����Ҵ����=[�m�jI� a�9�����$�C�қ��:{=8�D-ϑ����W��Lɘ�/��\�n��'jပ�����iӰ!+W�\�� #�h�UO��bS ��� ���^ի��P\(5�7�z�S�)� k"R�8x�,c��J�9�>�����|N��ks>�.X��<+��U�.-��4�x�Рx���%1����G�����U�8����n��0�f��&�h��(�����4o{ͮ��;�pr6��\���{��rX�[ 	=��9ɛ;�ݻ5�a��!�1��)r� Y.{��U�Hh&��`k�(4�{�`o���7���3��&;f�4��&�����od�b�w���g&��Iݰ�5D��M��YZ�>�&�Ug@��)�3ڬ��X��z��+y���x��!������)�s�c�Axo��\1�bx=�>������C�Q�� ����L����@
/��D=P��0�tH��p�y��/��E�{k��� Idlu�'&����v<�jZ�y,7��ye�x�c)�%���2S[�9��&�M#�v��F������u�v�b�[츂CMſW����Iֶ?��Y��T8M��y�1ꨄ�⯲g��Ȃ�u�0c�Ő'��w�����;��G9ƅ���QM��̱b�8a����/mO �l��OʄD��)��2+�x�.����}Vĥ=���-�i=��Vu1_�l9_po������C�r��O-�� �0.�U�|}�\o ���tѠ�/����-�4�I�X�& k���}h7� �l�4��X��n}��gM�'ɛ�5�+�ثX��po�
�Y��ai��
��0��G�i[�}Wp�n�û�n�H7+Go��=�A�	�%`�}M�e�$4�����9���3��y��Ĺ
ꢢ�M�����`��\���,��\�(��Y��f�!�I@�
�U��'� ���>�8���A�����Ԃ%o�����(�X^����ك M~V��ozڞ�O�?!yL�lB�������Dz�I5��Cu�ܬ��F�̒`>�ڃWQ�Hp�P����D΀;��d���_���u�ȣ�y�޽�\ ���nF���xuVt-<bp���|.^�L*��X���s�n��kH�<�k���gr<+j�54P'm�8_d��J�D�<�50�q�l���挄on��y\�y.������=�.�aAr/��z`�����s���$
����=�S0�50<�fC�iJ�,̫yd�%O��1PMs��w���&Uo���ݧ���7) ޾�� 5���P5y��mw�p���n��`	�r�1t�O�*��ȃjd�Ib����^����PY	*�=	�oG^��L���3��)��3�,.��s˗��.q���y�ё@>�a@�:$�8�_' s��ֳ�Z��(�8;$]�5�lm����U�#
z 7�@[�. Ԍ����qId^� d}�}�|+���A�3u~��٬�X�pb����G���G�Ǜ-���[,虅#��+=�<t�Օ(+��]��"�*�>�cWE_�ES�H�`Y�oH����k���Q�M�*�-8/*��eu%}�|�CX�a�S2�V=V�~Vר�G�TL�f	���z���NY!�?{|=���doUY�j�)+a>���Bz �Z+���cJEq@���U]�GI���3��3�Dn��o�_�a��v�;��YhZf̖�%rM��\�"U�p�R�wӁ��7$_���WK��s�������̠kk}�8D#<RE=alI�d^���VI^` ���K����1�k�3����z�|�������Η�<l�k(�-DrO͞�="R�y�u���E�����%�G���X�I��A1@R�4x��ZS�RT��+߃��Dm	�"�t��������a��J��-���հ���5��fV%��9o����Rs�Xְ�[��,V�x׸:jP�� ��)�|�ªJG�p<|��PT�*���A�P�ճ�C���a�͠�VxZ��	����ރ�D�}�O�wR��sa��o%r�cxW�ǲ�]����p��J�dLƯg`���E0��	Y�m�l�a����RZ]ՀA�9��	`���y�[5���
��|���=m�^ͼ��p���'m)ȴ�u�[��TY���m1�\S�Fɼ�&?r�������c"����奏3</��L����(}������_�d>+%�I3���i'k-�@��➠�f��P�,��M�v,���$ߙ�^|�T����{�م$e��cP�:�4;\���_Y��ٳE��Zm64�=~MZޡ���բ_�y�yp/?��nk�����=q�٦�=B}�~�8v�:o�N�=�e�Ȟ*��h[�}��VDZV���>���w|qOģy�$!��]�d��P�uăq���<`3<<6�ɧ��������xd�zM�q��;o���}���-��<ؚ��<Ӥ.E���,k��mF� y)i� M�m.V�����"6iK�7-؜ߥ�\�+����"@N�XZ���{��ꇼq���ۍp��aO/���\�����t�{�>Y}N�b�8�� G9���S����R��_���^�^7���_g���AX�hv=����בs[.�������m-�d���>*��q԰+�,4Q�6j%�����]�j����xT�
�M9d2g���r��"A��L (���~@Cp��2�J�@!G&{�]���#��-�/Η�����W����]v�
ؒP�=�ђ� ��/VX .'훧^@��NH�"��ܺnV�]ܓB��P%k�Yސ�i�1������O
%9�i�GkT��7���7k�*�E�d=w{X����2�<���u��=� 
Ϭﴷ+r�4����a��#H���R�I~���A�VY��:��H �� �`�$<Fѳ�`�,��r3J�: -��x������Y7�4��V ;�P�w#���!U/}�����7O�&|�K��x�M���/)�1�ou?M�I>�Z�&��#wH��Tc=��|ޣ��k��F�8{��$�RC۳�|���� M���~^
p�-��p#;����)E����N��ܱNpM	��Ɵ~��3�0p��w/�����.F��nd���=X*��s��{DG�{Q�gs��uh;�h8�B,��X�]:�:Y�����r�Zh[���3@�vǎ��h����U�Y׳��g���Һ�E���:�k�,=��f�<{�B�`o�ts�ʵ�?�5W��Q�8�H1�[L �a�H��Y>�٤�f\[X$@��=�g3�����Q��yCNt�K��`�sxj�4CȈu[rd�ɚ�g����Q�:ca	T�L}c�����HX���Sx�"ɯ�Ǖ.�v�Wڔnլ��+�}:���{���Յ��^�pTz�|h�x�6�}Ъ2v���3�IHQ����1b�S3�@�>r,���Xd>�}j�\�qJ�����b��j ��xZے��g�<*�	�� v��+)���:y�I"��N�{���2�j5�##�߼_�����
��������;>?��ּ��hJ^����ͣ�Xă`����������C�ܜ+�w^��돜}�h�i<'�\�Z]w4p9,�b��g��DPA����/�GSk"����GK�-e���<���?�G�?�{`o�N<y�؛y�@i���	J�&FW���(<(��㨉��.��U�7	'��c�{ x�CXS ��3%3e�(aw{�AZ-m� �
q�z���oS볭U���N����[�԰7�y���b;wY��S��dՕ���}�j�	U���2WGW��EP�IM�����H�g��t�p����b���_^�ӳ�K�fa� ��9d�b���y`��m���l_�f(j�(��}d�?����L�]�*� �Ae��Wެ�s ���*�_����`9��+E�U^Sq��c��
�-`J�em�+5W�v�ŀ�=_e~}1�n��*�k������4$^�:�s��#�I�T_M�MVt1�y���ط�֊�qԼ�I0W=�󏖞Uq��Ȏ&����S��
$;T�E���U,��,\�뾟����}^�*��<K|��F��z/����˹;R�p��F����������7F8�4�LB;�}hv�N�1��s��3������g
7fb�,�W�i�� `\B)�R�-�N�֤�����dW�!R�V-�~䐳��9�a�����bI�SW�mQ]:eD`a��@du_�1Y}��2# �`nn>:�8�
��7�=�����cŏ��� �*�B��w�(�#���,`XG�#�8:%�[}������)X?<>��,Jk�F�ؐ�Һ8;e��i�#���tv@7o0&`(�
��U#�Z�8�2����8�eZ�k��j�>>T��A�Q�-K4���u�*V��B�Ma�#��B��죦���N�ە�km<�cS�z`���`�l�+~V0[��򓵃���w���8X�u��Ue]��6��Bh��r�XcT��U���>#�H8�kͷ����^��i"���X�ۿ�
���B�<�Z�s�(s1��XƱ[�`����٭n"��% -��hFw��D������M�0m-X��6��$:���v�9��aS��a��vf��f @�do���Z5`��*L�b����!j:sC��x�Qcm��E�i���n�J�g�6�W`�Bf�2Ѓ�v|x��Y.�|jc���9nk)Ǘl��|0r�S��Ie�֔�FS���9 V�FuY�ƺ$tƀ�U�+Dyo��ִ�ݖ5�QE����3i+�N�����U�ǲ��^�ĝZu��E`��`�A����2�Vu,����Q�9	i�
�1%fYgP��p`�ّ-�~�Gg�Y��crB�9�A������8�����P���e�ǚ	� �x��kO��V/`\�L'�Cɠ 5tKY>�%��M�tcN�F�d��>��w;���d'�$0�����56f��Li��+v)�m&���t��� �$���Y�J�jk�v�4n��{���;�*�~�gIq��`�L�V&�*}���i�ɬJ�|�˼�y��v��ic�M�
0#dw�@k(b6E�~�2LVE��U��Ì��
�V)^�E��Qn����e[��z|���?m0�4�X���&P�Ɉ��^5�S������ �l2	����w�)��Soq�%�_�-L_�����^���/�re%	�����ps���l'�͎]�X�A�CJWS�x@�N���L�h�C�狃�L�)�U�������ff**�e�4U��q��`�����o	O}g%zP�O�X� +&p��`t�o��`��`�HO)e��4e�,� :�ST?$! �~���c�j��T���1q�Y���%d�,�e�y�g��ٲ �瀔M��u���Z��U�7;@�ө
�U{��S6��HN��S#< Ƅ��:��^S�;�T;hN��M�s��Ȯ�riN��4v��<����:�	/����k5�S���B*��1�X<g;4ј4Z!�Ժ�[�z#��`Eni�������h�[\�,M�;P��Ƀv�|W�P���`׫��1�g���YYX��0�ƺX�P���,�7���Y��h}������W4Kݣ&� �?�j�H�jd�㟙8�g�Ɔ�?��wޑ`6����UuVΐ���Uk�Y�|B2ۜY�B�8U.�S}���ʿ���k�fo���i�6�����?�.��9�Ǐ�d,�Ģ��`O\�_����N@��l;6i?Kj���=$����4��MTE�s�\L;`�t��Im�t�V�WtٞT��2�R�k��:g� +���qz	�gU]2 u��
U��(���٪�
i�	�$�l�49�LY	�M���'�����B���y��H����|�Rӂ���֓�o�Ne�x�7S���ug�Ij�ov�5�t���VZ}%�;
��j~�VS�������	���򮁋#Y2�B3��"b �|��E&���y:c?�&����<�ae&�q���
ɯ3f,��c'��$i��ٗ�积?���́��S[���-D��pʧ�N���&�6���U�V��96��LҊ�OO˴�-���9�S{�	�qc�I�f�'r��i���s����©�ڜ҃����R��ά�+[d,ǘ�nj5��߫����<�z`d�����R�,�Z�1&d0p�X��\ݘ/�{y�9PZp#�Eח�*3�?n?1��r�4tJ�4�0�/w�no�y�X����*����Y�$�y���C�_3X	�6�����B��t�Sy%��k�2q!�3�/˩�*Fȏp�
=�*�m`�X]]kCy؋�M���/n�Q����ʪ�YE��Fi>@F�T���$��w�{e����#M9*����z��t��_�VK�����`K_�'�
�{���v`E�\Ōt��=�k)]S�)+��7j/��|��w!n���m�.��W�)u�Q[Zu����j�3�����(��T�E#^hB��z��2�	�'�)����^
���.��
�P�=����9��@���x�ty�Ƙj�6O�ɕ���r�C�oó=����/�W��c��A��4���8'�Jc�`"xT9V����_8�DW̫�R�O���*=��A���L��J�	7�͖�IP�A��ZʡU����蟛�|��/^���w�����\�a��5�� ����Ԏc��h�9�
�Z;V`L:���^<���l�,�*����XL��*���e�iu�������KR���a�`Je�Ha��̨�5�� �O�q��A�#aDJ�LX)��$@��� � �k�!�A����=�1��q�y�ayg#���������r2o�償����Z3
�'�8z��2q�����DW��_�{��O*�����~�������i:[�G�d�&�X?�]�Y%�	N��"�4�#���^Y{���xd�J	�-O?S��[YO[n��I#�I���G�cp��T�&Ԡִ`�Ҝ�)���H�!�-oę�J�����>`褴�A�
�?R~{'k?EE����gkr� ���hs?U��@'��s��I�o�hU��|�f�m?�:(w�.�ٙ��l�g)�jTi�-�bZ�(��싓�Aa|@���<9�Ve�-��8>t�����w�s����`O���ռ׻.��n��߯I�*>t�Z�Tu��|\��ƸcF0��DɛxѼ��Qe����8.�����<��j�4%L�4�����:��3�Z��gmm�}XW��jč��A��A� ��7۟�g��p]�����ދ�+{�����ؿ�u3�D5m�,�$/�꼳C��}�uN��c��v���_�l]�1����)���}��c1����w�7ܧO[���`��`k]L��V:ƕ�=��j�L�o�:Nc�u+����!�����#>���W�?d���=9����` G��Q��Ȁ��Iۯ`)A�k�L�b��JY�j�� ���Ϙb�ѡ���,R����E�x���3�VO���U���z�{g}�W��	�`�T~o]_�V:^�tdf�Z�k4We�k�v� '������b�e>m�� ��
���f��}�v3�� kU��M@d���bf�T+�At��5����P5���b�.&���I���ߣh9~��ݠ���"f�Cj�)��Az�d`<|�B�4H�S���^bi3H��J/TU�O,�񕉹A͏���WYd�h��I�|#/��gg�����\,��}�A����� l�����bӰ���y7�y.s		�4�6=7a�۴)ߠ�����4���� �Ȟ�G�bަ��:D��-N!mp��<Tm�o��6}��`�P��J�!�i�n�"�D��2V�p�δ� �zp�~~�����H��Y�
�Re8n��t�t��*)B❲]��'C`�	�힪���MlYu���)���耞[���;�d�&���q�I�p���[cJ�]A洦��p�=�Z�@�kq7pgr�'ptV���~i�xֵ`���̏1h�����n��r��@)���׍S��_?�GkX����@�e�/�����V݈�M��S� '��T�s�I�AX�V�F�[�OY+!��$�Cn ��c��to�ta��d5�'4`�t`[q/��� E��� Y�RL9�qB����O�[C��ro��5�"\/��Œ��T�����z�Ɩ��ҹ�Ř���{���4��e@��&R�;^��}��ξ���XY��S��L����d����\�s�a�;7d0��D�v*�1Cdo�Ҏ�e{VcW}�U�-�
�wP�h��8bcW�#G�rǙ�ڗ;�r_tʳ
�b����7ON���k����sE�P�#�ڮY�`{�wM�l���,@X� \	�����\^�SS|�G��'�`bET9-l�YSVR�pĎ�3�6���:g��*>E�@ �����[��!XT�'w�k����N����_~�M޽��lxz]�?kErC�2- ;�*�uz4u
^�49X�`:��8��2@��))m�J��V�R�=7��'~�L� 7e-��H�VOK&� ����w�ӈB��;�4��j2z\�#��d�%�J�0��M��0���ʊ�t�I��ܲ$G,���R��s�秠��e��p@WN�ϗ�ݮ���_h_c���S�QS�M�h!	n��l%��萶5ňpW2?$T7���VCA[����`!T舯	�`�jJ��R��2M�`s�@��Co%�s/�D�ۧ�P����wM��B��r���V?�4'�#�@��+h�<6�P�� ;8S�"�N�դlg��|ʠc$;c�b�i�.����L��H^��>gn�UYW�>U^/��y�78��J�h��4X��f�5I.�w`�� �)6
�mc��J���{�s1�dc��E�4[�p�07|����� �3�w���O��8���E
��h�!�Κ5;#�>x��P�[*����ΌW��eP����Q��1��PO�㢈R�����{c*�3b�Զ8�4ςُ`n��=/U�>�����UWl�8U���L�Ʋ����N�����������'�ڲ�-�K��$�V�2fū!�������'
��X�����,8`�d%ٻr�F*G����ъ� ���g{�ٲh�ۆ��We�5E&�kh��(���[6ܼ���0�_e�F�����/^��_�cW!�tpnڞ��ٻ�h� �L0�i��H(,��-q0G�z��f��[''���'|����A���	����"m1�m�\z�)�A��g���۹Φn�qpD�b �6�P�.a�����of-�p �	�����	Y���*ž������cO����N�<�����	腇�P�������Ld6�Ǆk9�#�b��}��.ZlMj0�s��B���)������N��sm�O��=<,e��	��]
t�Y� ��v�ʗH)͝�AT�U7:���e��U8Q\�YR-���Fg��.� �S.Y�8j�J��'��ƘS��7al!�^��mh�g�*�9�܂�b��Q��R���=��A#c���5`û�oe�� �7����MEzA�� ���t�9<H'Ճ���V�V��F�h[s���go�������lc���n�&ǭ�a:M��&�E+��V�!(�'k���;�Q�B��~]�}I7���5N�c��:��ZO�sb�혊���Uec�*K��;��_�+
�-r�|M{�mCMM��3�N��� ���W��I��gL��ȜS+�&,�ǭg��Juc�p?���+�۩������(�Lg-�z:�7{s�J*m�:�'0z0���YĮ�!��g?���z^�"��7��w�+ ��2����H��L0k6��Q�n7�<�� ��+g�� �?�3���􏎏�`���,��mLо�
�5?�.+�Ll��H�tWd���bܼ:7��G���1v�9|��
�ߞr>Ao���)�s�z�6M�����Vۍz���a��=�@��Sb�
|�l.D�m,x�`Z�$}�|@�y��,y�T!IȚX���,���J��v�P���߲Q��>��3k7
>�����f���jv�qI��t�Lӡm�M�]��~�1y���*��L�_*�rу����5c���2��ߘ$#��|vm�W�/�D�/�}�Y�Q�{1�j�T�YİŖC����A
�k�f�NE���-���U� �\~����}�B^\����� �Q�fT�a�2J�`q�5�� �.b�����)kװٵG� ��â�6��%�[�����{�e>�3��zb{�H`�be�.*�{�ioᡓ&!����L.�^q�nW;� �ë��rIK�|�����	vqU�K[�
 s�OS"Eo�`#d�]��A�/+IGpzJ>ۥ$���R��:���ͽ�=�eE������8U�لb���)د��2W��S�ʊ{~���#j��ag޾�x�.����@z��
���s���{�?z������4X%�Z�"��?>:���C���0tL� ���$��ۣ�9/�.A�"j�lǄ�`>pr�(����S(
�	S��荡i�d���<���)��!,F��+RF�Ҵ�rIЁk�������������:kڻ��?�өA� L-Y,.�ތX{$6�?�BN���0ā�ߔ�m�H(q]�|h}�u0�ujIK�Fۧ̀yզX��kj�q�^�M93kCM���w����v��F�+��7��ͼ+������D*��� ������z�JOؚ���sZ ��J�:NX�����M�9f^FA[3)��m�.x������y�X=�<иQ$���O�z�N�)x x|Gcb0�84>>����]#^��~�0<��p��ެ�߬�1������Z�K�:@��C�7{�Q�����zʺ�{<�D�����wb(=k+RA������L��Ѵ�m�t`m���Gi�g��w#��}��)èA�l��^D�H-ցb�� '��3x.!����d��@|�ݶZ�ҥ1�jq������!�V��ue/;K���Z�a�~�.��H�B0��d��2�8!���U�m�
#�l�䘣�I�*�g���������O��F :@a����Ȯ)��9���6��&��Cy}u!��y� ��خc9N{(�cϰ���ǼQn0o��>�=O�ߴ���ጒ�rj�*�G�-�˾�z��A[�� 2I�`RQ��m�E"l���=&��d.�g� e+�v(pң�c���$mgrq�Z�^�N�� @gB�B�fh�f#�y�`��x+�Io'^��iݽW�&������#V���Ƀ[���c
��?\������_~���}J@l��8GG�v�@�B8
��Y���6��&�0�is�sxƂ�	��=_" ��ȗ@����%@{�z^��n���c���㰗�)����"�gv L��<�/W�L$�/;�`�f��^K�/.�Ӝ��}:}����:�^�wK��zʀsv�6��Rԓ&����7ě�;��=�� �	[Ơ�b����z/L!pB ����/^�˫K9�q�Y����sp-�w��G����G����3�a].�	��.��9��AG��qj;K�WW����jŴ���d��"k�GJ+
�L� �(�)�s/0�*D@�<>9&������� e��:���J���+��K�>;;c�J����� �|�=��zo�] ��R��+�X��j�Q���zq]��_`���T5�4!8^^^�?|��;�����)��|�����Y?6"���E ����i�����C��_�[ƣ���/�fg�_�P1fWW/�����#�������k-������i��䍛E�T�� ��<�'�NhGA�sCO<�6�X�����@WVQJ6�������P������V���& �	��}��}ü�࢏� ;+�p����u���{�kj�=���_�幾������-���^�q�����\f`|z�O��2�0Q��zpС�`f����t�ڥ�Fe$�*7��]U���� �������4-��<�[X��b>5�{=DC��c�F��Ӛ��$��p�0w+c��� `�w�*��0xel���^ǉEgGy��)�?�)9�^qL��1`/r��Z,z�A�/U��c ��m+����dwWd���2��W@!�n�^2K��թ��?��|��+꽎�^�޼mC��d��:b�lX�k��J
���3�S��7�l�4���4j����[���X|}���(���~�3`��i>L��D��?��2'�ve�{�W�x������rx|�b&[4��q��7vOX�Y�0Fa��D�j�1�A{�y�`�߃�aU~�}&F&�{$�����*��d�8;?��A:I�M���Ҧy��V�6:�7i�Lt@Y� �C��t-X��εb�`�����g�#O~�M�"dݛ��N�^K,�^y�iJj�E]�wt����'��B�l�P��7a�e�ROt�r�^60���t���Z��aWx+�E��Fwx�N=iG���q�j[T� - �m|���)<M{"e�R�,>���� ���A
��W�NZ�4'�O�Z��FI󜛷;�5A6���y��57���7���OJ c�#�n5����<���7o��i:i�
�TcM�;��7�`���O�����m`�m]NR�Lc�t��k�J@��������Mf�r�X/����Yqc��&�����~���b�z��z����W��9Y �S���L zl�W���/�y��_�|����O���� sj�V��׎�R����W�^��<& �Ё�<O����Qno��{��e2��r`�̣��L�a@�������{�O@�M.Q� 0$�ҵ\�=ҟϽ�ׯ_���o7�[��0 ����/���|j�(ʘ�%����_m� �Kٽ��o���Y��o�\�}@�B�����{����4�17�Vv&q��28@ŭ��-����s��o���<����5�h̎��� �s�.��=�7o�� ��cڣ�	��ݾFzt`��2��	�`�� �6�YO`�*�&����i��+^rQ��\��P4��xQ�oƾ/�p{PGto�s��T�d@���}$�<G۶�?��g�����ſ}��es��O����)��%�p��8ú� �	�Ct�}���q���k)M��<���W����o�����zq�*GvH1�K�a�cܙqqחJ�/}��2\�m�-��Q�+����XA�5��>3m�?�='��ݟ�㓬Og�zL�5*9�I�0�4�_t�aiN.�=����٤	Y-3���s9K����*����Z���%�[�9j)�jnSՅ��1�����ƥ9��7�[��1*0��:������#h�ˋ���כ7��۴���ן������o�_�mڌ���Xu�7��P��7���&pֵ9�g��s����ט)���W�����i���r_��P VgGw�ht���ֈB]�3�c�Y��q����$��Z�|��Kw;�ôy'�ˤR�/z�������o��:b�����;�W4��OR08�ڋc��1/7	�znڪ�@�um�W�4�S]s��,�'x��/^�bp��s8I��� 7ן,�C�xL�"��y
N`- J^&`��7oe�����;�.��x�&�f����`�"�o��.ܗ�#���ݲ��|���������	�`�$����0�~����Z�����AA�2]�Q�Ԏ�T[6gG�Q��)�?U�{X{ >?gP|��EZ�������� �ӯ��Jv�ifPj
L�����?������L��|��.  �g�'L1��j��P_$���U#a��x/�� |�p�½y��}���<���0�>m��}�����odan?�H��3� b�i�O�����JK� c�G� �M���� �XB�xx8'�d���}�K�.7���g>g�#vrr���U�w^�VJj��<�/�W�|�ǇG�7�AM~��:O���7z��-gi#�����)�W[+�Ҕ�ꕴ�)�Zz �s�?�(߇.�igc���N�Á���"]�k��b�9��k�o�7�f��"�����~Hs�*�����k �� k����G�[�`��8V`�����q���8?0�&��z]�;�����ZS���������ځx10G�&��2�4��\L�p�j��G0���J�TA%X���m���*m�������a����Ƈt��Y�[Sx���f�]FdR��,rɫdL�Y����d)#���C�� d,���ʶⓠ�j�
�t�_�ǝԁqv�&���@q-��F�}�B������߾R��Z��U�P�^�4*�;�Û���l��}!$�XY��\A+/�&��Q
(��,��h�S��<��{�c]Z���&�?`�q��2}�0��\����OuM�i6]�5���1;"[t��e
��t"�Iz��ҭ�,4-uR�fEE�~�z̪�0X�֨C�BC��ԣ65VC>�v2��W�( �j+����^J@�X��{�F���D�h�������ߥlB�ݒ�����<���ۖ����& �5[!1�"�$+"y$F�<�5����_��F��tP��Gz4��Y
d��B�1sW��!��>c����y6	[�Y�����z��	� �.Df���	��>����~b-&+R	Ե���e����
L_���k�X58z0+��pĚ�<�L%N�Q���B*r����q@��iڐ[�9v��UZ')p�p��N�9���i��yX=f�X XGǪ=(� ;�M�/�ϱ)�j�]
R �/_�`P���7����=���x��u3��%���\��	�;��ظ�Bc�tnը����҆#��Buc hT��@,��|}.)O��d�5���sMb����Zˉ
�3N�VP�3ά��	���3ڇ�OО>�4>��?�;�t��8��C
[�"v�MUq�p]�i���C�+��S��7LZ�����ԣ`�qϑzľ�q�ZԽ���&]��q��p�R0��|��G�\�i\P�5=,-K�O�t}a�:�}�zѢ̧��c����}֔1M�5�ۂLԁ1�gi�Dݦ�M��杤9��Em.R�[�7����6V�P�� py�VN�!������l�/�R��!1�cu�q�����J�V�*���z6���Z�[��X�#̛�df���e��"�<.L߅�c�7nl�oTw9֓���ؿ���$�1��A��&��L;s�fӐXOW�9,� <X�����$�í�U�a�ZX����J9�6�(�%�6���8eq�����,�K�R�S8^9M���d
�	�Z�z��`��5�������k价/�~�N~�����:����k���^>�Mg����i>��6��U5�z��b��
�OT�Ģ��}m8��H��1�>v���zM�y��� |P�*�#&�AZ�4��g���Q(���a/��ū�L`�ƭ����q����`c�� $���%nԠ7��,��1�<~8�G�	V��-f���_���%(�u� ���dUD���ZO�dP�<<:�F��-?�"w^���L~��\���u:-�����_�ۇ'R��CM�A<�KK�zQI[[*2�F�C5n�S4o~�J�~>�H�E��ZE}1;�r��xZ�}ȴ�A'S�����g�\!���Ҝ�4&1;��B룋��Nf�&�"�;bEJ��i�@X��*_L{���UՄ�d�ԡ[7!|,�d�80:��/A�m�+�2�zH���X	�4	��cxZ�)��	������JA>7��sq��Ҙ�A�4���xе_5h28������xr0��� �j�oJ� [۬��(7e5���}���������V�	A��Ǝ~�x/�@�
��r���x�,�OM$ 
��C����P�v1���APj*^/[}�h׍j<0S��`7Ўپ_'���ْ�A�h�=|���[6�n��p%��Y�M[���i���[��5�A�:o�k��hpa/9�;0��k���J�:ը&��RػP	�T�c���
Yp�����V�z��Uf�57|@"��:=�sF�}���HO��=�"�H�6~��B���7��i�� �g�оj跼���7X��v�
" 4�ru�
Kh�{�0��Pd�*�\լ
��a���g�����ឩ�)|����"s��Yz�%+�6*¾��,�59�l����0 c��s�utxzµ^#%���]�T�T�����_����C�>���l�k����59��zf�HW�34Wn��P_���R�S�>*���f��d�c���:a�����iQ
tvƪ��%��Lnǵ�bq����b��f�B����!�V�U��P�\���Y1���ɂ{����9�0�ʿ���Ʒ���Ǘt@��Cz1A�4_����(�}q1@�`O�v<:��wo.���_�"���72O��v��*��/<�k�I��׼H�����qc�\z⍊�Ӟ�{tlv�xv nU�_Y��P3:��Wɹa�Y0�FǢOsF���^����ƽ����xA��A3pnLA��*h�{�^\I;Sc��W�(�=���$�N C����`bU�M>Q&�1;� ��hg˛JN��M�,�f�Y�W6�h�t���p�&�7��M0�B����*�5�c�X9M�j<hV)�`"�ǟ���t��D�i�ki���EATcjm��+�R���{ �٤1+��c6{�1{j��8ٽw*q�m��u���#��9'�s���%-�_�>�F��H�����	mc�[Q[��~���z�EJL��p��K�P-�F�*/6�B��L�9�v�x���T����z������ˤMq�U�z�5V-�� 6!�2�X�0�'�h����Qec��9���oh�iD����U�)5�
�1�3h�4%�Z��T+���m�:�����^p��L��V<�yC�U��"o��`�x�fBX��P����B�n-n�� 4{�T����s[��(X0MƉ�v�
Ź��֦![VhqF��g����B50#x��[�@+����5#zB�J��G6��~����a����:�8�9�� ��0�ߍ���<��١�d�5��v.9�榾�ܓ�1F�Q�`ͮ�Lհ��ҾM�?�+���U�u^d��l�9��
NgG`�T�����S����+�����A��ӑk��Lek���̺��ZqA.��g������> ��@`\�u`��	�Ӣ�:6s�=e%����ʬ�3��=ġ�0��8��}z\j�U�֣�ܠ�mX3��w��b,����<�t�Sw�d��V$SY������oPĶ�i�tvwQ��Y�X��`�9Y�;
�!��7��_Ҁcg�ܲ"��g{�����>�;���������h ��k�!cL����i���#��k��-=9c��7/�������o���3�ϣ�GVk�0���A����S2eZo��y��C�:�~�\��H�my�̬!��]�qN��"��/�f��)g��#�CҾzx�b�1�����枋�j�Z��������z�i

���:���gjF���F�M*g\�!g��¬F���Y�Xr�]F�� ��w�6��%�A���6�/���+!gsz��Y>�9��(�/ ��j��������ك�~>�M�
����V�I)� ���.� �������Ƣ�����
`�"Ȭɒ��2r�^)��*m�G�^��C���W�O���ú�I�3w|���ߴ�$�\�]�S��ۛ�&rv�6�IM�2X�t�+v�S[z�G�0�)�E�q�',ۮ���dJ�s�����j ���rq;.r^2�d�w�+���Ȃ~k��iALۅ�&�'��Fյ�5��[k��@����f+��<n�V.��u�����2q�?E�\@w͌����PƃO�8pt�}=�I���@NOΨU���
J�Y衙��_]�+�.�R��)3	]۸h�������6p��Ȓ�i���c�mm�5�7\���Ֆ���~�Sa%������)�q7����c�����
8��S'7��ܽ2�5�z���s� �R"u���U�<���o�N}�ԄVT�������i�*�}Z;kz��4e�Nu4�~��*�5Os^&�x�5�Ui��2�T���I�~P���d�U�0��*��{��F
4=��[��Q�_���p��KB���D�6��M]�.[= ̨]�f`��Jh'%���z����~�{��Z�c���B����-S�d:{��{X��8V}��i�[�i�R������������K���v��ux ¼�Զ��ݓ���2V����-%��L�X�EV
���N��|�jԂ�ݐ�Uܜ��r��"�1c�!��ꍁ��6����N���00��^�'ڄ��O�_��?�?�􍜝.�F�iCP�5LTC�^?�4��'��2K`f����z�*�d��3��v��0n�5�[�
]S���Z��A祈�x+�tK����l�U��.��A���3'K� �-��!]����j޼���\�kuF��T�*U�@1�z�DJ�����]�,γv���?��6�{¹�CǓ	J�#�h�sV�Q.U��'��Ȉ��I ��p_k%E���\�bq�|q���x}Å�翿g��l�6�r	��j;��dU�6��x2T�(���<�?��M{��%��`�Wvi7�ܾk��y#Q���r�&�_^�����N@�ϧ�z{� 秇rt�N�����4�:�@�E�����l�U;�کtJh�i7��v��� �[;�JR�
P�}���of���B�٨hDʃ��,&6O,�6�a��*�����`�.IP�}@\����5=�6�6u�g��{ݼ�N�ގ�"y���T�T���u���7榬���EZ2}�9���Z�h��ߴ������T��Q{B�}2{�,f�*��� j,`[k
:'߃��S@� ��|+��B��n`��[ec�����-ҍ��kO�麃v=P�����O�����U�;H�	��� C�Wvۋ 0 }���%utM�E�4ӥ���gn�<h�]�Lq�ŭ�Ϭg�eV=�2��������O[�Y��{� cA�����J;�hJM�w�S��.��e,�}]:N�m�~`�j�Jx��UT]�9*)O�9�;��A��c�H��Z���W[gu��	eʢ5��W����Ւ�[�'k��7[��}H��S�m%d�$Z�<u��A`S+���ښh�}�B��7 d]3#s �1Ø/����AN3�g��=��ay�Ki`c;NC�|��[3A�aJ�S��H�4]�³|�{��^��ڵpA����w��nz2亟��Yz2��hȖ�(���VΏ�^�?����}s����.���N	jm������B��L5���� �B�
���:�7�t�yJ��S	T�G�2�\t:�q>Ln<G�2���K��,�N�cl��O
`j����,Vp-�r��^�`(f7q�8���'}z7Uec�I��L3)�RA2Sԙp���rȹv�CMA���AfBߕc�zq�����'�F?Tf���6�^�>����X���Oa"!���������k
�3��}���M�L�ؒ	� ,��:�C���MjV����<���8����V8^��
�q��2<��"�rz��W>�q���ǸR*�����TU� �G�'mP�u�Eܳ^�V;�Z�#l���7 o�SL?�1A#l����\�j��X	8�8�Z�v[6���yv�V�.͍{���\��R��S�L����F�W�k���\����L���at^U�X{ �^����ڧ�-�~���1=6�%O� &h���U��D�^7,nl�`a6�*A�wpcS$�\��U�*;WOf�za`{�t�2m�[ܴZ����V>& ���J�.��H/K�ai.���d������t�\��z:���?@č*�N�Np~zƍ����7'�'r�B�o�c��J7�8ݿ����OuU�Ԛ���䂥k���� ��t0׮G�-��8`���mڊf�Bn6���A��䉦c7w��f��O�D�Z�`���,��N��?����LK��|��'v���Q��p+�ɨL�1bL�N̼�׶?�ժ�	��δ6�����b��-7f|-�+�2C�f'����k���l��`筛�0u�Z���= ^$صjG�I��q�;M�[Am�j�����9���+yq~���^���'8؋�g�Z��{o�t�8XLճk:!#��s����A�S�U_ W��v38d� �j��R�a\;�������!�pxQ���2(���h�zeљ�4�qh�����]i7ƃ/8�����$ծ1�H�PhpK�H�?�	���H;�XP�}xf%[d��{c�=�5Zq��x������ l�����K��;z�L;b?f��"l��44�/������O?���)��g���Ɗ�	��e���`�Z���ɹLQ8�8r�h�ˉ1ͶjJ��ӳ��Y��ja�!+�M\�n_!W���֮̋h��~�NL�R�e��������
g	4VJ�� X���1�S�I�t���@4����R8hz[Ć��A����s2 �~���Rqѳف����Ʌ����M^,�L�7(�|��A�Ϻ����u#����T� @꿐��o�j���7�(�������fZE�n����;ǂ�=�٪��x>Y��*����4�����5��� ��R { ��)ji�7Oa( *>(�n��;� ;	�\ �i�e)���R68ٕ���z�桚��pcS'|(3�z���C,��[���bϣG�t�YnR�W e%�أgOnl��כ�&�O����cu�^�����&i3P�t�0��` ��S(��C�h`oG�~J�0-,P��,Jm���9��*������(�5����N�X�C6R�����x����I�E������! J�w2Шv1?�GZ[h8�55`�Z;���LBN{j�B[FH���TY�`��^#4:�<Y��M��Z6I��8X��e.�G�f[�^��X�v�@�&��U�ߋ7�VϬ�������@k�t�����փV�Vs~�9�,��U�����ڶ�spt��M��*Cf,���DUd�>F%�:�?UX�w`�P�b�F+l���Brk4�g�fV��5��2ͩa�ȮV��w2�}���'��b�i���v�ς=l���N���C���=��h�Z�v%�)��hy�E3&(�9L�}�����'_4�ŀ��`sM�ZM��dIįY�f>.d�&����?�*��b��VFX�GZ)�x����vY4u���;'���}����4K��<���p���C�qg�2f���/c�_��L�$��CN%<�M�Y����4� ax��2ypФ��r|0��˿��R~��m�gi�l�ߨ�\�~D "����*����X�`���6�Ͳ�7f��|���{�e�� f�7
��W���<�>�Lˊ�,<pt!-�EK鐗�(�%�_�&f���W�"�F�o'!�*hY����N�!}�iy�;�zI�T;ʎ���d�<jz����uNN.���XE��l��V�Z��,n)>-�х�b7b .K�!����8���}vv,o^]�m`7�V5�!AW4 V�Ņ�P��[�0qc`��nb<�Q���i�h���I�2Jl�8�����|eA�3C(�"b�<�������3s���~�"�9tz�7�)=��sH��FC�
,�eAo@tR�[U��պV�}�6��F>���t
��zmփ�'�w��.��hil�������f���ҽB��Ǐ�F�'��rڳTn�N�c�ڕ6!>�����I?4�'V�l6"�8M�~ �/�)����^�+Z�r����;zѫ1��IOV�ZӁ�|�9��x�`HP�^m��j�Ra���o �N���6L�WZ�=��]h؊��Z eR:VE���5�5R�n��4�\E���Ji�u��k�ֆf�Z��4����7���X*\ ��C���s����Fnn>������n�[�4TM��қ>�X��tY�挧�\���%�)�}zД�D3�����tiڈU��*���G�� X"�R�:n`7//.��<Η�H�h��Γ`� �R�-�>Ѝܗ�h�ksZ?��n�.7�� L�h�*s8�E
[��Gv����;�𔦺Yb���#����V�	��֏r�;��m�QA{rt�1�5���7C>CG�TkM��  �Nh�<O��Lp�L�b)r;488��p\�D�Z��L4Q�W�>Nv8�+��y
�t�qEۻ�'h�pH����aǲ���T��%\��/���ƅ\>��*;�K��<�R�{��*�GZ��L��Ew�A����q��ɮ؂b���Zϩ��:���?�wo/�h��w)
���'�=C����uՓ��,���吻pT!�����"+����lL8O`�3ӨF�E���trt�,4�(�Y0��AQ3c�l�55�f4[����N�G^�E��5<5(`m4_ZK>�R-Ft!�I�u*UL;�m���&��-D��K�\IX[�heFmXH�ő,��)b�W~���|e�'�4uʩې��h"�\��@�Z���ĺ��T޼~���r�N6	L�T�υ*��ͩ���P���0X���� (�5"N\AݲOS�k��a��g�̵㯲��b��F+vM#1O���¬@W�]dg��������)�U�����順X���I���Hţa4�'0�c������'��� %��B�=����g�A�ǓQEc��+J����������͊��s.:?��"��"r�< ��{"�����Q��6�v
`�*Tl�DUS�՜�:	�����˨�Pتs��8z�0�I+ڽ�Ze��!(�l(rW/�����.5VQ�Z_�% �Z��U�NR��o�,L�Y�
�z3��i�mq��ȇ�`�M�>�&j��N�i�F5�,<0`�y���t�2���R�OKP|,
魤�1���u�ן�~l��.�~��u������K�3������̘64�рLPn]Bnl���40G��i��w.�*S�5��6�9J���A��90a�Y��qzrªO�VR���d}�_�T�f��ܮ�5�\�0�A�J���=@�lhT��ϕ�1�U�A��L7j'�4XJ��=����m��k�gh ^��|+��
�S:^�U�UF*[���0��6�]������Lk������?|�K������JC�y5ڜ��r�*g�������d���!!W~�7����a���+��+K�P ����w���"�X�eed�{}���=+��N���MV߼L{y����Q2��v8���M@r�Ɂ4`�V�C��B��2-�����ڸp/��;��ב+E�K7^�^K)��8����
��MiC�R[V�cS��}��c0r�{�T��1q��*&Gr_(^�t.`�v�(׎�t��Hag��篡�I0T���m3�׌]`�jr�����I���:8�lBBC�x/��n�ٕ��*7�����������kh�R�UL���S��'L3�܋*>{H���5J�g�e�ʇ�ˆa�k,��#��l��WޣЩA\���15O}�ދD�N�����������E'?�˟���矾%����N#����iv�����`�$��.�I톍���]5c/�U:�����h�t$��*��S�3�=�阪���M=@6띓p2���`�j�5�D�+<�Ea5�� `!5�@x�q�W꜍�>=����4E�aol!��&�f�ZiY=5�@�~n *ʳ�
��Ό�X9���.S�u�2��4;�Ӡ��5�Z�A[-Ώr�x�J��n���e64nr�n�H�=-V|��z�U��y���u�G���vw�~J7���m]Z+6�ه:��]��l�ҳ)�����앶�I���r=C�D�ۘ�8��H9lv[j��~�}�A{U��`)������6ml��Sg-�tgL�bL��`~h������{�'3���8��|���F�n3U;k	�6�/��>[�`[��Y�`MNs! j�Ĕl-X�`�L-;�-�ĺj���`[����1��1���V�� �žS�uh�9��{oP��>��(V!iՆ�D.�0.���՝�:�=4����<}���}�?{�1���]P1Pv/��C��zY�9Zͬ��`qL5B�6NGF2c��	$�v+vWy��6�7g�Ff��B�������;������Pz���7��=s���Z�Q4,��݀�<
�4�Z�!�V�e��a�� J�mF��~�	�@�y|���o�RL���9��5%�ణ6�~��4�OV�вg��tgu>XD�!_س�ѕ��$z�>3���>	�waH��H�3����`H�$X+����C�B:=H����_��G��P>�ޤ��A����>B�L�y�PX�yrE��T�-kn�$�}^?`}���/9����V�W֣�b��,\�>X_��BU�"^_��$x���!0P�Ӗ基)�+�����/��<<��׍3`�b��l�>R��>�ڿ*]K�|����/R#����;Fo���^U���6���lVˋ�s
a'R�ńJ�(w�]�Ԧd��f��"Պ��T0]��
ZP��V�d�E�(��8G��%��Tj+��!��=[���ԟjJ;���i�` "�
����T��	�ߙ>�zu�ΠV�C�8�ɨ��*�LC�&*���]3Xg�P�@���̘����0�G�����,�4��,�f��5X3���WM$ �� �'�	��P��E�̡IH�[�.��+ع��D-Z��۫(��X����`�<5;i\0�k���@ �
�&�}k-�p*��~�U=iz���C� Mv
L�ڸ��Lg�5Z�Ё-��a�+���jZd@;�-�����LM�9��}�p=w�A<� �ދQ�oM�����2~԰�b�!b~ij抴��i���אL~��$8z�t�kJ��*��c�2Z�H��ͼY�y�EUe~]�[cq���SL��Ӂ�0�s/������D�� J�Ҿ���-��̵~ș>%�1���T��&�z�#�����,��x8�z<UL�_~������)]K�~ʰ���tu���0�8�<ގ��(���0d����9�<��������mR�i�cl�0@�,8�L�~;����,�XL�彑��4�i�  {yu!W��l1��d]iq��m�b(ѰB�� S�f�k�|C^��H�Q<�>R{����o�	���VV�Њ��\c�6R�&!Ke{τ�Mk6j��󪼊M2��y�:}��f�`��r4��c��wmHg<E� �������t�� ̦�8e����.� `�BDp�Sso�g��&��l*:�в�@R'E�Y���4B�Z�̞)R�WV[@8�`�999LT� C��ѻ5�6 �r��(&\*`I!���yx��"���	���r���:޺��O
~��X�J����>_���[X3`�R�ʫbm�K?4}��=ɦd�>|����o^��鑜c,�[lP�T%0;�~��#
�Qe��J`!�00��TY�Z����s��uC����F]����ʵ
�m�k5��[�U�+����"��郱�Q��bz]�-U}`�`Dyz~!��	��Չ��I�Ӣ�6��Z3t�Sm��f�h��"gBڠ��ڸ5�4��zɈH������[�J>�@'@�6`��>M��5%��\�9 @%�26�	,>bNfXE�^��0����4@Ņ�*�c��:L�nԠ3�k������Aգ�N̰2�i�tܭE˵�Bkt���8��"5���ސ)z@!e�" �F��x_��Df�׽AS)���=B<�+tQ (�P
|�0E3����!k&)^˖ ZK-�nba��Χ����m
�����H�[j�q)RØ;j�������t�^8w�*ǍYh�Բ�Xd���櫶VP(��h�V�t�[0�dCk@`o�e�.E��'v�o�wX`3�s�3�B�P�⒙q���H՟_^hUe;1+����iKd���S56�,p�����,-Az~n6.�Ne>Ӿ�ZQ۳�?���a�kk�-�
��*��#%U�+=���*�i���Z޽�,��=���گ.֜4鴸�����@:�\�A>�G��ʱ�ƪ�xa��\��� =b�9
����L��`��uq�Ê��&�H雭T��v�ek�9���\��� ��Z�)����ř�fJ͗t�CQ)�Y��C��1UT�W�
_{�0bP�rv!=��֜�b�bg&����ll^�ء<,���	�x��oUW{ȱ\F, ���[,/?z���i����K�q�Z)&ah�F�E*�����y�to�*�V�=���
����Wa�T>G���_Od+�g��RɰZ��.h�(i���L�%���Y���FF��?�ʚ�0F~z�$��+O%�ęy��>s����n��k䴱))м�G��{3K�8�⭗B����k7zӽ�6���Nxg�Vh��\u1��u͆�+ljd@A?�sj��W�HS�媓���,7p��J� 8�*�*�K--�S|:��Q�`Ƞ��)��f�ғ1
+�瘬Vs�SfDc����9�S�bVcBl�r�� ]����7���-�)��Fw]��;c��i��U�"`��cK愄8���?��`�Y���_�� 0V�M:�߱*U�2
��尙"��?���v�f��@�F, }��2լ��`=Ze��k�|{��zУ���%���Ӓz�N�nj��M<���&����Z�����%�e �Y��F������D�6 ��e�8j����)E���z�T/5�d�W��� �Nl<�n (D k�x�T6���Ě5�QSX`�zK&s��{�^��	C����G��C>�ܤy���� A�l̳�z
��g-@��<��hT�Sx�`ݟiab��v<����R��CE1�]���=R���=w��IV$��Z=�xA[Z����oP@���	BO�GZzt5cS�&qF�kM��w�ֻA���_p6�:"=���?(���Ԏ�n	��^yŧڠk�j�E��[`��d����yo��7x���9(p��K��݇������f_a��H��.V(���W&֎�]�l�X<��;C��8�-2m�M�=d���Zai���imB�ѨƳi�\`���ZA9�q�}�E{�V�V)��M�YE�]5<�*�HvB��f��);�j� ���G3�I,��>�Ĳ�f��VF��=Ğ�����b�a��Ӟ�v�-�Q��z��(͡�������,�m����f����5��(&G)��z��i&�É��"��Ӂʞ���i���v��IF��}c����đ�f��@#p��/G�`�)b7d�tv�V�M@�l�>��U{����vy�2�#�=^�ElBa񙇒3}1��Y٬�bu��/��� ��Zhg�f:>�����lW�P���OP��	���J߭�8�������ޓ����k
��D=�O�Au���qC�!I'�X=�"�<�=[oC
RO�~F_�u�ձ`F�	�9�������cz9��������I��|F�u��$�����^ִBz��Z�L�{��Vm1����7�|��ᑰ���U�� t?/^]�7߾�W�_0�����!�ϟ��<I�
��V�_�f�����O���(X��{�vH�q	�u�@��˗r~yI���~c����[�閕i��ܟ�o�DIw��H;�h����_~���!��%}� �qO,؇�G��]�H`)��!劃�C
���{����θn܂� ��>%��c@��`�36_�g�OϋrM � �|z�����Z� ��"%Y��3�����k �;��A	׉�\0M�� 7ޠ�@ ��&���}��9ݻ�,�S�&���v��	�}�7����l.4L�^YA�����@;�c��	����K+ V�왁���v��!�V�
�{�Adc��HT2�`Oq��g���R�ߟ���S�����M�In���5��Nρ��S��+ ���,6�:ߋe5�أQ��Ƥ�.�����Zh�ޮx/qmG<(D�z�^�t}�4�~w�7�66�� D�b}[�!�Z���,�	�T�����j�����N*l�� �{����.��ؕ0B��DK�*�W�Ѯ���S^��_�����g�_�t��M�r\�N�1�>ڹ0k�::8�LEΪpks��vч��<<ū�^�����,a���ӽ���UJ���R����0��a����v��P���;k97�mAsm�TLO�+/�"y�b�G��!��5�G��ENA�v��X����Z��`��<Am��^Ր���X�UИ2�4��N2��_�P�v�
9T@X������u�=4�_�2�j�-0 H�S ���C�G��*`V\�Q��4/����g����D7Y�-+M'���J��Y�����`:y����"���hw|3�<��?�O=������k�j�B[;=9|�Z={8]�x �1W�xMOG`�f5ߜa����]�S&�:[4%���F~;�(���� ��Wq6�OsF*Zg�M�`�ZmW\������q���^7��]�a�6�K+�#tTm�B�y��UOo��=g������t2P�- ��̴:H�D��f��E�fzb��i�/�Ŵ��`��@���y����Lg���zVm�:��L��S6Ϡ+�P�j��S$�1��Rp=<9M�u�6~m���`si40` -����*:��-з,>OI�4����y�XlC�����_%#5�-�J��b@��'��w�2n�g3q-ӑ�^i�7\���A`�&iS�
Rm�iϚMmm팀�)M���!�a(���FjV2i��>j�s��A��@��9�;0����5"b��ʂ�M��6g�%I��&�HW��UiNi���y4���8�����Vx��������w��V���"�B5��j-w�h�:k�^A@�V�i���t���	j��F��P�{�5+Z�,װ��4�eԴ��|Ě`!D�>�\���)f%�	�r�2A6pvo�ӝ�M#	p�@� �6dL����{�K��LT��ׁ}�6Z��s�s��2@�c�3Gj?L#�h#��M����7����������5��o��3�Z��_܏�bb/掶z�ς[~���^Ir�G����_0�5�/��um="�5%{Zi���^�H��͈��γ�WEI�
��gk;�k5�j�2����q�.�D���c�#���;t�^���(�:����o�&��{z��in��L$�[���*	hm66?��IF���k���X��_�E�Rv�����hD�h���)�o���:=Ye�R�ka�-r+	��R:��Y΄ʗrs]@a�s��W�1�v��5>#t-(�lk-g߻\I5�/�Q� í7�.�G��кdЛ'S&����h�9����0����?~eV��W��c�tK'�xY�Y�,Tf�A�5���L�����mB�K'���}���?�3���w�#�dGv�b5��1<u`l�`�"��AW���i�dBq��[���]�V1~}�`��+u��B�{��?ȟ��'�`�H�䓣c��O?���%O�>|H'�[���.��l�J<8��39?�bp�����|�S6ټ��1�HG��ӥ�:a�+�?��n���߃u;Ls
�./��"=P4 /5:�[cpT��B�0.8���|�F.�.��n�u�gHu���:���݇��wKA�S���Nz��|�����?���)��k�6�X<��}�S�.�Xa��7V���P�����7���� "�F�X?77w�ujۿ��6�����@uy�RNN��P�*��!yH�
��w�?��Ӛ�k�A%
#../�g�>]�	+��<~�� 
���{2u󧍜�\y��΋�|�����狅�y�RP�u}�)��Z�W�8��v�TC�5�=��ѩ��]�{�f0��H��`;�X��~���Gi���i@N�K����鷚���a���n����;��_i�6
uM��bƼ� 
��U�#�S'ggt���|�Lq'�5uydi{�*��s����,��57=]�{�4����+�t{"?���\\�ӳ��AׇT�qZ�`ݼhcޚ���W��>�׼M�m�,RWi�?̀��K�1ӂͼ�� J����g�����t�߾y��d1;��Z]� ;��)X�~x& �(XL��<ы����>}~�$Y0d��)����@� ɜ���7��Q��x;���^�}��7�m�m��2,�6
�M<'�U�&�жZSv��kŰb�	���QJ���)i"L*T����`�cuio%V�0��`��a�&��;li�B�n�*|5��L��F<�x�sS����jz���t*q�P���"���|��y��/���
҅�#o����W���7���	��^a�B�d�A��:aǕ�e��_0^R�%��\F;pb�;7],�'k��w�6���F�� ���J�Q)@*��ot46�_���:)��0!��F�\��P熡��J:M����F��6��5�Ĉ�i0����86?k��&�xŚH{����������D��6G{����@Kg��Ni1n��yX���.mp���l��fS�oSi�G'3Ք _��i,��h���\�l$j+���8�I�vƴ7 N�*e�.�����\a�	��y#0N�_��#�ҔM�&U`.��Ѫ�Y��2���5�6l�3g����������s2:U���0S=�Ī ~���y
�	 �{�� L��j�4��������7
����`��bq$'�=���Nb�xڜ+�'�b���n��8ī��
a�/..��7���Ɂ���^�g#�_(��H�&:��fѱH`�-�N�D��)����?��t�9��ag����o�����4�GǇL�~{���ۻ�L6�*����U��3���bڐucR���]иޚ�׌^#��s>�0��Q�8�a��9g � �����i�w�il��mЇ�7�&�,�F��)<��`A��ԼW���;h�T�I���߬>e�h=��L��@An���HX� ���c���\�>J�W1<�>S�;YQ
�4/`H ���w�"�0�:K� x���{p`F���t��RƎ����,�2&�j�
txpצ��]�3���� �g��'��\�R���Ր�M���z+1�t ��~F��4x��>���a$�c�W���u�/�0�����k�a|ԃ���(�A@��qNZ���S��!��*P�fͽī�9��!_�(�i����K���7.�M�\�=���PE�T�e��c$�1`Q��,�}>EJ8-������_��x��������o�uR�ZA��޲` Y
r�g -�^'�5��|Q#0] �FU^[�4�Gv�Í�;>�o�;��j����*�7���#��o�=~��By�}��weq���"���Zu����va��IM���6�犚��Q����,9�q`&Y_%y�2�㕡#t���;�cV��}�tQ�
��+��Z�ͥۼN�^��<-�v�����z�R�S�'$�Цf������ BL��E!z�H7�9�@�}�������߲g��}&x���c����>|�_~� �?ko�$ɑd��{�y_u���������+��P(��i]�:�"3.w���T�ܳ��ΐLttVeEz�a��T���w���-�ia�˲=�:�U���x���v+�ڧ��@��%!XV��UBC���k�R8�&�¹jc��%D8 -v���Y=cf zO p� �����T��^^�L):�p;;;��@� Q3�����Qr��C�%J���ұ[�E�+r�v���Ό��*�5��J"l�Q_�<�����qg�/��:9��d�?���&���f��- @��0d�Eǭ�`�@������qFl��P�#�h4��q�"zd$G$d�J���v��T���C��NIP ��{�5�♺�n����斥J�⢌|�;��m��<�?��_*)�f�Q�\G���E�|��x�lS�D����K����ew�8͓�@�(ҽ����81��Ժ�̘%����Z����TȒ[�T�l�y�������J�nҵaP�-������C�x,T�'�g?Mk��F	B��n�
RO�<�z�f�@����R�0eG�ʘhv�P(�c���"S�^�(��ǳI`3�/J!`䜍[R��"�L��J�X*@k��U9�Uq$�+��(�1�UY�������7r�����徿��.=tlO���3&��5��Ӛ��,�M.5��z��R˙�b)�l��X1��E����Cj�޻n[K��h:��lX�����ؽ%���{�R!��~6��0{�rN*�V���
�m�zOk���u��G�2%њ2p�ʍ�	�*7K�u?�dt��p�y_�/砗��s)_A�]�����|iVC��_�[_�3��x@\`S-���샰��¿�3��*��_�����.��֐����ɞ�#�������U$�����u��H]~ȿw��fyE2��X��h���` ұ���>��t�@�u(�w�=�)
�1?�2�fz�
�<s�K����Uv�.ksʷ�Ŏĩ��i��}n��S++:�Ys���H�1r �ReX�(��AW3@_h�WQM- }?O����rr|�2�v���iS�����A~�x*�N/�<E� �#�� ~鸐M#]�Z��8��*�����P�m2������2~�H4��t
�D��C�9㭃��b SG�Ȩ�8��P�|Ha���k��E�>�hU,SĿ���	���@��H j�7=nſW�~8�go' ���D]��P�QPb:|�l�&����26�]G
;��yo1jgai��8ߡ��������ڜ!ș�S�<�T�ų�1��&�P��KŹ�S1�1N�5%�����sݰ[E��|��cNT�	���p��� @�nXl���l�E8G ���P�n�`����a�	�ꔢHyF�>l9����&�I�������`<t���`>�<@:4�ʠ:u��d�Xg;n'@�� /2H**�ZUʭ��c�����ӹ�,9S��;��
��"��Hq��a�j%'�0{׶F�,w���+>;TR�5
cr��(y�����v>0mY�ct\��\Ҍf���e�� ���g�ӫ�ͼ���55�Ɨ��ߦ�3e�Ȅ{Y����f@u�㒍#w����RuM� ]� ^���������^����1�����=���?VWh~�s_Z~A0��h�NO(��B���vb}��Y>63�Q�nL.��3o�p
�7����a�Vl�RN�'a�),���"'c�E�����u��P���ҿ�ѨG�����[Կ{Y؞����pRW�z��$�3f�Ѱ� �G�~�&;-1���so%O?�CH��7k#E��b��pF_��O��s4F���,����4V���?
�q�JkNL#���+t4E����Q��tج:
��7���P�jG��J���X:�܎��U��[��g�HO��R�L#�E�hY0�2�j����BϹi9��|d�pc6��0~�i�Lg6`I�q�ȇ������Gy������䆰�.��d �ڂ�����'���D_LI@�*h*G�l����6t8*��i�cG��Xf�4�nKd3P^�"���/�R�f?�J���5k^c9Вi<cjcqr�^�ީ��� �cg��i��jC^�ы�/�
wa|1>3{��,G�D1��[0
	�mg{Ǯ�v�=g���s�I�5I�6hY3;TG�ȇ O�yð�\��ej��yHc�,�/M�ʮ�i�]���bG/5���#�|6;SCu�@i�rڮX.��k[,��#�����8v�(��a<���Z���f��hr!����\�G����D��n��6y��wH\����Jm�3<�h,��������]����ܗ�G;��7p砓���|���%��������>f�  |���kd��t/'�7M�?G�
�:l��`���v�0�(����|�y_�M��u�]���=NuX�<�I�ss���[���1TX��
ff�3Uֈ~��l��&�vS�@��z��z� ��i���⾈o���Z;<u�����*��h�gѶЅ�����._��:�&�U)&��º���=[���t]+�iC@�`n�Y�C�U�O>c��Ikbզ'�������Wf1a׃�hK�����FM5�����]E>�H$(6�^ѡ��B��U&}�\3O���H_��?�
O�1��<�ǝ�mX�4b���<��6,t������`�x�1����������o���~������xIͫ��ԮYP���.�CC��v�v��y4�?*�ѳ`O�t�	�O��_!V��dt#�s�z�������\��fZȭ����"ŘV��M��뛬P��s�������oԒ��yk����0�K3�UY;v]��4Br4�lRsݐs�⠨�Rۮ[Շ۴���P;�7�\s���=x-�Q�D��� \)�ǿ�����x�b@�ߢ���4�>	8q��Tհ�c�Cf�;ܴ���T�ͦk�✭j�!rGW� 'Ϊ�*����(jIk���"���
��M�m��nOL���U�؇�I&�g���}$Zh}-�����?���6�]�@u����:�
�R�k�h�����/b���6��z/���h��G9q4��=*ĕX��l?+=��LCe�:@��0��h��h�����ǃ�f}zTl���GK�G�{��NR�K'�7YP��c
+%R�C�c�Vu�saU���� 9[�-W<���b��`��p\�y� ��/���@gJ��/s�m!�7́|�u�`��< ^\Á����U;��Ui�$vk^XW������S�<�a����6���g�#�l���&��35ehT�C��Z������Ps�?`Y��M���ۜ_�*s{N{Ӛ�]���rb�T�{�.�+�G�,��m��w:P��߅��C~>}Q�iɘt�ƺ`5[��tjB�f���Z�3
�4���~�-�Sb+�S[��J�gJ�C0/��+�Vˢ^-�7*�N�aBkUp_T�π�Bk�Ճ����^��uջ<����~�A��g���>EE|��gc���}C{K��B�DP�ye\��驧�=� �����ד�����֪��Fǈ-�dK3��^�����}
��yr������_Ԡ�h�H4S�'�4E�vG9�2b�z`�ˮ����J"x�Et:��4Zb�� IB��k#��R�-F/�S���y��E����ֿ\<�e:>���t5����� {�f��F�Ũ<3�a��O����^e�����z�L�U�&�m	h�R����L?_0>Z�����MĈ|.�2;ĜS�ȭPa��``�J�3��{�����\aϷ$�����t[�-��m�l����#o732gv��̰>�v�?����JaQkӴ����0�F�o��S��l����0����Rn�.ٱ�� �;7  ���Dv�5m��� 
8�>h�lpsYj٦b�M.��g�Ɣă����6�FA��K]�X�J��9�����f���ݬ�t� �f��.���Q,U�]{�Aen������'[�����Ŝ
��P�\o|跈+|C^b��ԅ� �_t�w������X�26,AY|`��"�x�M��N'8m��=����6� ��t+�[�	����4����
:{� f�R�)5(-b�ZmG'�����
�rx::҂�r����
���r>�06����^ `��tʢ����2�%ߏ�Y����fD}
\K~��អ��wv�������D���!J�Cd\�rA]�E9e�{G`��FM�},�\9�(����P�
`���1�o,z	a������2U�<8qi
�jgy%�%�%l��f�Ħа��P|)k-���)m�e����@x:w�sH�4,�J��@h�y�z�����C��`o�u�k��6�Gi��	Յ#f��Q�#�cz�T�TST_L�7-o����R���/ݨ��'�?����N������d�5K�HF��rQ���FJ�a�G91��ӳ�*7���T	��Q{������\��l8�4�&g�=9��(���{�\ӓ_�����?3ޡ���m�E(��ݚРXYHED����L��v=���A�Ě.��ܜiqTgQfV���n�1�:�=���7J �앂�$��,C�(xD{�m�%�6*)�(����|̱h�nU�2�P�4��o@��cr���Z���4A����^��KF�;��A�����g-3Q(�P�eהNa0"|Y�Q�����s�cU`�ݟ�ٳa�:[��O��{ :�k�����<-_���J�P�����g�4��/�p�<>�)�s�d7a|��B��ϋ$f7b@k0��9Gs� +'�2�)c�(('���t��f��jm8P�� �	r72;�r���-�![��� G��DW"G"��ٍ��X�e���Խ���P���T���iw�ކ�|��X�yf�(s뾊7ʏ�'�KT։��1���bh�q����)	�}�G ��Q�df�J���V��,����t�s\�<H[��ByI���S#��a @�j��mՁX�]�y���:��r$O��_p���K���@��$���ު�Ԁz��gA)<p6a�u�p�RJ���w��B��ۃ�(�|��o�����"5�ށ,��>z.��d3H��Sș�.���AgDz,f[k�Qo5slFm��4�3նP�+�������&��d��wѩ@EE�];2w�3ޯ��D����M7s��>�e<�+�����K���pmw4�����օ/�������(�g|E���V=Z��M�BF��� ����C���V�U�zϼ{�������_ ��2X�d�����:b�h٤�rNˌBdtLȎW��_�M�[���;���;D�J9F�_�E �"t�w�x���ץsi�#Of�ll�,�-@��5I�/F)�N+��g4�z/d����h�=�Di
�ra������Qu�3AV+��@�n��I�0V$��o`cIԙ����C���ܡ�k~hm^��3�`Lc���2�dJ���x�9G��V����*��u�`��FD���Su�4��92� ��t��.��Hg�L\T��-��G�V^e�OP@��1�٧�l@�Y�<ZF��@��=�Xe�+�]�2;s�6з���� [0 LԖV��w�r������R�e��U���D�<)�y���B���-]P�w���[�f��6��E��z���V�M����W=3�,��A�nk�4x���*�c��<�R/3bO@�{B���\'���lLs�r�ā� 0nf�I�AG'
-����"�vp���`:\�<x�ôn@�Gwf�Q���6ZX�L�yŌ����֞[�xIZ���	f!�
��.=�{̀���Zې��s�3�.0�!��}����-�B��jv�j��U�pdf ����l�(�(���A�Z�oTD9`�6����������	@S@�z��R�h)s�&[cߢ���o��L"�	��}�Qff$BrFϯ�6W�xY&�ٖ��k�R�+^mm����s�U���߭i���~L�ͮ�^hi��)h�/t��4����H�`��5� s��5�`7k���a �����k���l@�	��ݭQ�,���*�?W�p?���vic6���6<ߢ��(,|
����]�T��7�������+;��U�E�U>�Vq�X� (�E}L4g�VбKkA� t������td������.~g��eq��n��#��v�sB{(������WY���uO��ί����I�ʯiT�1�h, æ6F@fx��n����m�1.��_�P����1qW�1�{��)��"�����; &v��L�]9k~�r]�(��l9E ��R��ж�����w+U^�x�]ya�1�YA}$���=�`u����rh����x�`�rT,9 �Zf�Ȍ���
�:�P_���l�f�<B�(�_�nD���� � ����TxZguc|����ћ�p'�����l�6�_�."--+1:�w��ٞ�{<�{�5�c��z�/6�����d��j�{f��L�%���r�q@.�F�<$0����t[�b{ N$�f�֙�.���/��ZTEz-����Q�ڢp#���B�wEʹ��,�Z![;�lÉ^�;�qxwwϹ�$q`��PU@w�c���l�Xޡ��i��#�0�>*-��Y�d��(
j��lP�����-�� ���a1��ކ���=�JAc#A�#5�m���S�W ��	T;�9���g�90���5�ϰ�C� �7�I�Z��jZ_�B	ɡ�A��6X�n+]G�ު	�!����\���'`�dc��t��>� ꋶS�Oָk"�3_F�S�,�x,c<�Z̝�js�~��l-�t:_N	�r9������^�uMG��&viV6��d�W^�Ժ���<\��43��I�|?�n��a1�v$r��fC͗�8����4\ں��8d�%7�>|~�n�⡐��k�ߙ���}��
ժ�(����zS�4��غN`%�k����g��P�Y�#�3w&N��Y,X�0��	�=�F2��'��3`��j�C�ݷ�������g:�U����9�(��)1U���>��J��#FuԊ�yi�~˂HN�g�����S��5�
���h �IS�:\�C��nM�ĵ�Dr�hY_M΄8��KʥI:m�M�d��n��{UZ[���!U�5�xv,�ə+3�A#T8���K�p^ќ;fZn0������XC�	 )|����=����-�����2}��g��2���T�^��� �0�g�(��"�' 	
Z��[�����:m��Z->9��F�m!;iSl�K��V~��b�ߠ;.\�%c����A@b��1î4"� ���W�t�Wk�"Cm���C� ��o�5_�/G����]D��OG�yh�\*[m��&�r4�5�陭�t�ٍ��n$r���HȚ�����I`
�mԥ������k�3�r�0�;}���}�y� ���Vij�qQ:�Z�ie�Xv���tdz
��>�S�# r0/��������r �?�qv���L��C�q���:����
ǅd���=��#:`x&h���::zV��-[1�C����p~��}0� \F����X�ϣR�(|,J���$�u'Wio����{I��Y�5I�
�j+a8���͍/�S�"[Y*P½Cf�E-'�m�3w?��`��V�ôf�������e>6��l�c�$W`��[f���%|���hD�ڠ�>��̶e��,�q���3��㠠�Z �s�庸���u��*� 4�]Ե6�hU��e��B����^hp�B��J��k�	�hH43f��Z�.��>ݻ��6Ѹ�e�Z������hR�ea ��u��>+X�)y ����ִ렁u�k( ���Bf�M`��q�,M�?-�.���z�
B@���E+8"b����;��E:Neԍ�����OX�Ǵ���#N�3� ��d���6,5:�����i��4�6�˷X2%>6��cy�;z��tM�X~Ҁ��@��K�JA�
�U�4kh L���+h���Wa�/��M	�"�Y� �-����qX�}�O�V®���}�p���
5,Ťi��� GwB�X�Sp��w��-E������+��2wY��g�@EC���y���!`mG�8���>�ʤXP��h���C;5���+�r2�JED+��(ʯ#g�:�����ݸ<0N��[ƣ7�32b�?��S̰�F�j���j���l2�����b-h�a��{���Q��#��*H�W]&׀5�1dP�;�͚ʘUa���B0R�l�sF
ˏ��E~z?c�DI?ʖ���^kd<[婕�K;bU�f �jI��V� �������单�@,^�V�MC�V"�d+t(2�Q�F	�^ߘ�f�8˶��j+.7�*�������	�����mU���YP.i��6���l�>=����[�|4�JN|��<�F��}���F��_Ȅ��
Kt: ��6��3��j�X�=|Ƽ �,���˙��e�q� 	C��Yz4^8k�^@Bu�R�; �1xn��	�r?*��z�IK�ps� �����+h�@��.>������{~��dc@y�vp}�λ�J�wr�ދ�tm�ǘL Јi7�s�T��&gY�o¸���>����s�@l�
�j�uuqu�L�����|&gײ�@,����N��a�K�,@l�f&�f�I��#�����-�-Əb�)�����y�>��l:�/x�?�Y"�A`��U�EΕ�����"��a��MDvo�v��Fy���tG���6��lkiY�'.D} A�h@��9`+C��d�
Nm6��bu)�_%ht�)8P!S����ZY�c���!`޹�=��|�\��2K��=�M�����ָ��i���ۘ�=���k*�*��>��B3dX�|6���9bma�]BkA�e��7j���a���lr>�����oo�����7V�ZA^���e��T�<�h� P\������+�,ד�Lp���� Qn�k�|6mm �隫ⓣؚiT�>�Z��rVZϿ���Տ�'K���	��-���jt f�i�	�!6ڥU���ۥ����^qm�>���xpUO�u���,Mݶ���p� 9.��� �g�l��s,�%]&��wt� ��mn����������*gŔ�L [�-�zʹ��55j�;Ⱥ��	��!����"��HZ��T7�&�G �jY�J�T=�e�2r 1Hׅ���{�2Z̼��2xd�~�N��-�j��}\�$�y��k-*{��g��&���QIڠ��Î�K������ ������E��:B��ǳQGH����L���A��%Į�"[�aD���;4!�<�[��1q�`���$ �UBi�Fx�P�L�ë��q���<��0�p,�$�� �~������9 �qCB�NA�)�������\������yP2[���Ò�5W	�`�1�����ë;^�����?��B����xk��ɩ{3Q#t� �d1�$�e�T�
?��L��/ӽ�tz�����Qn��r�@Fټ��\\�(�P����kf� 9zf���|��:,������$��V:#�l#>|!��ų#/��3!U�%%����s����eV+(��6� �+����@dg6�%�׌����3;������t��[�8ܫ_����۱��7iF/�ݦ����TΒ��?��,8 �����SJ/����O��l�;���O��R0�&��а�{�u��T��/������L��$@�3)���[j��f�+����mͬ#K�2H�`�&CPj�@bͮX6e4�	�@����*��3^����H��ME1b������z��*���tZ,�(����\b�v��Q�ۨ� �{Np�w�u��Y���8Fa�UJ�IDs�V[�N�=�M	�8@�h�R+*'V>t���3�������6mzOzV!��5&����%�1����+n��e�d1�T���.�h�V\G7{G��r�������n����6��aa�kU��E�<0�fD�eS6�uɢ��^2���ЍC����X�I�RvP�@���2`�01�n�d	���&g�����3��I��I����o���̗���j��	kkp��[�"�RNkQQnVƫ洣��H�yc���o�hiAi�\k��U���d��n�H��f��0�3`������k����E�lA���1�a�{,<�\21Phm�<�w��`�o�꨿�ܢF��SBYm-���%�r&�$}Py��R ]��k���H
�²�X3A����ݤ�[ ���j��k��}H��6��ɏ�gj$Q
B����@q$US]ܻˊ�D��Ƒ�yf�6J�EUw�l
��V�|�;N�@E)	�0��R3oQE:qI��E�Qp;�XZA�>��%� �u��*f� !)�;���ه3�n勵kw/  �X��O�K�G��{���Q;.1���R>~�����`Z���ҵ��.䗷����Љ�ظ�#fgg~H�������	�(����/�7,�_L�>X&�yIQNྐྵ_����������ށs���2���Sx���#�;WV������H޿����<��c��Q'0rFݠ���%>�s~X<��ߑ�5�\�Y`�8��S�]��C�' �A����C�g>�����<}��sF�*�Zt)�g����c]]\% R��fs�p8W7 #�rw�T�Ѱ塚����h����Zo~��گ�k�H/.n�ҩ���=�	����o	��R:q����C6�:���&�E&�#s�2�"�.Ι��M ��p����P����Tq�J�h���&�C�_�8����Y���/��Q,�<L��g�%��qPEE�iT�;ݚfU}dy�(��s�M ��L�7�5>�P� -�մ��#�d���	J�G	�Z_i}#@Z2[�5f�g��HP1 �1IvjȀ�JX��4c�$��k�/�? 0<��"K���O`9ك>LXG�3p(�|��{	R�ׁ{B���{��=�;�N�=K�w��`��h�	p�e��7�v�:��cˌ����ݽ�?�)�@��?�jNk �%�p�����A� nҚ��N�� �y:�L��h�}��Ç�j%af֐�Zr,����s�;����'��(v/,�I'�' p)Ӭ�����L�1w�]�-�#��(6bL�_���H���r<���΀��;v�b����M��D�5a)�T��NǇEjr�x�B�������w���{0�{����4qR��<�����wzv#�S��贰A���Z*�t5bs� ��@s� $�MEQM|����h���T�܈J�oyO*8�ɃjU���.a�t�YU��ƍ���j�pv��*n\L���D���3���Q�cCn��e�Y8p��qE��b�$A�P�h�l�i��������yzÒ���!��B5��f�|(%��ąu�!�G���NQT3I�l��ad$z��C�����IWƳ��Ua��|%�w7��M��A���/.��}�f���O9�Ϟ3��� �:�N4�/�P�B���O����.���PǠ�Ͻ����~w_���������sf�\�[��ˏ��FKk��
�����Y.a�f�!jP/����O�%9�b��R$��98'Y���Z'��J�Q��â����A�}�̬%��|~�NJr��&�UC�\�xJ_y3U���&�������Iw){�qT8Qdl���o \��0+)�b���g�0�9�s~\>��N��P�5����\���C�(V�m8�����o���@!�
n�<�(��6���!q=ݏ���
� ޻�-'��'� ��뭖H Bi>}G��K�%����ߛz� �vX�6�q��9/����`*�z����⃌>~N�1Pm�,�a#{PB_�ǛZ;�8pr.���\&���)��y��%����%A%��[���B�)�#iu�@ʤ�E�q<�k2s�hp�~��Z��;� ��/	��J�P����<��1����4�s�@���rעf�*�O��%�=���K�a .d��l�9Q�_�,��8��#D`y�������o4��.����>VF�p�-*��`���w�Y�}�IN7׼�!��۰���c9<ؕ�/���a�xA��)�o,}L�Yȇt�R�ί�����G�?;����j,#��A,�K�̓ţvg����g��vd�oSp#�9�V0}��˗���Me��F+Km��!�������Lvf��;��mz>���S��2��Z�yu"߾y���V�E�]��%g<�S0W��svMG&�lOTH�[�k�JWÌ���!�8�����_��W��M$e��m�F�jF�6dZK�T�V�ށ�M�E��YR*�wX���<��y�Y�F#���b�����[$kج�t���e}�ݿuZ�wo���?�,���iNd[@>G�U�Q&{��{F�hU�n�u�q�]e�;��.B"3�|a�K��� ��W+������P.Xa��*�����iC�`�Ul�xJZKj�V4��РѴ_-�C���t�)�<I�i�z�M�Ե�vYj�4 JcmkI3a�
��D�Fŭ�Æ�;�K�f��B��wwv5�fC �FBp�(m)ɹ�R�r ��Q��A��5���iFQ��7���c��Lfr��Ŝ��I���/�?��}���]����\�2֨���/7��m����G�v�3����[�{�0���F��A�	�$W�u2�#��]��������`�@Xv� ���X[�ӛ	(\\\�</�1P%E�,���.?�z8լ ڷ� _��Vk��*�f8]�-I�t�(�=��zI��n��Ŝ��̴5NP�Y'˞�?��w>O��R O�⃥�����p|h��OeA@�<��Λen�����[�\��R��p� �?�&����,7��ڥ���+�C1�$O MCp��j��l(EQ�D� J��K#���=�UX=$�v��F�,FCn\��k�14d�s-��%��[%��!p�
M��}��t t A�Ռ�4��ߖ�l�g�J���\�>q�h�V*�A�Z�Z��$J�?	��r1��	�p�u�'�C����i �^c��525����9��2�g ��ٔ6#X0��
	�����ݗ�t��طf���Z��h��#����_�oE�ղ72�ؿ��P�t4�gǻ��ٱ�iv�4�
� �s/�yi&)�=�QH*^
�җ�k9Kv�J�p N�U8F�;Syu�'��L��v�F�<�\Np��+�ӳKY?�K�jL4Yyy��"k_^<?J�<d�����J%�	}3{�jI����p$�S sz������,�f�&�'���L���@Y壔�s��r)�dS�r~vE[|������[J�,�R��� A�&qT�G�D�J��P���} ߊA�ξu(C���l�W�#��?k�UoV̙3e�W�E^nqQ*�r׬g=���-.�g8Wv�97R����4�eI���O,~����ܣ�����j!��l4 ��H[�JP����"K�q���x��p8eא���V�V�K���=��@��:{?S��Q	� �>��?�*���>E�?���U]~�Uģe/@0��Хq`��1y��8m��JΏ�Yn�W"��pH0D?��ڴȸ����}��W�tͦL��^3n�4R?h�� ���8�9@��W�^���hf�Tk��������Q��F���h.j64�X��~�NXe���Y5KF�8���=yv�>������QrD�I�,K\^^�H�"��Ψ��Ǧ�����N���d���<K羓-�!���Z�U��-�0b��\���/��,��[��29��k� C]���2�Ɏ�\B�-
���C�h
�N�TM�Q5�s���,%�3�c�%cچ/6ܠ�/�-jW�J��CQ��C#����|+���1�T �J6ϲ1@� ���Q��ĉv>^U�F�G�mzmU5a��nTo(���TvA3�J�.���D� �3!�wK��b�1�!T6�
6Z�_ԑ�k�Rj���X�<��&}ތ������̭k�
�آMJ�fVe�HNi�Y͢*s�8;�R�\���f[ҳi�u�D�M�۠���BrV�U�*F����Un�;,u6�,��YұT�6�v��X�/hGfYz;��>��Eh��`��h�`��}�����#��5�~�X\�(�4�`"���OҦd����C�� 8h���������y-��Q���`�_���hي�;t�
����C~�q�+?��g9>~fݺ��&��wR�	+ڐӽ7���)�lՓ�c���t$��}����rx�)#�0㾢6]���r����cp^Y�j%�������<uf�@����q5ώw���N�����*������}ؚ���ݰ�<֫�Sy��2S�]��l�Ky~�'�_��	�}QI�"v]��}B-l�f���mJ�n�����)�n�op�������,5�Sx���˲��Z���ѐ�	�#|'J�x���^\�u�y
Bo�������Y�W��C�j�l�&���&���{k{�t��ev�:�N��f��dH�R���N�V�y��wɢ�ܐIND/C����V�F��r D�Ǔ������,6�JĘ?�)��ʌ��3��8KB�� l�DJV�~���ҿ�tv��t&�	҄�I�̜@�d���������5�����������v%���ſ���� a�ίO��r���0�%?6��^@��rnr���P�N,���೴;�Q�v�d�@�^��9�4(~a8k��� (�6>	�Q�U�{yL���<��xS"Do��+ ���8���F���/�͛����30ͮ�|�����&�G7b��ϐ�ߐ���z^붵���L�})��+�g�D�;��"�7���7�_����`�l�E ��ζ�����	b� �c�:��BZ��o��?����{!S���'Њv��o�D4.i]p��|���vpݯү,��39�l��(,m���в�-�S'Ù��" �uS��h4`p�	~/=8����\��H3��h`y6uc��'j�k �c���^Bԙk�E{��ui��6p�P=S�W`p���*;ܘ��7l[ǵҐ[���"T���"�ֲn�@�A74����>l�v;V�
�	 �ҳŚܞN�^�=<�R�a�Ѯ���杂��'�q�m�1<�!�I܎1@)u�g5�6�LuP�M]�h�mԌ�f�4|ӽmov�t��i�m�Qb9{�f�]�T"x��Z�P��޵��+k�w.��+�9��K���	W�-4}/W��ϸpm��,ҳ)[m<ea��3�v�N0d�5Q�ZR T���`���qh� PRC*�l^a?�9b�Xr��n�Q3�YYA�rR��D���ŋ�6^�����}.�ʩ�M%-���t���f`��$J�w�]�-ӄ�@?>ܕ��)m�D� ��ae�\R���U6��,����RW���p���}y��ɗ��dwg�>��Ώ�$�ḃ�p�U��\ov�==I������%��RL�l�(ݟ	�_���T?L:�j�2�ډ� �9g[�{����wa�2`�
"�ȌZtޚ�e��xlmt,��w�u�nUI~�,d		��v���$g�q��JEV]C���V4�!s�F���MBx�Ff�]RE����B��������=��(t�ؤ�f��$�d�Ι�\2��x�D@�'�j�����r���J
������H�#��0�h���B
)DpX`�P @h�(���1�9��y+����3di��z�g�:?K�y�d2�ۻ��@��DN�����y�G�f[��(�3��h�_�f9p��.��"o?|���6Q#⒳�L}��N�_���9Y�f
�X��JnP4݋q�����勣�Y{tp(-��7�&���V��o/��	�����䘮e0�J�m��*��"�+��8C9J�r{2�Q���Ǉ�w���z��))Q�B9d	w'��dW�M��/?�*���Ȯ���BTy^���O�lZ�c�*d��+��Ry$��t�C�b�p�� �g=��$�'�wRt7�O�[���b�H��Ȏ�(��(�ʋ-�O.u_��ӗjZ���@�8Q����y�2M��K$w�~�$Y{2���:I���54��J��RC��Buv�|zNDL�-g��c���t`�j%�̴'���k��,@'�e�R"�2+$h�/�Ge��K��Y��:yè�#�lD\3:���ȺbB�0(��%��Im�cy�,kW �g�lGlY��I5-	r{�d	��$9���>��ճc9��%����~{'������'�[$C�T�R��PZf{�R����o^�H�}7َA�l�6�ۍ1��UZo��"3��"ff�<o &�Kɚ}j�79 m�ܢu�z3�[�ؙ�h&�-������
Ŧ���{��h]���C��B��,�ɵ���}e���޵��+>�2��S�`&U�i�%����Ո��U�8���R�YCs��u ���zT	
�k�Y�%��vw�ͫg�6=��(&�p�f��O^�LX~o���`���^Z����T��_~����"2��z8E�K���V���s����5AV��}΁ݖQnŻ�kVo����N')G �Q�.�[,��= �m�!G0�����=�Q�NOɟ$UݎЏDً�:+Z&���J�$����\u2�&�w�GJ/��X�s��q���,���k�m����]b�j����:�J�#�S�֐O��������?���\������}�O����J�� �U
�������>J-�Y�cE���x��*q.�4Od�Y� C�q�������ڼ�L,7 7`p��,������'�w��7���]�N�ρc�ө�Q!`�,����ͱ�P�&:�f6	|��@Nt�F�7��hs��ո����2ԋެ�k��e�n�~D�P9eh���tƋ ���H���M��Iu+ެ��&������r~��[���KJ4V�X�t
|͔P�h�D:�o�� ��EL���%���P�f��_�������H��˹s�J��h'Ek��H��6S�9O�mNT=�m'06� �D̝C��˫�{�)���w�{�4�
�="�<I�g=.eog��ۄ�x�rz)7P _�R8xF
8=�� �Qn;���w��#�c��ͫ�ߞ)!;��d�H;��	���!zK�]d ��&0�ݯ�!���c���h���:���Z�h�.l(�K2y���z��v����9�8dY�u8Us���|�����i�D�E5:�R<��y��������f�w��H�U�Y��H5B�~P3
 �-�A��J-r9�I�jp��4,#x�&�s�\/[����js�<�#�t���H�ln���I�;�d^:�-��7�_$ ����6[���C������="�F;oE��)J����ￓ?��MZ�3�׼�%~Y��$����g�vbl�#[p�i��^k�¾��f�<�e�w��,���#G��m�{���v�Mto����H�5d%�2��i�e�ܱVu�$�=�)���#�=��e�bQ��Ԋ���~5{i�5>�vh��zi���ь����(��䈩=׊�h���s��u+)K�j���A
^��A
b�v�S�����L��b�)6: 2]/��'���l��o�❵�{M>fLF�$z�ݤ�:R �h�\��J�ʩ̸���~�j�6L��ˇ�?{������G��.����Ȧ�l��{Z�މ6��dFh�u�lr)�d��w�xw��P�r#�I��|��{�^,�� "N!� ����/�����TN,�'x��HE������<����4j�ݟ�Wr�����lQ�@IK�e�,]?Բ�\�^"т�r��|)��d�,�������ңڄ�����;���΍pt���;�1e��9_�ϝ��q�`4*̀�J������]��)��|z������]�,�]:7_^�R=�;�|G����^��a
�b��CR�C�X�VG���/����Bwq!��t�a6�"I�i������t�d<��	�i9x5�((/�`�� ���̘�aT�*��\,���k���;���I�>�&$�7J�i0Ml� ߄)Cl��ˀ��ƴjht��$Q�.M����1��+�H
}�Z�j���F3<Lw+�o������]GH�Nj���d ?���.E�ߤh� E�	[ɨB�M�V��v[V1�hq��6�������������_���_�I��aQX7� P�c�yy"?��&Eu���<�s�Z���0���,M!"L�ut�#ۻ�����.��������̦�^BXV�$@�j8Q"�� �:)�b�K�0l �{{{���+f�nn�x�	5 ��-�g�fqTju.ka�ԝ���dT}^�S��g@$o�`\-�!�0v�#�kM������N�ٟ�v��d��F|ce�|O�d�e�=�ssia0��\�iG=퀂m��g/wEK�q܏�X%���ҎZ�Y.�� �?Mk��3 �o���Pf��2�.$���g;^\%g����V�\)t}-sF�/���/��[y��X3ԍKNr��=7���6.�܁²���K'��~[��%_6�\��������:��s:�u8�#�N�Y$��RI���>���4���CZN	Q�#�t��2f���#�C�ʞS��M"D�qJ��u)Ш�F�@�1FS�o[_n˄ZV�٦a���I/������(M�rE�U�hbV\�d[��`�͚�V	�\a}$�N>j������3�q
B�x��Lu����5/I���+��K6v�u2�&&����p������>&	"���ro�=?ry��b�mƳh���N����]��h����Pk�Э����Ǔ}o��߀�B����@�����	1(���ܒ���H'5h3P��I��N�E���r����#;=� ��`O�7��A�ส,nk%���{��Ç3������qop}�ހ6������صV�>}�I6�'�������<?�g��'G�_�@�x$�ɱ�,bH�4��1�)��O4P��6�Y3H���;�����.�h���^ų�c�I��2�?�= ��zΖ��=�6����N�3U�(��U�O�P1`E��ǹv4��+FÌ����&�'�舥C=]��#�k�N��9�aF#:�U���X�v��n�2׆�
l�hL���~����M��6�������w�嗷���UZ4+n�j ����J�k�L���Z{�ʥ.L*� 1{<Эc|�\V�5���qpV���c�ݴ�R:��J/�"]�.	|kt��s�ܗ7/���?%P�"�|(T쏒 �8�J?��:[��YrL���E��:K��[vHnt\J�;�����������-bhq6ΞQ�h�_jN`ob�Y���3!Ժ�����5��/.�׿�iD�*���1�t:$��$�Z�ek�����bUS�m��������!7�:٥h�Sc�%�~���=+�t/q�8b��ň��,tX`��;U�&���������`P�>t��J1�%%���"t �_3�^�Kg��m��yb����)��E)������;��}�R^�<&�H�\
H�+��n�@z
�f�JKT��.5̀N����^~��O��B�K��D�ǉ��G���!���!���i_R�u�X��4��t�(���su6d1J#�igT�|v�F���8�N�vlϖ��	��3��NK�;���qZ��-@�u�NA�����ks.�E0�|8���2 D�N6�� ��{�i�a|G	����-��K�F�XD��ʇl<�L�D�p��������珔e'�<����*��y>y��e��8j�	�#Q�*�7��l�,+�Ϲ8�B��R�ͥ��&�h(�Na#/�]��}�L�����K��Qe%�.�����k��|��2^�;���� 8�l9C�Ҳ](��_�)Yd�h���|� ��W	<��xX�5��_�NC�|�y���xL�����%�ɛ#�F�J��@�l�:���>}��l�o���Y��{j!�^���ú�����x_3gG�s�Or��H�}ò�"��"�C�}�`�b��@�f�qC ��Ym�W�@c2B�q��/z`ղҺ���n;����kcg>��Z��e�qs���c J�{��� a{��iZ��l��W����e�������]�*�7k�Q��X4]�o��Ƭ�i��w��.MmL�0�a��c��k4��" �i����A��,�4K͌��FK��	6���b�6���{�����Y�����?�(=����� jㅲ�q�ę�@�6z�!�h}Fd�2(e/L��И֚�>�(˴�{�� 	݃���lņaA���W/y�ۛ�t��k`��(�̳�`�m���FL��I��$\_]�ĉz9������XV��Q�"kO^�:a6cP�ҽ��:��=�ۑ	 P�|	 ���+�%(	Մ��@7���!Ql6zy6����h�O���3j)L���g'���~�^^&#ylF���Ez�y��_ȪAZ��hu�h�X���`)�_�
�z�)S^ސ�~�\6�lDG?4�%^�2~^�uh��8�ɮäU}Y�+�9���n�������W��Q�>�/^���ze��ˁu��ʝ=b$�X������w���^%��'y�옥����^�~=D�HV���mY��6�sFw�����g������߼�d˽f��0�����҃w� j 2""�&E�W�Y6a,?��I��@�{a`@���j���5y ��~@�Y��}Ϡ���:��~֍6	�i�m������g�rQ9��nʪ6��KǼv�����E�l�(�f�A9�ɢ|�`�u��6�Ӕ�4�#���^���غk,{�§�9f3lJm���JPރ���͍���An�o�:ڦ�.]=�ɳ�wr,Ӳ��(CN&� @������1A��x
�#��HwY�=<����i
/�F��j�Z�[�l���t�mV-�&{$ߣk��Gdh�1I8f�z��  ��IDAT��� ��Ǉ�N�^\�Nk����`E(ԣ��ri�N=8#?4�y
`o�o����5�1�|j�=h�!@E����w�B�W���E��ɞ"0ğaw7�9��)�d �{t"��>|x/o���]RTx]�j`[u�v4z��ǖ�Q�{jJb@���^���-o^�ο|~(�)��6zn�Z	����H%7pʢ�A��j|����b����v��Ս]�{��Y�.�ۻأ�^'���i�����,!&��Ky����󗯤ټX-�H�ݬ���E�9�C)�bUJ�|�i�8����A?Q<���bϊg^�[t���L;�D�F��B����r�� ��q.����ӡ�.U/�,�|� ����������^�:M�x�/�e(T#T��ި������ܸ������a�.G��W-��	�Б�������/�5<{~Bc�tʥ��������u �g�T뇞��dD��^����9�^� ږb��`"��SD7���d��ó#��2��8m�ݝ��NNY�E���?	i��YzMY�d��%7	��a��-g�!��#w6��@�L��o���
���#���_(/����K�!�-�����	I�H�Ci{��ӳ3y����.7ZN�Sf�6�\Pv������҂9\Y,K�;�3=_+}0c@+��"��WpGhr���{u�E���
�: �s�|�fɴ[/J�_�S`��{�z�,t6��� �w�=�� �����ٚx�^��]�>3�hPF������o�ẟ |�����[��jr@7V���3��u��E �*�㴞P�Bp��xе�N��#�K�:y����D �q
�vw��E2��w��_��n�	��z\]��ק�7��ݠ��b�ٮ+�Ղcϐ���9 ���B���a��o�u��g`CQ�,A p�Y��GS!o6ۿ�K��&��һ��L ���9���ma)΁��f�U���v�0�4�Ł�x/u6��5�85��3�O����A~Z!\�f�M>Ac��t+ʔ8��{
�%j���Z.g�538UV��u�H��A�)�N������1��\JNA�`j�������w�#p��AX�.�����6a�����<&�����+4��Hh&�8I@nw�T�B|����fL� T����x���6��M�v��Zk�w�,��)��8��v�0�	�B���C�a�Zu���0	��b���}!�07�
��pt�'�;�
�����Ge�Y5�4��T��c�(@�--1�-Y�����G�/�K�	�e����_?�Lk�u�|)*:(������sd�v�����s�{(R o4<J�h��eDRL}:���ؚH�\���'������3r�x��H��� 'G|�F�]a����!��O��;�E���<��|�z�����;��1"K^�eC�����ǖT�)��+���Ӈ��`�7؅�ƚڧ�}�:�4�ߤ�q&���Gj���_���L��%��4��cV~�.Y'Є)�G���C{M�8����@�۷�ɯ�����9��3ZN7�y�������oK٣�j�L:[_$�,dH.���GqR��58 �g���9=�dvQ�3�V�L&g���0s�MC��7��&�PƠ��1[�H��T	�~�B������Ä��|?�y��[�/Rq4	�]I>H�a�)���F��q_x_��}�x��k\k$d���@�ob]�iD��I�Eș�{[={ut%���p���5��g�|��Xפ�#����@��݊
�\��?8���	�@�r6c���\�M�y;��o^?��w?�M&vq�#Y�L	�stp8������g���Ǝ�Od'���ƫ=����Y��0�E�r����kUU9kYS{�d����6�,�1 ��K�Ys��-�KSKqɅ|z�/5�Oz K$W����{$�S�O$9'd��?'�l��8�̫
��e�jfZּ���N1���Sn���1!_����XP��w��$��������lj�q��[t0�gW�x��Ϛ���s;r�����nYt:��L,`"�b�t�L`ǆ��}Cfh�T|�#p�y�$��yǺC	�nPQ9����IBo��߿y)�8z�m�����ە�h"����~nH��$����������O�X�kH��n�!��6P���t0\��ONN(���7�K��[�^��:j���������>�&�(a�䖠`s��pz�jP�p��.�V���)�M�L��2�o�j�E��WW,�:XƜ�8��j��H|:��D�w>q���W���d_v��R?�m��O,t`95ٌ?�{�B��va��s�#��<�ؓȻ��|��[e����e}���dA��`έTn#ʩ^��n�N��31�C9Q"�l��9%����i�ea��x�"� k�����+�z���G�f<,���Q��?�J�qC�yK�3�ga��mr⒄���}/�~��3� >Z�Y��#ހ��`*�p�6ۈ�nT#J�?U�I}��`'��G���X�K��D:�˫X�n�`Т:K�ߡ� ����������L��`l'��7����/e6�d�3j͟O�X^�5�>&`��1,<��t���^��-s�YÙeȂ��" �M�ur|�6(�J���A������]`&�b�B0�ty;�<>:Jv&;,!VL��R4xtp�a���Q'�î!%�R�1��f�Z�A7���dKp2�V;�O��SQL�pL�j�ค2����k�]=�s&V^r�7�,hו�A��/�`'��V�m���TXJ�zN{Gs\��&�@�� *T�r�U��30���hγt�K�Dɿ�ߏ}�}�o=>��O�!���p>���! �NN����s�ƅP%�AЮg*��Q��Z�zNRj�Xk�|c)�Yrj�EI�T^�k0�!������S\��j�����H����9���3Z���|y�#���Q��$�~��E�goQg�b{��2�϶����z�߳�bb��#�OP9�6�@�նF�@G[��=+� Z|DKw/|Ԗ^�fy��<2�,<�]t�p0��,GCdA����od:��AR Y|d������af���m@f��ꜣp��pY��X���ʖ�,@zP�d2*�(Tl5T:n����M6�d���\'��ȷ ts�қ����&]XP��)x@	H�&-���EI�x�0�ߺ{|�ͣ.]�ݑ�j�j�TD+.��lM@����� TX1��:����t��^_����떜j<[�5�F&L%T��2��2@�{dA�k�Vȧ�4m%�)b���1��� ��9����G�fӞ�ٝ��� �����R�5����K��R�.I�ٲ�Lu�:�t�)��߅Xz��@2�T�5т�`z��g���=p���Ɩ9� ����:E�T�Υ��N�B�Sf´�7[�Q4$�9t�@�Yy#���"�@�Ѻ�.���rk]=v��4Gg�����v��}���έ[E�����"}D)�@�j��,9�F)�����-JP �L P+񲶨#�I��@B ���[��ڴxZ�;��~���ù�3���@����3y���l40��*�������0!>;9�����ß����L<2O��-8Q��H�Z���Z�퐪�(�@�1]���׋�'�IH��i]��S��]�!&������=F@�0�0��>��W-��r��ň@Hˣex�����;y��T�f[]�و�d'������u�.�@�Դi��Li��ZR�m�%c�GC�g�hp4�9�x��칛�ȸ��@ި�{���T�$dǷL�U@J�P�l<ɛו�sw��G�d�j �����]��,�q�"fE�+�a}��pc�@P�R׵�����ww���z`�Iݞ)�����{����E��#׺:�s�Ü�hYǝ�1߼�F޼~#��L�}Qņ���9�m�m�{2�T��1׮<�+���Q�At2����^V.� @\/OK/Γr��5Ǝ-���}A���KLR���g���X=�̎$[&�;���])�QXwl�����{{�8��������C�wk�;��Ѿt	>��%Λew�I����!J�Y��&s�3]�@�� L�yep �OT/��<G!Q}�!	?Yb���F��ve�����Gc��z��  8�v@W�TrH52�(��~� ޾��d?o/�y"�齏�~���L0�Nd�� (�;�E5o�<�л�dO':��e�
)(=e�7���(ٽi�.F��=��IcZ�a�����O8J���Z.�nR�~�.�
�iU�4�&�wr'K���r��:֌�F��
z����6�TQК
4 >R�վ@��4����Pj�JI��P+FV� /�Q�?l��]�D�r_��q�`�h$V
�?$ ��↝��Z�B?�L`�z:?<�!����Af	���\���#�F���ߏQcg{��Uv���9�!��� o�k��QqX�|�6��h5�>)(E�F�i�lȭku��d�E�E��b�����]���N,3���lhWM��/=�S����po�;���R#�2�;ҳmK"$"�n��	|]��م|>�JN�e���f	m;��h:BzbF>�'���U��6J����Irk�����o�a�,V'� [;��f/^������;�ã#9>>&S&k�an��Ņ����c_H7�K�r�癦�^��)f�]����7@�#ӹ�|E�5���+9����Zu�����j��r��ॳ�ts��j͌��ĝTӴ)�C�T�G e��F��]�����NǢq(�����#h�g��\@Ȯ6�UK����Y:���k� h�1����f ���$P��*@�u0N	89M m9��T՝ĺ#m��J��G3t�ma�9��jF٥m�X����J��᳧���z�qX�l#i��}H�;u7f(��Q0�0�;��B��(8w�O�����9\ұ�X��E�[r)5r}K��xح�l�9dBv�G�$9�`G�E��ܧVK��-�����\���+sV���*;�3 �$�'�Z3A��Z�t���SOԱ�p�e�rֱ���{��vu*�Fː��/�_��������0;��$&=����`^���So׮2��ۺ Y�R����ٍ��Px�]�gFt^ ��B�E�,��uh��΁c�0�nheOͼ���˹��Д�����r�-�H�.�V!=,�&kVrs-�-����k4#��
�k��b�B��v�U�:��9.NC(����������d��UY��~I~�N������x����K[Oe�>&)@�&�9�[�dw_�ۗ��Y�N]��P��9��(���ך�1OyjF���(�]`K�dvۣ]�(�B�Qǲi����|�O2IM��RY9N;�����u�s�����&��X��1*��0�oAb�Vp�� `*�1�9�!X3\�k �.Ȣ����ɶguy��Չ c.>j��*rѣp�;f�,�s�Ub��d����WD��|6y�"����C��Z334�!�P$,Z���|���������ںb$��J��q��֝H�bl<9�-օ�0e�nD�q���:�~]��e�W�u�h<�*�ME�_�.�;�2�ms������R8��sAZ��N�&i��/jzS	��){�$C�d!{��	�ΘQČ3D"���B%"��й�d�������z��:�$k,���<���EQj�L�g����>����g�|����"R\A���jI��U�z�>h���{UY�7"n�؂Ό���0��A�A�c�ؐ�Pw,0�l�&�dx��_���������&����`?��=n(�a:��j::�.�ә\�cp�Jf]�xS��M:�s�� O0\-ז�	���I�c� ��]0�ݬ��w�O`�1J�Fj��>��y����'��@�x���H�a�㯝sVB{;�5���M$�dj�UȎK���@K##�]aK���N	�
����,H�[��=
��w�c�i��5��u��F���*���<�� �	����+:�
^V�\�E�ҷ�d�g,h5�N��3>N���y�˟�`wF!D��r ���s����m�E�m�}�~x�������@�}����Lk�����˛��ɥ����9�L?��&=s������=�%fPK�(d�� �3�u���_��NxW��YAy1g_�����̲E7��_��$�Ѳ����߿�B0JaKk�6\UMW���G��h��`�ǃݲ�Z� �~����A3̔�~~�y�J�,���:<��B��e(���
�o~��|x��#�н��� ���`ǿ*�C���ƻU��^�l��A�,��8�'�K��j���<�(�'���� �ד��GlL�]��!K8��@�N�T�2٠��v1fkG���A޽}GZlg�2Sy�p�S]>� ��ZM�֔l�_ ��b~��d?GM����a�8k�WӯӶ���i�6d{0��d���K@�M�]�s�]��FDP*��&��ڠ��t�QՔ���gQ税�m´�lN�	�ˑ�l�ltodqc=Yz'�٦e`�,�{���������V����X�Fl�$�3���k��n#��M�+��WT���w��^	V��2@YȲIQl�NN2XW�k�2���U�6��H3�,�1�� ��I�h�3�\zB#3�>\H5��iZ�����N���u�\�`�l'�^� 3����Ȉ%���M뭮��pǤ��v�5�E��-Y��(U��n�� ��T5�<�W=������,)U8V�z��"��+�wэ��?�@��ح>���(�H��9+zX4�Ш���^��2��j�w%�0^V�� ��%ʜgS���4]Wc37Z��
$<���Z�} pj�Lm]��)��g»h� �1��|����YIWͤFIi���'���E�@�7�|#O�_�\C1����+��	ޑ�K�?(D�0�ۯLY���9v�rƨ?�Nj��1���g���P]�Ì�r����0���3s�;2/�%6	����Y0'�J�eÃw2DG���D���ӥ\_]��YԥkU�M/�Y����F���� &�\3��Z�C�VZlU�FN�~s{ˠ�3�T�8�ҹ���q{{J��"�S�m��xi3zR�zƟ�L���n/�s��]l��`=솔���d����d)��/������V��������$��u�Zm����i�*C���������|<�vG�@����x�\���XW|Os�hձ�d�@z��ta`���M~���"�d� pb筓�zl��>��<1�f�Lğ�/�$�*N�bݦ׭�גՒ�R���>Pb�$�_�\ɇO�^����1Y|W�������4hoR�~���?e�5v@s�:#���j�3d�"��S�H���jx�Uz헴&��+�Nr	�@i)(����%ƽ�'��|d� ��:p��Txܬ�pB�sT-��> SA�1ӓ�.h��N;j����)%�s&*���m�Z�ЭXd`d��vď��]O9�'z!���C��Ϟ��a��d�P��;��BPK�ܑU�*�_f���YS=o�6�h���MS��M-/�8x�@��~�r��C�5I�L�����z���Z�/F��#xi�d^����U�����;�t���J�}�7H�Sn�Q05J�yd�HM�HFD�dՈ=Р��Z
��N�v�lu����hxy�t=#a��o��ܸQ���ɤ�e�βnxOD" �$Py���ڈ�v_��d �l�"��{;{Lǿ�p.��&ۚ.��䘀�Hi!Wh2MTsQ#2��TA<s\��S⣕Uۨ��ps��~iA�x��gd�:Y�P�s*+j��&Q�ٵ�W�a0���~��h��c�a ��S�d�������xM&�JϺ��K%WO�fO9v�0-b�5p:(G�4�#�J�F�g�+:Bk��,�8R����짂CE�9l�m	G�����˓As4A��f�2�Tٚ�r �<�u�yy�2{�K�����d�9������h쏢a
-�	��	�r�V�3�0� ��� �4 �s����!!�?,����>JN�:P�m
��SQkji�L�qe���0� ��(��1�;W^��$��TY/,�UX�,�EFmJ�75��,B����2��������7�t�����t�y*V¾�/	��#3䋺�|&.�+�_�������ݳǬ��J��ã�|^�")u|�_�hP#a�Dj��B��`��`c� >
�o�:�Wp��o���;����|�����L^��Z�=}l��g�����)A�vI���� �r�s�내w����V�Ae�A������X5T~����g���Lf#�N�S��O�?ɇ�o)�2���|Gv�;l��pl�Ec�>s�rJ�G��;(��Շc��t$Ͽ\������ ��yd��wƟ���2����ӵ��-�����e����ny��(�$�XV*�^�� �+�ۃ�٢������h�D�G9�s�����J����� ϥd�j��������2N�� )*�=xP*�#�%щ�Vj�3�����w}�$T����Z�$���Z��Ҹ����F����1�l��]���C�n���M_B�m	C٥�ڕD� �Y�J� �Q:`�#�Ҕ��Uu҄R3^n]2љ��З9�3(W>��?��"Tx��hs��2�TxQ;4#�lϬY&K��K,�U�՗O�=;�Rq�,EY4�r����g������b������&��fW��25�ONN�q���;� iT�L��V���4tEΠ����jy�!�d�F�XBc2J����Z7.\�te�L�Zc}����G�)���f���S ��Dg�R�	 �LN�ȣGG��h�_�F��������ƨ�YHnu�=e6��hk�R�в]#ZB�J�5�Z���Q���;�h��0�E�=��b�ved�2�ۀ$ɻE�a	lN���@��`�]\����3.A{9ʇzتoS�̹)�@���ģ�=�;F>���]�]	����` x����@ 0�����aFb�%��!UU2L���r��Dg-�Ć�d�(��?v~��%�p$;�i����r@~��o�x�3i�6���(�� X�)�,4�b�1�� ������ŴL� I�&�5�����*#>_�̦�e��Ƽo6�.a�f<�(ڈ]Y�[z��VY����4�_�]�j�[�ﴖnM�Y�by�7\س/�2ng��4ki�@�\�9��7�[<�b�?x i7q�P���_9B���Rv��d���]���A����R'jW!!�����Y*�`9<k����7w��m4�'$%:��QmA��Aw�QAQ4T=:9H6{_���+�t�_ɇw���W��B� 6�J_	����$� ꁀ�i�����P�& ������Z>|��
'HD���;T�t
H�Z$ۀ!�u�9�YA|\'� �K��6�^��?�ȑL�)�^�xDr�tυ���y��~&Z)��]j �͇y���U��8�� �gK����bX�9s��_Yȿ��?��=|t�	��XSRtnóQ�ն�V� ����B�]���\ld3VkU伦�m��H��ᨒo0�ƛB�v��=�Qz��w_uE�sM�x˞����:�
���HQ�� ZW(�9���q�Om��d��H�!#�3�t�PWN4��c�������h�'��U	�:i�_٭��1bb.Y#l��F	?jr���/�7��.�u#z��$EA�K1�4c���/^XgM+��6�͵tR�dbb`��K =o �~��VT����O*��(��2R��`mooo���R��q��:=m� �A�8.F�Fii�����:?�����W/�o�@��N�chߠtِ�i� (k��7�d�Jf�Z��Բ�*r���a��L��u��&��d��T;�,�gQ�����D�H=�b�R�c�p�	čg��W�O�:�;���@�:���M��Bg2*."lJ>*��D�֚B�c;���FG'�W�Lkm�S�I���l]XCAv��-W���D�J&�@]鼰̵��֞��8�����e�7�,0D��%=�gC�)�;�4
*��s�Aͮ�L;�T1^�O8����)�����ic��L��Ѭ=�Dg`�c��$x�ʚݵ�Y*�#f��ǡ��������m�/���B�췺���AfS�P?��#�(^��,�f�43�,)���6���Y����'�K��:om��k���5���������0_*��e���Z�g9��N:寱�j��J�_y+��/�B�X:?~�P�J�L�R�~]~ 7��s�LW��<<g�_ǼҎs�R�����W���yA}Kۋ,�c���l6NA�|��c��F�:W�,n8�}������ʣ���t��rqq�%�tQ�jj����;��0��n�kj��Z��ސ��OA-|ƙ!����X�~���l@�b��#��F��om�	���0=�%\(�u+�zA�ٛ%���f��s�=K�Č�a%���XIir���`��m�kl��r"���g����-D���\�yӳ�
xi�Z�2BG�$yZ���X�Hl���.ֱ�ֵJ�T:"E��n�q�V����eZ�5�?:�m XK�]9t\�=���
�l<2 3SS8@��B�79�/fܰ���ck�H�wSjzCpș,�����"��c��y 1���P�!��Sߚ�ˉ}v�:�?��hNչA&���ԙw4�Q�B,�4��i���ײ�, 8X�sdF�Z1���S��� �jw!�+S(	��ʣ�U��-�]��͂�'}MdD-�	�XCԒ��J�م�H�7T8>==�V���n~>�����;��m\u�Qci¾�M댁�ON�R�w����a�U� ����h���d�@������ťԏ�す �[.��K�Kk���$�u颜�FtҰ�CKN!�o���8�*v���m㒹S�a�����p�F���������p�jT'��z�)�l�^�3�}��:��k���� �\��H�/r1���c��1�P�.x�'߻S�Mޝv��$��F�ʗ�6�~1((m�3u!�ڷkv`�vN��R��Ā��j�F�ԄɈ���ɳK�-:�JǏ�;^���k[;��Iݴ�&��o�vƩb^Sk�e�\���6�6P5tm:�3��W��*Z����~��������C�{A�m6�4���7q���gv�)� ��
�jô�o�f�7���3���u����ڐSXG'�3x>-��T��B����neЎr� ����=�ޒM[���3��f���_d?ټ"hg�z�o���mU���Tnnnigʲ췯]S���z�	�rAↂ�"o���Z��r֡( GS ?����U]8ם��}��,�Yu΁�˅R/T����WCF}���n������hՉ�(9�>���ѯ����?�U�hϲ��.Ĭ'��i�q�ZR��'���q+9�Q3��ߓ�Du�MkQÎ�.sh�k��+M���m�܄WH"�B<�a^�V��������{�s{�e��_�{�X~^%��^��*c�͜�`�7;wBɫχ��
���uT(=�k�HG%�Xd<�҆�Agi��[d�6h��H�u��ɡ��{��H1 �ϻJ��J��Gy>�`6~`�g�%HD����!�T�1S����Wa]�t���jךw��6�S���n���� #7Y��0�΍E[h�<(�������M���2������û����]|��s�*�	�%�s�Y��IMҁtt(�\g�a���с�^~��08�_?|��;��
�	Fa_���8���K�!b�P�O� ��_~!0�� %����[T��!x�&O��eWdg{�f,=��Gr�7���D�f�L���:X/o��U�0�{�_W�N��5�̅f��9�5,66 ���i�� �mV��J��cYt�B�c�Yk�k8� ��J��A��넝����g(�&�T�<���a(C>�H�k���`�`	Q�oF�4��Etax��� 5R�E�Q7�;f��S^��Q,�y�r�䌖�{�D�B�{Vë��?G����й�e`T��r0��U�𱔦r8ȇk
"��4ѐy�Z�z�N�Q�B��Du>.��wJv��h�}]�s�!��U��j73�H�p�Ȑؐ_��h�Ơ���̦!��ۧ�h�$�u��uj�e�+�.� ���Y�O��0������3�E	u\\�%�!jyV5�����gS��U�>R[�h�1(�����{V<� ��9��U5��M.R��^�R~v�r(f��-;���\��s@;��7O�e�2ҹ�Ԍ��d�����?��O���Z0�D0甆\�B0 {���ŭ\\]rtYU�*2#�U�<Uf!�Iv6�� ��PZH!P��ٓO���_��Uy��{���ڎPɇ�ľ��a�T"v  P@�9e�� �J 3k���i��_3�1�_f��B�]�]��ݞhNϦ�6]��m���)�2�9Ө��^��Ti)s��2鬢)�f%F+��Oeyߺuh� r-I`�ڽ�-���2W=�ɳ�2,��nFy�s(^���_����*M︣��h�ؽ	>łb�..؊i0̀U�ڻ�ט�#��@Z�v�"�[����uS�;��lv���r��j����`�{4ڃ�����?�%V'�Y��hܢr�j�(�cu؈� ����J����:=��'�s��}����U%5�����A�!�C���e�	��u��[���K��,��n�D�b����}Fo���̘�)��M�5�ȓGG����xq8�e�eխ�Nȣ�=�v�.2�.�=�A<VD��g�2�N�ۗ/�8�}:v�[�x},߾xFg���.�S��G5���9߽|.�~�þ�wY�P�Vˇ�C@ ��vp4U�⺝��[ ���e� L�5�Qb�B۶c3%<[�/�t��h�d�~o ��#r���gD�Bi۱�5��9���G8���Ur��X���;��% �r���\�҂��g��նjl�Q�W�u�e�7�WZqƱZJ�lL�@1��ޘh�'j��Y�"�cԄ��[7�6��X����?�-.�'2х�E���u�8�O�k����_��ZZWtK��'����2��/��=]+�0�
 l�����4�> ��k��>��y0�'.��,��U�ky���e����δ�l(?#�B�W���I�0���<G�D���?��$(<d(�"�*?���3��J5�*Hz�ژh�;�W,��Er�e� '�]�*w�L �
Yc�ձu.�~qus'�>a7$��s4f	�=�yB��q~y����k�;�Z����$��_���s���v$E�h�oBڨ����5���W3ٚ�)�Tҡ����i���H��}�=zt�/ ��f�gEyo�J׍�O�7�3�T�N���R�E�JA�a�wȷ`���ҿ�a7-�a{��X�ة���=�}칀b3?�����G�9�h>���@&i��O�kB�g9�p�	;�/���~���D�x��+V�-ə�|�7|�L�t���(z�4�7�=��o� O��]P.{��e¸�C��O��(*m�F;�Q�b�V1�����:+@xcM�2c�Ng�=*��$�D,e}E�c:�-Hg�Ʊ�wr��:��H,�7�Q�tU����xas��4P�����H���Yp�����G��}�~~׿FQ�E�7�����@@T�s�lBɟ�@?a6�7S��_�w����u�<h����ad���8:B��N�t*�ܮW/_���(��∭�s��?Ju/��9a���4*��(���pخttц�v��*�
��{c��T��3 �=y,/_~+��	��G,�\k9aI�\+6|����� 3���/72�҆�u�յi��2OZW����e�v�b /��JNFٳkt����:A�<�L�����F�le\�V;�$�:]pN�Аho��#�H� DTl���a�cZ�U2b���i�Э����  �X��y�]D���)�P�׍)��_�Kd	�0��,�{��Y��3I���Y�� �]�Y��0���3���x����NY�-�u�h��cۻ�ա�̞�7ߔ��m�.�������~Q��q/��9��:�q�����_�o�%N+� ���C��KS2 �����y�F�%٥@u��k�Q[)���0�j�GA\Pڠe�����b�5m��DeLXUM&d�{��C)��n�h��Y*�z����G�j�L" ����T)Nc���0��l���ƚ��dM�@o&6��G��?�Q5��?Y�)(۰�#sQn%J� P��%�o�q����i����˅�Cۥ�nI�����<}��`m���s�tת?��Xn��y���v���c���&�Mˬ��*}�&Q D� Mh�ٛOe'�
��XF�B9�m�`��W�t:�_�z���N<�r!7�az���i���!���cN	��b^ea��j�h ���+��w+y�}����z�]������9= �&P+8/U��XOH�|��lSuyO1h"b�/�>2C:I��X���H�wJ�!ۗ�ʈʭ�u�w�~��k3x��f?q�E���j���=������� �v�J+�k0])����)����u�$7Y���gVW���	5(�PV�yE�~vc����g�����2
h�i��t[g�� ���	9�CC��
�B��<D3�9@U+�?-�jG>�ƷH7_4uB K��� h���%��'�8�]�)~y�C�,׭����f����wr�@	�,������'O�*�>I�z\�uq���'g6Q�=<;%8 �����c:���9�RR��~%O/do�<E�[**��g���GG�uJ�$�A\�v2&�9���B�88;����9=�J�yN#�n�#EnE���h���c��������kJ��)��]/侴
P�R�Ò�YN8�8 B�ʈe�������fِ׀��Ȩj���0C�l�Z�o5��5�e�L���fA���������(��h5��~Aw�w=�k�����St�m41��x	:���r�s|\wg���iϔi�'��<J����n]Į��˕֧ I���)���D��0}&�S���Dtn�3�<3(AA#��KUfB�g[\H?S�זچl��._��zeg��\R�e\AL�SV��lA22y�N!�M�V���3��Zf�A'�TM�מ_��	5�Q������@_�mԍ�ou,	�w'#-+s������Q-Q��N5�1�S]J�@�Ԝ�hD ����Ip7��Ŝ]�:k|qi!vЦ�3>`! k,�������/r��yV����n�0�'��r��p�me՘�tK������~6�D  d6.�yA���O��}ͼ#@M���F��vl�uE;quM!�KV+N�؞���kۙM�,؁��<�{�N7�z��|v-?^ʗ�[
�:��u
���^�M�'F�t�F�E�,��F���	<��]'��L׾�T$�k'�ڐ"=���u��EZ�5�8h��Nk�\ic�W#���Y��DEN���ZZ�Z�����Xo?z_쩯�O=�h�����/���o^3�'<�������F��si� LB^Mp��T~H�D(Q:��)�-����.g@�����D{w�XKC�Du^�0����ː�<��������%*���w��ܢ�2d�U�M��2�i�>�1�Tc,n~8_=�Ч7���|��(J���b�a���X�iV���qw�w���G�q]k��P2?�x 1NX�uw$�T��nu���SD�5}t�,ם\�,�z��`�
�,��Z%j"k�����}S�0̶�t @���� qU|�0B����]'c�c��/Rt�o?����5���4�+'��A�8�8\���7����T�X�� :;������y�᳜���tP��%(6*��n��
L(@�c���VO���3��hR3#��&��"1��Z(賬X3
E�h3�D�^��h5n}DW�\ \�
�)�����C�ԑ���KE*H��J���R;�`���d�7��fPp�ˎݲ�B���*�m��!��{�֌Qi�3��Ap� �۴2�͈�s"E��%�.R�H���qw��ﺦް�4(��F���jÆe�Iv��n�.6鿷��U:�\�C�r$SU�.Ֆ,��ݥ�ߏ���u���qUL�X�`��4�����5 �!l��koo�u�vE�����(��:��"~/牊����*��HGGYyƬ�Y�C�)�ZJ��!�� e���.˧��L��kY��W��dɞ����|!�*�u�D�u�����8J��	�����J�mR�#M�S[[}0�*��u�>p���H����e3Dl�NM8��)�X#��d	V� LADA��ٲ�I�{���Qk�4���R�y���Ãz���ѐ��ҝ�6	D,X2�Jv��Ԑlɗ�M��w�u�l��`KO�#��EV�6�\�m�|�v(�E9=��?����l_�<�������4���3c��OQaaw���F���7��ʻ�)H���Q6	"���,�߭A�����̶'YG����[ʲdf�S�f� l�k�������� +� }
I�d�nӹ;�����my#��E��W�`�2ʚ���aS2�LH�	&�T����a�8�)���g�3���rL�0U��o?������-�	���=[-bэeG��}���>��]-E|�ATOT���MD�TUa79�8b{%#�κ �iD94��h�w����߳p���p��+u�����w��Ha��^�CI2����-�:-�Vo��k�V	B�~l�D2�r~���`��w��FG��:Y��i�nWɈW��U��='�{pD� R�O�r�z������օ�@
����r��, D/8DPbFsz~ͮDL�׮0u  �Ͷ��kiT�f�V��k��ݲ���$�~N����� *ZL	*�W���|A���w�}����lϸ_�ҡ�I 
ژ���9I�m�>Dt{zv%o�}����Y���la0�TAN�Dn�C��B�-4x�ؼJFb���NPP?j6I�)9��_K}�1�}=1�:����r��h�5!C
 �^�X���,�p��V2�h%G�9GAmM��:���g��!.LY��<vi��^�1V,붊Ţ��ƙ �"�3 �8L�S1U�(��)J4�����}��s���m��>���h,u�!a�f�ikx0�,=!.'`5
3H�a����;�ҾB�C�Ud3�\&#�3)���6Ӝ���`��%y4���J�}�����eIaw ��q��B:eoo������_��������]�ur�p�:2~.z�N1�V�@A�ɢ,��eh� ׸��,9�-� 1�|U��V�t�^[�J/�/*U���ydL�ϐt�'Pj�Y��mJI@�l���i����ٞR�f;�[ ����0��f��f�G,�f}�Y���` �#�? G:�+� Z{�#n9��5��hَ^�B3�zZ��2����O��J޿�����Հ���/_(C�F
M��SCj�R.��x��v�>:�e ��V	��Ò��c�U�ư��/&Obt�Φ;DK
����D���b
˽>#�5���$[zi�*������oUiy�5:Fi«5m�6�\^߳4�!�܋
�3�l�Ӌk��Ǔ��{����uC��I�.�����nŨA`�����o�%���iM����V������W�Ǽ��3��&B}�A����mT��3�r4�Ｑ��	��`Y[�}�]����������Djo���}t���[4�J��~�g���1K���y�F,�l9'+8���ܲa�����DgA�n��
Ě:d˵��(F�m��b�T�B�FD��Å�_d������[Hu�z����70̐�E�c�7S0�巳�^s��YÇ�y���W�}5����{.��
f� Ho����,��z;En\�y�&.Z+�)i ��c�A�(��`����s���'�����' �@��	@�Ȟ^�����h�`����x��-����������My���}>���ۣ1R�҂̾j���+����O4`E��#W*b�?�G)�@����!lD������_������7�@$@�&s6K����ő�ծ���Ka��
�ޥ����5?���\���%�p�{�,MhE�KWyWq�ݔ1�\��Cd'$���05�fk-�3��nrb���ׁ<9>Jk:�a�M��T'�#ɪ�κT>Ԫߧg���֒G�E�\�w��R��g����<E��	LO�I�����v�;3���o�hWk: �f��ޢ8
~��b����IxG �Y&Rt|V�RscG(�FK�0�L��X�@�Q˿Сc���6��T��Ǽw8Yt(j��j�k�%�3������&��3Ct�y�FW���	'�R���T΅|Ŏ����_��۷����:9�0b�7��lDZi��L�g�� 7�9�n��b3������8}���(t�"�����ӕe�J�Hk`d��5�6Fs�I�5����..�����%��xm0�'���aՐ���o�ȳ�'�a��9rM�BK읍tj�3m<<G��Xf[�|�* �M�K:{{���R9r&�Ia��A��~F������:���"�'�j����2':A�L e@p�p2ٕ*:S �.�˟���r��邍E;P+�/�ү���Ԏ=��<��|!��QBe�I�`��A�|�s1���M[Ӧ]c�}+7��R(����Ħ>e�8O{|:-�s��G�[�{����X��
� a��A� �3�ί��?�"��{��$��ҵ#𸽾!J��Ǩ#TR*���H���+5 ��?�>���F�(�귧c^�G � ����s���BT� ���U��;W���q�qzZMcr��S]Nv�o��7 E����(NI
YO d?�Kk_��x��a}Ƌ�ϧ%�,`�#��2�޺>1�}J��Xoة���߫ ��>��ˍ}�uA�?�T���`��ۓ{ 6̂I>�g�
y �����g�/F4R��?KC*h�E���C聚�����w�s�]� M#�u_˛���{�S8�8<D�0(���?�V&��z�#VD�����tz��ѝ�,�%��W�9�u���E�.Rt�;�f�O�����w�D�-[�m���b#>�ɛ��ɠ޲�A�k�G� ��@
M��m{pJ��oҡG��+���./6�0��`�& ������[Fw�w,�N�a��V� �G��U���~��i�!�Cڹחg�� )��bĎ,�)		�F �u���A��Ú���9�a���TG�Az���\�ʫ���,��G�a��n�4Ƒq`^hw�F��A�-t:�����e� �z���Z�鈘�? k�mU��d_?9����^�$�G��> 
��7�ᚖ��*�Ɂ���@p^�%ú��%�wY��Fi0�x�2R���*�}�D��PgD��蔛�?�L�V6�.�t���)k��P~�Uӳ���������U�I�ΒGnV��	 ń���h<Mk�^8S8�p>ggg�.9�_���v(?
��r�J���clY΄���BP�&�³����ҽb�����ﾑW/��7O%�8����3��]ړԻ��ܵ���/'�t|���J���{�nqO�l�g[8��TRƅ������W���sy��I%[�^*�`�0�"�a�nx�`cHj���gn��95��ͽ���:=74���\Ed\�̚l����R"�Ȱ��^�7)0\��$X�.m9a�&�.�N:�J��gЩp�� �ڭ9b��a��}���ܭ�kn�, VP�����b]~k�H0?cc����o5����{�C�s�w��iޮ�Cd:�HE@� �U�_R�ى@@��u�a6����R������
ϧ�3Mg���`��l�&	6<h���?�t}�� i��m�,Ȯ Spz8v���\��N~��~U�]�g�����yY׸�4S8n�=lM�2Tr�EH��U�C�ςeΕ������g���Y��.j�̇�S������J����17��Nr2������w�Y5f�z#���44�X��VU��l<���������x9og -��� ���d�*8��"mO]�"���C���=���#��Z���t���w`�~v<�QFj]#7�Կ��h5E�ӊ�ג�m��Β�&E�����̫V5���M�R��:�����E��uZ�O�)2N�	�OatAz��fy����	����3�����0d��F��W2�]2���N���C�n�t�C����oߝ&�u-;�P�Y�(s�$�a.PY�@���%'�L��g�3�X7�2W�7t6���WZ���"m��/��|z�����r�(
\����9 )8�ؓ��,3a�l�:� �l��P��!r,0ܶa����O�=�����<=�.,&��~
�v��i�i�v�r�K�6kY�i)g���>�ۨ��- �W�:ڙ�w�<�?���ͳ'x��t����N��� ��r�j�_i:w�M�����i�l�s}��1�Ñ��
�z7�(��D��UeXS�^B�'.��i�1et�B�&�����h�Ϛ��i� ����M{�~}M�FJ@w:#�K���"�����gٞ?!eht}�+Q�l	����)?��_��G� a,֓�ͦ�@��x��� ������0�1���tm��s�S�M���1:�dw,ӴO:���4cF���%����:�*�S/�^�x�@`'9�1A������$�������ȶ�9i�������( C�&��Q~T�s�D�bQ:����n�<'��/��3�?}:�U
* ��9���|��[�*`��{k�E�%]P[�od}��H���b鶍y�i���pu�8� ��>þ雪�;�C�#Ga�Ԧ��U�QH�� �d�7P0��`�ѐ#�J�X&����l:g�j������Z���r�4o~Vi=��\C)��B�����,L��(�w
�1�ràE�2]o���״xNȶ!Ajj�},���ؐ�kۛ:eD�@?���)��3@*q��7�X�6� ��6n�I�/��:���� ��]�B�m��ܑ��^A�}z�Ne���=h_��q�(��|���U鉩�Q�R��A3���/4���ʑ�{��5]�q.xy��k(#_�0/w�5[z�dËv�e�U�qJ�i�5�k_c��{`٧(�7��덿}A��aC��&�l ����j%�7���6(@��zy�,Q�cq`8�.F�Ҭ���f1w����x�|,��;�C*��dh�͂F dh0�{bܯ���~������%3 a��H6.t`h���q3{�lR�iW��ɨ�Kf��� �(S�5�싒���h	�R]���ł%�M�j�Z���mh�b��'"Q
�,��"�d,�vH23
])d�0�>p�8�+�n��<���������=V�R��P��&#�5ٖ�ޖ<=>�ׯ^���ȋ�XwӚԫֆ?�w����y�<^�&F���`�3Bp֬�q@jNg&��Y!
ƫ���G���@�A�(�(�;jW���*��H��Nu�$�S���FL�W���\3G� ��W�*U�ZY{��\��~Ng��"�`6I�PXjZ���ڨʂ��P�d9������-��-(d�>|�(�W:/o��������K�K�9��ɓ}_t|�r��a*\T_|�t������y��m:+�_�M�Ni���eD�dX#��|� �x�;��)�Lv����������zkf,6�3U!�5Ǚu�[N`�x���	�cK Ҝ�)��ξ�%�z��)�����V�3��Z�w�/a����L>m��J wK�\��0�����Ay�a �b��
KZ�9�F&��:kM3�]p˦#�W�3�,��΀M�1ܥ�S�3�y�??jMZ3����^%i�5��l4�:�3�h�Ɯekw�5XTY����o� {A�����&��]�b (6�
�2�c���d�Ag�@o��]��܌M� F�^:�[sǌ���~� :_\k��T}�@�^)x]-T���t�j��f]�܏

ʂC�H�̄���$'�� /6�,C�w�ͱ%�R;[w���:�z�J�M�,p�صN��˵v��q��Ri.���KqN�޻w�η���g�]��kY�������� �庌�<I�I�!��;�ۋ�^`��-��Y)��X�]�TL7��A^O=������7�{Ȁ�_��w��8	�ߧn�W���s�rY�=��Ix.�-Xo�٧:0}C���7�ע��r@��]��";���h�5m�qT�";��
:�S��PH7'G]G�N:<3�X��K'c�]I�4�d� q��I�Iè�����x��Ҿ�TlW���׌�Ӂ�[�(�����3v�;���>H{�)#�����`c�:�q����(c����	�R�{���)߲��z����v��=Xt�Ԥ&Z��GB ��uwR&�XMS$K��)#/ �v�Y�N�i�"�m`W2X(�� �Ff�ģ�}������|��D�v8�N� �����S�	 �Z�X"�G�Z5�h+y��@Q�S5�@2����Pg-�*]�=��M ��w�22�9����?�LgpZƸ�9u�Ո���}���5�I�J���ÅU �Er(;�~�RY��l���^�L%�0�1o�wXi�X��� �����g��@��?E��Ņ\^ ����N��R!��^\�ɿ�뿤�\��o�L�&�'����!@X2��9�7���.�Y@�7�ь�'�����c+�qm@9�ƣdI.�K�Y� ��u�zAUw�~B� xy}s���{�@<�^`2�L�)��P�_�&H�]A� �F�6�~��dk����E%�B>�9�]i�~N�ho>�ˎ�쥳 � �p�J�^` `ڝo'��X�?.�^}�A�+=h�v��P���J�v�e�;G����,��`!�=�E݆�Eh��A	��Rmr�,�s�ZӴcp+��]��>�����bW䈲rVn/����i{�a�P:���c�q��Q��k�i����D�lM
H�7����p��adܻ���ٝ 'w<�B�����Kv�c��Ǝ�66�]���4b@���ӧ��O,衹��˕�{���
���)��S�l����92X3��g\�$%� M�^������P�dT��f��F��_�`��v������=$���Ϡ���K���a�'�o�O�C���+�+b|ؘXE���Ė�/�Zt�y.��Hx������b���u��ړ�W�ǩ�1��P`-~��^������0�����B��=���DV+}JT#��Zk�˸��� �/F�	�t����}
���k�\�-՟�@��L�I����N;-`���'�,�u9|>)Zxmը~;�t��(h��R��G*��ƍ��`4��s*A`T�VcM�_��$±Uc8��>MGm=�L�s�Tb9�_���a�Y����jI�g��LI# �3�u�������?�3�4$gI�3!FQFJ�T��٣#y��Ic;����H�W���{vqEqHl��@H  ����DY#��'�^��������V̠���u�\%0�)���w�I���Y��Rm.�{v����9��j��wtٝ�"9�翞����^��D��Q��1����bE+���U�s�M�f�Vx�X���r��I�R�D��M���g���q�B��g��ֱ���X�7a`�g�`����씜�u�X'$P�̬K�6a�$(���l��L�����sH=%/�zb]�`PEm�)h�]^]ɛw���/o��/	^� LT�B�N�G�%Y4P,�[�*%$:���J}-�ՃK��~p\6Wr���Y(�C�} 6��!ɀi>B�{=��C����3��+4���^��1�V��k ���x�+I�&��̖�񡞛V�҆��6h�S���.Ȼ�������>^A�f`���0��v��R+��`�֌AQl`�vѰ$�g,6��ݩN��lvc��st2�Xv����XXQ��zyF��"jr� 0��QBl!�*=��%:��������<}����>�pDQ�_�ߦ3���[�����8e�MOV��c5�_D;�~/�L���:Ψ#5u�R��:�ӧV8�r��,1� �����{��8⡟�\A\�1���5��Q{���\�W|�kW$��8�VG<�&���.(p�H�ZS��J�Ik������z�Q�py���L�tp�Or*�7�V)��;�n,-�e�ˇ��}QT��!/�_�\�LD��
�8$
��eih�JC��f h��8��
�PV�V���#M���D��F��*��� �9K}c��wT/v"3<J�T�ǐ�Έ����H0��185Bp�nJNfǨ(�:�:�`YdgwW�f3�M�i�M��Y7
�a�*s ��űZ�+N t;�)�e���kYVthuk���� }M�f+����ۤJ}��~.�
�'���]N(03`J�Q��b��՛i�,"�"���;sF��\{�H���Z>�(��_R���"��h�w���4�'͂Yy��#�Yk)�৬Y���ܩ1/-k�L�����O ~��ǭu|�2֯5n&��
B��rDy�����?�,��ݩ<�49׻t=K�+�D��$D�ǜ�0���4���uϠ��~���*ك5��-�����Kr�B���Q���GT�Ǵ��݆2w��P.C$�,��	�*�:���r'	?Jmk?>9� lr� Հ�&� Zր"��'������)��X�1ҡi�J�Ť�w BU��QQ+ ��O����7o�/g�	�-8��M�^1�:�N�h�����}�A��Oi���N��*��B�+m� �f�c�l;�1`����$�Dt����I��8�+8=g+�or3֢d�Wx�[+���ӧٞ��뻵<B�W�,Q��@�>�����%���]���b�Bе�*u��OiPK\2���E=�9�U��nCJ�E��;��F4di�DT���wf�K��\�j����v�nT,`nh5����sϚL΅���Z��T��T�b��J`�V�/�_�L�X+f_��x:��T.,yYmK{�,W|�����,6��8/JA��6|ȏ�7O�ʓd0�@v�����=;KA���{�5�dK�%�	��h%I\x��{ ��s�t�)�o�Kچ���d2e�ǭ@���mT.cgv�v�+_2�U�i__�l����w2\�?�^~_�B~o��~Ʈ�ZI�E�X~O˂��%�/`���R'2�2dρ��y�5 ��!���7��/Z&�������O��i�B�}��	4;,��!o['���&B�l�;J΄��@�;3����~�Z�q�9R]#%|�n��5b�G�Qo+J"e�q<Ճ	QD�Z�}D�/�M��H�LB:H��}�J;;��"m�D���w�Si"xŬބ.���(�����S���X�'�8k��
ȰE�L����t���LAn��/��U�F�P�/t�(�X9�@a3G��C;�	=��T��H5��(/�������Y9�SA�Y����m9��&��3��d����^�嗿ɻ�ry�`t|�"S ��1��8��f`�2xp�Ś@�6�$�(�>h��	�����ZM�pլ�Δ�՘��l2(��:b�"��
���?�T�5O ��D�K��׶�=���O�P�knN 8�L�]5�N^����+��b)��c�C����4̞NF
��	�A<�q�	IT�a^���YV-4s�3�d/	�b̤"��'35�Υ�A�0��kNNN��n��&3\�,K� �7:��ׇl�E�~^`V���͆ �˗3m&H_?�rM �Pj"R9^	�Ƞ��@���O�뻏9�9�T7�~����y�q���f۩�:��Ȟ(8a9�6/�*̊���	,�Fˇ����Gьs�<������#qU}�A����������t(3ϭ�#��nGC�C,���Y]���W� L�̚��6��' �Sk�7��Z�݊��~M&�C���D��2�.�� �/p���Bѿ
��� �5ղ�;�<���*{�u��ӛӬܚ�oO�aA�U�l�WP��N��2_�\/}���3��00���K�3�)^<�o�y*���,G��TN'&�{�#O����=W(KBX��4G<�v�8��;�gE|&k�|M�LQg%��$�W]���#����[����}�=�+<�%^X���`$󥆿��?;g�2�+�zR�����hB����Tk-�i����d����XzM���m������0X����ɀ��]�|��,J��+�
��kƱ?���~WS�j���]G~��'"|�{�:{���;oyڻ	F�?Rula�>C7
�۬���Z�-�2^i#�B-e�=v�]|�Q�����i��y�.��Q.+Fu�i��п��Y\�R��t�����K��i���vm����8$ԋ���/��i �ց)�Qe�	6K��
7	�Zfjɋې�Qc�&���$Ԩ�p��s��'�XF61"'�XHMTS�0���h�v��#F)����O� ?�z�A��a4������������%�J�3%�+�+m�WӘ��R �b�3B9��u��%�Z>֥^�߫�HS���k��28�|����H��is���$5�:;%g�\0t��P�==a�����k}��Tvw���_���_|�����7N#98ضl�IY-��i�� ʷ�Ke��r0m��@�)%����8�?�Q�O�)5R�5(uL�&���������������SѪL�v���!*�lp�0J��UE����-k�P��k�}]���U��Sx�����9&L�~���ʾ�^����lU�_�Pk��9j��b��,t�qe3!k=1[�ya�NI�.���28f�����im���G`��@@ea\:�>��N�Q�#�l�'A(:EK՝=D�L��6�5��6�p�Q
�0G�R4/�n�w�M5�7�3��/���\���ח��W�s���%śWr�����"��Ƞ{565"���j��k��m ����P6��#�"�o���&�(r')�N:,܄l��>�E����I*�����\;��cf���#�tu6���z!�i���p���߿��~�^~��<{r"[[c��@i5*�{27�~��w������d���BC9Q
Bg\-�僙$())j�A|�Ih-ߢ"�!���&`��U�X:��u�/!�j���a@�7)3X�����i���hƳ3!c
���1��=(���Z��+U�E���R묚U5͛ml�q-<�em��
_���\~�������HON��>O�:�5y�	A�إ 
G�����5C�?X���2iu�q�����d�FI��cw{"����Va%S�5F@,���nW.//��o���NӒ�E�N�l,�����)�_U��5��jF�k�$U���:&إ$w��ƚEg�*�:�X*�ܔ�5*&����ۈkX�]^)��a��l�B����n����e�%�1�@��ꕣ�]#�I�T ��`xX�f��l�G �	�S��H�cEH؍��%[��pG~������jV���P���ЉBB�(�#��i�����щK$�:rm��s%π�o�dR7"٦�.;��c��x��bx�"��Y��\�Z�(N'�1[;��¬�u�\�,
#�L�`����O���oؙ{{I��G�=9"Y{b�M�T�B�,��l�mv�f�Y�I��g��9k+�0;��EK^�Pk�O�F�E�[S�.zm���@y��z�<ϫ	׭���r�iU�3A^��lIfKf�ʰK!�Ʃ:��(�P�# �|��,�#0R��G�6�ƚ$��6�Z�� ��m1(�QI�V>�v��H��q�!�_�^u�.�Y0�E����tֱh��=��~�oĲ`��c�mEڏ.���UY�G�3Lb�U�R~$З:kgA���G� |q�s\-4�6w?8�K�Ҟ�x��A��f� �l�c�o����C�@��B���t��	K�
�Zq�X��-T9�Y�"�y�"2c�@4�*L�V݈�� �c��ڼK��޳_�E��'|N��V&�k��Ùg��&*D{�N\ҢM놌��ޡ�x�T~��y��<~|";;s�4uz��V�nࣣ#�15����~��T.�n�*L%A�jpu��6 0�gg����9�3n/��`"!P�vj�����qm��rv|��,�N@��#Dze��_���S�_1�c<���	���)����}E�0̆���W��>aޗ��J\�t>_G��h�v�v�)>?`�G�;������6u?
S�τ�����<�ĥE�C��b��0��W+%k
�d���Lk������,�w��y\��	�,8�$�J!�������S�D�آ#�pȊ��?ȿ���W������B��e.�˱���@lP��uN�HޥҨ�dj�k���1Q0�a�k��1��h��^�Q�P��oR'�16ɑ�@C2�:��J���7�1�đ~��&��T7~�6��k^h{Yf�0�i�	Z����;�|y��,:�	fϝ�-�[ ��4dT*G���ه%} s�2�$�Ҁ�����<E���3�?�N@eƶr�� _sљW�G�eAv-�I�L붷M�YJgg u�+F�߿��B�,��*���O���UH�\��ԋ��� `G�:��n�U����M������|���svX���(H�lQ�� xJ�0�� �Xw�s�����}��[�S><�2�(���sC�ͅ���s����^�f]ۨ��fg�t��a�d�n-)O������0��wj���l���
�f���i�>�V�p�m��xf��y[�z?kV˜󂝍k��r��i2�[��
4P1}��r��v*:��H��DW�£�g�G���o��$Ω銱W�F9�c�T�'p��Z*��R��l��<@��3;��1�jNj��}xʱٚb��6˪S-��:b������w��|F�V�W6�zI"�m�8�(���4Zd���xW�����Y��_Am*���S5 꼳���"�����^��w��Ͻ���?��'���+y���������^�6��;bXHz�`���%࿾y'>�rl��3:e���C(��
>��ekH�ؗH�h�CG[R*)���T�s����DgɆau�0c�´�iĵiCK���e�ր�q`I�������O��{y��9����t�4H^�g�E��[)X����%x,Ǐ�ɟ~���?��J��Y7����$OͲ��>g��m@#��0)�{��	`�� u�i�*�M�*�7i�~�N�i�i�3 �� J��i���L]���� |O��r
�c����ƚ�
�7�qI���H��@-�EP���5"�pb��<��I�������4g����e��?_D�+���?�y�w���G;(�q�^�p�F+�𪦢���8�Cqn�(�[����O�ӣL��ڟO���z�D^~�(9�=3��P���h2[ӂ)wv��u��\����[H\�p�=���qg�<�H��Z	�|���U�G�s�҇�B�X#68#2��d�L�TAYzdÖ+է�r��G�hZ�kf��bB���6�Þ-��Љ����|J�QF��1ERAEd��9<1����χ3Ő���+���9�Y�d�R�D����"�Ih\&�����v��F#Q���u-�����0*�8=Sh�!R�(�TQ�����K�(�D-;E����/�	�2�g��L��� �N� d%���n�ߺ��0��eSp�,L ������eآv#>J������� �TD�2u�_>S�s�1�X�� |���Z��hl�q;a>���٠3%(�ic��9�D�aY,���:/O�yk`����q�TkB�̬I���zf�9[��l��.��ʓ0��r� 5�gY��֚v}�Py�9888��''r��LJt�"#��$2�]h!F�ز��<�ҨT�wЍ�^�u��' h��$�:�a��YE:Hݵ�3;��0�f���� �t>OXAF�`#v��|nww�r{��ɲ3.�J��6U�K����K1�v���,�Z��S)q�6]�g�h)5�� X �p6Va\dt�f%M
����5Kj�����ﾑ�'P�^���Q��S Ͳ*����%�m�;�� {a<�i!m󷴧�LkL�D��y�{�ܨ��bP�®*��O$OF*w��#1��.�D��5E-Gm�*M��
2*��}���m���l�+ϟ?!��ݏ�'�u@*�v�v���%U�������3:Ok��m��(���/j6iFK����׮b�ʩ�\7���mv��~���VdE �Aۀ�h啵�s}c�O/sY5�̹��g�\�ޫ/N9R|c^}P��Lbv���B�w�������&�Ln�pK����'䷩1Zk6N�8A�n�JŅ�Z��C��(o�\��MY8M�kb"\�Y-E����w�m�ACl�����7��Gч/��L��e��f���F4��HX����.���"Uj��ښ����@��x-ϟq��zq���*�k��F�����O�c�
2�z+?��by��!��W���LR�Ά�i+(
�2�3F�O��A0�M50 J��9�q��M��#�,��HVK#�k�|�dF6��~/hW��u��g��S�%�"d+�&�*g���g��o��<��|0�&�?2	��{|�7�NJ���n�B��$��?'�p����{S��׫vb2��).�͑>�ʣG���� ��j�*��n;N@����Rr8��'����g	d�3p��_�m)��<"�����zCǿ�RF�\ȩE��A�󢍔��ݕ�/����]k�����h���� fu/�_Xz8<<L��OЁ=����l�8�R���q����q�X-��5������_~yC�0��Eռ���'e`�DyU:,<��<������\�q��y$�9���x0�૵���C ֵY�������s�@��7�G�r����T#y�&x;>~$��?�M&[�J��Vf���X
^��³�c�'��>��Vg�6K� d����ؓI
�^�!�T@ ������~�YrɎ���������w����Qr�Sf1i�Ç̒,����y�(�0bdրe��^�Mh� 5�R8Ea��x2E��Q�1V��h�3������ .�j
��m����f �B{x���^ɏ?~'����w��A� ??�Uvְ-V�9	�(��99=�(5���ly�h6CF��-�!:!��A~�9]ާEg X4�J��KoD���3:�~���u�2��%SI�}���[�ޏ8���G������oI%W�M-�oبc��-[�YoVf���3�T�V���ٓ��[
po	�����TZ�m�bIQ�S��8?4X)�&>�_B҆�!�ֲ�JU`�dZSic�F�7�S��V|�b�2UMCm�[���(�	����B��>^��mMJ�m��B�8��5�k�!�J�||,�ʄ���Dޑ�����!=���z�"��\� 	�����=��͸)�f�le�����Z����/���aݷ�J$��x9³Ö�O��W�2q�*Wzљo a����Lɋg'��`����mx����QN�)(�`��aף	ˑ�JA�p�Ttms7�"g�P��T�HG`x������qëΌa��f(�stDa���cK�|h9Au��yFUī�.;�~�i����dA����m���~�����������j�@����^~Odh�I?������t�K"��ײ\5�6_�\����u���9p ��%�31� @��ސ���,�� 	��(E�pq��#��I`�������t_p���V��Z�cm���y���R<��~�/m��}	v�.Fp��5��.�@��d=v��8V1S-=���l5S�ٞS�L�^ ���y����O  +K�DkspE�sZ���k0���S��QI���ˮ���jЍg�ԛ]���J�-K����^2�Y�+Sb?c�iӞ��1J�M�C� �ՁS&�;�"�=�L�
݂��_���ҜF�`NK0�<@�¹ lß����霥uE�
�[���^}��Ϗ�B�@�߳S,��H��j�!�x!�R�ӓCy��Yr���^����[U����h3׮����:k�/4�l^dGo�"�Xg��5��ٯ�tKu�F
�pߍ�~�$ئڨ,�叁��b����� z�A������ ���y�6U��c(�'  ��!�hk=;:b��8_[��l�y��\]�RM�[n��F{�V)� �������eA$Wl�g�]��?ֲ>�&x	�|d���9���(3��`~��J�&��|+��	��b@���;]�@���V-4r��Z�ĳ��?��CI�$I3��8���L� ��;��� w���n��{�=Z�%�����GdU���%����n�f��f���[	���>��|�-G;�ūV�taԜ�m���l��U_R�t���h��v��$��[�Yz�L7�2Z�<:�K�JU�ӹ�����i6�(_X�;%Ca�7d_��M^�k��@�V�XO�f�`ql�3V[�b���؊�
�]��B$w ��T�KՅj����6D�9�� '�i����~����^��O�r�2�X����Sh�.���c��
��2��I��o{��[��Rb�}����
�ʍr""Wj�AZAVR����;�?"}s�b�O#�¹h[wxJ=(���ݕ��O���C��?����|��_��f�I20)��SUa�y�p_�L�������4�;��,����4J�,4�]�Kd��Ǣ�i~�����?��:��
���)�1>+~���O���?ɟ���;�x� ���Q��A��%H��뿹�EGs g���^����_�o���\0 7��6@ݒiCX���T�t�2�&#I�H����N����@Q�AvN��#~��H��:Lꌲk�w95ͲI�+�TZj4���\U���En~�c����f��V���5˒^�	>X�2�������&����KF��J��J#I�XQZ�R����E��<3�f�$k��r"���"CY��ʀ�n:���a�
R�G��M�r�m����ɿ�nK�q5W��WQ�3�Hi(�w&.M��|P��rb�kft�����D&�1�?��Ȣv�[�p*GưK.0sA�y�GG�|����,�S�1�����Ջg��������������_/���M��6H{�2⾖����	�0�
�h1�8|T�&P?M�/��{ruu� 4��@"K�l�E�M���������0�2�X������O�,.�A+��%�����Y 'LހGC���"��vS"%�
#t�r�w��
���dt�PB���G�*�nyl,��[��lE��0[�z{s+���Skk���éʩt:V���3/��/�$�V�&-���M���_�\�e�C~Mop��X��~'Z�ډN<��Na���{�����W鞀k���y���C`�
W�eP��(,d}i�K�%�cm" �Y��#�5�Y��{h�|�t����Q�!Q~���Z�.�/������ւz��Z����� #�he��̿(E
\8���K�a�lh�~���ڽ)<�N�"�f.��'_�����%5���|���t،��YI�2���ajx��/�_�*Pa���uY}�b�@XJX�!G*Q����b7 H���whqH�˖WdMo¾���.3āP�Fv�I��H!~�#�Z∼?�ug��qqY��s.���`NGT爋��l�gU42��=M�b_���hu�v(��	�ˑEr��Ѭ6[M�!A��U��LQǑu̃��� �s�!�����d�ς�ԇ��w ��S���_��WҌ�tN9�`0pcvލ�gc����M�{����.Fk���&��Y�w_!_~�3��O�#^XT�n���B7���X���N ���?���S&�d���VSU�D8\肩�����(��&E�/��Ӟ��cQ%@"E|��`�}����3NuȰ:MЬ�4v��5Ƹ(a�lc�B�#p;|ˡ|�����(k0�^�)B$g�R�3X皆�*�`�e��ڵX�Ho��������������_�5�ՙ��N�뵇�G���������(;�J2���|K�z\]_+-}.�]a��(5CE�2��������5������Y��z Ӈ=(����[�Am ?�K�%B<����2��Ud}Ѕ�L8pS��Tv�v�՛ײ�����%A�C�/����|�ի�X:F���E)hH�PD�ળN^��ivZ�5g�^m��Ƶ�ٞq���on�DH��B�����y�CcHȎG����_�u������V�'3� �B���
\`��c�~0-&τ��݂�^ ��J�,���	���"�|���^
J7S� ��Zvk���S(0,F�-v��fVU^����K�ڠ)�0igg�,��p*m?��6�Dg:�Ȧ��:���A��W� &9å��Y�?�X�k�}TN#��3�&��!���JrYw6�=ޢ|AEk�i��ߪ�-�JnM��5{��+���C���9#���آ�
�̫D�P�L2���{b`�����z��`�V�a��٥Tk0nG.�;�3Q�����iH~�h��~����{=L�x��r�
ޢ]�k;@
�՞Su:NrSE����<�>Ѧ��E�;n0�����v�d�9F�=>�5�9�U��xT��HQ��V�<#��cٷ����-�q)s��1����Y��.J(F �).d�$|��_��s�Au���*� ��f�t}��f��lB��J�hɹ��C(�n@i�ʈ,���4<��I�����|���0j�����Ӆ\�5��U*`�0:]�k�M�(�R���b��kل�Ƭ�c�n��ś1y��p2�N� ��a�"��AY��	�Ȉ��u=i����I�3����O������d�v�ewF�EEW�֮6dy?K�7��k�L�}���x��^,$G���'G���]���m���ez�[�Zi�grD����l��ag�/a���v���C����fS����Q~��x{��Wʅ+��=�N>d]�Vz?� ���Ś,s�w�YW�e� u�"E���T�V،��St���Ճ8��Y��ZCJ�@ɟ��!e�������W�S����J�}����'�;��O,K��1�m������嫯�b��kDm�1��S�-�nYSaO ���\޽}'��3:��-�zd��
kb�z{����_�^�|�\Ȍ�����;���q�(�I �b�N����Z�{�횀��Q���	��l��}�RU�K�C�48��jL�~��z��]�Rn�:�<��iM��׆��t�חruq���6�P���{�� M��,l�,��K�����-YJ �k�n�B��p]�s�ڒY�>h�@Y�����p���7���������-����$���=�b�F5U���3�/D�S�sEv�3pA��/��Ǐ�X3���1�cM!3�nP����=[�u���	�aF(�����38�����7����2�g�<3�)�[�f�A���#���'��Q��X��)Qџ�2rd��2h#YiOo�茮_B�$W8
�ӳ�DP���.�(���z0 ������U�L�r����\��݋NՇ� o�1��z�(dn���E|�6��߲�n�tO�a�ikRq���L���tR�&,������b�m?}ˈ�ؼA�S���������Q���[�o�J���7\X+%��`�j���f	!�%�8�R�KU�����E�V6��~��������G^�nu(p�8����Ȩ�x!l.�6�܉C��r��p.�����.v_��xy���5��RaՎ���t��B�
͛��|6Е�@Ѷ�eGEm��( Zh�NÝ[�̉#'�$���}���WD�+8��Zn�Gbj=�4,R� ��P>6��h�+%�:�Dy1w�5VV����1�ZPi�4
P�lX�38 �{tޥ�2j�����q����"�a��|)�gd�6鞡{���Y�4� E�F2G�5��l��K��ƚ���kp ��d�ĳ�
���!hrqT��R��xS�;����#	�U�#�L���`�)��M��*��2^��t�i*���b�K�.UF ����X��x��Y0���!���9����j`��+3�4�'�� ��/��R޼yMp���-���� ��������7���mo/	����o�XOC�.[h\d�ey+�AV���h���f& 3!qQ� ̀���~7G�f���\��T����<ɋ�3�,��Ψ�̴ ��q 1��Z*�-�˓Z]�˘�Ъ�D�Ǝ�fN7&pz�l!�F������l{� Y=��=�f�B0g,pU�|cN�e�\����5sρ�.�a�>d��	\�\�0c>��4M�Pж��/,�c��;��I��4���9�	kt:q�#�����}%s��
�U]p"�+�CR|�6���͵�����Ď�����,�h�����@�m�nU1�9���� d���W�N�2C��K� ,�S�n�<ū0n��b��8�[D�O���U�|�7P�BQhV��%�j6Β\��!J��R	�����W����J��&��RT���C&mB�\���8���)C��HY���<��(ب�踏��LA)/��NA ��	�3��+�w
�T�s� 0�E�Nf����9�W�s�zT��9�Q9 -ը��*.��X�����K��&�	/�ɧ�T2����@�P F�q���}����ɗ�|����g���@�[0F�j�2�Z�S
����V��P���e#�h6�Oi��ƍ�gg�qD0��K����-�N�(���2}7�}WX�����,EKas����H���X��������`�2�b �W��^����#MȕY�R�?쬀��4��S�<*�܉�[k�B���޸�-����%-��(dZiu�����Y�'H���6�W	��{�Pg�1�AUgoG�1��ӎl�sI�Ǝm���
����H-�����|8,Ʈ��S�$ul�䦑�e�:�Y�����O���QypTw.հ�$R��=����j�;�J#C�\��4��J��U�Sm3�9F#rtw�w����k��t�6��	 ��vF���~���,>�E���YB¾�`feČG�{K;��Yc�'�:���W?��R���iQ�>�:�e�� `�ɹ򹵽��� :hh���"H�SG''�)��j0vG����k���{+(�=�y�v,�/k�{�!���7t{w�����#���M��(\{�3de@T.��em�̫���5�B�"��֦�%����r5O@7��!ˈL
�|��ϭ����FK�m��R'��Z�k��� A��GV
f�i�E�3c�B,S�\<Ry�����+̯�t���}cS�D�O5&�Fm� ����!��gc�VԌ�d���b�KNX�MO|65G�b--ȣ����"�
ԦsZ�{��Q��m���sy����� k�#�v:�3���>?����{9;��{�u��wgw��ֵ�����t	\YH�@�E5�l�53���Y�
�j�U:<�&�vP��e%+
�� v~�����O�ã0������t[�$+x�u�v� �A΂�N� WкD��[	�3;�1���-y���v�<K��h�=�|�J��߮Z`��q�c�`�(��m�
�C���������T��ȠS�#Ŋ3��7f��ف�L~eQd�O?|����kY$�z?��f���<�!FSŘ�&o��~�1?��V�Aj_��7�d�V�F�QlD�t�a�c��j�!�F���4�-&4*d�*��Y1�Y!������"$�S��M�-h�D�j��%Cɋ�8�p�X5-��������rm*���ǖ{��*����
5-��4�K����13��pm��7-G��X�.EN��HH.�a֫4`15�����<;ؖ��5Dc��ѓ��p�v9/Xr����njm�U�"I��] �]Z����d$�V������.�P���M��R2�K�4ath��¼$�o��\�[� �NɻH���eSy}��Ȏ����>'e�TՒ ;M��N%jL�ՙf�\.����n:�[1�\Y�?��Ri��a+�U:;��\�������^ ��M<rk�@k$��kT��F�§�%�༨75���M�,�h�*���z�^ф����4�N��8؛� ͤ����>�%�ʬ��+]�Ӂ�b<.�Q1ӥC�UU��!?�<�1xf����Աp�|��/_���a`���P|����s7y}!c��5#��߇�:y G�`FL���up�'���YR��-C&.w�bvj��p2Գz��VrU\G���pк56�5��;��@X��=M�{�V �2���(C�;��j���W���%[(��4_qh6:�s��gZ�9Q�txp�yI,!�P3������|�Қ��B(������1��\;?�܉Z��hs���Rp�.�1}��:U�%gF*��n7P6��Tm�Rf�`@Z�;�\ ���
�M�D�3k��ܜ�)�R�j9�ٳA�a �(���ȱC6h��)����8c�Pm_tHx�]��̮!�O]M����y��5+f{{`#g�@i&�P�ղj��s�&v�G��*��>Q*�5��\�rW�\��T��ƺ�ΰE�*��t�Vn�A�)m8iJ:��5ώ��g�<H�彜-dݣn��A����0��s�Nٌ6���~�/G��~}� ��2��{���]��s^Kt&օ�6���)�uT�4���s��̇'��'I
��yg,k�	�=��t]Ng�VZk[څf�
f��M�dv�I��J']��/�"�ӋƘ:_c\@��]�N������9n|����'����=kf��0r.6!���Qh*��P�F��f���ce
�d$Z%�S,��85G/��,l��ޫ������![�_'&y����yĆ|/�U�xl�6���|~ �;3`�Z�\���cA�o9e�4��|.��½�i�A��p(Ӎ��6�I`E��m�����f�Ԓ/%6,��<�h�d	Y.�Bݾ�T�4�����w�Q�Ƈ�+r&�x�&%��_S����1�����O�!Ŝ�:�8���v���,�o8ND��U�ph�ܒ񸺺����U�� x#��W
(��\�<-eiD!�h��)M��27p�ggrz����pk�ܠ��ҡj�9Y�::����y����_�_��y�� t3G:�
G<� ��q!��(���ɷ�%>��k���������ɭ�t]ǞQ5�h���w+���o3"���qssE@�Ǌ��6+�k��|G�4������v����������ְ�(�a>�� �=�U�W��{_��4����_ij�z_͒�4ޭ�� �X�6b8��*;������9/�"��?2|(7��E����g�6�c:���5� �Y�r`�T�Gv�Nn%g��i����^��ȭ�}<�O/q��Mؔ��;��Kuњ��~��xx�}���P����$����kJ4�ݧ��x���_�Ç������ymo2��W:���� Р؏�!�u��B��TK��H�k��1J{�B$O4g�M������>���4S�}�`k���*SL��5!����$�٩�{�>�S��p{.0o�ՂRaԌ�2��DKA:	�K�MPO�f�"���M�e�'�2>�V:��0(iٞ��_�$���M̈́�A� Y�2�� e�-ȇ����6�ų��3>���b61j	�#Gt�����2 �^.�z�5��2�3�Rkyɀ ��4�&�3�b������T�
��)�4x�*���K0���^n���Gu��^p![�#9���-��n��SPssK�1�7�7�AE�لQ*W��A��0�ZV^|��K�9� �p�U0��e��Ul�Q�> -%)Z���,�H�9�� fO,��HF���6Sd�V��L�����F�V���#�.m]v���d���{�K?�Z}Jp1C��t�m���	9�
���BSq�P�JF`�=���������u�ZM:`�-� �9Fk7S�����-yq����$�#���#m��U�CQ��cp�_�2��0E\�``��Lsh,���	�lp4]���nM��;�Z� �L����#a@"�������h���y��������������-TN�UC���O,mx6������Y*�J�X6fc9��a
�E8:|�����D��=��Z��7Գ/D�t,t%XCi�"�
]iu?�������9�r9�
 ���.�������/2ѕ`�����₂�6����ۀ�w(���N��I����k���d�idD��~�w a0ݸf������hؒS����K�L�~v��&���G2� b#]t�_�5� � x�@����Ut�u�(�͝�맆���:X�S�����)+,;D��R] �~�<6qL��yBڢ̘��0{E�O�q��H��s���j��� ��s��E�ο3[C	�B�N]'�3`,ɭԙ��r��R�k� �uyD霯,ˍ{Xut4p|(Eߦ�����0��V˪	T\�{�i���f.ߟʻ��	ֺX�Kҕ:S���WFB�l��ŵ���;��Љ	W�� Y�c�h,�!a��<
����w�ޑ_�5"�0�vQi�@ǘi�6�a��:;�+�ؿө���9�3�(��V�f�VhvX@�,Ra�Lv��bFл�o�9�r��� �L��2�P�q��f{9� c��� YǆT��@9�oh{ЏzA�gI
��"�����3+�g��&Z�@5������{I߳!?�V*t��RM�Ǫ,x��%�MO_7̢vZ.c���bJ��Җ��ȑoK^�ګ]a�2�gsħ���jV�`����S=Ш��T�;�I�CJ�.�d3zhLc��?5{��6`b�~�+��V~l�k"���>�6w5,�ޤ����8�g��؆�l@<�����cV)h����)K~��*MR'h�E�k<z"�!=v�%�9�bt�JǗ�٦2s��̨��^�$V��% �N49�(>}=��Ҧā�{\1�Fہ��cH��\%�[�c�j�1!}�%��4F���ܱ֜���0m����_�ߴi�a�g��U��,9���<D��^�ثZ%V�u��Pr+}zQS�9�p_�趀`b���F��67�rt�+�;����r�F*��Q �ݻ�l�U��d:~*H�7��͒<�!���4�����90U��2*N�u��*�v��JF�}���N�E��3'��C;ʧmzJs�s Zj��1\p��=�Ʃ���-[�� i��Q�D��vD���/��Ay�M�|���ru5�N6J
0���ͫ��w�"���3oL�F�� �%Y�*���+��2Gz�-`Y/�s8�S�Ip{V���s��*9�@ JA�T��J��.9	 H0,Qz���C4�1v�����>sw�_e�/G����t6�ãc�QA�k �<���¡b#�l�q�m<0���eU�CqH����� ���	�@������%�3��kS#?M���t(K�(�%
��Z��f��3����c7Mh��R+��A<�^��M&'�2�� �����Di����:{�Y�4��J���)z�ҳz�ϊ��9���E����(��+��<=;%ge��Yp'��W�፪ʮS��Q��t{E� ����XA����5tw�@��=Axw�tL�L�qI�,��Y���o%����|<�`3
��U �^g`66B�ʊ���m�P�����0h�ٞ�Xו�'f�:oX����Kv'C"B?Kgs"K��h5���rI{	�tϦ���r2'���1a��|+�P�q}�ԿZ�{��Z���	���ځ.��CK�����2��N�p,�ࣉ4sN>��D�f`w�b�����(:��?'e
���}\���l˜�ۺ�K㠷����� �jUUE?�k���ޭ�ql�ә������ۯ��#�o�����{.VЫ���k�u��#�#8�JEl�Bps� Q9"�_�5ݯO�W�!�?�s? ���<v�Wk�f�mf�'r<�Q�>��s��$�:j	f�:��CԹ��&M������9���`y��ίD�s �~'��YH:OR�z�6��V�w��v��T���^��ք_����w�����mTY��F��D	����H
�Q�'�_X�XT���Y�"�u��&t��.}& ��2�'GEj=آdޑ��5��Ws����E=0Myf�E_�]H�!kE�y�TwL��:�?���2�0�v:��=�O���xS����G2��@�jwg�����R�Qؾj)M`�xoZ&R�ԕt�ݪ<]��S����u��G�t���i�a���%�7�~2��̠
��@ǒ��'���(,V.^�f1K��.fV!���/��^x8n8ݕ;q�m�HtF9 \l���m�Z�LS��B�]k�_U@g֣�(�1����s.n<T�=9�0֨�2_,�qM��h�s�$"���A	��ߥ�;���c�N�e�x��QbBI�m.5B.���
��ՀX}�t��v��&2�\*�:��ap�J7��7u��3�>>^�F�X|��b��csb9�"�Oʚٯ��K�kjY]�uc+E��?�u�{@�݃�#o�6Ά�m,	� ����l����Y��P�P���Z���+�3�@�م9��~�E��r�\p�j�@{���l�Ǳ�*a������z�9��x26�}��w�k˸�]�g�ץ;p���a���p=�����\�O	��RjȺ S����.�9z���R��}��VK~���Or>��ʴ���A��ŎH�O�-)�����{���_'0x���4�T���#��$;����[A0��D�h�(.�f0��5���%� 72� &}pH��`�	۴1�L6aLۇ�p}���<�����s�"s0���h��%����C�"�[-��X�D���$�:�`�)�q`P.3:�4'��+���-�v/��i�pw�g� �W]-�z�)%_���?_�6���"�>�LT�g�4[]XРC��b���L��xJ���S`�M�?-��ͼ�<�����P��%Ĥ�bg3��}��H"�Fa ���S��N�������2[�6� cw�i�Wڪ��b4M+{��8�/���kZ���.��'6@�	�ywwfr�|��U��~�����D������!�������S��J�WdN;V�_1fE�Z���%|H�oMKѺĉML�Y�t�wRЌky�L��S��UTT09�B��v��(����SA�d�N X�FA̚t6��҈n<�O�W��8@+%��tTߟx�]�Z��y�a�(�W��z��r�f:z�"�y�S�1Z�.�_gd�� �(�Y�3לuF�4f͔p>M�po�n�ώ�x��� Q�P�)j�U���$g�\rB�&k��1�V�_�N�)B:���ж��q�o�F1�A��?����LFSQI�Kk����6�5V*�����K��\��J�cr�>�̀�S�tb13�Ь�Th�o�p>}���N��w����˗�ZFFP0C�����fS�a�GNOSd6_��Zg !�O��A"���� {}r�-{;[\kP���?���^�����@н���=U�q=O��H��=u �Z��AY��e�mt���R��/�/Q2k�zr���Ҹh>�S� d ��L�����k�vpb>��?� ��_aɉd������A2��� s2	fZ�U� 1�I|D��u���,an>��ń9�5��r�$6����lF���B�M�4�;m~UX�A����D�R��;m�v��q�[u�����R+������ao�}���*؟�Ɩ��ѳ����y3#��P}09_��mhV�a柃=�u|}ugr1AϯS�fT% G�+kf�p(���]�����v19 �)�+����UV��Z�	�ϱfX��Hn
�Ԩ���-h&H{����b�5��ks4%_��?���R�W�\'����;������ў������oo��p|�� @a&�q��T�����ץa� ��*{��F'IL�� �foG~_|-�߼��j� �_FfL�լ�m]e�GQ�&��m'�� �����cT�"���u]��g�C�KV�#��;�yAm��昝����=�E��������ܷb�6��Iұ�>J��[�� e�gώ��/�������*�������D�I��("@��u�2 �9�ܹ�������O�@$��9lɳ��w���Ǭ��+�E8���t���_����S� l���
������/	�Z� ��
B�ȡ�T/Up:��zߤ��U���5������rA�8�c�C�|�a!��S�͋�>lmDZ(�4��r�Mދg�r�0�2�rY��Ѥ)gFk+�c]k�)3p�Ld#%��CZ�1A	��ު��Cӗ�
LT�g������ƚ<��EP�!�(�֦MRM��LPuz4����1��G�F�l�8��𔥺X��j�U��]����hd��-p��6<9��/�4~�KΈ<X�v�]_E���?�0��(���ጶ�`P��$�y��W�b�9̠��U�#���Ɖ�˂<��VK��_�����j0Co��0%���i6�&�ÆQ/M��� "��Р��ɍ��]����62~2��}�qg�<�=� `w�P�lȕ�Ey��#��*?���&�rc��ER���a�-xp�H���"��-�U?U�F0TW
r���Qu�jkL kLlu��&p�Q@Mc�l��-3bKM��J�R��Ǣ��4���DC�n10�tb�y����ﳡ��>���˟��ș0ə9_����=� Gsb��X[8αLpȚhb`?*�/s�Ei]ʚ5��[���Ѡ̋�9�-��.����W>�n�6&���MoAnX�bC�Чϛ"Ù@+�{�6l�f7�G��AǢ���9{�2�Z�_Z�X��?���,ى	J�e����6�v��]4NT��м�©�8y�@��{#E���i�+��o�jX����ę�X��D�����C�}!�7W촜�����}��|��e
~egd��Bc�x�Y��2��^�a૰`Nm
�UmA9�&��>��B��eAs�-��V��lR�r M�Yb�}^���z6�T���#W�&@��u�4f����	���A�1)�T�5���&(�6�C�ڄ8��<�N\NJ�Zi���� @Z���ݝd_�־��;
2S��4�4�Ҝk�F;�WL�,	�V�+*2�϶���S۲���@�fa�2��>����0��5��r�x�@�dw{Kp�K<�uձE����YY�eC� ld��àv���ew^�4��<��r\# 7��;�G	b]�fe��L3p1X�%?c��`s{���F]yI ���s>�	sFKm�1&Y�6�4�M]18�E�L�[�s��8f���Ѵz�:���$���a�����S�W7�/ȥXA��H���J=�4��`�U�ry7�nԒ�
߱��-_�R�|�B޼>�C, |b�_���!�!ˬ�|w��w �̩�SDgMcYB�0L�|� at
�Ls2`(��3�k�������w1��ހ��I�Y��!�s�hF�q�"O�)��YP�kP2C1�`�/�"��M�z�!֊aC+t���E���o�a�hY��?��������c*��������rҬD�{���j&Aa���S�G6�C��~I %t8ܯ4X����wN�1�L�KF��Ҳ��Dr���eU�$\����:�6��MXR3F\�N�f�b�:P��o���cű�}������	l~d$���p8�o~�;��]����g�ż���
Yv������d�Ţ��_`�8�\{Y/�54������u�R)\2}��vk��;V�oON��U+��Ep-g����65x�YL��h h�Pp�����W�	`�Ks?�����&����(ٚ9�	%st�b_�V��3�(&�� �/Ӛ}��B���(N/�b��;ĖI_C���x�Ex��v�"K�z楦�D���q}0�%P��"�zT�:@|����fU�������rI�wvVr|t��_��0��� ������\,�����?���&ߦ={��:'���A�X��U[Z��q��7Ǆ��g�<�:BM���F(tm�hp��s��."����m�l�{��R�>9z���>/����P�PH���[��d�y�JNa���N���i�*�j Q��}V>>��b�lxV���{PGF�6N�L�o"w�)�t6p�3��2|������6��ki7��3���/�H���I\����¤س�$!\\��'r�B>O�(�pJG��5��%*��> ��7�L��~�&'WR���fQrm��.]��US���;���=66n�3̣����o�Z*� !m?�dooON��dZ�Ð;��ц�Q.�E5�K\u�.���)��"��4�b#�U�Z=-L�#�s꼼&���ڥ�ՌSi ���+9><���s���tv-�N����`{�B��tb�`�{P��2Tr:���~�L�����pa�2$�$�!�	���wh��m&虵{��_��D�\�[��z18��Ţ�7�p'�:L����vڂ�õ�n�={�g�k3{�^#�Z���'b7�d���*�X��f�pC`��Aw�`I�e�i\�`&����G�U	Zg�v9�U�Q�v���r�aė4 <�<���H���~��Sؔ l2�� �	� Wi�l�������Or~u+�rz�}��Z.�O��4�T��/�m�@OR���fr��)��y��,�Ԣ�Lm#1pM���h�7x��8�������~��x�|'����u�
%�NLP6��2�.�D���uϦ�������A꜇|�\�N~� b �-Ϝ�RCi%�%�E/�_�����e���#��8�Z��q�~�e�1�:_2�[��si�u:'p
w�3H�I6��hb��
����ٜm���N��

��˴&�ݧK���(~��RZ�\�h��@2H��RIߣq��	t=K�����p0n��~\�.�5��4<^dOg*����y_G��,�}:��M๠����Cb����������{������o��B��Q
{�e�[yJ��V�R���5�`�����]��(�l߀a#��v)�4K��aJ�Fd�}��.���'�}��^{������6�O����b�ol�'�����'$�c��9���o����: ��lB���,ٲkv
c�m����C�":�i��t��5��YZ_�H��W18>����#�Ub���
Bc�B�*��^j����N\�>�^�ź���Iؼʚ��r�+����I45�(>�ύ�v	{��xJ��5VqBQ������@�@S�RO��@4��u(�4���a���&4�AM/��s�D��:�.@v�E�~sXF�Jf%k�J�C��,��I*�a�R��Y"�����,C^]�ʻ����"?��N~M__߂���E����Ä�&9�ŕ�Q+��ܟ�ț�G�</�A(yIM��5��6�g�N��F����̼o�w˪�>-މ��Wb�<��OA',���{<>C����snA����"o��� 뱁Z{[��ix����� ޼~�u2�|qA��H�T�g%QZ ����|>tnB�}�����Qr�[����i�����/&�4V�v����;<���s���'�5xvuG�����ls��{�0Ub��joal�ɳc�����/^��:N�K��í�:��q-t�6����"9@-A �L�'��ʸ�n<
 @�˲��_�J��!QՖ�㭉9JJ�D<��N^m8Fi�F��T��0ù����4���k��>���Y0`����
/��>8�<�І�������+�}$j6d:�L�t�
��i���u�;[�λۛԦ����N�5�h���d��2�-�G�z�>�R��h�MP�0�B�6�IV��w)�O�p�.������g��w_%�vr$��1V�cWW�1�K[�6�������!���ڕU/�8l�{�drA�1A<d3�˙�v���q�Q�M[k\h�ay{�ڱ&"p�6F�mJ1̄��l�վ�%���m.��@@?����y���=}ʖ>|�:�����w��8������Ï��R@�Ў>��0��	�w�87�*����k���w�}�S�D�k�KӋ,[9H���'�e�N��dcV+KC���UҞY�L�z��^�}���r���
��zo]7"2��8����ƭf�4�����e�J���$>ے7[��9��>l*��m��-d�4^��5�����c�m�%G0��zd���F9.LhPk�E��!�H��i�~R�&wy��j����u����r�!�z	!/����U�k2��mU3k#^X�o���L�D����Ù��_�����K�U�X���W��^2V�{;�=�x��
4�Y����p#�(�S�}��و�����	����)?�e�l�5+��#>�U\ϐ����΃�;҆F��.
�s�6o��5+��A��!���u^b��F�Y3@㽉\�,��x~y�,�>�kY��e�JNOO�	����� ��6���s��Z�S���(mG�=x�)N�iZc�AF�m��X��4?��&\S��t]�(�1A�v*/w��_��o���|��e������a.�m2/O����#W��{I�S�UѴ侀3���fcf����"�c`�����s�:S0_�7��������E�ֽ��LY���օ��4�����={O�N4��#Kb��`��s�XfC����=;�"G!����39><�J����[#4����Y���Q�#� V����*��еY����&B�N�����<�B;�! Z��![{��+��5�DI�J�����Ե
A F`�����n]`�7t>�^6l�
\'�����z��1��A>G�|E���T��ڜ�J�+m��,�d�``�A@a��u�3�)k��ǽ)�AW| ��pz��k����8���<~<|]�����/��G迠�������b�G���Xv#v����� #��GG�v��\���$V=S3�a�h:Y��W�� �H���y��X��m>a(>�Yed�'AKjT�Sa�����}b+�l���Q�Z����JK�yY���؃0���/��}�УǞ�}I�ߨ��i���B��cP�0�\3��2B\o�e��_2���9|�\6��x ��_]�C۪3���,f@%�$�wz��3��[̓ݭ)It�7���އ7&��S�;���/�qZ�E�i����R��Ï�����䗷���q$���WA��(/�/X���2i��k�����b͈�~?k/,n��X���X��g�9ˣ�k��o���?��@��p�c|����D6n����y�?�߃��~iZ;�\���\9j�mPF�nު�v����� ���hHs���l����;{��� �0��&��y�)���ӌ.� ��Txs��~=��l�h*�����n���X����_d%�Z���G��ӟ䏿�B^��'�6�����O�����z#��?E�-��W�vrrL��s�YQ"B�d����)�����Kfc�
ηd:��@��	�vs�} ��ñ�Q� ����0ҷq�b�C �+�2��Q]g�!=�0��,7�;j߹�kN8;hX1����ۢҲg(�Q���
���z���47���"��o~���y�Bvw6�zI��H='hHhǿ <Ʋcp5p�) ��9�amt��6�Q��39��(�ɦ�[#9JΌ�.K���dV�n$�G-�Һ���T��m��7�@�p9�
�M�~no�M�ێ����f&G�fN)�bK_�N7�fd��3������UzG�jH��c��`?�ǚ�3�����c[�n��zh���u���9�^W��C��}�������QE!9=��M���r~{�	;���>����y��LU>��Xs��m��������.hbX͓���f
L@���_�W_>��]d���Nݖz�W��~C;*%dЕ9$ѩ�bu�]��v	1׻���i0:1@�c���G�uVI��`E���+��욹ڂ6V�;�a��C> ��	pv�����d�r �2�&�PO`��h��ɼ	WkUw�rd$�R4u�D�/��,��@���Z/[87�Ua��L���c�D���	!�\j�e.h��&��.>���1D�JkBA�����If��)�<9ؓ��t'���_��S��y*[3�7(ǢZ���y�[�+���k���S ���xk?�����>�Ɂ���Z�ќ-��%��ư�L|�<=F/{}�>j���Cj���������f�@'h�G�MH`dwsJ�ѹh
��ɑ�*ڸ��!����m�MT͵���S��]e�C"c;��+�1����0���l�5�1�M@�ɗGa�^/΍�ΐl���/_��d ����������cn�@��q+�IZ)H�ȸ.vw���k#�B��Ӷ
\���T���ˆ�=2���zB��/!wap�{4p�qpl:sR�߷�,[tM�v@;�S�lE�&��!�	 ���nr0(�]��r�A�C��Ō%��mĦDd ו: ~�g���&:���Gٕ3�p���ֲR�1����k�䎝�*��}̎X�rg�) ��V���c�Dˌ��wٓ�O���9e%���Z����r�%e6�#����u�.�"Ӽ��v�]����ѥ|ߛk�,�yq� ��ӛ�'m�C+�۰�������ߧĵ���q����0������h�}����O�3�B�0����i�T��#� K���>�^����/6�!�	�d��q�pM!��M���LjS��R��Ǭ�Zq?����$���A6�� �o�Zo�|
�_��:�_멚�{�4J��yO�Khq"8W�1W*tU!_�x��J��Є���_���C )���t!o��|�bD�$��l�`� ����@��M��<�M�gĆ'D�{e|�?��U ��	5eS�f�D�y Ə:E�$|������5���i����@&J��������d5�e��,-"��d�г3�������O-�!�XOZW�d��1�?�����������91������Z�J�F]O���1|���Q���p�i�e\V ���x�9U򥜘�6�NT���X<;�g	zgk�e��4QbҲvK��"��w�P�yԉ
��{��1Fd�M`�ݧ�ή���3Ӑ]�4B�0K2J�m:�d#ۻi=o��QB��Zk���?�^�6�hi�ɠG�rJvD�~���Fc6ۤ�>���c9<<ҙ��Y�e����j�e}9'��@{�-R=��Y�>�m�7f���c�7܂/m�V�	��nKt�9/(�^�K̝�0sJ���݃�^x�C˳.ڄ��o�O�"֜���u���K���u��ە��{��(#���\�D����Q5@��J�n/ӿ��Ð�&y�3Q5�]�nb�&`,f�#�d�7�Q�����~����&�~�������&_.��V�(0�K^���Eh��l��db�����֌�-t	ƣ��+iO����(�ɨpR����V>�{��nh/�C�����߯���}��W��>�s���q��������!���$��}�:�e/�����.�5[ݥ�Nv��|����z-'�1xL79���Z4T^8>9L��p���*��9�YnC�(� 4~��'�S(a�˙����_9����}�Z�(�ћ/������ �Q`
햵��t<�u� �a��P͝uy?6g�8_A�?=�AS��j��[ޑ�U��������,��k!���^�q�aʺiM�Q�+5�^�,L���w"D����@���M#��� j�����)o������������u|�������q}���F�
�9�8HG��� ���"��۟�0���?�|8�����@s�A�c�0w8���c�EA�rh��y�� %F�m>���F6 �(㛗�d����D���r�,3W���r����ʟ����{��Eh���w��/o���K��KF��8�"�0�:Id,F��\ty2'��mݺa��"˗1g�^2ȕd�^.5�<�md0pN�窂���K�������Ɯi`����*-�gɀ�� Lo�Q����eE���,�O�~ϔk�@}�>b�M1�c$�z���9'l����ڷN��ڕ�^�*_����$ �U��L<��ݽ ��@����Z��v����f��TT�*���L|�H�Y-����5h!�L8�+��0%�ݗ�&�K0mݎ���:_�b-Bf��&Go�S��ޫH��h���%[{'	�Tvŵ�Z[k%A�Z5�i	��&�c������?i$����J����W����|<�m������ZA��������ӿΒk��`}p�za�>���ogE������r�XA���1)
���lom��_�`���p�Y3�P]Q4xE�Z�=G�hcs[�Odcc[��IqY�#J��6�>K_q1��a��U�Xsag\�px�!��g��N�Z�E#*gh������8���M,em{�W2`$T�[����MM���K �,�D���w2
>%QT�rT�k��l��w"�/��(J���cV�+v���<���]���ZNI���Cj3�����}B���)Ժ=�vq�4&��(mwwS���uq@L����a0,J�.���4\�Czf�ֶB^���Y���M2p a(�����u�o����m^�H�^g�N_|B>>�'�w"�|~������7��Џ������yS�0_:ҥ�j��9<*<�1I��@��U
&�y�(�Tu�n���s1���������8yT������'��?q8���B��a�c��J�I:�N۴��D,��.�;�j������	�uym��2���Ɣ�uе\ ���#�?|�2di�!p{;c���;�T�VQ`(7�v��l�D#�_W
Y�2���H˺e�߻�p����#����B8Xg���s�}��Fk/.C/)���jV6���a�\\]r8:��㑭��V,yk'��4�\O�2�C��GÖڲ�Fv�}YW}�doG�x����1� @m����\pOA�t3w6� �Ã�my��$��@�<D�V��#�9�������C`P���Q��T�G0qy}�r�\���Y�h�ȭ����קl:K����Bu��S�s�������@>�X�c���ff=ff�ۭ��|�����?㩰��f����X������H�!��� #��1�V:�(�*�V5��9�ߔo~�F�x�b��.|�H �:��a�x�|4�Tës��`\�B���*O�P��j4e�J�N��6a�)��^�sW$� )SZ`X�(?��h<�Ó]6〾�%e/��%���N�Y��.�Ƈ���u`5��-	�:k.JA��"nQm'�N����8��@v�Q������F�D�Bf a���d���V�X\�
8�&م�����F2�"���ר`ܹ�D��	�%vz������~!7��B��4cg{-B�3z�W�U5Ϸt3����I_By����[3 vo���p���L���^�޸���7�c�4<�]{<�x�G׎��>'���:ML�,0�T�rn�N��f�AV�R䴸����K(��8�	����� e��.�U����UKɓ_ ú��*rXr��Q��83�wj��FV���[��l�gI�Z0�`m���=5:X�8p��}�N>]� S
�Nxũ�V_�A$q��J�Cm��8��*��׸<���J��`��m[����a�I�WߣE��a��f�{�����+|��sh**���2�juO ������{������=K�y'����4�}ڡ��f��~�-�/��^�x�A�Џ�����B�/����S���Ɂ챥���U�t,(�R�������g���Ѕ��|2�
����L6�v�.P�>�����Rݩ�.#��q"1��8�e�⥚���n����Iȳv��Ԅ �ױw����g�к��Ͻ,<z��x<eaŬ�Ъ=����6�3�Ǚ�a�r?�y��x���e���r@x_��W��Vjъ�/ tI�����SP�DP��6K��(F<��n4��������FB/�nƿ,u��S3暁Z.�c���*K�����v�y����m��C0I�p:���C��SV��s�v�z��|U}�j��Z~i;K횠`J���bƱv�D�pAy��0�M���f�y׊ �6�?AKr1��ۿMיx�n�����sd��#�Ѹ�`�2�~A��Z]���or�SAi�q�C��ev8Y�:�����:2��C��'��:*Bp�ք3��wg���q��r +��k��3a�m���!
�����ֺ ����{<��S�����S/��9��|ks�vrC��f�E\kF]XQ5~	::��s��U\�(�'�ʺ�w����"�@��z��G a�Ŝ��B9��&7�͖�}��5v����Mc@�?�W�J����kD��0A�=D[?}��C�f4*�	"s�Y~��q��<D���#���I^�zI�/d�5�&�0�C��D�%��j���WG^��=C�u}2{p���}1�x�O\G=u�Q �A��!�6����fX��~޹<*HY���l?�{�$\X�����A6�"} pU�UAه����ﾑׯ_��R2ȹ�~`T������Ⱦ�psڦ.f��2�?4I<;:��}�:B�V��?$���>���o�bV�$�QŬ��D�e�pȣƠ�����Q�	�|���3ClØ�E�2���R����v%g�K�� h�lݢ5��@��CZ͎��AxT a
�*$\�ST���c��ك"W]��CO�����p��c��uD���2>��z��%��_�����7��u=#8����=�+�<l�Q0F��9
��h'�ɿ��*7�����:���)�G�:Y��І4��*o^y������x3eƱq�=��0T��,�3�����1�SG�LA�8�0$���Dʇ��N4{��q�3�t��H|�j$�(O%�S[����sޘyH5amk�T,5H"�hf�'t~��@�:}d*ʼ\)2���Q�8)l|
A�uμ�������d膘�(�������ZpQ?܌H%�&�d�����1K�P	���5a�X�`ѕv�=[4����l�È/ZK��[߈��
����
��������r~a�ʆ��s��o=�7�ߌ���A�ܣW^���%�+�Z;K�,���dS�����79�(h&Y��XG�p��+�����{�����|ц*� %(I!{�5�Vz�M����u3�����`�)�c�`�G�XP�rz`Mw-�1�P}�-���V�aD4�^�����1b|ثWoR�y���M68�҆,�JA��������t$�Z���e�EK�����s�7a����WD���#��mv��Q�2�̥e��z�r���ϲ�[?����p��ǎ�9�y�r����s�SM�R�XQ�Mc���,9��cy��x�B��=�Y�5pqy#�7w��]RК�@�|T: oP#����gt�)�J:��6�	��i:�v~�5�������Б�΀t�����{�Oum��Qj|�����ZyX0��p��[V�3F7�Hkf�r:
���PT��&+t��B��O+�8m��ӻ�	��7=X�1F3����]Gp���Z37�e��
��/���=j	דrn�ڣx�^y��O��'�_2�����.>�9�wC�5|��+<$�
:��}��2= �#�6�1C۩$�rt���`90��h#�����~2[7��v�&b�����V�8Ǘ:cKi8�c;f��kf�C�?�0�V�&�Jgk����y���v����|��4g4a�������hf;�v� 7TY��$W�v�Q@��vL�M�DAY��w;�y�3`K"gtL�|��Q[���W��f�Z3��j��6t�5�c\s(�j�B3O�f�4�� Pk�tww[�m>nΜ��<��7��Mu���p�v�3xw�֛��'�������Z[a���3����6Q&����� r���}��|���׍�g��7|x	C$d�:x/��W\� ���X�e����LYps6ʊ�6̅D�LӪ����X�X�Ř�j
UG�s��"��|����zt=�Ѻ��:��ɦϧ�[��捎��ʫ4UTfN��\�m��f:��=�v�]t�((@�h�p<���K�1�>��jTP��b e�1�s	�������*�~���+���a�^�
��VVMߖ
v�� j�%ds�X�|�&�x�G�$8�/��:��u��э��l೏4����/U�egw�9u�|��X���?rn���yO� B����1?tN`�`F"��K69�0%���MfSʇ`�Գ����F���y;ݧ��� �h�����������Y�u`q 2����
�o�$Ǩ��=y���Q��v�p׽��\��\od���VMEm���d��B8�#�$�KX[�w���z ׳nE�u�!�^;��q�w����3��l�w�yg��C��ݜ�����Ap���#��{<.������+P���`V*���׊v���HE���9�k�h����>`�|YM��ٰ�,[(���?3<<�! ��ڑH:���g����J;�q�
�O]t�aocb�%FeR���d
2����Ad0�[��*�e�W�U���U@��AT���m<��:S�fE�+��Y2��t����͇��:͔)/�6��-��x�
OMkk:O�T����A�	�>�~�-5r�m�*-;�LJ8% �H�@t\ґ�J�n����~�p��ukOm���7�4�U�@f=�l� ��|-D���P�u�x������mV�`Xv߭&f5�Дy�o��ȏ ���Y�[����ӟ��آ�շR,��{S�-����Tm�筨�Z�at���ʝu����8<�'k;�2�RO�G�y��%BJ���J���;� ����5���0(B3g�(�&>���0{�q4)���Ĥ�zu4Xe��4Rߋ4WU/��CK*4�,#�/D�ѵ�ܙ��1�;�-��F�ryo8j�7T�qF�U5n�� �9Ȫ��o�5���e��×:y�V�p�+��^2M ���_�"�:99I���r/�n��w�����}�����=�W���+��ҸH0.�J�R��3YΗ������A����ƛ��EP�|���K����ʏ?�$���^nn���uaHU�QC#��N &{xuM��1/�	�����!��T:�p� Hu�6��V��k�˪�U4SD-.�';�Hv��k˅D���C�5X�g�y=��
�׬rmR|�ݧ\f�=s�m�e���C*m$���q�_��k�f��x��v�P�P_Q_�6l�tF��H�z���~�C�#�1� �fc�	."8��I:n��,EIkЍf��b>3����P��#ة���S����N�d��e֐+��$�S+��T_f�ߋ�3�	 �4IČ���?mh�TK�vPq����f ���tqr^Q�H�4�?;�����M!g��7�^�`ݸ�9Bw"[��H�^W�`
RLS���`�b��_|��>(8؆� ��[V��8��D��ZXQ�9<<d=�@%K/�m$E��'f|��I ��E�O��:�z
�t���z9�Zt����v:����X�3�Z�	e0+j(�*i����JK,��E_&���󍖵U�7qp������qE�G9��s�;A;k��Jf6qeU@Ry8���jwn� ��3;�zX�hA
����`��	���҈պ(f��{(!B��[��i-W��t\�!�I�bGЈF�ԑ��ã�̍�B��r/�*����5�ЮG�A �Xw7,?�완�D�Z(>wϳ�}��?�o~�B�ga�o�֓Y|i���@�^�Íu��*{�Q4����'מ~=�d'W��ut( �TٞNST���[ыRɷiuvN	��I>|<#M�%h̨�y2Έ5��`���5�R�	M'���eoik��ʴ)�f~�>�B���'���7���_���ȅ�:7c~����Zgw(_^���_~!ϟ�<����;9=��h+��ҕ����"T���[��˨�<Q�)�>�ъ�
�zC�����V��Y��i+����o���(�CP7����n?���J�@�7Z�g4:@��{a�2�/2[���l���q��ע%���!�}���:o�q����y��|ޞ��)琓GT�&��
2�Ʌ.Ix�d`<Ò�;#��8�LTY�ˍ�#ȗ婣~�J�_������Agus��1��=����9H.8�v����0�����$�'w�ڱ�Z��gC�K�5:�`$D����nD�_5:Ëc7lP��+��o�A!�U� =K'�h,ˈʑ�/µ�z�i�S��W'f�y'Ȱ8/rrH~�Aû���H�S�yY��io��`�D�6�goBȆ2Gk��?�����C���D�dݝ'�n����U�6}Z��ꆥ`��>Fy-�5� ,�KV@��*��p0���%;��C��f���vC��.C�a���v^0�u���}}.b��N���J{ډ�Y��F^7�!��>W����W�Ih�\��oUgdP���=< �U���%@}�R"���=Q(������ߨԬ�6Fjԛ��������)9?�K�u�Fjɵ_���)�3���Qm���,tTWTa��_����σ��o��Kc�&�ۦH;�`"@��ЇZ=|���ǘ�yj 7 �y�>8ޜA3���i�ϩNkj#ݯ��M������F���ا��[F�l�Xi��.�1�5 unb�z��jCf���t��q��m�a�Ɔ����_���~�5�O	�wY<�����}.6�S�OKY�F�a\�#��  �Y��0�K�FF�k��Y|��Ҳ�3��܄�+U9�����_o�<
}�c�u�� ���}0|�!��_?(#F��1��U�q��N��/1 �_����ЊK�&8 �g��ܲ�- .������F �*�Q[=�2����VZEj���N[�z���������}�[�6�d:Vi4�����qԲ��+�M�-��%1L�<<��}YCC×�5!���*��F
`URG{>��0�jPy�q/����R�% ��u��eV}�w�{�3</%�����a�y:!p9��9tqE���A�%%���ٮ~���|��|1l����r{�f��A�/_��V�s��#���"�	�Z�k8����;�r�1 �:^�o���N���y��|�£߲-W�E�x��\����&mr���|�n��s%w7���"����k����eM�9��l��J5��Sv�Lf����l&�+�Ƣ;Iwp�i�n���_��o�d�hi}��nѴ�_�5� ͛?��/��P$j� �EL�Ό���J�juK�I��Z�f[2Y�r�As����M)��ƤT8���ĩvpus�e�J�e�Q�T;"��\H���c��ؔ��zI�t�>}�(���S��7�L�Q����S����L��_�%��+r-�4�Q/P:LOdT+G�rӨ�\��i����>�ԋ^�%�J a����@�د�c�;���SX�=��)���L����%�=�I�dA��P�-fV����w��wܻ�U#��K��%Df\��{D$H��ٛEh�@ ��a�nnΨxh驭uZKm���鲨b�C��[�(jD,w�-�d������h��/���D�����܂*}�6k�qy��!X
�`�֣���wVq�B����;$�w�o׳�O\�H-4�����|Ǫ�<ب��#6���l����Z�1�i���+;���8�oX|e��m�����ZԵSЫ��BY
���v/b4����e 6,�C9Dw
:�+>��[O�~F���PR�9������}�6����T�S��^�M�U�[\[�����_��mS��
������J�i;�C�jn���͔0��&���m:=/��N[����� �dX|��.E�f�b��R�5�8�ЪZ�W����Q���2GS�Z�v�c`����	tm�vd��OD�"ڬv��������B��J�r\O�?��K}��$!�@�o�آ,��6����@�H�<�>��bچ�h�;����3*Ϋ�z���q��4�H���|16hP��ir�i0�;�Xy`�Q%�S���s���
��x��ε@+�(�G��-C��1� ��௡M�K	 ^�B�X����R��C(?���g0�m��Q��?����z�5�k�d�Y+l�||!:�� ���-u�4�����Z�p����sO�8��d1Sx/�b@��� >��	�A�Xt�8��ژ���Pޞ�����l�5{�v2�'��f͛��ksVoE�B{�끥��cگW92�K9`K�D��<��C�b��4���F����4�]�3*8��$�n'��t��h�"b��a�p�^v;�\X�ْyãt�o����a���LY�v��H��!����]z�~��V���I� Wח�H�@=7I/��c���׎Wz��UI
��{O�h�?m�l��3�������Q2f�0Yy���U���6>+�I��� 7s٬ԣEň�J�"r�l��٦$��4�{�gCZ�G�u�Xmͬ��q!� �k��p^+S�ױ� oT�a4.XרdS���*OB�l��Kd(�Sk4 ���/����i�h`:�k���w��iY������N��hվ!�3�M��4w��V��'�9p�;�HXX�� �s��% m��4�p�n#s�5���5�zz�͏L6�\8�ߙw��w���U���xYt�]4�֦_��ee��@R(i������9�6����� �Em�B�/����O��b��Hc?����d��3H��d�M{뎸�[�g}�L��,�.V�_�<jm@�
��.QCa*�=ܚ�\�q��yb�<�s�*٠�|�+.��!�xQY�uFY
���= L��DMi6�Z�%�OA�1��LF'cӒ�B'���It٨�y�����*Ȃ��z?EF�$�O�|��?~~�3�oo�p�EP���\x7�F7���c�q/2�!�%���=-�"��
GU�.S�)k)8��ző����%F#����Jn�/���J9:���X��`ͷZv�)z*�Q���n:��z��K��B�vY��Y3�u�<���i\��xu�JE�f:��J�N�1��3Ή���րL��gm�a]Q����,|��[��S�r�"��"���hZ�����?.T�k�>�����Ѿ�&�9�k�����ݜ'Cy-�����o��V���Q^��;�������?0MD�g�%d�ZX� U�T�o�����}u�h���<�������`�A��\�@���������w�O���f�]E�)ׅy�):���J�x�F���0=��|��H��[c�/?���߳����F��j��	�ײ%��Y����t��.#ؑ���ք�Ԉ;�U�S'K[��-L�tn�~�S{�ָ}�ƙ�԰V���l#g��w������Ȟ���%��5���49HUani����{�����UL����� �#j�@��F�h[�3]�	ro��3F@��A�X�U��6��0���1Zt�w�2��9C4}7�T�~��XN����F���_�� �q��=I]V��C��x�W*�ү8� G�  %�@��{��X�)����$ǌ�i��m@���m�^�<DWm_����@���E5*R���@�}���F��g����h�5��9SP���b!�Q��)K��H�yT�Z�x�5�ZtP��=���q���P7�}���<��D�پ��������R���Im����tͶ���'��~�7�?)A��Q��yԞ���) �/��y�YډңR> m9(Ҏ�C����U��-�G�������Mw�bC���] ����0~�h:Gs�(yE��/�tU�L�̢�N����j_ю�ц�{�wo��Q³p��,J�𺔻�s����Ǉ;N�����)���I��J:�Ǽ��G���<� �w�-��	fPÝ����K(��(��=V���ED�9}~Wo�*��ǧ̡���Xڰ��´f{e�t��{�@#���Ki ���K ^�h�(ٚ?i-r��\C�E�A��pw�<�Gy����Hp6��q|�����������?�;����wryy���\^`]J�ku*��{œ6�`.�O���p'mL{��H ���,��6�gk�t� e��	;��|���|����[6�s�m(�Sr��v�\�K�8 
����A���2�i휲y���/�������PG���7H�_�ƞUp>��ۊo��z��Ί)TR��0{�T�DB�6����M\p�3�>^��������,�n�8kH���4Y� =�nF�~ϊ�Ѷ.kΝ6*�cT��&���|E���>fk��S��ٲk�#q��m����`����08<Hmw]�%�����Q���=h�xȟ����oN�(�/	v�OUa7�>'^�sc�U[���.�����j�����r�t�R;]��]ڿՖhjiA�p�(c35�l�>�ԛg�k��z�<,���mo�+E�9tov��ǇG��]�l��&�p�rr����Vq�QN=�k�8�R��`�,4�X?�Bc!����l��h�;<D�p�x6M+��%xf�~�Lu�)�2 �+p�1a��`����\��Re�6�����C	1�JҗrvN�Ҋ8�(l�,��|�gF�^���*_<�Ϊ�&�b:�T$���ߤ�ׄq��>�|�)�������6է4��An%�[��	-3"n��c\�^��Q�ˍ̐��s�H��\Jl��F,s��J��V����0�+�v �uqv&W�_�F|J�5��NoT�
�mK��%��������}t|�9˛e!f��լ�8�1��R���b�v9��S�K9<:���Wl��v�25iMϭ�`���33�~�|Hōe(y����]wke��} �W��77o��yRjb�<:�V��;Mo̫[$����AnE����+� x�������_�Z�����q�y�V�Կ�|:���s k��
""���gۭ�z�J�'' >��e��	��e��M������kn�H7Cߍ��͛7{�Я��h��å�/d�i4�1�&Y �'�wL�]���[����>�P�q$�<��L�B���/�a�|\XJ��L�}A�W�@6m�Ih��њ�_�����aw�9�.�R�2�"]�����~膱?mr�5Ɔ�Mi$|��.��6P���iu���:J�G��t,\/�0G���3Dl�x��6��v�t�]�i�6)N��Yp�L3�+c�0�v��)�ۓ����y̫���x��Z
	@np�훱�.��Zd�9|�����u���=mh��`�Kȿ=?��\,�"nc�{B��Փ�{M{-��m�����m���s��^��J��!%xE\5�kU(,B>W��pX��G��������"o<�!F�..���*�ǹ����DU�L�V��11n�h,�*M$���|f7��|&��lȎ�멼�>mm� �@<N��;�R�9��ܼl�C� ⁌:=-������B#��+p���J�@�J���Fs^}���t,�h����	 {Y���hD=�l��&?�Uj�x!P2t�(�jBI�59G�-� ��uX����N�7������?Lzm�di@�L�
��~��?Ƭ��'����m��)�S�$�K$��oc��z�0ڏ�7	t�E��T�.�� @�����f���$�-Q�Sn,h4�  ��IDAT��|�,�ʹ��p�ޛ��	�M.J�ZL�%Ʋ ����fi��J�`���I�԰�����N���1H\Q5}�@��
Y��-���6�Hŗ�pa�����Pf��N��P���ô!j ����])7����?8:�O߄�H���R�M�7;3�wҘ���@H?'��wp����״�~����t�ư� �&�z) l�"[��{�T�:y�vY��;Ӕ����z��a���k�%p�����}RH0¢ykܣ���W�vDI�WX��5��h�)t~��T;���_e�*|�������ұ2iH�5!���zco��%+ڏR���9X�T��q�JX�Zv�짵)Y[t
�ӊFt<���<[M��������:L�K�Q�����^?��p�q< 0�㩥�q�+Kca����p��ۯ�2R�X�q Lr����i�u����G�o�1��WaM׼��Q0�Jڠ�����D�%n[J�X�׆9z���0��Ã}�ĵ�$��d{�[B�9��L�@�DU�n��j�\*�@�4B	n-�1:�e�̧Y:G�:�����7O���/�o]�S��DΆV ��n�\f��o��$9�ͭF� �a�H��>��{g����Na���C���64�[I��S�E������H�/`��zhG�&h�]�z�{�y2غшi[EH�5X�c,��`b��9�W@W���c��GW�ʃB��_��l��I���uTܖ.w�R�'�:z����{4ZϾ;C$��-?�F���LRe�#��b���h�����|!��'�ԝ��Ǟl���Ͷ!���Q`dC��yC>7���j
JΕ�1�
I�����X��(w�����;9??M��:�{������g(���ѤvW[�+�˰���K���6&Y�re�DeF��A��P�$ý�\3́� \�٣��x~������ۗ��oe��Dv�5*0h*EI��`��{g=Va�P�٦Hk]��C��u�,��A$`���9�Wo��C2d_�����I��a�D���s�|=x�hM����ps)���Ҧ�Q��8�/D�����k�Xhj��B4�eQ����Ac��"����7C�Vv����d!�ux ����)X�ô]F����׹��|�>���^�hT��ߩ`.J�n[I�J����2?�����sr����kR3����SuFLF�*��;miƔ����D�C�mV~�ꭟ�F+�"S���SC 3��oI��j��E��Q6dB�������,����F������`	`�:�l�{O!#�(Art犈~η��|�}�������i'�ο��{�M�����{�aH�EE�d._N�������\^^ѡh�������Q4P
�e�]� a�Ru	��!���nb �<N����w��^ЖF�\����������^5�<E�Y�!ϑ����[��W����{K9��G����uk>���#�El�kM��0+B������� ��ѫ&ُ�Q���mr��iJ`x�#���Є;�8c�r�����$�s�^��9�v��yd5.�P�#`�N��M�`l� �):�$U�l;h2�q�/�F7q�<�Sk�K�6t.�I� 6��z�����T?�����\�0VA��1޿��X���S�8���~�[Q���H+'%hՏ�d��I�_W��ʇ�ۑx���<n՟�?eWbn�`���J3�0lr qMȽ�r>�&]�Q��T��(1=WKq�76 �<����F�N?�gZ�>TDUvv�_0��V'�B���fs��E) Q�ܽ�魚G��Dc�(�^S����7��w�\���:���-������wHy���:&��;��e�g���-.��"�Q�2�07>��Gӡ�N��8Zw5Fb�1�b��}�W�+r�ZT+��3�p@@XxkKuW�!�XC��3�e�ctTGbs\,�:�*MK�xB��� � <���z���΢�u�ڴʴ���%Fo,J-,O�`��;EJZm��q�1/�\2���� �g�����Y���P|=�5vq�(@����|~9���U-���:G!����M{-UG��9��ŷ&�^+O��N$x^7���aPaݠ�8]lI�����D	� ]�y���GyD*s�dQ�����xd� �`79{����v�im ۆ�% ��0
-�]�,�O���s������Ś]�2[�ϥ4/nl�±Aۦ�/���_~_#�9*}�_���Nkٰ�}/ ~lyK�܁!���k��ibV�&'k�i��EY�����}�v*��I��5��O�M#��3W�����o6[�)	������U�����t����|�ɶ>Z\����T�zt<2U/�q���`�nb�_FK�cH'Q/��HcB�J�Țq~�eSc�kπ��K>�F���c�j�W�YL8zw���؃q6y6j�˙�Hm5<�h=g� �&���K��p�s^Ԉke���7/���tS&�i2���<ۂ:��k�&�O�ϲ��Ԡg�88 ���˱O��wx��R3
�4�?_R0h:Bܒt��߱p��zq�I޿�^��������Dɫ�����>�ot�KNJ��ǻ��k��,�	����i$1hA ":q���
ӹh��{����ϟ>�M� ���'�{x@YTϪ��m�����1�K;	�__�Ia��w�3�afE�8�����AY[*be�Y%$�Z*�7��cL`�Av��o��d�R��㒆g9[jE�tMc���l�UB^����a� p� ��&w��J������U�]4p=�AI�(�"mЁ?#�\�Z���iW�-C�8}k}�;iCq?�)�P��6���g?�c���.�r���BI�ե�/{�m(�R���l���j�d#�ٴ6P)�M!�Kr��r���[�����=X��)ӎDu�xq�}�0�noy����\��QYG�p�V{�<z҇��5�&L?�����ݝ�-�8??���V�{�GyHl�1��'��q6����� y?N�yN Fčk 0��\5��UT��f��1x���x�Nu���z,1fl��1���.ڂˣHR9�R �4�r��1L�|/p��W��3S�s�"��i�5N����rp'lWםA}����ٜ��z��@[v�1����2�
t�����MZ��Nkb�����k�	Z��Z�vl61;D~�ڳ� y����{�F�<sS�g��Ojk�%�4��Y�I���d3;D1��T{�3^��?�ើ��, �R�{zYΆ`����GPn�d~
x�ߺ������B�|�b6�������I�(� ��A�ڍ����={���/FN9"�R�L���yWM�'Hވ\֡q��ӎͳ�����kˠ�<�]���g9��I.�|�go�{ ����� e���F-h0ݡ�np	�S�'ϥ,2�ʱM�=	x�}"ɽK�Ǥ�ռ��Ŕ-k T8\$냻�ɴs���>8Ysk��<7���ѻ��<�PF/�9���F,��4v߶�R�;�DC2 �_#Ճ������J�ÆE)p 
pFV|>�?tAl�3������f�^���Z��A����Z*H�"��>��qǔ��n���s�XY!�XLcz���G�ֹ�Pm�]���H}o�����Q/v���[�Qǻc����[��}���}�ȿ�1s�m|�o�1�u�����_�:A�Z��e�xjM[0�2�l��q|���ZrY��y���#�Ţ@8DN���ye�nިXź�����}�+^�`mWuـ�.����L�k����G�P�&��1�Nh����9�D{�֌��
#p��:B{���K�N� � �¸���t���O2��(���`4C��D�F+
�BK�"� �b�g9V��Z���jN�l�˞�{
�n�W:������j���V�t&Qō��ʬ= R��T^#�a�WF�6np��C9�}��R��#�+�A��I���+n���z�8�NP�M�f����m�2T���WU����5�U5J'D�j�\���wMi��L��+[���a��sR$�.�?�Fe^��_�3|������Ww@��0�a`���9��V�)�~�����kt��㨏�'Re���s��7�r���/~�˯�3��k��,9
��o5/ P����G�H�3/J(��RG�~����@��%#���ݵ\^����?P�mVf�8�k��!�8�pᤳ�E�Rk]�����h<ep�e����?_����W�ظ���"��6�fp����/_�r/�?�gE+�փ���f�YU�U�X��<bQ&{����>�����k�dċ��`��%�H���1ڀ���3GZ�0
a��eN����.��t�Ua{{��x����	�.��V�:DǮ�n�D�<H.�F�'2���Ann�3��>Ru��o��-�]^\�Z�ãD��*���Bd�3����L�S�<g��Wʋ�yf��\�:0�
��mKu���s��<�ݠ�m�~�M�"X��F-X]۸�`���)����%��FK� �0���n#�(���'�@T'��Qr�,%��$x:X+(��8�^�\I],Y؁����tӜ���_(��ϛ��F ���mM�"[�1�3��9�	\*)qN f�<�������\ruy���er0y��1��#� �Ohz$߳rQ�}�=���\���b�k�؞�?��Y�"�u�K�u���5����o������Wξs��S	�+K;�߰.�����d@uj�N�7���v�&�ݬ"d>�<��q[=��`F��H3��d:ם䔣  ��ҫ�3���J�%3ֱZ�F&sU��6���F�#av��0�a��BY�8�>f0�E<J���33�L��A�X;z�E���N��˞RFo���������������ҡ��v����3/���~�KHj����k����|�7$�1��X�v��*G5��Je���	�y9����Ԙ�[�C^_q/��n�ע;/�FI�ݚ�3��c�<Fy�U���ԉ���򁑯˳��%y�g���  ��z	x��`�TPW��2?Jz� �r.��[T��ȻȂ.����H)3�b�]m�Ug����A*�x��;�l����ne?�	�[-���D��U�Y��2��7^�ٔ{߲�A�� G`���M�N���zM�||�S]U,|�@�?R5� GF)noo�2m0���4~��7���������K��@��&�dl����rH�������d���Znot���ݻ4?>3B�{�6el���@�%	�"LMb�U�,�u�� �	�NҳJ�p�4��@>Ј:���ࠎ������_r���k'��Z��I�,��W�FH��6Eyd�UY�ʎ��yS�᳂ ���2�WZw�ZE lH`��y,1�p�@��}B�c��E��������W�$�~}��v��r��5:���R�P�L�-�T�~�&Z���4���*����I����eMЂ���v]��^� �4��ۏ��s�}#.�;�����b�� ��`z��A�ǵ���)�P���fw}�w�z��� ��{7�T����Jc Ȱ ū\�4(p�[�P��Q6?!5���6D��G�#��Gh1���7[5�X5�r`�4�z�whKw�O�K?���l�������̙*�������D6"I���^)���9�F�U�VJ�K�/�⠕�^�8)S��E��BH?�QR�~���RJ������}�)�aWD��z�VX_��o@�
����܈��t�?�ؖ��LGQ�|�u��ч7�ּ��B4�O���kkmղ��"5u���((�pP�|S,Κ����u�%��7W����{9G���Ҫ޶���@^}���U���~��5 d��r�Fr*#�*���q�9<pӗ�i��7z=� ZMM������:;�F��$l����E���\���^NO?'��Guh��{��}�����S�b��k��Qu�]R�����XġZT��A�&�<�]S��d�A�:���Ǒ<,~Gô	�x�EK���c��)b�����c����Z~���	��܃V�1�tA�?�/hq<�\�	��ɻ�?�I� `�$��������==���>��W��GvM�4� ���Z����������K�E(�LP�`�h�]�D��kn�8�y�Q8���S�Vy4#h�q����Q0DM�B����چ����\�i�����vX_O��|7��B�,,Z�j1�C��>��	� ��,�3�[:�������IO�l�h5��"�֣l!�����T�/.Ҽ�~4�Ua��:|K�+����.([�Э5Z�D�Q�!E�;� �	�OhM�uy��D~.�N5�HHkz=h#�[!��f�&�R��ȶ��h C�r��A��-�	�V�>{�Dє<��A���>�/�Ӥ`ws��a�L;����#_=��93
YfE#F��ʅ0��Å6mm�+ �s7���ϻ�-��"�W@���z�nc.���Am�G���'�����P).�����E���*Q��5h�H����ґRMpq�Mo1�נ6ծ��U�7sj��v��Z��k��(��N5����areuLE n�c=����i�0�E��Wo����a�x\���Ni�xO<(Q�� y�������ϛԧ����Xh:o�t]���d����U�ih8X�?l�8xn(���3����^P�@�����^�$ש�$�T@K7��LϸAH~.W��������.������D����ձ�l��)4��\���_S&�ߡ|6ͳ��^T��ܨ6nD���P�͘�SΡ:�y�[i���f7��~v�6�d�|�����I�C���������	�5J���%nL�h:tM9]�����g�*�sSK���E�_��������2��˗FipM��Z���y@�1=��>WB�sZ��4}��#�,7�e���Jk�'9zMRw`$�ѕ�y���H�'�%�
��G�8�#%�U�-��ks�NV�<@xB `���L焧�2�^�[yğ�{y�]�8�Z���u�p'B�9�G��̓����z�
(��BY�(1���(� ��Jc=ee�Z��/h��F�Cv5�b�{�:�����HǺ���8#��6���;�2�&�U*p!R�>� g G8TK�~9�mj�1}g"\g
 �5��b�#�}�b�k����l��I�6��4'oXCW�!ZŬ[c]Ц�V���"�3�Y�KrAͩ��^X�Uن,	*��s��H��J~ƈ�V��[&����h��i7U��Q��;����{$#�
uĨNu��c�QNկx�:���|;�wA����MH��C�kagO�s�
��,��{���X�a����~PE�<���F�}�c�/���J�L5j�(nz�(����rq/��s?���>Д*�P�8ss���L���q��&��5 Wm@�w�`dǍ���T��~�C7�8�ߞ����E�w�VV�ݛdC}�G�VfA��R^c~���%?��\�LgU�s���r�1V@�Ȟq�3�z0��=�o����/�a��������͕�k��ە�ׯ�_KEyMEՔ��i0r�G�B��Q�6��@���MΧ���&��WӘ����ǈ1������O(L�>���Z�9!��H�lQJ��O~��?�����͍2��o�9�Q@M7����ɏZ�yVc��5�b���Iϵ��U"� h0o��1mN������#�K���H��-��ӈ��\��ѯɏ�Rg"��ȷm��[ !�u�6H�F�'p��xG�Γ�^ DG�)E0���)ثb�b�P�WNb�L��w -�"����<����޷9����lI5O,��$�I�Q)s�?T�N��R=@3���'���Q�c��e�"��JF���r�0s/��rz�M�	���Z������t�T �퍁_�n<�q���#m�� �1��v� �Y`h�N��t�{�{���_�׿�6�\yO�9^L�߽{O��wქ>{v�h��@ܧ����e���Ks���IW���r�4Z�@��9I�-��2:8f�A�ihd��&�;��(=��ٙ�����S$SL`o!9A����ɅE�k�a7�:ӈT��3i���ݘ�5*G\�U?V�&^�����IP�2��|G��z��B�(�:=�$��k�@Ӷ��Te����~gv���Y'��_�ͺ��΃�����lɑn���Kߨ=mڵE�/s�����������`��t�ԩ�ޚ����^Wz��+��L�&�tY3-o�yO��s���]�}��&nD9���3\̺*��K`kE�#c�����ަ���B7�V#e�`m,C��z���Pun*�ŀ���Bh:Z
R���3<�4���V�H���Dշ����y��mF(���׏L5^�N�4ثd�V�X�^���^'�u(��7h���l��rS��Pn��{X�_�@�����dfWޭ�D`�{4e]4� ���U:� G�iS�M�~&{�;��Y&К���]}�O�n|5z����\k9�-�l%,E����#�:���-�Ǯ��t�=��� E��%7d�(�]�!Z2%L�Y��Mu~k����ն��@�gP5th�M4��?�[����U��_�����ki���'ֻN�B�,څk�+G ��^�*o��VM}�� �f��z�����CԠ�~o(�^3Y�����s��>d�ѣ$�{��W�Xے��oo�ɓ����V��^\�����9�+7	,a^�i���5�c��\_�0B��G��s�H�W}0��I&�������v:@
����ݣ��"�s��~y~Ţ����O ��M���կ�|������p�]ؘ����L>�48x�#�9�c�>,��*m� �ﾾK�y���q�m���ą���i����4x�����@�>l�����t`P|���{����ת������ĪRv�U��"��N��<����3��ʑ��|]���o!/�V<��c��>9��h<:�4�z��^1��6P;s�]���
&����R�ZA�/��Yr�~�f*0T�'.YS�@ا4��%d��M����wl�%��yl�&jԶ�(����9K�0�j@\����i<Έ�*��,�Ѵd��Տ8�{��~hե��!�PI\gq�y�zЇ��$����o�5�{j�1�"|k)��ʧWhဦ���)�et�
�25)B���` b��."s���c��O�կ����/�E3tAj�keO� �����V�F����ͱ�
ݩ[V�8���m���'��r�����`����9���;�m���_��W�-��H���<�q���GKļ�q,����}e��쐾��[�=����}p�%��֡gٷ�t$�/W�qs���;nj�mMϰ��zK Uw�H��u�|���C�ǒ"��D��deEd����H�hJ���~������L�u�0��_΍�z�y��hB�W�7�?��/is\�7��U�=XHt�
��B􊕤�ZJ�d?�_��k9>�c۩�ل�h��h��QY�>0�Ҵ�g��5�����*c���7�Ƙ��BU����fYe����p�Y6�c����lz��,oQ����(Y��u�����3a�X�"#��4�''G����LI���\{�ܝ����/)C��Q́y����I<�,�5F�@¼Y�o���6E��U��3��o��
���`�_����g�ַ3ͷ4o���F&�w�[f'TBbIҹ?��9A(&���A�Q
F�`�Ҝ���]z.֑"�g��	|% �Rg��-Y��;� QEt +Bk�ZFCp�6_R#2p��8�rh�̛������m
�WŠW��δ�uR�����I�|^s7G�σ����Q6?Yg�F�N�Vp�� @p@��'Hwԧ��RU�rUQi����YQ�
��x�ސ��G�&M��h˥���.l�c)P��w?|��|*o�>��vO4�T�ST�7̈́�v���V v(�>Rv���z/��R>1��A�����A�G��%�*^��]o��贏Z�	��oi"���:2trОh�H{7�L�-S��U.��#׆H79���1uܢ�m�[x��C�Z�6k`8��~6����P6c&守ML|go���7q�>_-on�o��v>��P�#D�>�9L��%5'�J�!�x����J���>�F	��O(5AΗϨ6d���C�y���|�^Ɵ�9� 5�,Q��z�ζ����C F�5X��߼a�`[��]x9���SF��S����u�,�e��RDJ��HSȄܯ��zC�^�/�nMg����Pߘ@$ˮ�33�-�n �N��6�������.���p�D}=3;����wp ������W�e�ѯ�"�6zVM#l2р��w<��:�(����!�űmTr�<��E: ���c��O����R��lL��u���t�F/t�^���{�ߪ)��$����{�VO�v��N�@�#;�����_q����1P�j�j�{-�o{��ｍ?��QI��X���A�j��YS+�Hm^�_��l�#t�@b6�{oi��E�Ru8!_���g�_d;�c�g�t4����b���/�0������TS�!���F��)�%x�Qu��>k����`/���ڽ�VO�i��߭���v��\���s�s1�����kU`n�߳����g�n��c>e�8��#��z���#K/��~`��o,m%г��{����hε��ͥ��'�NZ3QBs��X���� �c.[]N�e\�c�XСi#H�|٣�\*����a�ނ:�%�C�ث1)5I��ϗj-��?� �U�� ��^۾����j�,>�}�� �FsH�sH�A;d��4�`ϧj�C��$*�n�w��2���ټV�RM��[�imr�4�?�N9\U'vbr�X��;�R���|b5�U���	���-������ɺ87ԗ���|��d�@.};ݱsh��	�z���h=�-M��v���oo.�iǛ�dT�輕Û��	��p���ϱ'?6�����l��?��r:6Y��ydm~�2����*.\�w�����\�O?�"i��N��R���`'R�>2D2��7+��K��f���z�=-�Az��0U���1�v^���$���l�D�փ�Q��0lں���.�m��ٓ���oi;�|���P�~D��=6���T���v�����+�̋����������=�T`#$>m�`�EE%�C�#Y�P���������.��-6�)�`�d�mlr	�g�����~�o?�a������جq<8�c[��zIF���M؞((����Y`��BJ} �l}���}�N&1�-��p���1"=k:�*a��[�c
�`��ܧ�|��T����-��i�=29���	������զ�����[s:�tZinO�I��,z�?��!;h�&��������4�ޘ]�9�]��Z�0�9�{�8������v�K�m�q�@�16"�v�`~�8��sE�S�/�0D竞K0#̶��Lfs9::&``J��@72������pf��^�Ԣڴ6fC��m�� _��M�K��v �k5(ZBD����rp�G��Ez|)�g�5�V�`W�3� C���ES]ױ�w?!REx�G^?�����e��֪l�����,ޔ�3�y.�5���!X�'��>9�i��l�VR��*`���Vz�1��6�ь��hF 4�f��-^11�r3�Q3`��T���	)W�t�HE"L���R"L~�bȣ�c�P��	T���֒�1ڒE+��@S�r课o�F��;G�j�v�*L��C�d �V���<#�	�/ld�9�K~��0m�{E�*�E4w����wϓ�K���lV?nUB����J��E��-��E�쮞đ�===�.���)7�Y2�Z=�V��8^�S}溪{#�rcY1/QO�S�nȇc�=I�=�n��KC�!M�,Tב��:�hO���Ui�}���r�������- �2��<-X̕{e��vf����wҼ�fJ����E
����F�֚Ηaz�L0�����k�2RB��5Z�=��{u��p���3�� ߌ'V� ��#��G��fzh󽵼L��ͮ)�T�E��-m���N�
h���Gz�Á��2��Lx��`YϤ�z�z�7� #��ER�o׺ƙ4������ �#+��>�^|�")=Z���&[���HA�nL�L�G�v��CZ ��M�$�_�9�b�fDJu��X�>�����ھ��a��mz�_���|�8  ���9��25'�2�2સ_�;ݮ���_Ρ��S������s�b,�qf�j��!D��KD���"	M���dke��u`��MI��=���]ʎ`c}c��ҝ�u�"�n��wH����7�����v��H-��b��*��]�J�`��x|#�{;:Vc��Z0=���F�"�:����5i��tDk6ʰO��>/��:,8 ��L��[$�kx���wn�m���|	���
є�Aj4 03�3^p8��[�����'i���ǀ�I�o(2�P�L��7�p0A-YM���%0��n�8�ix�J��V,��=����ap��@����O����V� i�����`i߲Pl��3�|��/<�|��}�ۻ���z|u"��:(��B�6�ya�v�?�
���_O�禷6~M]?w?6~M׌{������8]�1{С�ކ����C��z���a_���hDo�>�5���UpT�a~�" ��8��T����-����U��=�?��@'i��B�mrqw��dO�w�^m�2^82i�wH�`׵&��g;	��7���mٚw�ѠQ0b�[��W&6���#R�4�S��g��ގM �|j�M;-P@!�t��4b�ɡt��gss�T l3:�#2����ɔg>X�۟3��8��f���]�޺���t�dM(����P���s��Nl�u�hsT@���*+c{���V;�s�UU�LvT�
�M(��7��/l]��z�H'{��fM���%6��SL�[��R���c�S�Ϡr�|U��� �9�AS�l:�'�����j����)(�oC�c6c7�Uq�}h��=�\��R��߈Hhz�4�Cd�5
IE���b�e��g��3��/�0#�mac�we/��������'�`�����;���c��-�E�J��ƺ��(l���)�L;��O8�ا�o����㷴i�����Spl�$t���:�XU�&)�4X���xn��s�YhBՇu�,��Qg�p�G�)\TT��H�G��k�0X�MGD��eS��Ф��1ET�[�(2@�?]$���t�+f�|Ev�l�zr�  X� �M���9T�}�'!/ZR� b`�Y��b�&(uO�o��C�dӬ[b�"χʐ�K��x J����i�#��Q����@ ���₨���3��"J�@�#`�Y����N�����A�"�"�P����'�����1��NX�F�F/��ʯ����C�ӄP=�?�8�����ya���1C�F��S���}�����߽���3�M���^�$��G�ޱ�Ft���������/F�/�����ͼ�F��u��F���[:����	���0[6�ޡ�����+ݰ)�ȯQ��#�PО~mc��P������i�RPNB^�QAM�HG���h���V3�IV{���4�	�z:So�����3?c����/�Չ��(�.ӴX����M�X���z�<�\�W��5�A��-�2���q��ê��A�jk�ւ��$Zm��ZNm�9xe�V��}��Z����[˨w�V�H�T��D��|�M��U�N_��X"�2M��d�Lo��� �s��{�f���Ls�\���O�[F����+���
�B=Hs+0���}'׽��Z_�VI���6s�WUY��ㅗ�;`X>���Ǝ& v�y�PќNv`���D�cr>g�]T0o�)v2����J(�ų���X��U��%ߕّ�,�~���"�N�$�@ur�/�i'Zq�B�1�W�s[M����=G��JŶ�v41�M2��F���%.M��GM��(��ך�����ô�!�E&�Q�.Fz�(/��"��h��<j5���X�/��Z3�� 	He�_��x5�7������7�YȘ=	��ƞ�x[	���$4pf	��1�
�۲G�E��!Q������[9,�8;���0(@����ō����V����C�|��7_͙F��!kkA)#���6`P'e!��|��\������~�_�!Q��x�z�3�w�.����ke�/}��)��G� �n��E��6�k�`�Q���W_q�~���dg���o��`kۃ`��nr���O�t��!W�S�g�y�p5�6�y0�3-�	���2� �.�6J�1��4Pɉ��,]��������b�|��]КMF���a��Kt@�NƲ��z��;�k�6�`����od*��sD���{DE��Ž<˹JF�X3sO_>�j|:�O�>�fs$���Ǟ9v�Sq����%�U}�;3�&'�oh�ڊ-�)�����l�-F�<j��l@w��n�O�0(c�^.y:�#��p�3������q�(X��"=�$���� |mM��ԤӪ]-���]�M�3,��U��@}:q�R�V�6��';�
J\3^�Z�J7/�Y4���e��l�A?�����`Oi�4��qaWg/��[Y��s�U ��^V�b���F�st���/�O~�Ν�������2U�2�^	vmTG���S"��ftK@��G>��r{O��:�%&��B�K�������j��L�up;b�R'i]�:����C������O2{�ڤAҊ��0"�(��~�� "yw�����bw
�V�':�g���,ZZ����k>=c��X��cjBޢ�?����۔�#x�r��m\K���C�zx˴Ṱ�P�04��X/1��F��p�V>
ȿ���{me�UJa����×&�[N�iu�
���G��z�P56�"a>�^���aE������?�q�(m.l�|w/?��$����é<<��Yz9nr7�y����A���Z$���y�KV&\��c�ek�����V�"� ��s{���]2{�>h��}�?��zdz�my�uZ�vu��1a��3;::b�b�H"D~~v.�ݣ4.���қ���'gf�R�s��b�ʍ(��~~K�r陖S��
	"]��*�COi���
�ʜ�œ �ø���1��luis��Tt���I��ND{"�mm�������c����(��	�� 	��QJ���>��c�5Ut���_���-���Tȷ4���OU��	9��D�uY�/l\?�ȑ���Y��rdJ�dx�]��">Y&���⛣�UoK#��0�� �X-	�����q���p2&�FLEJ����w6���#�Jn��EN�?7�r�W������#�h]�!+ˋ�<݉��E)�����j	��_Y�J�@�=3KT`G�"�T�`�6ΕW"�k�	�&J��6@t������`v��T���3��n�UE[�ϳ�&)��K�
�c���431�E6>��j������#���������坦��oo�k��%'�#���P�t�[�aݧ�s$��ߤ!H: �cU�gH�ݢ�>|�<��٥Y<L��b���`jOwQN5+�Qոr�:��:�X��D�Ggu^��	��o;l��AqjC����$��ӱ9.�R=�d�p�w���)��&G�CI��iXsC��m�96��A�NNg��(�:��i�x�OPa�:(/�|-�=97ð�E���8*�(�T͛��k��x3ڊKa��VD��\��ޥj*u4h��-xV�q��_�o~�;���� >�������zӫQcX @��.��z�{IJ������^�K��%��P����kyu��t�Ts'|F���lp�\�wk��ss!n���Vl>���͏�fXc��K3>��LQrO?���Xt|�o��V�$���'D(�O����>������}���W|ᕘ=#O봱4�� I�=7�ζ���<���+��iYS�뢱qPw�{�Q���~AO���!�MiPz� @󿔡�F���)���-��m��..��ǫ�Y��
��i. "�Mb�����6�:��?K��l���V��њ4�̩ZY����<���)Ą�Jץ�7�7��oZ7�G����Ҫ��ɟ���k�k����Bn�4����.�$В�f�Fv�@�3'4dV�%� �b:U�K�$���a��~uq	��/-bP�i ��"�AM0^";xvF�<�=ҳ���ݥ���Mx.���n�;u����B�5�8Ɉ臞���T5*/��=[MbqÄ�e�RD��Ŧ��u֔S�|Pe���'�&��ޑ��9�@A����"DT0���t��9�"��)�9�6�ky_Mk��y�	�W���!�I��k��6�� O�l���������[���؜
���Xt-J���3�e�z�Ec ��1( �-�f��YI�g��/���<}����٥�����|���l�xߜs��Z�8�^��nÖ���4��U�z���vk�ݟ��8���d����։&��ch��W�;W����n�#Ah�He��K{^���Ń饄�1�(ߠ�
�v�^��y�X��W�d�5tL��hQ$�({F~4�VH���������R7]��!;?X_�>�Fx��oY�}�.+��j���"��ѿ���������"Ip�h���ڱ�䜘ڰ�!�`��T���^_1
 5��������r�r:�{���`��0�~���c�z
�6#_/q�<E�c��Wv����
Tc-�d��F,2�0/�����p� ��4���utY�w���WF3���b�ʸ^��PgFD@DK�=�'�����ե|B3�V5jD��>�ֶ�u�����4i��{��[(�/Lv�����L�sM��t�B��h�����,�y��$ �j	���Ed�:^���'X�������ImZ�M��hO��m�y��I���k��>�#]ߗ2K���an�#��x������=�P������WΪ��b�%
F��(8���"�,�J;�@�-%�c��{  �Y3t]���C�)��EO�M1�0�=�q��6Zv2�(`�3���d� 64Z'���w�~�`�Z*b{o�⑱,Ni�Hh�����F���[Q�4PRXm�~EOS�M�|�@�Xa<��	v����1�odiܼ�Q��QF��µ���i;��ټ�H\qݐՓף�qs��㳿������S4���S	��������=yؾO������-d>_1��JW�����M�\y�����P�v2< �+p%W�����2H=&;�6����F��?D?PR�����+p(;�H���ݩ�VLC��A qn[|������",MŚ�]��n�e���)�A�A @�H|=�;x"3��.$x�0�C҃��d>��o)9ꪬ�&��~J�ae���U���_��)�
IGF_H�DC`D}�����X(	Tw��Ua(��nM���"�Tx�P�M)\��ɿ��o�7��A�����`*׆�S��!�����±���|E9��щdT1��Eda���q̶wD`�;�-��������~i�^6�g�*��?y_��X
i�̓e�m=<<b��i�t��ig;��ZCu�B�-Nq�D7�f����J|ª�	\���"9өj���* ��������{���0�X��!"Mʹ�J{�yD��Uj���h�����U����+]�h����w?����"��h/�I�`�55�:|0P�GGLۣ��ָ0xmk����ܸ^��w�v��k��v�k�T��1��+�,�߳��ד�i��|B�cy֙��E7ia��6y�0�o(�T�n���5�d�� �.�Qm�4�F�ڼ|Q`ww/��k9�@ �"7�[c@`0�r��_]]SU\X��oQ]����T���=�" ���Z�GӨ�Q���D�d���@��:�#Ae�B��|v��w�+��d�&��\���E���{�y���UTd"���9Ȉ@_Zv���\Cd��m��qе�S�M޵�[��6f�(nB4A[մc�oFMK1�v7��ۖ�����ʁ����O���������}`���Qoui?��ٗ��#���7��y��!�:�y��C��	m��YD-�P}��b�&h������{>P���ŕ�%�۴��I���^���߲J~gwN� �M8�9��՟� ��QZ���`Lx�pt���$I��+��i,���S�[�i�YaB�|Ӌ�jS[�؞g�S�{�����߽c�������F��\_ʂ��5�`P��0���֬�q!�`%��M��/s��zo�ڰ<�J��plp/Fɔ����+�U�U��Ս�vE�p�1�AW�\<Ԥon������iP>%CwOÄ4&��_ ޺2��o6��=�ͻ@�m���=�_�#��l�Cc>�fp��s�qb�O��U���g9]?�����M9o~��jBrM�Ə�R#i��H��W	A�6��|�P��R����g���5��+T��0�}߻����./o�����r�6��d�P�C�`����OԊ�Ϊ˴x0Ϩ��R�=�Djm����$da*�c��;p͌w�h�e�yؚ�d���Ή�i>I`�h�Ql��W��,	�eʫ$���қһ��
��!Z�<�jJd)WeF�^�9ǩɜ@���׀���Nu�4ˀQ*o]�3�S�`2f��)�sB��V�K��-Ϗ��5���-m���(�988����_͞�;�s�M�����Y�6�nM���u�B�Ix�H���9��%�Q��*��w<��%�s|r��ζ� �ϭq�h���bI��t	T>���BS����㽬�~�x/g�m����/����[����F���q�����<����6��>�ֵ�c�6��Ȣ��r"x��P�����)�)����\�K,�s�����_b	��~�hֽ+���4�fr��(ٵU�����\�+�*Zģjk�хE�b)"�LN�4(%��uح�o=,s�.�TD�Au� ���lªIr�8�
m�Y����s�+VR`��N�	���ʹ�Ql2���f�3�k�6�β�w� }��M�6b��}H?!���6����>���6��j����$�p|t,���L�m��Q傁��3��k��>��rk�h[)j���ȯ[�`�#����HY��"�ؕ�ɨ��VC�ʴ��.V���g����H�=�ĠIih�ڙ��w��`s���}�F��E	�襬���"^\i��!�'0��{�p�m@^0�-�0R�t�oje��xEj��?mI�\sQ�l�=|S�b��x)�����يv|�^�.�n���}G]���
>Y�����|tU�5�MW�M�:(4�h�9}k�#�+|��fΝ\^\�?\8�IZ�f�j���(�
�޹ՠE*��`�ڐWuOnX��D-�˵f���ո���ʢg��7��6��e������3"���ZS�j� 9z�~2]������7��#U�M�����zH�E{���N����1�69��\jA�~�؉2i��و7��s������WF����-�A(�M�-�L����`���8���o~C�+���7x���� A�z �T`߿�w���2٪��=�J���gM�5���͛W��W����ɛW�C�T����|��Q�����d��N�������W"��UҲWC�� �d�->�%�t�#�L��>؝��o��o��[ve���L�����+���x�]hi��DP�W�/m�֣x�W� N
��7;[�༗����6�XA��Z�-G+3�p´
b��'�K�Q�+��Ge3B=W��眹jۘW�G}F����s��C,(t�a�@�� ��h�C�~�2w��,����Qm<�toُ����OA�>��Ê��� :@8���s��91�in��*������˩�� ]B���x��Ǜ7�Ӝܑ	x��%�E_����V��2G�
���*�ԋ�)��#j�����i���Z��N�kU9��ziɾ�k� ����r>vחi!\��F�Hp�fh�LH�]K����ⲍ��-#�Y�q��# �V	X��#N9��{uO��
�j�dȓ�6�*�K	L�~��_�k~>���}����{����Q����C�=�&�ps-��:�&y��bb���칗��}�.�!����8�]4LF���l�D�[b����g��c&��)�:��H�|�#�H�s� ڈ����~�$"���[�r�(aX�`���wc|�er�56"����₥Ö�yXh�xDM���(]��2n���|Y����ж��B5s*yE�Z?���Z��[@(�_'����<��m]�\��%?+�G����)1H 0-�+1|e
�MYS�H��mg�X����%ݧ��%�OY���Ab=���`	b޺^D�5�Q0}�W���ߍ�a֤�M�Uj�b>��s#(�Źca�=���O�9>�H�
�6�	 ��7�ț�o��i�+��v�f�5�����GeQ��aKs��I�s�;D��e�{��x�^QA���c�88y D �g�������hP���[��W���5{�e�"ͱ]F��vE�	>M繟���O�v��F�V���"���3����L��$����%��5�0�VX��d
���Ǡ�<|#tGױ�V晫��`���ך��[Y��1+�R6��h������g��_�qM���4�8�M��<|�kA8�~$x��S�a�9]�M�ǃ ₻M��Y�&�(�ժ%�@d(��Q����`�l]V�MP�V�Q8���#2������' ���˫����4]Ǵ��F��%sr�@4 &Y�@r˱h\mQ���ޮ��01�.�Aw�G��x J�O��т�����-i�j��z�Hq1U���t��)K�Ռ����,Ň	P6���猷4X��C�9�LR�Ps: �j?'��J��G���k5��HB���}:=���+����/�������R�b)!|-g�Ï�fpk&���I���*닥`��<^I��\�m���k�8B� L6��w��E�X5��lL�x�� ���G��QS�M!���4�/8�u;l� ��p NA�����NM���;?g���c��ńYUfl���b��>i���wiL��Q�㜞�Bn�_��@��&�Rh�Ԣ��ʟJ��*�J�9����X.��@Z@�vN�ݞ�����N����.AX�*�"�y�׵5��N��?� ��	$)!�B���)>�v$w�0iO@�N!��z�Nc^4��e:'jف3�&����Q�f]�J�pv$G�t~(Aڍ��0w�����
����V�s�'&yp]'^�Ɠ��r�T�c�(�@Q�5e7������a�*�u�_�祥�����&f_ lv�[���.���_P(�31hoND&�M���i�W<�^K̺�>;� ��_�ӈr�$7lW�e�����F�@��	O�n:��y`:�����\�}Iϳ��<H��B�t:F� ���vi}�ɑ�uu��&�X6�&�n�QK���u�ɪ�3��醿V�Z��߫&A�~|�p���x�^��_���S4YʯE��P��r�)�M����91-��R�{O�K� ��ҝVy�����I�s�^f4	+ p鳮]'�+��xHN P�l��:U^9�L�a[$�6ܡZ�BN�.������&N���g����t�A�e;'-��O�$-����/z4I�4�/P�L:�P���ƺv�<b1ϷƜd;���
q��D6�z�V�����<���Z�&@ȍHU��M���MOqp�00F�L��|>E��H�_[�Z\��ڷ��y	�tW��hm3zy\�H�����ϧ�ÇO	|]�P(
��9�� "��4Y��m�h#۴Y����	e��lxg��MrҨF��Le=��s� �no+��:������u��|�ά�̦�_�xn��|D�FM�H��9�V��X�w���vI�E���5kJK)��iv�l&F�Q�R�ȖE�F��f��!��N�׶εu�ݯ���L(x@D�a{�����eh���o
���6�hh岆�K_�f��������4��bD���T����#yu|Ȓ�I��f�6�=DŶ����__�=�{Ͼ|���f\�珹6�+_&�g	�`@�6�A�Z�ח9��۸`�f����Y ����$��V�G$��lө�W��Gy������v^�H�����3_q�\'n����S#���X>I�QG��������0� L�Y�gӉ	�*��{ў'{�7a��E؁��<�\��y6��C�E��<(����\]_�zrb�>��o�za���~ݦ���M5��`�|�S��	%uVv'Gi����~��i�n�Ö�%��5��H���l`�ZD�;?4��<?bw�hk�NT
�Z���m����5���Q��3��J����apsH��v�zN�/�0���AS�W�XM��}�s� �}K�$�2�������OhJ��0(X�t�X� �g(,ːhFL�V�8Q�է�!�X���#S�HhN�^t��*R�2�;F ���65{�m@��E�쓚���7g����h'���jHo$����I��$8��Q	T��%�Y.�'4��5!�\���Y�_&�j��T9I�q$h��x!�9��6��,�`zu֠x��~G� ��?Ҡ�/Tb`ݥN�z�������'���\�\���K�Sӆ������LH�Z�D֍�F�N#�]�2��[S�(>!�(�aȆ)�����,�/���r�-n~��ʛ'njS9�e��^恸^��������v������ǭ��<1����|��*��Ť������|�
̍Fb��Z�y���bɨ*�N��X�;�����B޿�6��8�\8k��7̿��ñƨ/~�M��᫻t��@�ف|�4ӷ_˯�yK"��ř����x�&{��D�z��i/ș ���`WN����}�����4u�>g	V
�H�;;��m+���n����@9!�פ��b�lQ��y�e�B���0X`�8+�g�r�4-� ���;���L9tdQ�3��3��b�-d��g�Q���z��������.�����sY	���0=e�k{k.}����\�hn��������'���a��=/� �шtLD���nX� ���hQ����WuA�V���C.�ױ�	� ���}�M�K�	�O 5��[��n��'r���хn!"T8绛k���#5�X��} j�PϿ����"�ɞ��J�uwJ 	�9D���̶ b+F�ǭ�	�G5��4��/����0!so�=��w��*�Y�A���l�����ص���!?=����6��l���{�TTc��:����|��%ZD0���(����<��������e�_���^�l����x�#��K�� ���Yz�`۲JBv�,��m�5�1E��'.S�?M�.�+��A��w�NT��F����z��
yE�!Ʈ����	�r�5jk?[-��9D�pj�� `&���@e8 $b��a�'�߽�k-��_}�>h���a�ĖꅭՓ�V��Π>�NȐ�L�d��Py�^j?`jc�f�4�4��F+`G��A�3!'p�ԍ <�{�h������0� 1 ݋�@І�Q	ɮ�S�B砗O�j�kpW�id�Խ���H�%h���wDfV��=+]���1���##�"�U�g�~_��`k頻��N���̪�A��I0ء��z
+�J�.��l<JD�eن�R`�E�A���K ��*x2������ &�>�:
�u���jP^�0#��f�0�$�[SP�8qš�_u=x�M�˴��W�'[�b;q�j� �~���J۰R�<�h�,��������,��y�p��oW*�������i���]�ʨ��؇*��iLO�w�����ﾎ@�dˡ|��E���e�˛��"��qӨ]�Da�ۈǼ�8c��--�G�th'�����J�Y�nF^,}�I��؛M[U�s����$�X!o�<J�0�0��h�+ܙNC�;q`t*mj�Qzx�٩���ק���ηd�:(#��iZѼl�XX:gw���H��a��k2�gX��Z�T�;j�"F��~zr�~�ղr�Y��=�Y�V2cX+0�6¬a,����Ժ�N�Г���%�p˲3��s���J&H���c	�N��E��$��2X�{��3�h��$,�T��,J]�\��������BBI�V�m��$��ZK��x�,
�ʗ�ߙP��-�,#/��J{��ޅBT��;�Ng}(?�p:���Ϡ��Wa���aͪt?�Ƀ8�|�|2��H�rgV�X����&��W��ĵW<�e����~ǉ;�
�R3T]���"�{�� ް�0��5.[]���nnM~S��}��}=)(�Ͳ�f!�\��~v�%~�Zß�8Q
k�K
f%S���p"Ta��(�� ��0�_͇��lʒ/X�<,(0��hX8���E��w���k�~A@y��I
���)p�j�f9	Eƕ���N���+0�v�R�� 1�5���v��ų#���m�3��H�k�|��J��6�,8yf	h�Iq1eC�.ⴖl���}K�}�9�p��r������)��o~���eK{�K|�Ĺ8-}"5�<�WB]^��Q$�]�V�����j���H�hjZ������7�c������=y|7���ߋsf��������^����p�����N������/���wv��WUV
�1�ο����?�_����ޞ2(����=}�'����`?���z�[� YD���'��"x;9=�`o�^aQ�x�U0�P��cR��kj@�� s�S%B�sL�V�`}�i��Ȩ2
U�(	d��aN���6ႅg���3'VuX��[jѼU%�!��
��{[R�3�U�%��VK�@S�e��E$V�[e�7M��X"����Q����=�o1 X]��72��l4�%	�0���Mk�Ɩ�*I����ɝ`�<y�~A����+>�s6��.l� �,�qMR�ͽ��"�G���q�q��.at	i�F�Q�IJ��Pp � .�i|-����X�J͘kI����Bad�u	��������D��-}n
z��1��>˒a�c�m��*K��1a�~�?�HM���栖)S�n?�❖q�ʓ��J�m��.)d���F�Z��i⌆<��5K�)$�P�������Yo����3&��S��D���(��[��7�2wV
�&�xu�%?�^�7Ӹ�ڧ�fV�I��gY��B䮚�y-�`%���֠@��mZ�V˨?>�B�V  ��|ş4)�%4
.�>�����<�s��K`#C���4M����+)��& 8���Ɵ.ܮ��3���:���_i���.5�BZ̪{�p��6o�I�:{��qN�QӉ�9�����X���*8��
^�A���#$�O[�Z�;�.Ċ�����Ԛ�Ak-`�u��u6�� ���
��ieBJ��33���]��~9��vIK�y^�M�}D� �]���MԶ|�����W���̶��޹��tIy�]��R�?�3�"���������g��N�}����qͶlo�I�p$](&�J���L1?9[I���K,DF�<�Pid�sZ��J��wt�� T �BVH��69��H0W-�w>Y��rP��u�lT�*u�Qp�Z��,;��	�DnBq�����*Ȅ��J��)��^op���`|%X]�7�t�z?�,qo����[��X�X��"dذvM�w�J~���ďD��N�X)8�_c��^ijV�s���c�èP`������,����$/U�X*�[`#�1ԯM��T6�e|o*1�tv�ć,�JW�CH}-��r�T�0yoځd˧��;w�g9hwD�lЃ,�O9�i� L���,2��}�kk���wo'��ȴ}}`,+(�0)�݉8Oe���xp�,Cl�5�ܯ��$��ߵYe0�ij�%v6hB�}�Żx��f�I�I�6�<GK��C�0����|����r]��vdO�P��b�2�ҫXVu��}�D3����*^u������K�sK�"0k��i��������N�l�� }�Įm ��WZXb9	k�c���O7O<?�7o��A|�r��H�/��gSG�1ގ�d���L��i�0�PnN���J�Q(,d�{!h�PǍYu���*��s����b�X�^�ַ� f��>&��x�Y��>K�K)��g�tb.Bf��fdE>|���)��2�?�p;bl|�V��ٙ��	�M�;S����n���X�d��s�C\؄�+c��3�f�R��ڵ=Af�X�T�6��kݐ�h����:܃5��:x(لk`��7a���آ @������#� `H؟�ENמRN�u�( ���aQ�bcC�Jx�$��:�Fu@	�@2kH|�uZɊ��i�p�v+	@��hR���9��@�8�f�I�!b� �H�c�Yǈ_:�p�泙D�' ��������dyG0���|ā{vvFVz�AW��| ��w�(3F��2lE����H���
�t�s�nP�Pc
	XΞ?{�?Fy����ymp	�bm�rV}ԖM��\W�D�]�z�Z�<C��"C�"@4sHn� ���Sƃ]D��V_ ����� K9��6&���Qv�Zr�¢S�4c���>+��]\�5װq
�	�qϥ�J���u#�j@�l캤-�)Y1�
�� ��@(��pmV�,�{�����ɤ'ٰS[U�JˑO�&ʛ��4&N�������\�7��(��B�
Q��"�o+Z�;�B(�r�e��+�2�X�]�0OVR
E1�,N��^GP�{sOf|Ǥ�L&��"�Bv�r7�B�A�?@�S\(���;._���%����1*�G ��%�j[)iq��$���okZb:t��UC� W�?��cy`3J��"g�^ X�N�5
�Iy��/&W����F!�o&��	���4�\�;�C]�)�b��º�"�c�����е�~J�링���5U��Y/T��YG��J�z��' ��ﶽ�Ŧ'�3��*
�E���.�0kYd��o��r/��u���Ȼ����ѣ=j��;�pM��O�*�Ui�x?���ۉn/yV��RN<]�ԢqTZ;�ې�~{����$��B��0[ְi�BB[yW%RZ�u֢� x��V��U���\YIiY�pA���n]F���C�J�����ҒBf3H�9��-AZ��:�5̈́(����ѱ;��ӓS�2n ��!�Yg��6�%�4i�4Oz��z���{_�� ���������N^����wwo���q�|�e����q~�r#!?�V�mĽ�}
��߹��Kj̤�I<��^��Ab���0��q���B��p�f�:u	�ʻ�b�B7tی{a�	�i� ����n�[��k���Ҁ+�:X6N9�J�d����r��-VwJ�(�o�����cx� k�D��֥�����y|LH�+�m?�HSا�*�M��@��b�M��ˁI�P6p��B����F�C�E-a���<�{]�$�+������J~Z(�:��2[;�&��
!*o38_����kU����0�$�	 �F_��H���Sz#F�+H�)f
�00s��hD���-�x��b���|\L�ҷq�n�F�X���*��@�4&Rg� f�f�H.�dQҁ-�V�ʳ2 3�yZ���]�b�^�`jeBn4�Y7J�>�H:(Da��VH ���L����6��2��!�?iZ��s�`�EqM�I����86[�~��g�ؤ�ɨ����af�Ė�F���S��̮n1w��C0���\~ba!O���N��R*.)��,n�F:�����b���!7OR/���ֈ�V��x9��!�2N�Z�%��k/~6S)e���,
�>�1 ��mʓ��n�ur*x;j�h���H����T�8��.7��D��4�ċC�����l]G vvz�NOOX�}�5���i
\t{�n��+2���'Ɣ�ȽF�g���N(ndp��_�_����[w��Hx��f-B���j����~xD����G������i=.ܟ�����oH���Ŷ��
n⪫�ǎ����a�|�⥖�h��G|�ԝ�����@oN+,X���2��c'��AS�>��Z��Z�-(j?������8��}�H�ȾKP~/VP�S|e��|V�t$3!P��lSX(0��{����(0�h���_���1h0 �YZF�FN�����7�rL���C�/E��ф�A}�;�����C�'�����>���֜ϗ݃=�k���� Q���f�ZY|���(�D�^K5b-1��1<��P�t5���6d4e���T��׽��BI(��~c}�\f-�.3�Wʘ���) teV�[�N�H+�]W��㿈?�(S��a��crQK��纫`�,��^|�nl{��_	�[(y���/"�YP��R@���2雺��� \9���`�6�E��%�UBzq��o�%s��#uc5���~�q-e�J3-4c��T�R"��3~m�-���ɢ�em�<����� ������y���p�ֳK�?���#m�x���;�����-�e;�A�tq�"�`�f�.�ȍ(2h�Q���۹���� �o���Ӯ�V\WR�Ä�ȾxY��Q��Ab��6�R,4���$&���A��m�v}E+D�6�����x��1�!��́*�q*{�1H3n,����A<H�"-ͣV�D��(�@���y^'�wC���9]M�9�z5�.���&�(sG��Cr��>��h2�^�-W���Œu����������w߻��c��B����%��Q�E��7p�	�k�Kl�P���$Ŷ��ZѤNk5��F#�,��G���Z[�W�+;������Y��'��&t��U�xt�?y��>z���S��kק�J���6���J����pk>~�D@p<��v}ǹ����}��Z	����q��/��w+w�<���E�%dnF���5\� L(�v�e�HZ�XQ�+�6d3��,��i}���+�k�Wm&���_˞-@�F��??*R�����Os�����m�D��}6�9m\O+��L�z�.�9���AI��! �8Z��MA��2eHv3g{X�ˠ�Qf"r��@h'�Nb���g����D��^�J]��'�M �*6���Q�	��eP,�A�~���Ҷ�A
:a�	t�1B�9�f)����[r !	-�}�e*���4vx��f����eS2�բ��M/ue�ڰ��Pm����;��^2*�j�� �Z/<L!d����v����x�kJ�+f�]
�]}�Yu��H����.E�l�w~�Qm��ez�ƻ$��ۑ���^��u�M��RHK���څ7��R }��*�0�������p_�˄xd!b�u$�]�+�\L�׼���T�j��A ��i|�sy}CІ�'�#q�Ȝ��׌ �&�� �<�#)�����G�xsv7�+w7�G�����W����	�-�����u�f��&|ta�fpw9?��8��QM6���J#n�7�3wrrL�+�0XN�>D���`�j/�+�Z���l�m��w�y��a}��N�iHj��i�K����ڸ��{�'c{,v?so߼u�F v�28
�=6}Z�i�B��kZ�P��c�:�E8"`P+j���_@tmJ��Kݨ�d<��*='�x�_��+wxx�/���0���nV콃����m�֡���K,��ZJ9Uj2�_��	ٔ����+ܡ ��vB	�Vq,�Lt �������}��ߘ��qÿ����r���˴�V�۸v⼸��u痳8��2~P���a�D�[��x>Z�Z��*�=7^д����^��=�'+����{A�<ÿm��3ܬ83)�a�����0���v����Wt�ɀ�t��$���}!�����ܹ!���83�EJ��Ī�H��w���`��Z~�)��n�R�:QO��%?�%;�Z?�@�06L��*=��{Z�3K�ƍ��1���PY�=�hɯ�MF�`��j=�n=VZ PX `AjQ���u�*�Qq��N������v�Aj���f>���U��5�:�D�)�"��ȗ���:FO��by[ڡ� ��b���>G6�&�4�U��i�a ֮���e��t���)ƥO8�{p����>�E�ک}��L9ȲyX%�uo����>]4�J3ۜOq(L�XJ�C����� ��q�iW2�Y�'n��4�l[�Z.�76t㥻AU��@��Jn(ٺf��׫$�NN�?�!�A�=� ~}�� %r�=�EA���ml��*3�����#�����17��-���� �Q�!7C���6N�ՈD��>�d���^��`� j�����#wA�U�ȶ�j�/,R��R�{�Zh��swv�bT��K
1Y��+M��ړ�������~�r���w���גqxU��)h5P�1�- ���]����u�v�_\0LCOEi3�x�׵OBF?'�XO@ŀxk�ٰ���z㲯Y)֨��ڽ����x�rQȠe�k%5�pm �Y�O ��o:Ƙ-�q��cp�-���h�Ï?) kh����{������^�{�����
y�څ[�Zh?�����ml
µ�@} cQ`PIb�%���2ċ$��^Z�m34�0U%s}~����������W���Z�6}o��l�
���2[��4�����g
�Z�۰w�@IlE	/���<������ ��ޡ����Jz���ُ�a�x�sZ���ܶ"�+���^d{�s�׀iȄ�����w1q�3��*�TJE՘��R�3�t'Ĥ��:���n H�Z5��=,"X��:�� Xi�sX�$�ς��l���W⸼��0����.��+ K�+P);ߪ����~�L��G�������@Y�����LV0o�Q��	��酪h:�K�6�����B���Q�	�����O�� ��ԭT@��@�I+���,s�H���1���2�����������Y@,;4+K9VxC�7ޕg�\av`�wQ��n���<��k�]]��&�J�����i��^�h].�n�O�ߺ���t�޿s[ V�<	}o����C�_�_���.����	����̽?�@��1�z��߇%�!q��R���oȺ��x�%����F��C�J�>���������ߘ����>�����]ӝ���[h=�����X/�[�6^޺�TR�%�%k(���j����*=ic$��k��| �B6;��D�,�=����慫#X��&0���űK@��~M��3���@y'�c��P �>?������� �.:ԈwrC3���]�XJ���o�3-�����	#zߋ���	�Ў���.�O�sb\������k�"���0������(�0�2afﻝ�-&�0g��FX?�X�Y�xv�cwI-1w��롯	ٍ�G��c��p�e����*2��J��DX"L $Y�>���������6�b�at��l]?���{ow�H�g}v\8Cdo\]N�S�I���=M�W".^��3D�V�����s�_t�9J0:�/�o�l8�#9kc�`N�.�䛓�X	�hk�%��Kn�4�Ѵi 0��ʈ=ʑ�KQn!�Dڨ�QK:d�V$�!����L�)rԼN�?oZ1|��0mw��6�[ ��7v�4�4H���
V��6O���M�F�%�2����u/��@�|����{�lyy���+"(����
땜���z��vP��������w�pR4_2�$.�#��`r\���V�f]�F�6>��/.���dX���F?�]%��Y�!��	K��W<���o�X��J�xd�B��'�r �$.ƃ�״�=}�B���w��w���M��6ϣZ)(�$q�k�	����4KR�C�Z-N�����~Ѐ����߰� @�����Pm�%I�'��;$`E��r�rap���s.T�TX��N�N�j���V ��wU��^��Z�Ρ�g���8�BH2'Ϟ��
�J���܌t�ip��8T� �-�@L�(�rE�)�Ǭn�ׯ��`��8?��3*��[�[҂���ZL��iO ߦ���q���-�ʈ��H��9t���
J�M+ގ��{��WKi $�0�d<!��OݓǏhy3��c6_D@y��x�`#�+*r-V�'��  ��&�j�5+�<y����)�'��㗁+�q��{�*���uG������q^�n���L5�R٪��<��`��[0s/�i�%��}���K.�d�0ޯ��ej ��4C��Ml����ǿ���uoS	�e�kU��A*��g`�S�Ss��3��7����p�妨)�82S����~�e�/Z���4�F�M�p�NLO�e��Rn��md�Yٵ���@ΪV�)`�7�Zc>]��B�*,Wz��DN4�EfQ�����M�fP�H��ap�/Ј�̽���C��u����\Λ����3\X��'l6z�a����q���_ 	z_0ū����΄�k,�|��>�J�[e�W��X�����?D�3�rFq]������V*H ^�8�F#�V�-���QpWn7n���Z�W�(lm�����������Ҋr��Hx�����"[�n&���젊4S/��,�ˑ +tş;;��|}3wWW3Z�zM�F?�5紒@G�  !k���z��F}��R7\i��`U�{Q��%�='��e�S�dld�5����B�F�+����癦�������K6_K`��%�f��N)@�a�' ��_�%�����.0��R��ruN�P[�11��D�R"��*Z�VK򰤑[l*�(a�a���dIC�4�w��3�2�\� ۖ���(�
�]Y�c*	 /_�p_~�ea��$O�/�t�͸`|�J�\(��<��d�q�ǌW���P<ޏϲ�K7g��̊"W��[�&YJ�,>(��J��9S�?E��{~�?��X��C�+~������z����F�^��z�-�+B�1D�+��8�!(J��!���_O9�k����C�m�!4�Te葃߭~����FC�J���d˓������v/��	8�n�Ul�xN�\�W�/�ol��9��TD���Y�} (Rb$fD����r���qK�jiǴAW���H�����^�;/#Q�^���'U�	���pi�.n��i�d��9�F��/&{�ĵ 7��ژLTp��l(��� ���6w纂����2�X{3���d�]�^�4lO�KZ�6/�f�X�;���/��#�N��hW�K%����4uNEгg��~���kK��^�U��Y 4\��l��@r�N��ѩB�*F�Ƙ4�I9��;�F.HF(k�!���-jn��O�F�p'������(Y�������81fY���$���hQIn�" ������׸PZ?{���R�=
D���T��K| �֜V�B+�䏚��!�d��~æ��{���Da旤t*���ܑ�B�ca C(A��2��������iҁ�Љe�I��������3kLb��E�88$U\^�0)ckYג� K����D�U�ILⰐI����k<]x$��`�-Ђ��k�}������A�%3Y�!��'O�rn��rlia��}������d�1� �`/�l۽��8���gڡ������o�3�l� H�%y�֗XZ{O��V);Ewe�
�Ϙt�af!J�K�r�G׼�I�+ ������)��0��?׿עb��FJ9�7��ZU�e)<$}�P�kX���>��*�RIG���!Ҳ��#�1[��2Xrv��� �����)�����ΰ+�M<��$`*�=a���b����w9����UK�8�ztZ�A�,%�$�X�x���E}UO Ac�P��YSq�%� �� ���
��`�I�MVcm\9arB�h$7T�ٗ����+I�R���N�L_t �,�+��&uZ'�=W���+b�SR�p���[J �&���Q��u|P��ᇿ~�%C��+;�'j�F{��=Ѕ	�y������s��FJ[`@���R	��Ұ`m��p��$��1HpKª�j�<�b�I̐�;�fڲ�"��k&�i�겓q�������&#�e�h5�]v�Hq��%{$��� l�܁� 6,�͢�A�@^O	&� ��;;�tǧ�nw��a;;��˯�v���oŲ��@qS���b�E�~=9=��]��;SZNП�� �����-f�aӽ��t׳r�<:�"�W�R{|g� ��q>��V���=
xd[�|XhH�����������;Er �]k�,33�Ia�, d�=���	`�V���{�߅+�X��<��͛w��F�6r[(����ix���V��+(*C�1��{��	�M H��_�q�'ǜ�O�<v�Ͽ��}�� m�s�ɓGt?x�8�V�ԃ܏c�O�����W3Zw�	�D������X�rb��v�� �8�@����%�K��ñ�����7���]|�z,�[�sf��ă5�k+�X��jɄ�Vk ����ѣ�Vq�g�EH���p��\�������?���VS
����==Rr��M)k���������Q��'�\Sb8W}�}���U䒆z���<��qNhIv�x�ƠD(�A�{+�$3��ɥw���@�}a��p&�]��3Xl���)Ɍe(ݾR�#�Wc&l|I(T�r�/�Y��b�V�2h�4k|����R׭6����z�@�=�:�_�"(��͆*O�d�
����j�[:>Xi���YO�%���ݝ��)�(*�/�;��bXmָ>&�T��a0��??��q�,�:�`l�2ESzq/q�AA�&7�F4��en*����������2�1�]���a��R�s'Aа�t�������v�'��,n�7��[���&apc	C������j��ػ��-���3��Ѿ����������_��Ȇ���f��m�X�!ۏ�CX� �����nC�e�6z����]�-&�%!(E�$2	��wi�A_��M���ZJ�/ ��hE�*-l�ۻ����4>'�
�#`�-)G ����k~��K��I���swy}ō�ի�  �V�Z@���`퀋ĩ�>!����#Z��6�2Q,����gO9O>��Ѫł�T8A֜��ӂg�V
��c ���s ���p�i���yuJ��dd��"�y��]��k���ߦy��"����+d��UcR2<�mC-���3Ho{Ώ��G��/�뒎�/.�	P�r��[�y��Qs��#��"�H���2D��a.7,��=�������d� �;�s������t{_ݠ�X��Z�տ ߧ�R(LX�2H�)N�
p\�{&����R�~1�hӦ_���DR��w_ZA8>&V�uf�_x|<���Y9/��?�:�-g��F�Z��k�����cs�Ouf�q?e���kk�>�Q�$f���Z���lo��[��9JJ�-�����O>D�/>�nqi�3���!���2a`� i�����[C�5��Y(����`i��f$9	��d�.�ESکh(��̒JZe�K�����	�6lu�zm�ؾ�1i'�Vѵ����W�6��\o����U�Đ[���q���m���<��k����(u�R������̯����B���m~w;ٔ�d�b���X�S&�|7)��s>�"�j8�cN�����bK�x12 w"0 S/V�%��[�l��	N0
:셫�d��> K�_���}���q�z��D`U�b �S5f���d 6Jh��Q�؛��O����%kI"��8�����u�`�\S�ᎻaO�*��й�q#𒘥	�0�[XK..n܏?�v?"~�\a����(�#�
�ۉ�>b��55f��.,���V\x����t���e6���*t���ZH ����೪F+��RG�c�F��l��J�V�� /l�mKk6��J�T�..	d �����h�_^�����){nA 6#T䘶K����:��V< ��w��=�$�Ep�r��;��QT?9=#xƗ��k�Z]�B��6\�{�������{����9�# f�!��c?#��������n؇�k*���S�Q�K�Z�k�k�������I������;��������ot?�;qGg7����X5]����E�3{��X�ǜ&_qd�^��k�>mV9~k(i2�ڠ��l�����t���C ��/��b|W��Зb�����`fqW��w���<}�\/�M�Ypy�7o�.\�E�SbP��\�YQTP�&��]���W�b�.�%�V �w�������<[�Ǘ��ޯa������!��Q�>h�z��d�� Yܵ┦��*ۜ�ĀGE.ҩ{ȕMCRN��r���ؠ%9�&��@����	���/�a焀t��#�g����:YSGK�4@[�̎J�2���ؗg�]��jH��y~|��B�0��r$�h�[�y�#v��v�y��z�R����`[YR�94Y����2��l�g`%bd�k��P W7F봦$� �� ��wr��w��{{|���2b+!:��9!B�w&ZyaŶ������={E��$��� .�H�
W#6H��	i-��`3����ٹ{��=��X�������?��l��|�,ؙ���2mhpK�@�� �k�	X#h;9>e��5)���<������&��G�X��֮��r�J.������%��n��׳�5��������|] �e���OO0~��kA���5\ld�{�N�)��H퀾��X۰��0�"���:�WC������!(�g�g�(2�	�yZ �u�k���D��Ņ��L�;����7ĝ��-��@{1c��,��q�g�����q `�+��g�����]\��6�[�j<n�,( �j�݉E�Ӧ�*���p<��!�	 ؇�S�.���z���?�� �9V5��4%,���%A�rϷX-���_�L���H�Vzy�����үy)�d_����293x{MC���������,_i����w?k���L�`�Z��T_�O�i{V�69��n�wZil-��%��,&|�>X�Ե�����1�e��:&ɠl=�َ<
#Jjk9�r|����Cg��0�9!t�h��/a��{�?,����y!)~� N�M9B��
"���B��tY��VN��N�Ԧ?�|�P:=O���{2�✳�`�yΪ�)�1�^��@�!:�C�F{�|�dhړJ�ߠ�SwR��ʹ3X/i����+���@(�·I��.}[�ܢ9�9F�g���#T|�8 �5���d�TS`�LU�䒅�k�<׻�;��s��@��"�R ��Ta@1ָN�ʛ��Mi�3��'�H�ǿ+7��튛$�����^��u:ZW޾=r>����B���ތ��J{��-y�޼�)n�[n<�ښ��@��e�Zh��$�n �����ܕ����HƠu\�ZH<�eq�Md�-������ �=�G�� <j�!���,�%�ooM-H~��\�V�����3C1�BH�R.J� )X��jɶ��V�7 �E�8'e��R*�,�)�F��p�ڃq	U����>�tu+��-��RKn������6�k�$���]���`e��j�u-������gu �N`�V3ԉh�j�����_�z��Gv~�$�&C�c˹/ֆ�������}���N���-3c8���s{~�D���.��j	T�D ¬��_U��myf03p%%̣tw�3��՞I_z@>��='�m��7�'ɻ�qW��9������d�*2�+��O��)`�$���[�{zˈD�Z"�&��2�ƤO[l1���܂{�`�PĘ�ߵn1�UVP�Oo�t�ڜ+�S�u�;Q�� �WóD�5M��6�g�,m��E[NhI��i�S�Z�N�&��"������@v$��}�w�>�sy���-wNF���4�ѝ�:�DK��������!�qګr�+oGF���sf��/7h''AQ*G�-ĵ�����]�����C\	SK߃ǯ��jb� �i��^�5�	�ڭ��	�de���Zs-��A�}*B�W�Y�%c��%������k�oQ��@J.���������76�&n�q:���Y��Q����6U��/tj�Z��iM���p9wrvI������;2����FwY�&�4�v����kRc\�~��t3��e]���$R�������D�k(�D1��x_T�`�5
�"��D��(-��r��Lb�=�7c� ���q��@ V@�l�j�q�E)�Jƫa,]Vp��|T=�BFj�ɱ..�	�/��1,��b::�^CX6$��L.�O�Z�im]XYq�nQ�-��	@�lF�c`}�"P��EM˫�Ki�[����RC/h�[	v�x��"��v���q�����$Q��k�bIV��(��p���p���;o]�X��
n&[n��2��J[֦Z�̪:)L6��l����s��� I���ҥ�Iv��{�W�����_Y�&K�����_y	�O��ޛ�F([��5��h'c�ؿ2����B2}E	ry�uJ�Q�;Z�\qv�G�Tפ�)���m��C�e��i�Se8���k��O�[���p����Zˆ5��z��5,Y�7�☾J�B2�p�A-e>h��$�� q8��4�Y��'�����5�S3d����\��Z$ ���)��e�ѦSH ,7����B#$ fЀn���%�J����r�P#�W;~	@�k?�?�$|~���.`�d�c��Sj�j{���c���,+������ M73��K����S+�L��R�]�v%>#ZmpXZT���#'����.o��:u׷��dgύ��P�̒����,������~p?���ٗ��͛7,����ʋH,D��+��Ѷ��m��Q��Y)WO�b�@��o�V�ǲP��/��f��8�[ݸ	lI�"� I��J��w3�v�-!YU7���	��
|b�pY�����8q٦��ڕR�H���񜰜zQ���x���rQ޺V
Ը4BX����U\��*��*�3��T�/�i�^�t/^>�X��x~q�
/^��%�?��O�u��>���rv9��!HV���+��g]=��,N�0��<ܜ�9C������#H� ����SK�`���u�Vj�ަ:����스�V;�Un7�{�E��b����o�p9n����UxL|y�A�Q���5qdѱ�ib��5������޿�qO; ��_��L7:UB\ѧ��&˱�7�JW�HSkI���	�-��2ր�* ޴�Բs8����%�m�q2�������w���	���z�JdE���-�|1��Vd^J9
>d_'�aA��I��
��
�.�7�V�7,nZo�Ng�-M�2'q������4�?����e�
���嚒�)B SCX�Z���0̵�.[(,�^&F�S�����[���E��A��q���3AX��	�{Glp���m���H��,`���ep�]��V]զ�Y�4�7TNK⬤�Nדw��ѱ��]�E(Y�r=nƽ C�Yw�Z�pJ� c��]���pG �y	VzǸ/�۲�/��i13�f<����<N���aҿa�EX��u�k�5�Nun��M�!58H�T".��uɍW4a��u�ੲ:fT̬͝3��b&Ev.e$i��JX K�MSqܚ P܎9d�L_����]U��j��4)kO9#J�v�O�&�:e&��'���'eC��$A�B�
 ,|f>=�F:c�G��cwx(�a������k��12�����sㄺ�������Ge�8� �f����[�֔l,+m�X�"�Z���f��mMF�;8�cܛ l��5Q2;�M�޶n�lY��� �a'�[Z��Z�1���(.�J�h �����2c5HALI��&�|�a\�P�59��S׏{O�{�?TJ�[�ܯ}躵�k�������|�Q%���� �%WX�2+�;̱L;K�tϔ�Zj��ie����;fV7WwL�|:�#�}9{H��!��ڪu�j%������I�Q�d��Q@�N�h�����hY�G��8��SʖH��졂ˮ�P�E8Yg���영�X�U���}�w�b������<�
 �ڭup0�%���9Ju+�۲�w��k�y���_U�or��&5K���ƪ�(�����{�6� ~MR�8��<I+-�Q��$[m��m����\D��m$ɬ߄�����h�Q�b�A6Cb��;�,�r�DH���^�nQmb���,3+Z�p=�n\����X�:e��0�i*�A�����c�^	g%6�f�����5��נsq��~$mT+n�Fh�%���z��U��>!S�[t�aXѼ*Uz�Ţc�3�xAV�����h�m��
��I�Q����ͻrզ%�C\ V���
�-�Vdh)p]��g�IQ��yPW4���[�.W^�yvv~�g@.�o�7��N,��5��%�7�rߋet _��<v/^<c2�b�����$�}z���בkɳ���s�jT�7��r�M�D���%��g��6_���á���fz���k%���Zʒ{ Xʍ������$C	��ۭ8lbe�g��b�����v�tm�ms���˶8[W�������G��O|<���2EK-��/ ��#.U�9�nv$ut�ZP�İ�+j��8[1���`� �pL��6��w�[�G����|��bx�R܁7�}���^�S����Q��;S%����3Dc�#o�c_et�6M�:´IS1���t� hHi�^��>�����[i�2X$1�G|W�ͱ��S���R{Ҁ>7 ���f��iA�����U2�f��+���n�����=8�=��b4��~|���;���gEDc�,˶���bs�4I'����Y���L�*ae7AW�-#�5%\d�*��l�N
OǟcNV�[Y�l����:ՍL���\0�>��V���������6,��t'�P�t%�͘��2E��W����j/~�e]W���{#����t'~>r�El��Q�ڳ�JP����� ��?a]jX�:��z
�����[}Y��Xwr2�e��e����V�TdAk�O��1U���j���K֡K6-i.(Ȩ�b)d��Z�X�������j���"a�Ӈd7�$)��yN�uP� `V�ɸv{{[L~ ��b��������u��87�.˾�>@x˾��IX��v��P��;�t/�,f�����\�T�dmOt˚��$�4a���UŁ��3���-�C6�^�NIg�ڤ�m²�J�f��:&J�+�������oM@+_���,������%���a�2�3��������ß����3ֹR��r~;��RA�C�󂌻�r朏ټ}�B��5�{{Q�f0����5��Fzn0$���!�x�{�C9gR�\K���K��W�����x�e\�-�Y�h߶�y[� 0)�mG3�`���#���j�����._�R��b�SP9�ʧM$hb{�)�a�u�=hr�Ej�q�=�[�����@X��0�R���+�D��Bs�TڷUўr6�����E�|�I	>g�)�>�,J�;�B�O��K��*�)�<�n�����à��� W_R�4���%��V`%�#��o4�Zb���o��*�3�?Ω�OU_��(㷔 �G/H 7S�+q�	xr�OB��e[�΋-�� ���uDm J��:e^�,OK���&�ߤ͐����x��V,j�8I坨�������ۥ��:>1,:`���^��U`< 
�����g kG+%@������&�lv���@D�����nwg/
�5)���
2C�pQ4����d?���
��(p~}uM@��d�(�l<������}S�+2La�Y2�����s{�p oZ�<"pB6"�Ad{�_\���ߓ?%� @��ʵ �1\������_�?��"{��V宧�6���ͥ��<u��uƷ��B,��Ȱ���vO��kc�q9�n�Niֲ�KIɢ}����y�����@O�xM\���6ɠ�^!$�W�MJ�ܴ����*�>�&$L`�$7����G�x���$��
�	�����{��?�X���~��?�>>�贿��l\d��!YȜ�^+c=,�$������xf�WU��~{ǔ+��Tp���1ǰ�w�Or#��k{�M�!��|mZ���T����Ib귶-�j��L�fdT2@�-��f�Y̅�IIXY��/� �f�������D��j.�H�VU�	�oepdv�y=J�ȴ���@M�ɲy��h�i��)͎�����������T��LX�4��W���L�h��YJ�e�.�2��1 ��p�;�����?�z�e2c�2 ��;�B+$�m���r�X� �03�A�9X8�Z_�BZ�!4�6��t��n���-Q�l���H��4x��ۈ�%�J���� A��ChW��^�`��#��:4َ@E��C�Ȳ&�`����)���4Xa�����V���K�c�PW�s�>��N�D,K{�`��~���j/�C�d�MX�Ɩ�r΂�2��+�� �+ Xt@: �|�^_�)�A��L8����llOk,X� �FZ�=ޮ�u"�5)�F{%Htn����"��5&G����s�@�茰Z,��� <}���������f6!�܎|�jY��hu�6�Ș|�����s����$�ë�]��zv}���N�E�c�0��ƨ+�E+]SK�Yp��{�Wg��T�\�VH���[#��-�6k��U��>(�Ql7���ʳSKB�Ö ���ؗ=��.�����hS�Ӟ��{����d{� �I`���%V�9d�����o��'��>���6��ÑI���EK�S���uU�E9PuG+�q�G�q���\�7A߫�J
Y�SEcz������.?-+2z�`��yT<U�g�o�J�Qh8��a��Ţq����m~'F�V䧤Lb���})��~���Qu�����T���ு�ܯ��Tʋ�v�>�D��:�,���Q0�n��H>�c��i�U*�PF��Y}zN]{ijF�M���ks�N�KCU,��b}�C����L�d!���kg��~���>�v|��XO���A��Bg���mw�è�h�$��Jؤ*�hUq�:��v�@�$A�J��  �e��Uv��o ��7�b��8i40��=�yW�K�<`A�n�"�f���i ��eϩz��8`-�=~����?�޽x�� �G�.��H4#X9;��_�G�K�m�T%�;ɆÆ�ŗ�	^����Ϡ,R����R�X��	�?�@�7�j�C�C��\��u}}�\O�u]H���J��~����-	�b�`������V�--��<�(\��k���s�/���"�y"r��r= q=::"�-�>��݉�C���tB�PF<�� �����;=]1���S�I��p}-�<j�o����~A�A,{( � ` y��2�R��0���{(�pK*4����;;��E��t��/���{��1�@=8�DV�J���h;�\������f��ŵ{��=�)$п�K��)��u�k��Ŋ��w�Vyґ�noG��C��-|��V��	x6�B��cp��B4���幟�ݿ߱�>���WR�T�j\��4�n����h�I�S"^G��>��;e)��/�,�9[a�Ù������r�mr ˼O4/vN��Ce������j%�d��A�G��`]D�Թ�݊�`U%9x.���d��k���f �����*n>�b�WXŅ�V�ǩ���'�Q�f2wOH�Œ����;f�I,��A�Y�h:�d-�r0-eM$��ق�b��DMg M� ��nf��k�W���feb�W%13�L��Z�}l���v��o���_*~���3���t�(�R���5Q(�E�����i���9��mdI�d\�|c�g?�vWϊ�r��Wk ,�P�iP�y����!���������die��teZ�rJuE�
S�n7�f�v�dbD�t3����<��Gq�Ś�@�w�)Q�ѓ�!�Z���ވI 8܍���_~�?�X2��_�Ķ�uG�	8 d��2����Z�x��=AǁX���`�?==� �2��;?���JZ�e<�V���ՇB�_}�2�gKb�h�������X�c�-����� -������O�X]ƶ������ij�+�$q������^|�$��xM�"���OxH��w�H4�b��=ڏ�h�`K���Zl`��-J�B�P	��*�\���TZ�H�h�� ��{;üXh!��im�����˗��I��[鶼 ����,�u����P�U��W���:'�����&JI�(��i݅�,�E_�:,�X�|���u�3)b2��[�N�%&�\)~5 �QԄ;?m�~��1eo�6�y������P�����خ�h�]1z���ǔ8�ap�ϗא�e��U��M��f��Rů0�8�y�r� ��B��%2�����kֻl��^�����n0����͓�A	IJ��ͨV���2f��{�-�T$�sѓ6��Cƀ���H<H�R�8Z�5��`	��m|�Dm|FM�G��Jx��1���NK�8g\-L��1��ai�{'�j�J X��i�R�-U_�kv��]5��aY�:0���`1a./�4ՂY�xn��he�U�%\�gj��DKA�.�Xq��s���jm�n��p�����u����Ђ���?�	$��aM�9�R!H��� ��]3�c�Ҭ����0�rW9G���"����@,K��:�;әu�?��JkF�5�ݳ����������q' ��<ަ͉KT�0PLkI8h-c�b�@!�8n# �9u��򻸐�n��7Sw}y�no"�:܍��w�q����f0�%�_�̑̢���%­5�4nwo�����'�l!�Nb�����NYxh��������k�h�+�ѣG$������'܄��ҋe��y��B�_ǾPs<J��vqq�>�ci����"��x�K�cdF�+�Z�M 0�,a��3��;����~��ߺ'Oi��X�:�5�c{nܟ��\�J�������L\F��V� �"�u� 6ZE�ZcGU�krE]X�	v��kf�z'�[���=y�ޗ��/�L��t-��]�ޣr�;���2����<ltP��n'AX2\�K)�J*�u:����$�BA��8PN�͋�{���]�ƗM�j��� !-ƌ�ӵ�\�����9=���J�@:���R��e�s��p[���ϺŃ_�����A���`�x�ĕo%z�<��/M���nI� �f�^AC����ɶ��5�x�ԕ��2�U<b����k]�|Y�njC�HJ��fz{�¨���x"$�,Fj#T�p���r^���Ȍ�b�~���� ��4Z�k)��j�5s�1�����K�oEm�ʟx5���7����.t�>�`(�{॔���­��X��*2�����
p� =>ޯ�y_�89��P13�|ȋF�$$X��/�_�zӜ��ip��/��y��1�2	kڼ�вI�O 1<��O�6mҩ�I9��o����u��CM� �9
f�`v�k�ȗW�j��u3�Se��}⧢�5�^0̯��$fE֝d�u

5x�V-�r�+��W�0nj_�z����/��=��-��<��U*�����&�B�i6.-��É�k:�sȯ�\�/��b��j�[��0 J�*$܄K)���S���^X�Ro�}��zhb#�%  �!kj҅F.��%US3�>,K-[p��5�$l̚�[өl�L͓x���@&��1�`��+��x�5�@^�bV_k�U�Nb�F�Z��(���=���貖mb�GW!��# ݚ�9� �=\��*֠�%��<b�[�k�be��NǼ' D�Idx����䏜�5���B�p��|���;�/mw}�a���sgk�g犱*�p#|�8$�n����A=V��Ǹ��aQx�QE!o�\O�O��2�9�Jvh2肌si,s2�}Z�Y��t.]��q����Ȉԓe�Y��I�Ja,C�����A�\Lv��s�5Yu����q[ب�~�0SHb�,PX9���:pIj|��5�C�sO���]���}v9��t���b����l����v�EU�� ���axR1|Ƚ��i�-�`LÖ��"$�#�@<qE��ܙ/�&���D����5-��I��8�Q�s4L�t TKW�ŧ�Q!�)���A1ݫk�D��Ƞ�ₕ�q���xaя��͎��.�Ы�	נ�Q75jj+!l��J� �6M�^���!~�b(�aҏ���#�lfZ̎Ƽy%���W��x��!�ɐTQu��8�s)i"Ŝ-,�6�శ����r�������u���O�f�ơ8���m))M�Vd3� /��%[_��DgRj���8��s�"�*�)�CHM@��(!�Gt1-���(4� ��z��c\V\Q�;S���孖��eM6"hNmۥk�I�ba�G�"��n�������ş8c ��^�!��c��-}*d��-����Vx����^݇����[I����Y̙I��f�Q�-��Jp-Xk����؛"kr<J�l\��O^�9�5�[ɝZ 6h��,6Bz:"����mE9��Y=����Ge�:9���o�//����u ����K�^e��2FhC'֫�K�������F�����be�����,��l&�ׯ���kwt|�z��B/A_qL��9�s������؟�,o�����w�}���;_�}l3x��v}u����#���SR4���+/�R�`N���'�;���Y�wIa�)%��;��L� j�b��.}
ʌ�@���P�dW�%�P�W 0_��$�P�� �\{ʻp�w_�J��sQ�����������OÝ\���hf�J2�bJ�"�-^�!�Zu%M��2\���\��k�X�̢��Wv� �(r���K�.�_��I=�FP�`������V	E������a"�yl�ꚡ$�@��A��r��O)X�G�o���p�X|��F�&��z��-�Y�\o0
3rɃ�- ؒ��/����(.6)%�u�s��Pn�Z'�m.uo&{a��X<�!L�|6Rٳ@8Z<���~:�r���G�`��V{6ݦ��	�B�D��H�qg�JQ6���6� OX��@s�*�v�3�V��lR�ʃDy�5!0y���Rg����׿�j�l��V�T3�XI�B��9N[��6q�xV�����"˰�l�]�q��.bb���ȼ��q4ԴL����
"T�ħ�k���E0� ������dZ�m�`����G6A�*`f@��x�nBMʷ��F v���')i���-t-�f������Շ�8?��`�4n�W{�)rw
�Z�V}x7�oپ��]-h����	)�q �֢ ă��a����A`h�۷�| R�4�Ӊ�X����>�ׇ�,.�yP��6~���cj��Qh�����������6A|�~����ױ�N	���y��=�x}����{�s�
f�kwrrD
���"+��p�}��~�ߣ��5�2����;X��I@��ߦy��g�r�^��#-P���� F۾��{����G�6��y~~��������i��򌴖�*a	N��"��S���)�����*I��t.�"t.Ke
Y�l�^܏f���R `�2�ﳷ@�T���\1Uk(?�6��SiR� �l�ț~!7l���>��51�L�4y>_�����e����a��,/S/�æ}�\�����j}J]�������k�Y����3�!���k��D��i�hJ���0� s�%zØ�+V[�C-֯
J<T:)V�Zes?K� �);�>i
��D_�č�U��
h�0Z
��n$��U	�#``���
Jq�ѻ�0+Z�l_Ǉ�Z�دH��x� @�W��AW=i��K:�1��)�}�|�]�@����n����+��Hy�\����b�T�v`��kP~/�R��;���9.|��=�!�����c�ؑ�;iS֨4�C�5L:��F��Ϡ�����=e�-�@^&Y�Kh;i]�_R�
�w�ؼ`�8m����ֿ_L��)z
 Y|?X����M���L��.o�H^}�:ы�����8	�B(Z�|pVC���,�����~$��Z���W��f�u�{)�Q�8>�I�ї�=
�z��5�u��3��
�h�x]���?��D�"���C��We�M�����g���Z���!E�yķ߽;r��:;���a�=�+d/~����8��I��:� �\<y�Ľx��]���/�.�D����`�[HN�������p?���po!�)>��>�8��R9��А ���"X@[2�Շ����������u�p��f���u��Yl�����V�h/! r����b_��:��^A���������={F���%�.8��3��K�\���v=�ݷ��]]\�7��PN 1�lxH��P0����1[�?�9>�;�@�F``�b��T)�QrO�g��?�]Ku)$BjY*)���^hS�.F�����O�ًW�y���S$1��qō�ѳ0��5�_�8�2�O����*�z�ʹf��M�1�7ZPc@�'Ŝm����7~��q����ְ���N�ם���G9����P�h��N������G����C�����u�������}�Q��8IFq��>������_ڿ�%��I�@�tk�mE��}�<²u�$�f�$���B%�Z���nA �6�Ҭ���@��.b�ʊzP��H��Ȫ23�D-��]�[d��.>S���|J��`&��{I�!K<$�^�JA*�'�lEqe�(�F�������*������ş~�Y���(>���F���V�fsjj��j?ŋ����x�҄?�̌6��v �R"�``�E�Y�@˛���)L�Yc�3��H���	PS�E�'^�& f�*ɂ5<m�g�Rߵ
_C�!�k��]?-D��h//���w�+��`˗/�QX�LSL_+�חW-h����Ӹ*�%��t�r��� Ұ3ĕml�w�f�v�f�H�V#��R���u�$�yX��r���Z�!��x�9��n����n��N\����)n�o޾�1� k���{�VJ �ֵ��`}Q�b�66�L n���x��l\�_ -H!�f���-L�_'����>��a�1�t��R+�v
P��#P:f�����OON�~�ҥ�#t4�pÊp���)��@`�wdў͵&�ϑ��g���"p���ry��z.�kT#AlV�L���G��V�7d<�9PX{Id'�V���8ՌK�	����}�dU���l���t��hI;b�)X�F(%����t���p5����\�l��ᦡ��VK:-R^J%ᚇ��^���s�x����\�a�uil�����ԊOG۩��eBݘ� ^��7��`�D���B����r��x�|������
u�]1��BQs�"��c�ά�I�Q��۠쥋�r�#�l  ?vް�~-.'+#�$k�$dcV%�ƪ3:&)�$=f��^Y��\��z�R	���$��c�,Zǵ�K��\�X[�N^��cI��j�>k(b�2�=hn���5YBm,�I�b@*��l�49o���끒$eh��Z�
����O���$����%�]�3U��,|&��NX0�e\�nk5�-�v&c2pc�"j����)�(���t�<��G����KB!( Z/��͝՟�,������N�v%�U�FI��v����-�YfM**΃sq"3������{���1;���ZNE����zqs�y�R�M#��pn��a��4��x�i���u�
T(��.$�f���D�6-�͋9�d���w�)�����ߧ\�w���N'"�V�A8���^�-�aI<`A Z�|��l`����` _IY��b�%0��x�I����>�lE����*��:*.���k��-}��n�ؐ��Z��+�bE��-�W ���,6�z���j�>H��l�sw��,�p�eN��p-1;g%�(ߑM�; T��H��NH�F�~]��]��b���3��4�x*hU�>�sI�-1`b�\�.e�2�>Y�d\{�6�Nkٖ���48����5X�ҍH �&.x��r��c�Y��+��
�^c[��ꒀ��� ���p��������H٨\x6�R��b�:]R�:���CMő�ދ��H�Y���~d;?}�v� ƶ$�3��3�]�댙�jL��4��t-�P���\����7:�6B�5ܺ��Χ���h�'e��>�J��so��:��rc(�� ���Qy��?��6�E��N�׀���,�zz��>�f:��&7��ـ�]GW���0��i�ʊ,G�|�s1���A� �_% ^�	8���X�Gr��OF�ۙ6�Ԥ���#�ME��GS2��^j�!wm���<[���� �a\��I�'���_�Y<uۻ�L�8�/o����%� 㦦u{C#�J�q@t�&��&��$++���l�5�zXp`۫ ﵈��ҋEL \��� ɲA�&-_����d:����xo$v�op7US6�o�\�,����P�T0��a)���TlGW@`-_�E�sI��'n9ͽK�H1���H�\6��ˮ���_?��K��M���l�L����Qj��:�-_�ӫZ��X9�!�g˴���x��Ok�I=�%�f1���AI\��d6u%R��k��J1S�QL"��B�P9HL��� laC����$ �d���aI���>�<kK�������ܑQ��5����Y88�E:	�d-���d�ʼ���\��׺�ƾO]D�"��!���\{�W�?+,^���.a�/��� n����bs���`C1kn�x6O+,��Z%�qZ�t��l�d ��������ˋ~�\G�Z�ޡl�QI�P_YhI��l�q�^������.p^�
 T��i�����	�k������h�I�Gh�3r%�&����fj�K6C�Pq_��pI!��e�dc㭵�{�^J }�>(iq���a�x$Y�Q��Tu�&�v���S6���I@���	�&yk߳�4�(�TI'7dp"�d`"(ڔ�ۖ^R�ղua�bv7�(kG��5r��Q�6��z)&�t(ǣ�va�*N#��B���q,jx�s����[��Z�$�R�Y�n�g���� �`HRAv4Bp �>�àv��;�� ;:>%��,�6X��
fp�17����0��͠��/l�rN���J0��(�*�V�;��F�p����1
)�	���4W�vr)�2ņ"�(k��%3�+�Y{�ѐ�#䞋�/��#-n�5���Щ��Pkv�׺~xi�&����g�Xh���q��(�����c����"����c#p.����gf�.ϭ|:�i閐���M�6��U�R�s��D�|�B��Y4;ՒDy �ͭ�C�c�R���Fk���<�sX�p݇�j	����o��t�y������w�XT�܇!���k$sx��K��^7L%�T�s����� N�0x�,+%H2���P_c��]��hM��a-s��E�	H�����u.�jBt��X�m¦yo�d[���)�3���%2MdQ���:0�c�	���:�*�a�x�?�z��3\H��Z��3ߗ1�j5���j�q#�MQ)3�� �A+I4�	Cl$��Ӥ�n��N;M��4,]�����?��Cɑ$�Ts@���U�]C��W�dD���d�v��Lwɬ$���Δ<55"�zw[֫�8�͍�=eO�3Yob��jfi���}�VH<:`��d���p�y#2 g_��^�D�f��Y9=t|M����d�?M�裱��=!\���L�*\���C��M�H�)���5U�Vb����'\.]�_���-}���yqZ�{�6o����Wخ1�V�f���^-x����<^��am��%��%�{��s**�]��e.����1��ޣ��꥛�_~����
5�Ta�DL��V7D�����
B=;���?܋[H6����΄W6_�� Gl*A{ɮ٘`��GN���$�b���� ÛL̀��� M�fFꧧ� ��N�[��9���c�|�x+1?���%��8�a!�r�pΰ�~�fmֵ&��V�FL�f*�'#�8��ӣ�z��u�U����ơ67�~qF���s��=�^t͎��>��kV3H۠Sr��k��b*C��u;��H����B�BF��;C9�=�F�]oesZ?�)y�֦���3������ŏ��B��|Q��9���LQ!%�=�8�D ����9 }:*��D�n�� �ٵq��� JTbjm�M9���Ol����X���~ނ�xm})�P���k?t�n|��Z�F���hm�������q�{��&��v�W�u��uYT-u��ڜ��6�?[�X�+ J�ugM�3YY+_��f�6w9�:�V�����/��ӆ�F��':�~l���"c+�TZ{��2�>x��q�k������xn���3W�6�����}tQ$(1#��ɓA��=N��&o� H��Rw�LdrL�J�ˆ��昨n�Ų���+�y�����G߽{E�g+:�d�d���)g�05��,~��v#�'X�|���3Yי�k1�^�:[֤)2���t�����u��u����]�<�z!V�]c��Xuv�(��\G��n���j��ll߬尦���k�����ru,e/�* �B>�[NW��Y�P����Z���7�y��$��^�jG"�4�H�A/�.�L����0?�@?��sA�?���)��aMm�t�f+K}%!tF~f>y#�W$N�)[{�g����H�|�9{���T��~j+d�4���!\���c�3@��Tst�̤?�7Q��@&��õd�m<�����80X���ƥ A�-���Q���( ƬY@�^��ZG��W6fyg�?�)<M���5}��==��QW��,�O�)@L�J��+���(Uw���+��eȮ�`<G6ٙ}� z�{���@@9��d�'��7f����J�n�n�,��|�M�_h��Ϟ p��C׊ m
�F�W�3}��ωv��2̮7��`ݮy�`e#
���S�Xu!릦�]���|5V>B�C
]v�]�pG3���%�x#��=׋�k��q' l��H-@�j�.[��mT6_�KY�j������o����S��*8]�K������V�xYu��4yQ������;a�)����ĦXfЖ�r�0Ģ�NO�C�GPk��&W@�[� |�\Ac�y��pͲ�//N����w�{Go__���L���� 8.|�:4����1c蚵#�}�@|��-`rf�y�����M�%����#�x��6%qb�t.:��ׯ^�sb�1�%�1`Q ��Y�si�����}R6&0�³5���>�?Vu�dj��'�*p�^�3gW���
q`\A�w �5��ʔ��F����zyN/��U��~aN��o��ӗ;	P��L�4r@6��)1c<97�_S-�Ţ�2`T� ���~g�X)L3�J��n��d�lo�㏜QM��cOƄ�������KӍ�����1h@�D&�2�*ń�j��N��w׶}��e���Ĩ����Q����$-��R,_�y�Ϣ���Q(n
�g����'�uuq)��`�*���Ī �@�ʻܴ�~#̽���o��^c+�& �9������A�(����n��(�L�����z%l�e[^9Ǿ��}�dI�Z�9<s״+�r�{D��N�/�`:V�Qs�p����ZtK���#�fSRyՙ�AX7D�`�5�S�Rh�0%ɕ�K|K��2I���u��D塖���T�;����&��@S9�q������Aj�8M~�
:]k)���
H;����ߜJ9����6�a� lPV�$I�v2!c_ XW�s�{��������@oJ�q��&��=�ڵ/�zK߾{E�E���<Ú�V���/�5$�/[m���S
a��VT@���T_�	��2�g�̻���'amhX��gMP�ڲV����W4?Z�c����F��>��/.� ���L��N�T��-t�q�`����twh���,�>\N��F8z�^�K�S���e�����Z���;$��i�s��+�/�����_>~��������J?��I\�Z�lN� ԣ~U&�����A��3"�P �y�d3�Xy5}���O!���lr�ř�O�V��F�ϻ �r���_�(K�E�k�IMkL@={��|�9���`�0~9:LJ��F���|3-����4����Ղ��cО�D�P����J:'�4����E�{IPY���p/��,x9)�D/Űo�\�$ě�(u��"���� �"��s��
l��7�,���rm��63�ڏ���1�	�Xž�?q�)pܳ��MA�n��������c�p^��=G�om�2����}�[@�d�ܭ�cO�_ӟ ��[rY5z��	"��	X��c�����ƍ&q,V�@��Խ��TC�B�����3���$�LC���_�Z���2�Z2�
'H�w69�}W�Yꁱ�sA3�c)�VE�^�9 ���Y��+ܺ~��v���4�!
�}A��>�^��&(+�R��x7p�l��������}��$�!i,�oִ}*��tI�}S����Ы�3Idw���X�
!�P4��%��Y�67"'�HU��.�7��k7_,$~��2��-���ϫ�}��/�W
}��%s�HLXya��l����ܐtZ^O��p�q���y���h��m�d���9]��t�YT���t�(�}�U�j�\d�J���ө���)ŷe�o�
!��kl�,XČPMS�5 ��L�2нg�p��j9���i��zMo^�[*Ύ�B���k.����ayW��B�"]@���c�壹�<Ƿ18d�t��h��3���}!�abEj�z� ]����ߨ�:򁿣�x���2s��ęH��q�v}3 �fMLc1z*n�h�a�����rU��P�u���`��@���:�ѓůx�Mo��2I�[X�RN)����E���JϦ��&�����73�g�=\��O� ��?Zg���K5l�<<���.�2�����XOϙ���#��k������mH��߁E�5�=�h
����6�l�oc�i"���[������.�@[�U�F�`J��@���%D��&#�0Y�WҾ��yo.L�p&�d�H
����+�]6_ӭ�m�L~-��� L�sA��@R���=q�0��\~ڍ��-��+yc���0 T���U��w�]zR+T�%rF��-�M�8�*���Ȇ�6��0(��p�6-��JjGg�}�楼�O8��̉�Z��Wm"����T�$ː�96��d?�m��wke��Fbw�6��օUE��v�mŀwW�3�z��w����PW��nҍ����Q��⨣��#)���q�R�;em�M����fZXmO���ū7�\�$.l#�L����H	YhP;Sj�� M��F�Jƚ��2������ 齳��3��8���~��N���~I������o�?��/��/��Ki͛l��Ril�i�p\��3d�d�زr�$˂`2�v���w����"LItP0�9m���o4n�cMX;R7�!�v3n���K✞�i��d��{c<x9t��Rx�Mg&uWe�/55~��e.d՛��y�t�Rl[�TR�(�Z2�8�ر�]��h\\�E�� ��^4�\���<���p�~T��8(v�Ym�QH�LCX{S��=m��I��DK��y�םZ�bP���O�	��xL�����9�U���Z����[����C�|�iB�E�N�5�X��N��O ���d�`�.;#ԅ��:��VJ2I�Lsѳ�˪7[�Ă�� �������k�Z�fA0*��z����S���X������Q�B�K��j���:^��P�4)l�qO:$;��'K��+��;ܯ8 �#X��%T�f] ����7j6�f_H)�x�`�b䊇�v�0o�;!��ˋ�I�z|yyJ�^_��חtuq\��`��-�L�匧q49�{;�D�?�%�N�{aN��\��]�h����N	��A�/p{���]�<����2�j���Z݌	{K�#�m�	w�zDx�1����C��T1����r��tVr+�au�gg�Wtz���e��=b�EsZor&�_�mld���ҟa2��D��F�!F���J2	�B��J̈́DV��G�贔�b1��x�WmՈ���ߴ���i��/�b�\�	�����蛑?�?���� �jJ/����yw'j�dڳ����N@��RO���
��iOܷ����c�8)��Z�����!�h����$5�rM�\�O����P�wz�f█��`� 7i�#������kv����)��_��BRr��{\֦�Dޘ��Z6�2�ΎW��ŋ"$����mwf-�tn��W�1��@�f��z���Qj7n|z�L��kO�� (`-:��!��^�8����O��\{둼��y��T��mC����UkW��r%�} �4Z��h�� ������q@��h�E����E�J�h�!���֣�z���a�����宂�N�^N��mI��r���֋��:��º��d�۹XAQ�9����Qk�&����X��[t�����Ӕ���#�N?d�����Ϯ�Elm��w�t��Y���6�yz0 ��;R�� �Pk�0��P��*���Rq6�kӼ���\���^����3��A���'��A2k��jt9�;�Ǐ��pL'��nt�i̚�Rm����?t�2�:%\g��f��H{�[W�������㔽g�� �G�~1��a��[���~��q~$�J���U�y���T���L��v-d$�}Y[��n]���j�R���0�~SF�wm0�0���>x�Hl�)�"� y�<g�q��P�c�v��γl`�99d`�ߗ;�cƆ�����������e�yvrL����;���)H���^
�4e���cG�BTGW��≽�Z�?���k�D;Ʃn���YTE������S2má?U�e_�yf��
"y\o�o�x��Ó�qW�t$/J&HX-�I4�^t�b��Se+��V��FH!����Κ�1�H�Ta

�\�^�ָ� �<�����Wtʟ�Q\��b���Y7r������e�6���9��h�9��|������4�*��y�l�Դ�'$�8 ��L-e8���\�b�N��L]�SK�!�[�uW��s�-e�Sc�T���Z�^!(1�����+�h�>�T�|���o\B�{h���]���򇫛E�C����ZrY��1+��|�{�n����$ل�T�mjY��1��I�fNh,��d�(�,˞��<�1�պݼd�h�sd��'U�jY��h�[�<�~��o�C�/J���$W��q@6���l�jk��KD���o�1v�E�b��$(��n�7�
���� X�~���o�0�mo�ۑ��g�x�'0������GE��8;�3NҐ���\b�Y	~|z��!le]��y�.�/�	o�̳�&��}N5T���s=[�S%�����@�X��~��ی�����&q_�	[ڸ�z^�zM��td�3��	��Ii&)�Ŀ���,�v]7i�պm�h� R3�d���_5�!�0Ysa�`@�H��)�b�����l$Ў$>kF�-X�����Jb�e6�l-���y��,"��V\*������M�d��)B��idA�x "/�3���w��2��֠4	Vo��$��D4�"������I[ǿB*�q�Ӂ��
U]P�	��Z굲���.��ق�����Th�]�s�l-E���P���l���U���y�(M�P�z'���q6�+�ǓՊ�/.D���K��I�IJ��Y�p/�p���ڠ�:#��յغ%�.?� .��P:��i��}b߷��ڰ�kN�]ߟ��?6�95� �4�-�J ���<:wZ
S�,�D�?�-dm�B��R���j?��~f}��G.k��S�hj�b�3h����<g�sh��͵��p������u������v���|�>�(~1{��>{�c(��puaǐ1wY;y� ��%�pU��c*��Z��چ�4
�ղS%n8/;�V��E��Ș��W��{6� �ڇ�"^+�6�U.��u9��t`J&�m���=] `s�4F��[�0�0��d�Z�Օ=
�cݙ�l�b�M'��A���'��R]����|^����.�Y~q�R#Jb�]��5�{�>�s'�%\���(�
 �RX%�	������@�X��`񾣀���.^���/h�\	6|1*y�(xna�x���,.6�q���z	~�P��fk�eb�� �ߌr��4��SD�6�����w�������N���b T`J{.N/�l��2�dk��f��^|�R4w7<
�_���n�g�!y�7п��{y��+�=it�X�� P�DX��2x�H�7{��xr-�#�����R�S�����T�����|���������Å��~�_U,�
����cu7��ȋkY�g�p2�lq$وR�z�97�+
��R�Z�����Ա�͂)&�1#q!�NR@u0"Jބ�t�y*@눎ˋ�1MK'�|0KA/��LS���Z�X��/�#-�љ5� tt�����@c��3X���-Ma�e�vG|�hY��\��H抸�$ ^�Φ��>�=��s�PjU�
�����JsA��&�'W�/�����5��]>�|Z,�6�,��Vn�:]�=ާ����s<W�>2Q	��E��@�d��P?�y���Q^�����l^L5����t��VM2S��N�R9�D���e�5�MJu�����-��U���L�9)eB��d<tC�ކ���d` ˞P-bUqIAR5�^��?tYwh꓁Ō��A,_�vZP�IL|1@���ue�����1�U�0A�������%�a,��$q�ٖ��ʋ��$�ˑ-,�e�n+�l���xA��S:?���Y�����4UR��2㹰Ȳ��������\c�t/.X	���ɖځ�)�ըT&cRW�F���6;q7�~��Y�b}�~D�����?�6�|i#?/�~Р4++�ПI��0�L},��Q�\���䬍��k���d��p2��s���L�3������ �Λ/�����DxȎ�d��F!0dC�I�D������?ܓ��ɏI���Q]�Vb=X!pyqN�|������1�����ZcK��ʬ�ɷ�h��,2�o��̣V�9��� ��&���r���T!���@cY��uL�'�I��!����*�z�/ 7��)�[�/.�@����3�,��{�9,J�	��:|u��(��H�*��V�5���&M�ފ�1s\��RڊN�b��5��m���F�%7�7���%P�fH|2,�a_M� �X�l|�({Œ�8�v��ϩk�k@�!KTuc����r������v�տ'�v�F{��A���:�n�`a9��($�5���ˮCl��W�`�e�}�'�k�z h��`��{�&�w�_��"�
�xS�	5*���O3�x��ƽ�O��Q�_��RX�p�U �����Q��Zcϴ���������A� s(�����l�̹D� ��=�U���g1�	}i��y��>��,k�i����<�~�M�+i�]̡�J�h-F����x���Q�^;���1�\���j�i��Z't�l��x�~؇2�T�H��V�'|S�$�G�nm�p:-����W���Gc�j:h��
�:s��F�"!@�־d9�J6g�ZC��5�K�O��G��9[���+:;;��oºNf�uk��ĳ�+:.���t�'���2���@wtl<I�\m.qL�l%3,����k����P+��F}q-n���>���F8OO/Ō�A��6Sn���u�UH�#)�yrv.]��;-� ��d��);�-xX�����?�y��5+��?&$�̅3wA�@@�on3��9���O��$�j0*�H����d�M�pc0m��6�b4��AZm�ފ�@P�L������u�Q»D4�G�����`��\!-��2����|)LZ�_�99�l��@P��1�m�ɺɈK¬��%g̤>ݬSm��n�;���5�h�E��ű�<+8�`�y������
�&J�#M2	ϐm!�[>*��nY���t_U�X��|X������I�z���n;��;.�hɉםZv�抛Z�b;�� 0�h�ڟ�c�@/��^w��n�ܛ��0���bl-���뼇�Ly�*�{�;��P���������e��s��k��Ȳ���h�p�,�Z#�SQ�0n�3=@V�S��b�8fs�s�q��,���|!�7�yY?}21��%kmk.�lrn�=b.�+	gEZ�%@�XR��d���oT�#~���x��%�v|����Y�S
{[�c��ٺ�9+Y��Dak���������.f���lf0M�
�� �˓_��G� �|)���>B�<rپ���ޗy��1g��	ǧ���w��C9�� �>P&A0�O�|��R�5n��b2�{\JZk��ɷ�җ�9Z�Xv���n
�!~U�	B]�n%nM�#�4<�]�]Q�UN�E�0�tJ<'${G/���hN�#`�ӓ�I�����mˡ�l�����
{��9k-pY��Q�������2�k����οbqZr�\7D`I�7(=�E���OZ�N�������5y�³�W�0~�+C��X���..GǱ�P��z/° �W�^�P���3-�'$W'y�Ç#2��L�^̑\�[�i�"���U� ���M���y�s0|�y'�-��?n�_����!�[2�$%�F�����q�=K�fY�bؒ�[�����..�a�U�{}>`���t��s����*`�}�����w6��=��uD��f����O���7�A�^��1�݊	��Jd@��po��y�:7[��xL-Jp9�U�g8�%�R�6f�?-x��5_�`M�fP4 ���T���}��s�<���Y~sk��;�����d�V7��<�`	�k��s��
Tjb�����,�?��ЋU��F�>���<�#ȴjy��p0EE�u"�,��UVK
W�fQ��Ļ��74c}�E��*�L���FA��vU2�dWЬk�3ʐZ�ހ���
��d���l.>h_�2ęʪ�覜�և1g�r��	dq�s�� ��9*��������=�aJب\��CTu�}���$�n#_��8��-ǀ� Yɽ�vq�j�H�����`{�RGRa��I�2Me�)	�J 1Yv���� Z�x��(Onz ?ןb�@Q���ͩ}w/�H<�6�r���j &s�p<z�]����ޕx�h~��ιn��ެ5�i��jm}.}ÿHY�Yi�B3�A��(���?l���q4�����O�D~2?:���7ᬛ��{1y/��鬀/q=����C&36�a���
�L^�����v��|6�I���$�E��t�S����1�;_\���H��9�J�	�eo-&�| ��9�[\�VvM�V۩v)�f�n�D��񜽺;jM�+G�����j2`�wVj	U�YK�;�f���=���q~we����,�,֯�/^`=N�;T��!��iM�|�XdH-+���(���\FL�K��P�O:r���1`���� G028��H,��:��ڑA�����b�{�j �l�y���ѽx(�(Z� �Pj�a0����p�}�c��ϵ���5Z)��_|����	�@}3� �[79T��J	EN1���驌=���ZR�����9MR �^�<:g����3e�3�ղT�B���Y���`����`�`��wu+��lBy�d"I.�D\E$[���T������[�n�K��W��y�X� ^]�����]����fc�Q*�"�%T@�BV�6���ip.��x%�xsH�ݵ�#����3=�������W%L�Mf�2�(Y\�����^�S����M�sOϨ�yf��U��d�F�jmO�bMڦ����C�P�
~F�[(�������CO22@��~��08�����K9�i�XJV��4��'�T�4⟝0��i�ޙ#�K��RP����x0%����ԜqN���t���Y��=�S�gY4���,��	�V�5x`7�|a�"��pvB��Z����f���Z��}��9���K�4�Z��W�Mʹ���d��+�/E�3�h�4(���K��`M��"��q�d�l!�M�S����)A�3�)��F9Ȑ�����
�UCc������� ���9�͈�~L]A�F�@�e,Y�Ə(��7���hB˞k�|_���f�	h�̑��t�c�ژY?9�/��.j_�4F.1Ç `��I7�M��GXm�Q��	B�AU��!���ZgV�}h��L�,aE�GNuc����.�����V�1� ,Z���:$S�ʉ���O-\���Xh��з1�)����]x�L�>!�z�F��^����f��K뾜Z�Ϟ-���ې��B��Z�����M�z�=b��L�)`V�@��k\^�l�`�Cٝ��Y�,}��QS׈����*O�H����֥�EQV���lb���/Ǎ18�&WU!�>��"�Y��H�Z��H��	��Q0 ��	��������d�]Bk�wzzBr���]k�S�.,'}�u3�=�V��>���l���_<��F��>�������)j��?=���A�9ޚ��e���SIvZ*�
\� <޿���" �֯�������[���],�� 0.;�^�~����Iz�}�?=�_�&mOur,��q�oi{��[���+�&/rPc	�U�f��T�M��p)4��\@j:oT���aB�c�.�7W�ؓ�J�X�(���z��oإ���e�D��oHM�r�5�L*v�*�=Z��䈎�Ex�;���l�T���mBX_�Y�qi�L�.曑�?q�u�b��67̵h�v#4\��-o���l}1_�0���Lа�<��흟_�㚮�ot.O�鈟ň�\0$�W�Ko/��1�	���WY�����M�h�q�z_25:�|%sA�����Q�_�}E�����g`��I	�+:g$3�@7�T�~C[�uY��7(}w�O��7V|���@Fʬ$�+%�4�ר5Rk�{�aݕ�g�21����U��1j�ղ�t|P���M�pY�
��V*��JBj�hW�#�<V�W̲L�i|�/k� x�Z����`�Oiʲ��)h��2�j�B���~B�1�.��f\g�J���pc|,Mlݖ��r�O�����=���΍ָ;�r,������H�!����ov�F S)5�:���ٺ��:Y�^��2�5Z:+�Sy���I�[L�r��J6���{zz\��3���/ZlL��K�<0��X[<b3{�X�q�8ޓ�9K�ūI\�J�77��WG���մ$3hR�*��P��As�`�ο񘊫��y��wG?�kn��?�� 2���_*�h�~�������y'_�tq���٥��*M�c+rU��]�F�D�>A��xV ��Yx���-/CB;*Y}d���~ϓ���n}�.�KK����K6�r�d�p& l!��
��!&Z�� ,�������5�0��kof;b4��R�R4(�y0A���uJ@�����%�l�Nk)6YW�QA��Cj7�N<g�ԫV�VK9q��L�����X��QbC��'�r�#˶<ԁ�#T���9L0�Ƹ����|�$�5�.s����8�v��փ?�t��c<~#�jc�~�;��G�P� ���w:��k���t�@��\�C��V���I�._�Q�,���5@�����ld��l�2+�0.ow�BMD�\�B�^ޞqxE�@�<��  ��IDAT��[`��X7A @�(�AQ;��%�̭ŷ=�@�=��3^A� _�
�E�G�תւ
��R j��ȧAp�=n[���>}J�N���-�6��&C4���Vݺ�X�N]i/0�����|�Y�&�vmD��=q;ڳm���l���Ꜩ�u7�^�$�T�ީq�ά�P]/�:	g������:/���� �~�Ϥőu�#�V��W�����<�AQ�ʽɁ��XϓNk\KK�)r����S*��.0�tH�3��Ý��尅h�8�]���eg���ϧ��'��u.Q����Q	���$9�f[���#� z��>;�ts�4�:�N.$�J �|�O�ﻱI�>���>�HzS~����Ř�dq�=@����0y��0d��g��Ж��e�778
v�'�?ҭ-��:���V�_A���!<)�Å�j{ִ}���v[��+�x�����Ah$Y��%3�<�tI]~�<�B�2��Y�����	�J�������e�n�ڝ��j�0����p'�B�Uڲ�>I�-[�?�k@̰�z����W9�A|���Z�c�x��=��Ӓ�v3�0�d��@���A���ފ2:ئ4�pݧ���<~`kV���J
��S�]6K��3 %Y�wb������&o߼���|G�T����Jې�"�9��ܧM�<,t-?�++�=��(����J��4�i�5 Kc��s�rO��<<<ێ�"�k�	�K�	�O�u�qX� 7��vM��Z�\�<4�{��4lj��5��xm �}���-�������=Ԟ�����Ek����B����~�ңŭ��}b�E���)2�	'x���3���~��h�~�L{}� ��d�q5�s'��k�'ǰ��i��Q�a�^���/����n�~��-���ӬS�$lwIc߸�.9��.f��e�s٠�~7;�� w2�+�j�uU��f� ��v�Dw׷Z�����eM10a�[����L��-c�l'�Jnݰ�����A���(�ɿS-F�S�_F�:��i���������첸�gF�T����)�G���1ρ��=>�^`�צ!5*ն����e<`���-����y�%��ZU�Q�0��=��n�W�cna+!�.�X��)s)���%/ޔr���x�I6foW4�>���4Ha���.Vr2D�V��P:{mq>;E����ͯ͋��w�j4�~&��!`�,D-;#�D��>3�w;��T7*� i����'�TW��ɯU�{�k� ���<�\
sj�.��>�?3i�E ����g�U-�pA���x.���w������_�+�h��'�{��� ^"�d��5f�f��ӧ�����|\�V�� �Wo���� �}u� p����,<ާ�X���h�|�qH�hG�|.��Ak��p�_'˦�ᦦr��B�q%˨|E9�ْ:P0`�jU�nL�ܞ�=n�PD��rn���CM�O���nlGlK�s%����x��3^g��0���O�#6(������Y���-Ʀ�g��3�ԌSt��vo���h-�ƪ���ذ莔��cv�/�V�z�,]=|� $uL9L���o�����N����)�0H�,��\�m^�[&�d��c\c����q�ڳ��K��v-�/Ys�9����z{���"�j9� xc����uB'`<����r�@߭�g	K��.���H���U��{F����������c=��u��T��o�f�sV[u��.�5�����|����%�]�ly*��<S�߮���I���lx�(�!�O�Y�/�%l7����Ќn��k���ɼ��p��)��-�������kg�zPa�P7�ɽa����q���Y�9�*��[^��������'p"��v�(�q^9�1���p1�Pw۲��C��`黂�9�MG��mv�N��:o�D�h~�b�`�Q��xM-yĖ	�!9WF`,n�t���-77�5Ygϔw����[���Dן?Ѯhf\��7n7�6��$ F3\zu�B��Y������{ט�g �A����@%JR�D����2�|���~~O�
 ������]�yG/_J���`K�n�?{Zr��s�щ�; dR���ҲB�e�q<#�v���,�A\4��U�̞��ʂ���3�}wqyA������/_詌/ߗ)H�������d����F��,���E� �Ckm�=�^�s�@����^t3�6��C���r4m���L�v�C>��5l��H�0i�i��h�� ����#~g�U�a,G�>��S8������?fh"�+�	i��S6��ƫviZZ��z�|�s�7�?�x�:*��5��?���2���/0�FF�dɟ�o�/?�L?�����y>g��W׭�K���S��Kao^G۶P�͹�[��xd��L�Y涉*p�G�O�h,V�t��d_~���TIY��s9��f������A�.029볥&>X�Hr7�3G�� Z�WNl���q*s��&1_��6�1b�҂����E�eO'"p|�$���*cuvvEg�J߯��`���65�9���bY�e�ϡ�e�:�G���^�I���K����5G�^���'��%-�R���m1~hc��$��Ww�5�uX���??@����3���54Hj��h+���2����Y+$QΥ�`l���Ԗcg��6ɻ��
![��lSIe�j��1r%s��N �l|;��P��<"0����rv��Ņl�7e�^�����%0�߻���\g���8�a����Cj���}��7��w7�i�.`�t/�Wbv�FU˽ư��r'�?s���X�8����wS¬��y�PdU��~s�gl�#3�-��~gZC��9v0�L@���<?./���Hk�2�b���wo��:>9.�y+EeY�gK��ǟ��W:6�����2QkR7����r~�DP���Z������#j��_w�?�E'~Ǉ�0�� ,|wڞ:���~�]7�~?-؊�}��o@^ �p��g�����Mi1ಌ|`����t횹#�f�.���B���x�l[ۥ�}��޽{G�}��Zu�D�L]�k)�|C?����g�����D=>>�� L�խ�V2�.p�}?׭F�p1ǅ�kt�Xoqg�,̡`i��_���e�W͊BϤ��L�tZ���F�N�Y�B*[����awz�@qj7XW�[�v�ş!��5�x��o �jqE?X�ϝt�n9�����#=��4?��z��|���ruA'��\��_���5w��2�>Qģ+��j1�V+���7���d�K(��z�:L@]5�Ð��%ٞkV?�s�N�c�ά ��V���X�=zLǉL���YuΡ3C�6À��'�+�6ͮ�Ŋ��V*���z�f��f�- ���D9�T�
p���FdMuf*v����l]ه��L���e��<A$��dH����"Y�D;�mY�		�EK *��>Զb����k�)B���˗/J[V�|��n�e���E�5���f���
n"$4׃ 4�C����` ���9fe�f���O���/�����ɩ�<��������h�B1�?!��y��-��'����g:��^_6�đ�]��H�g�����<�����V�}��AR���_�H����b=8-`����c?п���?�(�.K�[�Z�Dg&M�8+ϗ�ِ�����nh@�f�N??D�0�K�#2�����nz����M�?E8�٫�{M�ۇ����s���H��	p}a�V����+��h���r/Vl-�@M�L�J����U-�M�(8�7�*������W\�������"��П���o������(�l5����s��r8�(�LT�]+����!����k!E�k��W��������c�Rqz�B�-�N����qS�t�tl�񝕬+��\�r��nb�������l�6n��kgd�'��{��F��4,�L�2��<=�񺗠���ۢ�mDn������� ����)-��v��Dϋ�{"n�� �Q��?][S6���N�>2p&w����q��V<w���t%Sq��q���qu��qH>�|Zg�1�C[�Q9A�C�V��~.�ő:Bڪ�S}X\�7�Yc��@��739��̿)@���pUdo�uRTf����}�X`���}_ a����Yeе��"KTM�
>Y��Rl.���,��O��R����n�@�e|,�NM���9��C'�$�+���gBO��������	H�ge�����f����ýf$}��QHWŊ���|��.^�f�cJBC�{�n
<Wnޭ�]cw��Mg�^3�Rg�����Φ�v2~�L�rѩ�䅜�\��Ynd<��u|�R�i&�Jt��L�v�͕�[���I���#B�"�5K�C�}��d-�s��m�;ټ�fn>�9�ύ��N�}
آu���Z�ة�r�V����-y�8E� �	 |M_��ٔ����i%�,��U+�&�F�[�Yǣ�Yn������5��/?���t,%�z���R��_�������?�D777B����Fa���5��-_��{{ؕvIA��Or��)?|��P��>�?�@�W�DX��kaSQ�-��U/�}7t{���noi�ZP.}��Js�hQ��;�j,���a����2�̓�*���{��s�&W fʙMT��IM�_��6%�U��q_����_�'.�Gw|r^d�k`G��e�^Y>v�T�l}r���3�3&*����S}N<��6Q��:֙%)U9�����XA����q���S��!$"�b-�^0�����No3��ۯ�2�]0Um f����f�`�T&��̉���c"����t��R��;����Dm��l,�]�fI�@^b]�u���]/�/�L%a!m$i���l4>Ok��\;�{�2�X�%j�˙D����;��`s1�h�A�R��Ġm��,J ��"4uO���G@u`��z=�u1Q��:�@���dfI�GsmI��'������y�{��5���;:g����s�r�����"e�ɉ������nJ�U ���8 ���~�����D3�8	�g���Γ`���ap�b9{����O
��{��ݖMꚾ��Sy�����=$]�v��s;Q-�3>�d�"ZJ�ق���Z�"��׀�^���@�y?|��E�X]�Gd��x�S���>�އ@� �W�����<birOX%<�k+4����;��My�p=P4 �����9Z�9�\" ,x?���Zzn��R�]�"F$q@c�qS��#���:-
g.�R���cʘ�~z/��fU�t�>���V�՞:/�%�;� 6OR�r)���~�"�����wh�7Q��EW�Y�*�&.~y�����{zx��������ݻoh�\j�1[i1M8�lyI
@�[h�?J��0��A���RȚ}��q��>7�
Ʋ�C$�Y�;�C\no�~����#��q����YT��3:�|I����WE���~,�02��n$Ӡ�: �s����� ���X���+��yu��T�����=�@��Q��`Qt�Jj�F��F b��Ҿܚ*���ͼ>�9b���E5#}0���)�x&;Kt7�'��ݏ���Z@��!�y����NW-|�Ԯ�~>��%�`��ƈ |��1વ���C�/��48�K,�s?�ވK���ǻc`G�"v��*R{�y�}Q��
[�����'n$��3��R��
M+�;X�`�l�N\�ys��>|�H�7wjN�/��7����o���c߄��uK7�ڤ=�����g�� PJ .VAʁ�|�S(��b	�*f} �kf!����Ef<n,��g�~:=9�2F�?�us{��e��Ȗ�(��a��E�<FK�=0�4�g*j����i���/��OL�����?�0:�Y������"���j}�i�R�vNAY�/ܾBb�|�	�������!�8}�)P�7wN�a-H
B<�H�D{�غy����0 �����2_9��cR9�d!5vI�x������V�W��hk;:��`�b�~�)�x�J�Dx���u���hn�d.�����2��/y�䚻��x��t~)�����\�+�7�;<�l�3qM����Z��zC��oF�L��^�ͅo�r85| ֜��c���%Ŵwr�n���/��Z?���Z�Z�X��Wtrv)�_�4?B���T�W������5u����T���6�(�_��x}�=�{Uc���������hO(V���`���踺��A��?X{T�)� � �F�!{aI�Ŭ��}>�jZ�����%;�2��a�l���JA�������=��R��`~~f�\J�`?�Kɐ���k٥��',pȔ��+��:�mӊE3M��˓����t]6�?�H�E ���ۙ	B�q��)�*l#�'��~��Сж�~V5M{b]Y\Z�Ae�v�O�X�l��|x����������|�{z󻿣�WZ��y�f*��,,�h�a�㏘� 5Ϫ �� ��s[�>y�Dg4!�7�ҧ"��ڤ�:����N�xN�^�{���u��Sk���������+)7QG5�Y�DL�BL��y,2� ������C�?��fj�I���M���q���5���Z�TY9|T!APH n��.!}�=�e)����Bc��=�R�.��1^1�����`E�A:x��}�%.��������pr�N���C������yvf6�<X����sP2ǀq&�%[�%�l��DB>�vB�ݫKQ�W�2�Y�1���{>�^j�MX�����
pCKd���@�1`[��<.�����e����Ï?
�?ן==��D ^��keJf�V��a!I*����l��vtO5Y����e�^\��:Z�m��#�>;������
����f���\���<ۋ��'�/���{,syO��(�ch�l?��i<n�@���o��}R�3�"W��#PQe�F;�;`�������X.�!���kۣ�ff)�.�*��ۑC�9 _;��)����k �nl���,�$�c�?��qk�f�:��T���$j&����O}��*]�ˋS93F\�aS��V���.i�g@����O�lө��m0�	ћ�۲(��q����,��}���%��4(7�Sh?�s �ge5!��{8��? ,�8�[-:3�Yؖ�7[������/7w���z��w����|��Qnbӻ`�c�]A�Dp�V�*��!$���׹���I���KـT����_�Q(6�eC�b���?t��(���b|� Ѯ�t�T&�@A^D�\�+؄U�����*�V�{ h�G "q~탯�̺�{[�-{(N�����1T[N��S���r�{p�@A��j
ھf}C�Bs��Cֽ�� e��ѽ	��p��F��Vp}&��+p6�Ws�����.��m����-{��}ʽ��<朱<l�H�б촔�����;67��حO��6~ZO����ٲ�eɌ8�������Ky����sG��^�,�����Y��[==m�u-��,.���Q�����ڐ�V~��M��h
��ϰ�;�!r�Jo��us1�}f4�5�y�x/VE�T &��O���5�c1���N.^H���啐\'㜬�J"8'LO�>i-��P�kvV�Y�xb����>(ֵʠQc ��ǽ��=�����v�>Ρ�7KW�,�����^���P�8��aZ�y�Ȏ
�W,`��F�"G1ǥq���2Ӷ��EAa�PO�lu��ng�\M؈�Oڞ��7��1����Ó�!��lVk�\�3x�j66JbYP^>].8�f�p�9xB�9������z<��%~C5׬\��L7_N���_�h3�9��E���\\`�P��R}� ��ds�@B�F�y�]����@v��Ŷm^�����In�$������yp������7��������i.��LyUd�����	W���>e��  �<''��X���ƽ�����;&������������X���bq�PF�2��*`sT�-!Һr��>�T�)��1����s9�o�Ĭ��k�n�����5��$��x�R�y��hׯ�G��-D]�+Ǝa���iA�n�m���H��v���/U@'�B� 
����:�C�Jy)��1�*Z��X�0& ���)��(�eY�,Y��Y�a��$`���PQ 
�V9J�������L��w;%+�:�k��ӢٝX�s[�#'�����8Y�[��xXY������dRJfgO��}��V��-��w%���h�+Zl9[����t��!�RW�ƅ�b�����A�@>La��$.��39@�6�����RH����˜9�~����?	o�X������Ǒ�
�S���;͒ո��m������_9�:�T0��4e���3	�N�ĖJ���p[-+�����q=΋��fs�g����$bO��@q�n|Й�R�u��b��q�7�e_����Y'��U�/L����WG�[3�����ܫ���/���|�I� +;�ҡQ��6�a���@ /��j 0S�_,��;- �����U�b�,��M�:��me�[�^��F�M`�M�:����C:&+Ze�O�̔�K9�f�^�!�����]�&��ϢE�#��Q�����M�ёb�Lt��cez�鉳�n��g�	᧥tKOga�	��� X��\�C%s�"|�!�%;��4���+k�� XrYhE����_n������⪧�/���~O���]_o�&vJ:�V{̳JHGm�>���Ӷ�9�}*�k��y�H�b���쬁I�HA�����Q�.V��[�<�
��9e�F���`ZWK���|i���[��G�'������ܘ�s��쁃�פ�#B�Y�4��.��ς�(�C.J��٣:�rMʮ�R�#j�.Q��N��U��z���k����>b�rc%���
�PGׂ�nCp}�����Z�"A+o�(97�Z�BP��;ps9�fks.J�gS5�C3��1@�~S`��<s�	H����kԹ�����T5:����;�ϸ_��Ǽf6[Y�,gh�V����GX0q!��<�*(���)�<�LN��z�����8��d����� ~�	 ��[�Ebƪ��Z�TB�{��ֵ���/�,�P�,�|g��\���(?5�{T�')����ʧ�/���N/^��z, [��� ���iw��S߬� Jr
����ds����k`�77�Y�� ��(�~G=��Lu.M�=�`�LuJ�i��ߦ��9���b��N�٘%���0�QCP���^e;/�ԛx�G��oĿ���n�뭽,t0��8
+h���_��F!�V#�QO���;��X5���ߘ(I���y!��5�D
�Fj��Ԉ �6���&����hF���v�LV;N-5ٟ#A�b����'��f�-�nV�������|�ӓ}��x�,�0K�8���d]Pj�Q�1-��� aɹ���խ�5V�Z��n��ǟދ���ቖE�|��^�~O��~'a��B���kTN������(��l�ٲ�{.[T��f����eb:��bA�@Z4ޫ>$��8О�s֫`@6��������g��T���X���
�B�X�:	���e�b�\`�YIP~�L�gLA�<����D��!��(幼-"�E7��p��c���i���2s�/P��c*���!@��O��2se#5�M���Bmq	�B�1 ��o�0)fY�h��Z����v#2x���ub�#�>�-yC݊p;����;����5+�TT A��-��eㄷ�L�47~?Sm��]³��Q����1��������Y����3�����N���K&'j���y��#����/����V�s��� ���T^���t4�D�v��1/Tj^�9L T01CN������	Ml�boQw:����ɹ,���(�\YD���V����\�iŕ%p]�>�]�x�sR��hnz�u�a��/����˫+: ��l�(���k����'Z���:F�6���4����86"��j	蚔*���c��lIRɧWk\Ù�s�M�w
��M����9��\;Uk[@�^)^�Y7t
_�u���e���>��f��s%c~v��)�V��Z��j��;K������	mM8��|lX��Fa��v��&o�-��%��)w;�S`ޝ�����ґ�a�C����09ExV��v�}�ᅴ�jn3��h�f�vbcE|������=s}-�IN.����5����ћw�����/��0�gs�l>x_a~y�5#�{B�>QDY7w7�M���V�/�Q!�Y2R���9D��$�w� B]�V� ����\���D�;7mi��f�֙����Ū��Ϟ̶�8��Okf�����f;A=�Օ��<o΍l ���r��\�~����㈹�w��j�~t�NK"E+����s���|�}`!���,k|�F$n�)�^;`58�@M�
���U�Zh\����X&n�P"�0wj�b�C��<��J:7I0�Ô�q���q4e�W� 8�N�A��\�6�����7��>H�q=K(P~q���E��Y�*o�?-ǈ	�V��X��R6N�i�Z��#>Pb�l��
��'{m6w�AJAS����q��
�3gT��,�IH�L�깰6W9�z)�_˓3!ʕ�c1ej���^q
�a�����i�����ogc�vUV�b���5}�tM��� }=���a<(�6����Ӏk�Z;SH�:7����'&��;C�4_jL��ԍZ�����]��5V���$8$ካ|�nw3�c�>��{]\ X��&�d/��L��e��
�M�s43O�2�(�1j��4�P ĨMD�Մ�s�J�{Bj~�P�`��iB�G���
�?,[�i���k�.�%,)3QH5N�o��bP1�����LP6�G�~��-������|��hf���tR^3��1
�$��,�n@Q���� ���@�s�b�ö+��i3З����,�ϒQzv~Io�+����/_�i��V��H���W6�>Y��=̦�[�B����ھD:Ȱ��]o�j�?2x���=��`q)�`��9�%9g���EP�엲	����n�5&E�����{a-TM+l6x�����/�����אn����R�������&O�nBD~�њT�'��i�'�*�}ؐMP�Y'/�V������ԥ�
��K��=�����ಋ������ݜтq�{�N�=�7c;bF#��sx�O�\o�f��4yBc� $k����e���t<�p��A�9���Fq?vҕ "�`�A7�aDܬ����-T�7O�g2z�8o��ImLHj6��̏2��k��<I���NN�������/����>]�d���U�������h��Ĳ?Ɍ
֫D��+}�v���=iu�O�~ۙkV�]�L���גeI��y�8�x!�/�x<.�K�I��d|�9�d�ɲsh��l)�K�� 8��d�r٧���2PᤀO�n�_>�#gh �>�֧��I���AwXF�"�$�\��ֽHw9�<bOK(���rP���h$�d����n� L�Wè��<��-4_����y�n�ԕF�pF��㤗M�Yg�c�p���p��0�U�q6Z
��{�K�yg���_���h����N[��๱N"��Tܽ+�&�� Q�588n0�irAk��,�bT�o9i���.�"����zG���z8��vE�KP�
�Y,��VgM�p��cZ܏A@UW�>�`�����z�L��HOE�~xZ�-�[��`Y�1�z����7�r��K����
�V�4�Mh��M��%�3(�ڃMo��p�"(�3QM��kr4�G�{k������,C�wީj6�\����R#]8������'Ԝ_��|��[�pXMLN�/ Z6�mz�$6� �5�6��J��F�EG�� ������!����� ��),�1�+R= >k
����;��EK�vg��UK��3��7`�{�c��<G�
�`#!�_?CLYo\ZC�G\��2x rN��,����ֲ�wX�dp�ese#i�m�*ZF�V��,q�w�(��}d1��C.w�x� 0�]s�БA�5U(8�c��sh�#gǿ�*%w7��D��X����cÎfK聅����9=�Р �ب�)�p��B���n��N2w�Fm��~�����Y�'Vp	���Z�]h���[�-�\����ޚ݇_����BaM�0�y�����{���}�|G_���c-sW�┪"V��/�s��j��	h��vAw X�GoY��j��V� C̰����i����]�w!�j���B�@A�I<�V��
��������ӱ�����#�?�@�
l�n��`[ S.�����Kfe��.N�.���M-�f���3h{|���M�1�?��k8�<�NP�������*�q���,�dz����Y��^l���0a+kfw7���������BL��/��ha��F�3�Y�\�UW��d�f�R�Y���p�s\=0���Z�������Y�gW����^J�����Ӳ_i��^=�+׻����	��c�����@AbiJ��K-`�m�te�Z��4��TP7����:q3�]���t�5i��(�	(�Qm��̉�O##d�J;�h� ��Dz��u�7��F}�C�Y-�.�'V>,��@Kk��*M34�~�Zj�֩���W{ع9��kf��L-��׾�kO�[�g���FȤ��[������ɪV���2$�ðk�ْ�~$d���z5�l��� {r�j��`Q�z����ݦ�����^;��;+��X��]dx?��Eni60"��tZhF�Ν�.���d$0�F�G;����ڼ�~�*�?���Aס$/���(�EW</oH����
���ϟ~���t{}M_�$C����e-g�&囓W�*�{.XS>�r�:�l�'el��<�KV��y�=�����9�uR@[��%����$i�Qa�e�Ȍuw���o��hzd�ϻɵ�=�Ӛ3[G��.	�������Kz�����J�h��\Aso�ӭHma�8��t��T���zԩ3�Y�X�I�^�u���SE�%� �;�֥?�������0-�r�0T#^^��f� !� ���{>jp�b*=��3���I/q�x*�Ҷ�Mr��I��dopu���pP�j[){'V�ET;$K[�!vޞ��Kz��J	4��O1���kU#�v��s�&�\����e����/��*�l��2y�L���KNȤ��F?�1[�9�������Xj���7���f���pW���v�)2�z�����GW/_KOH��r�e,o��Ԍc���>��:�ا�0qm#%K��f��Kȸ��ͨ��o�X�sM�"X8�X�Ac�X8�6�%��|��L@�*l��nEǶ�'6��'��Ǎ�C��*���r�Q7���N-,eS �~w@�K
C�L��*�DE��������U,`�yNA�L*
r#H��-a���Z��g��U����ش���q��ێS��UZ�M��%V�ypAg��b�J�.Օ�Kb 3೵�-�GBĺ���sm����#q��zg�_yCDi��``��y�n��*�f�L]G��V>T���D���I1|��t5M�=F��if�	z�,���i5���(w�q(���(��y�6��ã�w5#�{�g
:a̓y������|�?�)EV�17���M��RQ�y$|u�#s�i��/�$�=�.	�:1��������0��?�8	m�n�p��ġ��6��>�����T,�����l(X`����H�yɞ�d�^�`�<���
$o�W��5�q�Ry��� �`�F^3[��h9S�v�!��;��Z�MNa��X��<�S�%ָ�@l�sV�c�"���wA�u	��\A��۵XF �ق�/w&kkm�rƆ-sKe�׳uRf�0q�m���ff�'��A����ʚN�m�����r2dF�Q��Y�v�D��7|͢D\�U9����@xH�w���5ȊP(}ԯN�Xo��������R������d���{0f�e�J��el$[�2����f�ՠύ����=�l&�#������\^	��j��.bѳ*��l.���FS�W�0�G*4zI�
�&n�K�3v(v������䛘f��h٩�����n	�,�gy4��E=9�rZ�8�ɔ�+��Zfj�&e�d�sU7T�=�A���8��LF�t OA���t`�m�V:\t���@���־�L�5 ?m�
���X�c L��L�z�!T���K�s���)/*o�$�/����g/F:�i�=b�⫺%�-]��bZ�v��%V���U]U;X����V����e�ʣ�I�ON����.�l�ٹp�1 ce�闏�/���M�磀/.˕�E���")��҆N�ue4�D׌~���M���]�U�T�f#���%5O~K �&}Ρͪhq�ꋫ9�NυO����n�|��������3�sA�h�t�K��]��*U��I �S�ʐV����k�56ONhU���^��J�(��q��u�n�V��w�������m���ɧQ��� R�%���3��Q�SF�Ͽ�,nӫ�/��������=��lHi�`��>�ߋ�j�Τ��c�%B0o�}�#���\��Gb]&1�Шq_n���?ֳ�����x�Ї-WF�\l��yLx}u�=�B�lޚ�kj��@��;�S T�keK�e��l쒑׸5ӟ��8�eթُ��C�ڣB^Y<�{�.o[����P�E�a�{�o>����"���9qɄ� �yQKPF�гg\ ���@�W���2ʌ��ؗ���~A+������Ni�xAw�_h~s;@ʳ�ҏ����`��n��n������qz1Oy�s�����䥬sJ3�L;�xI��p!��E8��pp���5R��� db;p�u��/�b�;�ࣙK�q�9d͑p�,;��q$�<K]Jms��4ӑ]�ge�z��J
�UQ �L��Ge1�f��ǹ����S��@(7��֩�\�Ʉ���*a!�+�5ֿ�^?�{�;)��h�Q!<��6�pz�u�\54��:�� H��X�Z&H��ngE�'@&Z���V��6�}� �Mf������a�xU�n��p_3߶���<K�����&�dU�H�Q���q��Kݏ3_���o����`�X��������?�������H_��Ǖ;�e�J� ki�.�WkU���>�,e{���
V �b+@�=�W��b�l:�mѸ]2�k�.�Dˢ�����Z��s���B��m�ܥ���(��&kмdƛ�(�5�B6!�s)�!(��לk92���߉<�`�
�#����8O]'R�]�3i�N׹�����u^+��k� ۖ7>~����z#@lQ��y���^4�LY��s/k�Klu�V�>]�fe����LjX{��S�$�syzT�Di�����d���`:�g��3K����n)6^��]��}^y�OW����T	�%}�w3�*�h��kDY_�R9�,��P�hEL��<Q��qV`3L6�ɣ�H�9��8�޷,��yRM�3���Ӧ�`�_4�i\��h&G&�Dc��=R�fZ:(��M\Yx,l��&���4a��s�
%���S%d/e1b�F=��_K�̊�s2����]�]���M����&ɋ-Y�#�Ϸ<HZ3bf*AdA�����º���qpgW  ���0h�f�$b&M�WY���u.ֹ�Rj����͎�Tb!0����];��r��	_]����}����}}I/.���xi�ic�+z��]^�ͫ�����~*��{����n����[��9���
��Q(|��������T-K�Bk=O^|T�U��P�Ri����G����vѽ�C_�F��`���@��I����ž��`m?O�Ej�� �px���;s�������*�v�!��Rr�hVW\�b�;�}����~�Zһw���#}������G���o��������?�@��/�^~�H�|�B��k�d�{Vtp�a���	�$mkg�Õn�rğ�5�3��!SY�j�����z���� @������c�Ҫ[�P��+���<���J�ƣ�~�l���ҵT���3�4�I��r��.r�]�l%b�[`U�L]]z]�����XJn��=31<���=~H&�U�w�Tx�e�"�k ΎDYx�<��2g�����pU�?��U�K׏��J<b�2��	�){֗�s�C\�o�G�Gank�����7�9�� �WFfVfU�I�gzf��������>H�*�8�`k"�jf@Du��7^F�p�`�&�**z�}@V����H�
R�Kzt��]I�6{r�Ÿ���":_���f㣶�:= K�/u k�-�9b�'�}��z��=G{Y�h(1S����<"�x>j�������zH�o$�J.�u��c�:D\�Z����ҳ�+�����@�E�'����8��4��(�g<�Y���X�YxN�x�b�1�e�����ץ���|W�*��X�l%�don�Q�����1��
�AJ�׿�h��s�(r�ōɼ^��_S�fm�/�B8-$]�Zn�|���^���]͵'�az��Q��i
.Z�_[�J�l|7.d�u랣�Gi���>��MD�ݻ����{��)7���훴Q�����v����������k��M<�c)�{��f[L��/�Oy���u��7����x5pQӐ!S�����c�`�p��00K9J���xyl����,j�U�ḶV5@�s���W��Fs@=}�G�R����;k��k�\8[%�V ��I�wn�D�jY�2�.ƪ��*��mn����m#@�G�����(�����v��pO�ގ&��](B4ӯEi-��UM�l�ɀF�mx��� ���BM?�@�[/�q��6Ӎ��J��ytjO��x ��P*$��H���S�X-���ޥ��d�#Z��}��TV0ު�-�V{�s[��1�����33�6��)�a,c�v��,VXf�Wa@AS� �I���O*�߿�e-�~�hC��=\�0���5�l���a���k�]`>����m���s�-�t�U�z5-n�z������~�6���1�6`Og}i��gboi�3ϣe!Ί���r�v	�w��?
��f2�>�ѭ���e�s���77(m*��^���A<���X�|L5����P	��ʣ�+�$�>�` Q���m�=��F�K(�$z� ���+@fd��F@N ��Ji���4!�Xy���5.�4f�){Q'~1����^�4ʏ��
�r���t��5���!�t:���Yu��X_�2]����Ղ�=J�?7�M�����z�+P�Q��B,�u����*��߉z�g�����6�l�:,��^w&J3����AI�b?���R��M��n������{������f�!���0}�N<�8M1�~g�C�V��J��X��;	����E��M�����虈�:G��0�+b������ɓkkl��u�uSG��T�6��</U��z���rݵ.G{��i�li���\W=���u�$�*�'e|<�\�5��n������U���C�R�5�s��u�hYNUz%w�����-=���mڴ0�hD�h�r���9���
m�ǧ��Z�9�ax?A[<[HϹ�\�VEB+q�L��UE����V$����(s���j����\�?Q���<�肎p��!W�E�1P��kZ��^���\�ͼZ��&3��E��1���SkM��6�B+�p�����Q��v~�wZ�,z�͜�Lį�[����v��[q�r5.�Z��!�p�!���c�C���������������U:��ޙο�NVQ�˞�r�vV}
�� ^T�zs��Ev�����W1�}��!�&��G��Y����Y)��L����%�����4�5�)͑�,���λ[�	�D�֭t@�6�l3��i��R�c|�V��4���	�9a�c�Ѵcc$xm\l�ÅW���1 �4C�˞`x���'��
aX��Ff�n��5��P�D�)�2f~OoU;h����$�2��=E:�Hk�2�¡D�tF7�b��y	:uouƹɟ.E�B�����}s�g8e!*��C�!�b��7����k� �K��g�3Q(�$L�C�(�=�N+c���
�NS�.?�������<2�"�ڞ��̻���P1��`��rp�V�����y��"��y�����ӣ|��M��m ��\�x~9=d2'���{��y�p�f���|$� �q�����s��|浨�L�����U��L��ud���[5]Sz2z��ys��������ꈩ�악�<����g����u�"� �>�ߏY���(m��!�:65���[,���S�}o�%���>��#�Ln ޴|/@�n�3%	�9��1�B:Z�ͦ7%�Ʊ��3m�H7�?̖Dy�D\�XրTV������k�,�L���G}��/D�̱�2[�X���n�6k�@T�q�,�*_��ޯ����U��Tvy��\Pe+ѯ��;˟ِ�������$NG�qK5�Y��Жa ك��kC��q/�ן8o6�!Ǐru��������j�&Z�ў�*�nՠ{`��.�c��5mL[����T#�umO��kb\I�o�S95f�������H��3e+F�~$����7���??i��C香Q�A>ģ�8�v5͗�/  %�i�hT��c4�R��C�6�U 3�b%c�q�J�>����WN��b�z������Y12GT��b�3NSN�?�f�� ��Y?g�1�TO*h�ˆu��Wgל7M�*Pr�b�\�ɧmA߃W[���m#�^�j�;�g��[e���F�bvH�*G�*���j�|D2��Fi%}P}���	�}���Y���+����W�EQ�/i!��)��fR�Z�0�[���)HU=憗A��������p�H���[�o�9������}#� CZap��w�=�@�[�n>dS0T�y�5`��Rg�{�=�����gǮ?�Ꝁ��L�E�}/�N���#Q��=O����U��s���3	���G-��ǚ�G8��V@��4�F.�}�G��T���?/U��~�LǪN�:���H �p�T�;�k�����o=+\=��=���D��_77�U�m��&d����@�����*�vA�x"��;�E�!0��ѵ̩�%4ENs 9_���lI|Ŝ�t窷��w��0s��!�_y�b4�Cn6��f�Xcv^�B�X��aF�*ɧN��<V�IuM:X2�ffYᘭ3��|}��o��z1Z�Q�Z�"�h�n)��i!ը��H�qTm��<�g�v�M�������{�o��_��[��9z�B��.//y>N����]�摊�][<���~fY���/w6_��(�e�%��I����%q�ɍ�}��f:�=�����\\ݰmT��>��	�z��kI�N����@ Rj��I2��:U$M�;�k�%��bh���*����Х`�J��)���\4��ے4֒GA�0��6��4|K��G~��dy��KP�L4��ԯ�Lr-7慳'}��SL1�7"� 5L�h�J�0�(^F��5F.�}b�#z�e�����:��C��.�g� 8��p�
$��K�|k(ǝz�*�<��ٸJ��M��0;�"z夏��)���I�L9��7�6h��qWHط�v��j D{w/�� D�Ҧ����_~�ǇrA����\�&/��F�c�*�.)#������2�<"�NJ��e//��c>v9�z��~��>��1��y�x�Z&��|k��y�����:5W�3O��@L��X�W�y8К���s���ծ����ÿ���5 ���4�Zx�u�;�r�����qX.;ާ�n/"c�y����)c���8jqDk�jwO ��B�䅁��!�����Μ)��[��i�.�l�9Dќ�ހe�v�8nJlv��>_���~�
0d�[�P���eN�g�"���(�j�wv��d�����V;�b�_s4�J��� ^(v[�|�}(�q�~��z��W�Y�N ��>֛�eg�"�|��Y,$�P$u����ߘ��W"~{s%��ܘh��sp.�\r��\��蕠nbu\�������ׯήQ���q4!虝����
��~w� �O[v�M�Ǵ����Q�� T���r:�do`^&�;T0�2�i3j���0C�e�h�$�a�Z=��E
O<���_����`5������3ꬠ�1y���&�E"U�J(�m���5���\��J*X�0h�,���������9����}ͼ��IM�2Y��C���W�ʺ�!5a�4s�#Zї�< ��#TL]
f��k!+8��7���Ҹ��~�=�w�ş7CG\��*��6 �8��֟(�
Zt3V�DN�c���x���'�OOr��6�]/�\`�B_�р[c�ª�\�·��G��v=*�*9�Y$C�}Ѽ-�mh�����v���-�'\7j��Ƞ�/���؏����>�v��/�\q=����L�I�w�t�1O: Aħ���H�� �t$�E�#Hx�8�5������=x�Vܞ2qݫ���y]��"�ZSk �� ���6�EF������sL����XIr�8��s@Ǳh�����}\y�\���дmh��M�Z��.,�o��
��9�5�c�{9����D|1�`�93�0scc1/>7y-Mm�C�yee�;w |A����4��p@��)JQ�#:{����U;����Y�u�(�(/l�x��2Yl6;��)Ų�'�W
���;?���&����,�  ٜ�^q���-Ó���Z�x����ӿ�$ߒc�������� ���G�������$��R,6�LW*�uT!ۋ2���mL����s�^&�ɩD1�#����H���{��.��Q︀�H�n����?����rT�wh�p���w�O`�YBM���B+sc�v f�H�!1a���*%��eJ�8z3L؜@�g�����]��9_�\����J���`�ME�u�Eۆ��}Ǵ)�=�6y���+�z�A�qh�:�/���d����7u����sd��u(��nT�aڞ�4KjM%�q�_6��:j���2��+���X|��ab�&�h�3S21f��c�vf��+/�q[yg}e���8����o_p�U'�Ҹ/L�PE���|x��5�b$WnpQr�F�Vq�b>!M�j�݁�J��~{���該�Jc���fQ�7�ʣ�k:ʠ��_ޣ��h�,�{����Q'�� g���dc7���TYQ@U�1}��%�,R����ѡ���eHL�4R��*ڟ��U��:��E?���4%�G��T!uu�߼7��O�d}�A��s4��ő��)�
�<�#��Y;���[��-H�c���<\ثN��ƺ^%]��0qL�<-&b����\��Z܊H��G�*�y��c�&{�乖相���gs� �|��e&��e�<?�/���������������\��r��e�78�g 쥕�:C�R�$-pPq�E�e-�Q`�{�R1��������B�O��<����R&��]�>���N��^�A����Sl���r5��k�ն6l�12z�\�s�҇���:ѡ8��_$_�[FF�����Y��6��|��<?��q���d��;r}u#�����m) p hy$h@O'����,Oۨz�OJ���S�t`N���F�7CI��1BARt�JG h�ԅ���B�S{��#�>��J�b����Y�0��{�o�r����;y��o��@O�"�W����C�U\_�=ݠ���'~���Ѱ��M�GVq`\�V���[��Ek�
 ��ӷ�eU� �zrM��za�Ӱ��kf,�q���W� ���<�^�����[�����M&E�f=�ߐ7�ƆR�bߍs�9���V��xR��Y�m������H�K�͂�6AT����~83��'�N�8^x|~�0R��Z��0��R^n|ӟ�5������1NH5|��y��� �$��Rէ�=�ҕcO�����5�﹜����T�L�{s~^�����*TZu����Ǳ��y�d�����?[_c}_�Ƞ�=��A���_���&��q�k� �u�<�7?'���3��r��R��j� ��h���Z���9bJ�C4G�aN_ё/�汐2}|zN��%��zWM�ϭ���88rP-�2�8��^����ņ���f���-ǚڹ��kz����g�#ϟ��������s�_e�'�TR>x���8ZļD$���q�y�,wδon��d[����b�5�H���E{,�C���X����1ʟ��Y>}�?��_���Rnn����޿{'7W��I�e�
� Z��*娵�De )�ς�ن�*@�8�q�Τ8F�9�gM�6j�
O6���Q�3�_At�9�G䁼��-[�!��ց�i�v��|��[+��^	����$\���6�ju���Ϭ���o��֣���r`�h`�#/�曤�-`).�S�?��U"�|�tR0 Vy�=Cv`�{>�Xy���,�|���Iv��|�6��YUu�H�尩�$�hzb���S��[ɪ�u�/�����m�,?�sz�I��@�	�UX&�Ƴ�x]jp_B����'QeO^{��iRSf��������,����l;_y�x:T���^�2�DK�Y�d_�[�h�����6y�'ٝ.�54���k���^f�"!5a�}k� �bK����t���1/�b���w<Z��l���|v����@���
���z*���E^Aն�XZn�,�,cB"x�|ڍq�P��͔X΢\�s5߫\s��h?M(Ͷ=2�.`N֯#Y�c�Q)?��89�U;>�b��5�)�:��������WB:�DQɲ6<�Z ��52'O�c�j���<ߢe�}�W>�^�A��Q���6�L�p�mNOv���	r2����6$a�SG�����Z6�?w']_�Ղ��(�3�����0��������r�}n�T���3�9(�wޙ�l�q�W�����D/�/�r�A���Wv�?��s>OPQ.����:P��&��*F#X#��4oi/���0D/��,��o?���j���y��A�}{�H ă��9�Q�	 �9���(>]��3���Ӣ��b�=�-b��2��
f�,K�׌�p`[��{�jD����Ϩm�4 Zn���$��>y&O��=����l0��E#�K��~�'��;sepS�s�<���H�����Br�d�4�p�{Bf�{� ^��YުE��N���k�X��3�h<&��[py}-�~�k�65UϏ�vD�1�q�A��5���a�j(��u�x�1V�
 wi�W�-y$__koĉ�m��^]�B�Lɘ9?��ʯ�ߜf_���W>��{�����A�2��8P��}���d��ӿ%���z�.Y�&���)��a�������at_Z]�y0h?;�V*)@l�����!{�`���M�S6���ԑ��x����8��4�{���96"�"�$t�D�Ʒ70�7#G��>��l�X �_G6u���9Nv��ȯ��1�Ѕ�"m}��Ov��:N.w~V�
ȣbt<��#S2W�¸_%+=�z�_G�'�k�4�����ùk"��i[g��6Z���������:×h�(���<r`�y�P�n��}�n:`b������a�s�NQr�����-���>�2�d`hq)���'ӹ%2��������4E��'wk��[�$;N��a��S�XFS����H��>��#�|0w�b����U��f ,'�|������<v�Y�,�� `ph�	Cva)+���#��Y"�ɦ�N�=Z��
����3ґ����x��1B�P4�w�zB���*�l�u��&vʷ~�ot�>4F���!bvA��]D8��K����k~��@�4ʕĄ� 2`SP<��ɘ9pw�~�����Ŧ�Rxd���f�K���?�6�<�\��*z:�B���|�"�
��)'�Q��
�%@s8�5��ݝ|�� �/������ ���ay����U��qS��8#��-���Z�uP`?�Ӱ!���
��&��U�vQ�c���97'�:���+���߯k�\�ȫ��?>���:4��K7;��$�.U�kU#��Rr�o��H3~���ҧ9��#��{��C�D5y��ɖ��������+$�"� &�dM'Zwm;��rO��k��`�ۯ(��䱰��=���V6+m����֬��CI���J�K��泥f��9�V9>ql��P���_����W=�Qb����{^����Kz�&�ב�Z^�ǹ�
xR05А�5������{5?�:E\�e�y_�)��6�+9ujd{\z��|�����ȉ�R�Q���T�s-`�z#����d�К_e���V�d���$\����5���߿��'gz��M�W��b�9����Q�3?�L�2���;�8;�����3>��'�s�W�����W�?]A�b('����8?;�wVq�;|ww�s���z��~w82���p���ٜU���u�p�ҲȮѽ-��ߦ4;����Q�������t��t��Ѡ�%��)���MMp��v�6��P��mN��}Iy��6Qm�p$6�3�d�g�(�A0�Q�Z�;d��	 �J��- Ɠ���ث�$H�lf4�:�Λ	���]�U<�>N�B�p������za\����e�ϣL>����t��z�D����j��ait����B��Dln�c����.Le�u�����c�0���ȯS*#)�g�9���'\���+NLy�ڻt>LY:�D����z��y����yd Y?�WT�����/H6��dxu����쟽�%s Z?z��#��\�EG�n`��W ϻ��X?P|R6C��cZ2z���a�O����G'�Z]�㳓��Q�b>���EK��+�9�R�+1��jS�S�uZ�>�(��;K�l�_+��Yj����W�A%!��И�NA�HU	�;���&��le�Uuo��:��r�_u��� �F�Y���N�Hy�*�Ƶh-w�VDu$����װ�]?WWO�Ǩ���կk��?�T?�����j�el�Q�S�n��S��E���t�Xsy��� {�)��������9l�w�h��ŨE��S����3��7���aā�G����bM�=�� �2�-x�z~�נP,D���S�=~�8Dԏ�d���B�~��䐝*�*�_Gb�(��nc����zQZi�Ύ6��(/��c�Q��)ݱ�h�߿���FA�������n�;[ˤ1(�"Y$���{hM�^�;0Ta�r��D��1����ұ��4���.~��3}�z���V�F�ap]����.WP�Xj��Ф��|}`��|(�D�����἗��z$0�=>���#*$s��O�Bv��7SD4.��T��\�ֺ���e=����J�u��h]�lf�h�L�
b��k�a��f�R�<)�CV�g���Hm3�v�I��ix�!���b3��3C䎅r�M�׆�Z�q�y�iҡ�b�TD���!��
��]'kp�X�iI�>:���������+�U8�B� �fvm6K[�������n�P�wd���T�g /�)r7����!9y#G�~U�G����(w`��(u0z�+s�	`���FZ��K֪k�L�����Ʀ@��H�u�o���3�Befת4<04
_.���l��֢�Z����a6�����"���l���U�e![�Wv��,������+��`�D��?�@#Ld\.����5�k�j�	M3��Tl�G��Q�:�U��l~��ϼV`�G�Bi�*)Fo+T�v:�q���^
У8~�sw�6ZV*#��K~�������0��M��l�"���/dk��{�Zԑ\ɞTD&�Й0Z��Q���*첳m��� �	@�O�)��Ϧ:�U9Q��)��� �_<p�i��U�{�Vs��e��D�&���vKB�v�]lS���:N���S�$<m��v���!�k:L���׭\r{�Q� H�xB��z� P�?&GPH��H:ڢql5��r`Z2�
D9�VM!Z� ?�ªqw�$ح#�G1=@�j �"�pm����	bcO�.=F�b.c#H�B�Y�e�.���0Я:D�q�Rr���*\���,'�^�l��z�\�J�!ku-=����+2�6��D��9 ��f��֍\��+�Fy�kAxs52B��9�[�8�kY���tlpڱ��G4�=93�8�0�*�&cq�+5$z��F�*��m&m��fd�-Ej�j���K�yD�/̼k"9+�:E0���M�^]ԯ=�/4��T,��9��c��)�YE�\>�p{^~���{\��ÿ��W��F�ν/�7��B�����O�`�%'�G禱6 ����wsY��G-��!Y-r� �bi�l��F�}�A;��3H��>L�����W��F=��QQ�3�("n ~�po�H��<�~(B8�֤>�Kk��c}����Y�����q:��#��uE)��tf檥�XD���lԼz��fU�$R��Ȋ�)�~(�����Y-��Z��E-��M��Yۯ�b�k�������#b�<"�~�%�q����o��sp�m#n�d@����~l]^m���=M���x�1�l(�-�����`U������H�O�!$sr�e���؂���p��e���`�-S�)RR��U{u�Q��Ve`_��b툖���H���=�l���ȣں��0�ա�9������ZfG��ֿTd�^d�;f@|_Ҧ��������Ŏ�9�\�d0��6��?e�F�d@@w���E�"a�ȹ�\�C����t��/�zO˽�=OM����TbS���cZ��h@���g٦���Y�����:�}�y܁E�tV-M����gt�� ���\$�uA}I����c�TV���OD� cX0���@'	����A��6 �^#W�|(�����3F'}Ɯ^qC�{�hX';Z��W�P��o\=����E�*��Í��˒ 
Zg��wG������O�β�唍��^������fe%f$hu���F0xٺE�M?��ua걷��>(zԴdh��f�!�XQ��֍G�̛�ι49tꞳ|������Y�I,ϗCNf}��-�#����L��Gu��r��DBYb��0�#_��r��9��u�!�� ���(��v�j�Ki����ۘ#5�g����4���"Z�r��r�T��M����ao�F<B�N�4�_�?nk��8��u��)&��N�٬(�)OT�z��f��,��Ϩ�H��
@Za��~.y�:*S�ni��|�F+��>G7j{�D�&��kFX��c)^m��Kʜ6���b�ύ�T��Sy���O�"��$
U�yZr�����N����z-�׏�#T��V�Vx8p!x�y�"�i�d(��S9?���E_�������;y��-�
�E	�o�b�����N�PU|�����s@),9p��NB�S �F ��l��A�u�v\/p�I�E �)��kf����]����XN�57ux��A�VA����HR�����Η�iz���lp���v�컸s��)��~����[㜗�>��"<��+Wr�@�M7�̥�W!�ۊ5۲M�����Q�C�:�^<ƓP�w���j
x��?*Y�0�c4���n���k�Mё�Q#�u,�ejs��S����`�ȉg5�5��"��RJs��q!��g�a2!#@�,�J?cGXF�5j�/�o�6�3ى"i9��!0��\2xjT����	\t�I���kD�{�58��<���4z�A=T�щ����ߨؕ�L`o��|� ?�"�|�*7o.��j-k�5�F�2Qc�n H�,��ҷ�ǆ���ݼ�2�UWznk��8蝑�LƧD�:��U���ǡ�\.����T+�Yxip��@b��tAY�h(O��-_���Ҕ�e����à��~�y1R�C����� ��ԡ�K���* �D�\#�@a�˗/�)�kl0�l���L^@Ҙ5�|1c!��TJ6N��r�M����F޽����pϘ��\�U��=������C>�߾�wdʉ�\�]��2��-�a������L�(bldo�{Og �ϢC'�#�|�C�2��gkՆ�Z�K���L�⺺(�dh�F+85�{d�fD�{Aߊ.L��WUϋ���9׆�9F�ش9]'R����iW�"U� ����,�"m1?Ǭ]B�����4�\c�S�~z�9V��p�;�����$*��H]�tv=7�it���&���?�A�������`X{@rv���Q���_�����ϟ���{��j�.��Z�v�c
gR+20�JnW�^�Ѐ
�U�-�d���{�n��Ҥ5D�쾢�T ��-1؆ٴ@�s�s9cU��W���HL���Z�[��q)�
�ٲ�� ���Z��uP�u.��U9 �G�[g�qb!�~Fk�ǧ¶�*��øb$���p2�>�)>����P�Ȯn�A�h7�:�C� 2g�s��q�������u�8*�,�UF��,��I�{�9��y���Ë�x�bc#]����xz7���P,�~�lR���U�����NK��ι����4�p>;ǖ@u�|��u@�a�ްT��eg�Z :r` �r���"�Ht�7j:r����6Ci�<I7�E��U�ft�� ,N�	��= ��FM��ڦ�G�Q%�ҿw'a������[ys��E3R��U�~�7f�tӈQSV� y��"+A��|�0�E�N��<��B��7&�s2n��ʁSpT����� ���$70����ϹD��Mܘj!m���pS�O*^Qm�"�iy������A���-c�?ߘ6�䅅�T�P9�aZQU*�>�':^�`�������JX6Ⱦ�4��@�aA~R���@���(-
Q�6�QV#ߌh���W��J�g�`�	т��knd��}C`��O�?����/���`!`]<��(��%�)��	�qS�גD��I��jt��	`��W#^�R����*�z���K��6')#�P5��d}C(�ȼ4�u����tʃ�	3L�;�1�ظ�ZG�^�P�Z�W&��j;���Ԥ��V�S�����눹x��Wk�:uY�2�]���J����y��x\dN��5�i$���c�8��Q���~��0?�;m��k�����_�֔�Qa�46�$f&D+#�����B�m�
�-d�ਙ�����Bgr0��Oi--����\^������u&�ɞ�ve�x��x����ˌ�T�MK� s�(6[�'3���*���Z�/((B�Nd�����lӡ}8p e��q��W^So�y��� أ� h�t9t�,��K�ӹ�} `6МeDT�`��uo�=�u�<RjM�[�ޟ��do��
��J�䱲51�G^jK��0�� >*{Ei!|G4�����"pL���@i2�q���q�r{�}��cW�^`XVE�}.DK=v��.N)#]�aDZ)H R�>�OP�x��.f��[Q�e[z��q�.��V@����$G}�r����ӟS �[d�i$�=�F�w*��[?���N��u�ۼJguP�K73������X/�_2P����Y��������o����ʏn�j���"�&Rn)AlR%f��x��B*��'Q��*C��{bjk���[f� /��!2J�Q�9QY�ڙ�z��7��^w��,�o��5
�c�5jx��J�ί���@�	��?>���}N����6�FR�P�r����.P1e��Os��N���Se��X���.�X�1d�x��?"_�w��O?��o���>���;Y]�����."r��F��[�\��Z��.����+����e�3��_ ��w����&m\?��#zC�^�{���B�}��6����|��y�a�e�֜��{E��|)��7m)^q�4��������Q��&� _P*�Q|0=�:��wi4)���Ȯ��Tc�">p(%m�e=D&���1f���^%-+�Kd��+#kN�^V!��kL���	}~���ѯ���Wi�Y���j�KN��
��9�h��Cدs�i轿�����XzBj4��a�EOƇ�{�ӫ��_���M�w�}{K"�h�ݥk6i���"J�R�O��jU9ČU.��������?��Ԡ���_(K�$V�.d�Z2���Ⱥ���5�����ٞ�c�Z��Ta��|\:!*� ۰X��xn�� ���W9ȷ*���"6Ж]��sQ���f:`d�yA˨������(��ڐ�������r}u�q�������Cl~GO�y�4_�w`�mO�ud�[sDe#�T�~�21 0Y2�v�<� ��(O�	'�5Cfl<����-�h;�4�FӚ��7�-"tg�Z���������w�3}��w�(��2�	��;�x�B��9�v����q	aS�T��F���@����_�O]-�D�ū�0��O.d@zU	͙Z@(������G�6Y�d�c�2L�(�GZ���=����N�~�����%ۙ�52`h�����Aw5U�G��t�Y�����eC���3�[�^Ӂ�4���/	��Vӑ2Z��š 0'O�(�w f����ּQc^c��w�da��0��&�jĠ���UhJ�;,���v%�m�V9�S�g�|żert\�����6z����a
�T%��i �2�bm����t~���@$H�ca��3�k�u^���fDOr�Z=� �k���A>}�*�|�Ĵ��nǟCp�f}�� �aa͘��5�\��Z�ˉ�:��{��}Z�YwL�}���|��A޽{�+�ކ�����	R�Jy�r��N�/���jm�ͥ�qg�+=d�{��p:���i�$�j,�ҙN�o<�M��;��W�:	ڀ_��� F�4�R��*���-�AScQ�!7�cc��D�܁�#n5�J�Ǣ��ʬ�j<�XG�j��׸Z��b���S�u4�轅���bt � �7,֜J/F8�'W��5�ȬLl�4(R��?���"e�E%k���i�a�߳o߉�ƢJ��mP�Jc�{�qgMA�v�/�S;:f�n��	m��҆~�X����K�'H�鈞�vDQ9��m�^45r��1�W+>�� 5�h��,ЦZ$0�Xlԑm5D[ՙ�-G/ci�̥:�0�Ǳr�D�8@��~��5 F����G�>o���`@3���u4PT:�i����g��~!�B3�8*V�d�XҶ����*Z��E���7 !.��]�.�qڟ"ES��a,�&��9��^���<�I5f'��-�Q�<�l�H��n+}��̩�����Ų���1V�� l� N0P�� ""��6jdX�W��>�*C�ZD�����|�����4�;%�!ڂ��\ڤ#���Dn��*�$=���T��r�K�I�v'��Vb��$q���;s�mqT#$��r|ъYXȘe�����
�ҏр��Iv)��?�����||w-�4�O���Dg��6){��V�0z����o4~w�̍P�]x�C:��O�A��<ӐA+�u�:k�[mH*���	ahM�ǍN�;��M�g]6�F+F�'�b ɍw�.w0�tG�6U�&�]C
�7��oq#&�Rpa�.߷дW�a'*΁��1�A0���1yx��y �r8�r�Ϸ�Vl�"�6�n��G��*�
�� ����l,}��K=O�}�UkIڤ.���q#���;�^���1�� _>�}:�
( <��(�Z�9WEO�:������V$���`ʰ��r�*cof<�t��ŝm3�H,����Ѧ-z6s9��VN��Rx/���@l?��	 #79��IJ����A%�
8�ﺺя���_�x_�#B <\�����G#\�Տ��z�˕��}޾�����rP�2���["���j������ U�7�>7n3�z��4���h��n{� pJ �_����b*s��#��=���Y>�����N�GDFML�m<����@>�RZjF)K���E���F��C�0D�QP�����\]]q}�;����O����}O��ޢ��D�-�Gy�:fZ��BV�#�*i�Cz @��֢?^��-���U���ګ������I�4g��E�/u�ȝ��S��� Ο��4W����0:ed�9��WX����}}���:��V7]Ɲ='0�-Y=锪��a�ļ@3�_Ҹ{|N��gƘ XH`u��I�bC����r��ޝO�JF�>�P3Xq�f@ZNخ��݇��c�F���`0�|�R��A��\�=*]E�-ؾ���x就�[�h*��@��-#���POh���ɵk��=栟�*��v����M�6��g|�HҘ�F�M�X��x@Y"AS\�(".����Րc��E���gX��m�ўN:�����[ؘ�6�M̏�4*t�4�Mv��߾� >�F�^��8$	@p8X�UD{��MTނ�)Y ��XnH=ot��dt��p��l�95i��Ȱ`���&�!J�Mo��6)����;�3I�������ij�OV[ �FO?����q��xe���qc���Z��<7!�\����&q@�҈���lt��@���w���&���
�^���Ö�Ǉd,�	����p�|<[bлUÅ��H�ba��#<:gX4����o�G���_�߿I�"$�}'�	���?==�/?����ݩ4#g���F�k<GeW�L騣fZ���׊���*����d�'����|������z6�a(Q-),	�y��_㨍�H�Ѫ��]l��ԛ��>��<x��`�Ү�գ�>p�(֔/�B4s�Xo�SM�k*c�XJ��\���?"E7�#]��-a
����_��P�0_p�Z�܄�Z_�C�ά����I�|\�97�n0�0�iD��R8jV��q'�?}Kk�9�Q}m8ٯS�h߭@K����,����
���ֈZ��2�˴Y��;�DҮ�Һ~�����FJs@�;;�Ƒ
b����-L^FnDuϑ���5�(5-�\�h�T�N%�-�ZM�e��N��}���*�* ��l5O����@5ױE�P����m�Lw��B���� �����P�^a,�-�v'K��[ӯ��c	���*a?�=�����d��-/eu9�b}N�[�qX���-Z�[qBQcF�"��,����#���
¢F����r��A��;�]e^�b����x�>��<�/4cT
�5�FV�O�ѴM��b8��T��5�C�ܹ��4!\:��l�J�C�6�"s@P\��&;�ڴ���m�W��D3���*��כ��7��y5�P"%~ў2R��m4�G Ҵq-�d�������4&�a�����ΌF` ZuH�`��
�&���Z��Σ����/N���/4q|����4��z��di@1^^�J�޿��I4�D��*;F͝�z9��
o�0��� [�7z�-f�r�Z���������<&ck�#k)!��f]�7<�ބli�{+O���(>��H�<�ХϜ:�DM��cQ�e������s`H!0�NU�R)�x��,�8�P$��L1'�C��N
��W���l���B���}�x������}�*���o���h*�`���'���w�Y�qF�w�#����xZhM�	.��2y��������e눁rz������w;U8p[/s�f�Z�4l�Ѭ�y	z�0��h��M���Z!u�K�_����<K�^m�4�m;4J�Dc�[v�t~蘘<��J_�V[S�}�}k`T���Ú<Y�����͝�U�A�=霳ќ4��Rx�¼
 4:5����������tag@�^. ����_��x6J@,�M�_�y(P�	�p� �o����E%��pϗ˵\]�P���G�7|��bF�X�n�E�MhT�0�QM=��8��}�c K�r��u�`�e�l�S/�"J��,.���`A�a_�=�|�	�m��+���;��p��@�Hv*0dI���ؠy�	_>W�b/��.e�,@dӺ(�q#�9V��'�Q�㴪&O�g�0��m?�
A:���|{x�`���Ն�A��7oe��`�����BU��������ܩB�qvX[u�E�xBD|�O?i�<"s48rJ��*h�X�2�����Z�(�4���N�A��UG*'tAۥ�`�9��"��<B��������cl��J�{v�Z0Jn!����"��q]OO�tr*�-&�$X�mm[�E��"�]�Mc�+Z�
�c�`KQ~Un��C����^������^�Xv��k��Q��~�
����j7PӔ�+{6��!�̟�a�Y�0��Cu���V��������vqa�	и��R�]�i{����jL��7��7�Vu�C�tp�1��5��XnĆz��8joN�i��(k��]'�b�b���5��SH�xK�NF�i��%4�R$�I��XXT
�]�0t#"A��^�nq��~���3y~�M�ŀYO�mNΊ� Zmˠ�k�s�:3��y��^Kd��x���|������]���乡CB���
b>�h�S���Ϊ1�z6(:����� ���
1�i���Hz�V����/c\�t^y�c�:��C�9s���$!�:\_�1/My�ۼ ��L�K��F3ߋd{��+03X6c�d{��s*M�G4�mKJ�(C�A�SEbx�px��3L�K��H����T�Ъ��Λ�$_G�r��=_ҫ9H.��c��+Buu�\�ˣ�����</�h�	�[!�i\�ڠT�ҳ�{WZtn��Kp�T�� �W�����z���s��������h��Q7DK�Xݤ��i��4�`Q#�Cl]�`�$�����F�}���+��%2*wbZ�FD�J�U�FQ!�.��Č���B����v97m3T�M"+u����h:ysqiѯ�\���ĠXs�r-��>�&�e�{$�c�I
?̫/��ع�.�m���$�d����%�5��ĵ.舢���..��߶N���Y���#��H'�k�R�����УW&Ȏ{>��9 �י 4�V��L��8R�7y��
vN��u��}��@ ��6f!���9����G9?gߕ�Eh�|�&����G�^��ف1l�4k(Q��"��>5���1�nbҰD%�1�>	���z�>{t}�s��XGS�#F� _V��U���Y�^q��I�0@��V�yy��`���vԱzM�H����O�J~�z�j�7鞟��͠5���	e{!������*N�����*�9h�d@(��͸&xE�
9��[똴�)Lث�a�.��7H��|@���Qɦ�]�q����F߽qn,,�~�uh4-�� %SP���HɆ��EK*���4�F�!��H�il��H�q��p俱.Q�Pt�/g:$��)�J|2v+]gFeʟ��A��͂R�Г�Q?/��Wwqu-��=An�HhGqr+#���h��٨�F����t����=�U:���\�"A�J�L��>�8d��`iMq��q��l1D#�����59��\�1 ]� ��J;���s;׏��K�Ś���D�Z��0�H-A��lťrJS�<F����MӒ|��4�M���t��j���x��ZKLe��+m�
��k��G�ӎ1sM��E1�>��A?�
�N�����޺Ր���A�֩S�^o���8�f�ƍ~���+0]����:�6�"IK������#%lM1��߯��v�z�~�HFu�t�-#ٽѴ����� ��j������)4�����5�2#l����r� ��:Gk���F����Z|6���P�Jõ\A��Gys���+���WƵh-�-0����4�.5��@B�k�������0�yB'�.=�����Xm��t� �*f�/�D��͵r�@]��ڌ-% ���Q�S�M���>�8;�8���̒{jh���?F�󮞣�.��D����+S�`�s��"���1z���%�Ls���[���`�X���9�7Z��@,G�2Tţ�Q\Q��w�>�-mTHl	|J�=���R^�1*=� �K(x�z�����Ee#��j������P�*�;���J�û��$����+A���SFr�j���K�Xw*�)�|���J�;0��$�dU�B	�����h5z�s�(G��W��(��Ơ���2��Y��ڏ\'-�����q�6���\�̹y[K��R��^.�;���g�<���(���7(�� ���w
C�@Uf��]��ճL�j���b$5UH�#��+����Z�������₢�kx��5�8R�в[��v`qpP/.W����X:��r|�7=8_�.�h��4}�?j{ �~첣Q6��xU!/��ي�p���=|�vUg����v��#�b��ȗ��E&�g��gHd�grp�\>�ќ�"k]i2�P��T�|M6���j��L�����m�g��v1S�Ss��d�	�.�㕆�7�AX�c�m�\֡���y�sޘ��F�$����F���������e:+ �4��fԖ8�)G}0����:X� �]��������p,�1ܬ�s���BS��g!2���¢ΐ�Y]\8hd�z�F^4��*ϭAzp#77�V���(�kE�Ѩe�$i�$�P��t�H��d�@c��GSr�X�ț�����
Զx��{�b�+&@�����2�m�}�nfOBk��Qv�z ���m[ m��d1_܃�R��FQ58���-������y����wy�Q �S��8o�3ǶRM���h:�ʑk�B�	�ςhЅ�X#�:��3�)�-m�*��i��H���o#�S��x���<C�2Tى��P��#nN�����8�7��*�)u��0Kp5�0z,O�L>��Ơ�E��EZ�˗�b+��@>r����#�qg	a��Ɇ��6y�_�5�w��U�ɰ����.�g�0���ʔ�V�`�N� ����g��M�Aל�û��������n�i��ë�l�6��.mr0��r#�o��a�ލ�\9AR��� �"����H�Zth4A����rQ�m$i�eM�5���!����L �����!�U�U�ԛ��4~�� ����$+���_[G�c�bVþ�>08+��yn𢡋rV������:�S+V!�FE xB�a�_%�us�����:��w,��V���XY������� �n���	6��4�\ˉe�QE^�˺�;���h�~S"�O
�V웸��0��b��J�Ǧ,jK�aAK�5��Y1����=���Vޱ��^LA{���/Ogy�l�ޮ�����`l��д���x�r�7�1T����6��o)�%�ޖ+oB�4��%�綡<H�"~�Yos��`�� "WM�����W��~�=���jͰ\�` Gu���>�H���
 ����>zu��:Y���pZ�\J����Xҝ�}�+I Mw�5�ٚ*F7�U��l����Ҕ���LoCAl�����q�	f�NO����ڿ�����urn�s\��� r�շ�!Z5����;�r>��E>�mH��޾O -9����ڑb�m���m���&�k��=�,>~w��l�_�pV����M�7�������ڒ3��wk`���Z�g5��>2cB�9���tm4FҮ�
κu�Ud�X�m!7sA�ߐ��ٲ3x �B�9 �.�o��@�>#� O��I���8ǁ]Y�m��WZV���<<���?����`7�F.]�6�F�^�%_���g�iB(L�1g&ڬm���c�b�t��J�.W��q����I%��W4@��!v���Xr��� �G�b�sM�?���]9��܈Ao�3xO�x�9^�_y�����[��hћ�:��7T�Z_>��R�PUHI	wS\��MKׁ	~��`���*i#��a����%�D�F�ߩ��p�
<����8(J�[˙P��_=g��������*H��w��7E�I�_P|��{���s�F��Z��7��"��U�`��d̛�h�B�X��D%ֳ�������6���W�R'�� �Ϛ�!@-^�ak]#��|G�$����g��Ũf���b�I�fs�F~��Gy��r����Ӎٟ�!n9��o-]�� �������}I�^)u!����r��xȿa������I'R��<�dռ��9���M�ejՄy�ji7*��}�tOCA΀R
��Fx�raª��^WlՒH������9�Tm�8ӼHD$�b��CT���@X�Ō�<�tZ�^70W�+S;2���@���[�~-����������9��N���X�����=#�H�Ԥb�����Y9�ȁ����1c�MO�����\�^?=>% &F�W;�dCb��A��R	�LNT�WbN!�/�^P\␋Rjki�!�i�� ��s$#��pGg�D3t�P�uu}����M;�'X�����v^��9�H˜Ӽۢ`'�O�#ϥK�E<m������>���z�z����R�M��{�R5����9��cت�k��3��s��Љ��h����JM�g'�?vAU��Rtyy%;Q��>.x�&���p�5'��
P����ݝ��ݳ�?�X1���V�;ޚ�/T	:���"1�� 8���MM�H{:6en{�[y6�m�l�Vĳ�mlV�?V�Om�ϳPE��2D�B�B�����F�E��9Ds���^.TE�������֠��%��fŐ�YSU� ��Ȇ$�|�~�� ���
�7~��A���!_~ 5���z1�>ZѤ�aL�Ң�r/W�%-��������m�^����X�f�f���8*Qs��`iĉdt���]!�1U�Y`�.�ْ@��E6z�I�aۨ`�_� T5]Bt��6�4~�@������	z�a4���M��0�
��Մ�=�E�,����z��dp��`��˫wܨчlI ��] ������I�#Y��Ʒ�#fD�#d�~V�	��dD��L��l��1��f:=�%G5"��
��M��е�d^p�n<lO1X.��NLKl�<YVm\͎�n����\�1��)���t��Lp�P��F���Si��5N��p�]c�`�k0�|�x��PE�2��b3���5�i9��mgDr�ʥ
��|�2������ZJ5pzi"���@�����x��8֟��k�X]�5��CM��_�jT��Ttf{l�QW���G�6멘=wB��é3��UDv �K���Q�Bӽ��Ee�5!(:�,��<�G#����d}�ɳq��C�n���
������m��-v�hts'(A$
��F~���H� ���@Κ:tu
U���=NW؇-~���垺f��I�7r�p�iX��񠶣UB
��¤q�f'z�T�����Ӟ��R2�3y8�{Wl-eE&�e��R7�9�T�E�l��B0ՠ�H{L Q�]���� M'P��`٭���-���ϟؚU�����a�s;����h:l s��e��;�A���|�trm���ڗyT ����k�,%����۲]�T�����Qi/���~o�
�+߬Zo�'�E�܁z�������>S�zu���=��2e*�NP����+�(��+�/ځ�L���~�p�Gm��d������s-9�r՟R���&���/��y�3��Ioh6%��S()M-���1G�ZF)O���S���(��Y�/���.�������!�k9p�`]�R�����2�&>�Yko.MW����@��
7#,w"����}6E�.�!(c���~l��εx�3��,����W0t�2@@{V3ᣕ*[��!�7ԏ�g��h�{�Fb��ld�Vzm���2�&�^�ų�Sԋ��L�(1A9���T.�il1N�����ꚜV/U��7�.h׌&! ���[�/X�Ir�Ƅ��Uo���@�91�C���E�K�F��lܪ<5�՚�-ؼ8��>�%�Dwbm�DӐA��&�Bz���BL!۹J�5Ϯ�]�&t�3ɝ�zF�'�3B�wZX[�q-��LI�q���O;w�F���D�w0���Q�a,<��ᩊ�+�g�e�&t���:mX�߫�Ȓ�ԉs8�X�k��E#C�X_�7�a/�p"�#58m9����ű}-+��3N�8г�O�?r��l����y*�HSY�e�Ja?x�8�@�W?j���5���(�إ9I:9S�9ڟ�K���47v���?�?��Y�����ajK\7M�\nr?O� v�vN@g�UB�u� _���qT6b.����ן~��?}���I[�[9�;���j�U�:a��S$S��sc�z?�ՓG��ZP���<w�V�h,eר��Rh�L[/�9�gr�NJ1@���-�R��vʇi�S'�q]?o���{ޱ9��d�T|��~ �0jJ}�J n����&��Y��$̵�6������xO4�9�G�c��lO�Е����XTɧ�:5>��L	��p��
n�ݾv�����g���5�p�G���k|��%�ڠm�췼u� ��؂�i��on�����Ǜ�9��Y�9VyᾔL�I,f?��b�*��>~���t�!�P����1S���z<ǓQwd�
�: X��l��K��>?�������|���ۛ+�n�@ֱS9n=K��{�6 ���w���7�rq}#W���d�}���(NJm��R�dV��Oq�j�'�����zw{èB˪-$����a�"�
�%�EJ��u�8w[����\��W�'�IXD��ȇ�a�'������Q�M૱{rLv�)W�<���F��Xt;$��|I�2y�Pž�ژ��뮤�fu�B �ܤq����d ��FS���\jԪ��q{_��i,�)�`�mJ�FR�Ʋ��,	kG��,�7߿��o.y��tM�ӟ����4u���C��/�F�Y�������me��\���!��G%ݻd���{�gޜ��O��(:K,X%�&+^hOs����GN�0��7�K�2΍w�ȍj����ʋ.�=�m���E�vr���*7��:�q��q9�q�堌�)��0j�1��G�Q{��:5XR�V�T�8��/�Z�Q"|�I~,Uu�5,20*�<���t���`1��Y[J7z��&�`W�,Og�e���E�"5E��V�2��E*�ot�Ϻ�o� �Y!�Az������VP�ST�]\b�]��u�Ay@�r��F�N{��v��B
����\@�Q޿�N>�𽴫K��?�$	�Pk���=����gM:O/D�0/-R��W�#�&�W��J��ӧ_(`�1�c	ΛvxK.��'yzު�4"��2��b	���#&Xg:=Z�W����kN�l5�N��(���r����@��J����k��Ï�����^��O�>�����K(5e<H��Yv$��+p3�B��$!��G�,��M�\�������%��1��F���Կ=�ndqr�V�����y��=uj�� m�6�Vv�ޙ�3d)�ӷMw��	Ina�����S06�� ���RЩ��!G�����Th��������2�70��^�8�{�x\}�x)�}���Oi2�,�O'y�暲	�yg�F�X�-u`�X��,�8���^�r%��H��3O5�B�e��~�����ɋFTHR үd��? l L +-��=���aZ���{���k�*��ՠ3Adj޵:fܘϪ}�냁y���&���@{ 4�zj�:�����!G� 4q�߾|b 0�|�J`k�^p0N���t��t�ɻ]/t��M�܍4��Dy����soQ#�_D*�S�c�v"�:-" g*���yR����s6��eb�o�w�ㇷ�����M�ᴸ(*ck0�'�������0J��>�y4DLI���+�-�h�˵��?���EnBd���ϻg��������׎�<������(�s�A�UO��֒�S�G������*	���U7j5�غ,���d������j�{EuԬx���|���=���h�i筽|�7O��ڏ�?��X{��|�1��HOTт��d��#�AJ�7�P��^�����R�-�,r���n�a��{�Ӈ�'ꮼ� �V/�f�.���]�^r�r�P�Ҫ*[��.��4�1���wC��;9t�΂O�RZq	!WlY����2��䴽��{�횑�3�A?��{@�?�7λ�N������a]��|����M�.��(x��VpB�6ޥ�uh\A�g�l���������ı��qL�f�隀�r�� qt�Y���Et��_�A/G����[@p���l���ƛ��������?������~8ȧo;	����F��[�t����B�"��2|N�z��Eb��1�<GsOM)����J�ڿ@�~�K�y=�%.1!ˢ�d���B���W,k��E��-�k,ZjG2ax��R��e�x0*�f���[b@,������
EG�V(2�2(��g�	��W�>�d�u���u/;uca�һPD%)�RP��0 i]ֵ�-�>�D¾=��'OkP�mV��بXy��K�Ӑ�D*�r��Dd(��l5Q "m��L�l!���=� �<!tD2���GQ���ӱg�<��=w����0��ń�l��G���F����FC��T�����Y��"H~�v�V5�kj؎�  螽�"�L
��|�VQ�B��T9A�Lf]֋��/A�gD���3��^���\�T����0��zލg����1���Y������8O���N�A��k�X�uŜhsD������|��V��g~�۷oY)Ɣ�B�����; $��֖D���Y��6d�O�!�dh��ۦ��gJ���Y�
o�S�=e�4.;��+z�]���%����QRq%=W�f�Ϸ&�m"I�t���wt����݊�W�#�V���4Ku�������c���ﭥ�����L�Y�vҹ�z��U���{�29�߯yZRA�2�Ϊ��G���=ɕ�Y��-�4�:=�����Mr���1B��gk�'��ׯr�l���m��N����u#�(��r
�8�27&����@�&�IQ��l<�鼠=�9>��BqPl̃n�h^�e�'p:�2�Ni�]�t�noߥu��ܾ� ��[�!]��=�����U6e��8P4� �F���o�Ez`��=�|�Q%V=��wu���F�GW7o��xC�&�<4�ܡ���J=��dEB^@ƿ��������+�����(��޼����!�	Zu��\�����\���3;w��q��\�DMZ� �}�]�K���=�k���t-�O�=&�?tTEhL�Qy�l��ӂDj"�X$��RU0�urLl�V���j�5���v2����*�����{��̞�?����a���k$��0��|�l�]([5W�yK7/#Z;k�7',v�*�rGV�L�rwn���-D����g���V���k���}�����C��V��&F���lFŰ��O�sQ�t8�l׫H���!|�.�[%P�I�g�	��4pSeR�h���X4�h������^�w�D\$��fI����1�<��4�� l/�۞^�`$Ox�+F���OF�ƭ��g��ӭ8Z 
J�3�ξ`H�.T@��G��DMI���p.�-EƘ��ݤ%����|�����$ct!����2�~(6C�
B� `C�2�s��� �^��h��	�������{Vݘ���<M��:	��-U���4�$�"�}�ء_ &��`�>=>�С)7Z��x���GN���vu]e�|��=B䢄=��Ɉ�*���iIƮs�W ))��ϩGO�1Z
Q��ܻJ�V¦&<��"/�^��a�UQO�*���8c�q ��T�c�&��HKN���StM��R�ܯE��q��9���
�s.^S� *pWn�|�`��P����}a�Y/F��42=Z��ܓZ��'sqq�L����J�_��>$�����o����p��>����ow����I���_ɛ��&�P+���T���$��^���"�{�ȉEJhἽ³�~���>fпB�u:��ye�_A���t����ț$ Լ~�%@q-�>�	"�Y�KM�v$G�5�
���𜓨�\����(����KF��1i�v�R,<^Dp�i�ά�$�=���=��u�����/�w��֨{˂���x"� .�M�H!�f��[�t�ו9��c�@DN���Y�[����dK �b(�/����=�j�qng�e!���bnu��9�x�E�!d1o�\����RPli�ת���M5C2�@Cj$Q�t�猽�m\�$_=��[%��4�pi�4}p���F�B�{�����d�]��P��wRi��n����FYW:j�����_��U������j�#I���#"y��*i��}����=ޏ��{�۝[6��YuP�$�,�������z�;@�'�j�����]����˹��Ҍ�]����_M9D�ީH���!׶R]0ͨ�yc��/vpŗX��%D��{�A��ddw
�~����_tS�3�a{���'�<�GO���O�ڇ����_��^�l�S����x��)�����t��%(�6F��vM�����{i��ֳS	<���a�k 0�]wKs��Y�^Kƈ��-MU7�.���~������g�]_������do��8,�������|���-�r��Qp�u{�
������^�ަ�Lc��e��MN�`x$��e#����X��������������v�ׯ_�S������������\��<ij��><\��(�Y
��`��9�X!/�yd_r�Ⱪ6��-7���F�1X�~�NewHX���t�����̹��C�0��� �Q;�S}�(ua,VSn��z���3��*�	P�3i��ޗ`�}����S��w}���[mX�k0�ת��0�|��]��'g{7��������9M�2�/�m2p�����������ﾷ�O�jNb��)���p�y�����g�K���/��ǋ�'��8	$I���2y��6� ��'�}@%K=w7zhB�P,�!�^�ܖSBFg�|B+ʶ�b��bq@������d	�������3�yy�S'"�l#�6��{r�k�)G�sZ����1��p���r�^�}o�>~�ɓُ�?psG6�#��%�@󸣏┢���qa>UJ�7��ѕ9���c<4����$35ʄK����D��AZA����3�<�>��iCI����Q�N2a���ɟ�Xz�$����wr���܁��1#���6�،�������f;�H����d�k� ��0N��Ԟ��Y���&�t�dr��@k����)<3��ȅ�����O�.+�,�)�QJs�����y��"��	�s�����ݷ��D�h���z��~V��;vr�}�q��geYe�T��!�+�����F�`
��y��y�Ú�����;l�a����n��lM�ɱ�U6s	���8����_��g���o���%����;z��0��g�aӺ�jb�vJ���#��EI�T���%�U����خ�LC'g���J�v=��2���;��3���.8Ͷ��Ʃy>����n��ի�ږB��#�W�)�)��xH���L�1o�-��yl�A_Y�1ו�t�sg�_u �߬dr�3��C�_���ާ�3�=����)�`����G��Eb����B�>�w�ƺ�5q��00N9�O�S9�0�M>�Ds�	�W
t��� ^���A[0�0;��^0�?/�L9(���(�3:�[)po.�0�oBm��(��H���p�R��'�c�2do �� e}i������
pz=Y��~��^��Iu��:�����}���	��x�~�e��!�m=/�Iq���h,�B����׿����9�r_�|��ڻ�.�1a0=�h�:�A!��NS:!�Bk;��w�䌮��GM1=�}G��hm�����Ѓ霡D�̬�1�qv�A��$��=
A�l ���Y�~������ߺ'���
C�KXBj����8(s�f�D?�n���^��]�V�=�۾�u�������6��U$�� �zR�'�_N�<�eg��a46�:���|��b
��n����0�/t����ku�p���'�@XD�$0��=Xj=2~���Z@���b�D��ƅ��?_6>#Θ��T�(^�!G���ݬ����6�*pLxi�>�l��iW�_�
��Y���;��C�=$�Ѿ1Z�x����Z	�@+n�߂$�9Щ?4�]����Jaz��u���%?ǚr�[�Us�ʻI��}YR�u��d�}>,�pZP3���h��Q������e�{�n]�r(�0سC{�pi��00S[����dN�]�jC��Q�s��F��	��\�w~��$��&��]@i� $Y{�&��\��S�k���P���P=m= /�! +=8��-��s��o~S2�G�kdɎ@`Ki  C�{��h��>i���4-h�q���v��b�5���:���5��1�排̫Õ�|�ڞ<z`_=yĵ�Q] ��X f���wO�Hn\��(���X3�을�,�,�� �6���FX�a�� �� \�Q��WF�itPF	���\c(=�0����VEw3vV<Om|P�0iL�'�v|��Kz����6�1u����{\����(�߳^��kߥ�:j< X_�����Žş ¡�������8���ƺ�a�fm�n�����;j�޾}O@���/�<���ݷ��P��b�~o��
�����
����� x �X�(5sr����RH^+�m�莝�j��|Y\�X�J���;�k:/y=�k]���b��Wp���xkݬ7�;�M1$Q�-�y1��$dfb��kX�hvA������:��=��\aS�� ��ܫ�c?�L�j���X��y�;�M�h=b0g�3�%�����)�MW�Ƶf=�DlFv�W���2X�1�r���z 	NEzk���8��Mr���I��U%!5{6�F,�$���^�K��҈E��&���u�t�LV@\�͝��ZR��H�o�k��_�m`D�ȿs�A.:�Yـ�g"�5d��T��_��L�����l����?'��5��Cj%����$�t�js��"�z���y�u�@/9��O]���߆���!A~k�W�c��c�8{���LOc��_�(�$_hꀐ�ODԸ�l�P����&'�i{��z��!��N�&~l	]�����ͼzA9(`f�Ȫ4E1�y\S,j�nbRh.��+l@*�{5��3�i��a|���� ��4-5�3��e���~R����|��m��d�00������۬u�(��Z�0��	����-��[R�y����4H#��׃k C؁\|����?���S/��vc�>}�wo�ڧ�n]\kMS��eT�8:�3x�i0/�+X,��R�����	�+��C�M���A�'����gk�vl�s��-u�\m���s�+(���g�Hw*�T��0y؈�TL�Xz�@_b�Kqq�������u�?�����e�Z��:*��Y�^<���e>ۻ昙Mx� `�����j���Ĺ�9fƚ��u�6���>�'4�p����cZ%@��rt�,���r��~ �K0�`���1��ks�Nq�����7_��|�7�5�m;�
iv6�RӾE��5S>x�TL�N�3u�f#��]�akD����`ٷF��X�K�w���K��,.�d��c�( ج���0]1��b�v;M�[�������P7W%>"�z;`�l�,`�}Ge;�F���N�e-�1iD=z�I�<�:���V��c�z�([t��5����_)~��gy�V:F��@��.�$�E�7�{��T_[���ds�C�V���0}l"��l�����#'��h![�+�u�C�� _��,=�ONh`�#��^t�N� YS%@nJ`E;��[��P�����j�D��˿h�jo�������3=2��R;�����\\�$ve�)2Q�'��<m�}�_8���h!$��x�b��dJ����v� C��PceHg���48z��xJBi�V��98���fX(1���7�	�� �m M�������y�|��I c������؂�2	x)���?PM���H=��f1��|͚9�1���`Z�q�ܦ�@>������{��y�M2W�\ @�ũ�C��� G�Cf���,���c���H���p��X��6�=s�b�����%�E9��ť��/�y�����~|������{:L_~�l�WW�L��D��@�.6kw��}� ��muw�.����Cv����5�6�����9C��1��w,X�n������%�ʧz�ܞshѠa�'K�a�"���~+�g����*��>�k�_�-B�1�׹��zWo�zW���`�/�E�a?������">Ã-��ЀU[�Γ�~ne�����	������X�(BH�N�M_�8��.G���g�M%��3
F�Tem����h/��
ރ0���*��׶�N�K��af���Q�D�w)�G����If��}�='�����:��{�������w͢�1"�LA�*��(��~!�l]�)P%�+��zr�2ͭR2t�eٴr�$����9���$�x�� Zi'�N�@�5[��l��ܐ�����k<�$�'w��`~�`�b������1��VC��;����~�`�A����pe	ڵw(��Y��Mh���e������4�������J�X+GV@>Ismn.�kr{6ɗ�������1ݖ�ٰIj��E��"����`�����6���ث�B��:x���9`�ۊ}2:&L45�5�r��ۻ���� ]Ʃ�\�#�A��,�5	��B�;�/lpe�!(I�e����ݧI_
��/le�.��8B�W�P�x�Tg�MC.�C5�k��B9�h��I�t����ue���j�z&W����z;3@��Wb9trه7���y���林d�H��-�ōKcmL�ZI5�WЛD��0�t�����\�%DI�5��Rd����f�������<��M���-O����. �J���R1" V�MZs����$���5����&vp�g' ۀR6�-���Ĩ��eK���?_�6�ʛuO�f�5~��g�9������s���;m"c�����8��>U6��-����	+Iз4�� 
|t���� s���#��c3������g��E5�0��������C�/�������Iq����,7F�"�κ�o5�'t�8�s �^���ˈ_�(�u�gc�:�����7L`��Z&tp�y����7����9�n�Hvr��q����se���,p~��(G�����}��8r���gvj��͚q�j�F�:�)�DZ�`})F,}]��>UV$�cܿ�j��a�3t~�u:��\�k1�c��{�Ϫqf<_!5��Q�5�]��I���e (����rl�]���D���J ̽�uĵ�q���qH׷k2�)ع�%Gw�?�Hؼ��	��꽜�f�$ :S0�mz�d g�YW�l�`uCJ���^D&l�.�g�������.���"~,��
�����5!i�;	�NHʾd��.W.5K�9�
�:\4Hь��5>�{�n/1%CH��>�hHA��%�JRD[�&\`���Ŏ�!���F�0އ�5h��2�_po��R�+�p�ɱ�����-�m�<1�"vZ���K��*}�UBW�A�-u�o���e��M��h�h	Ye�V����,T�eq-����'�l-��kK��d�Fc�}5[0^s���"��[ci�91(a�����Ζ�I��x�jb����,�(��`\���ye�:��|e��"��4[�C�9�L�'�56�-�6C+�Y�{9"�um�D�KS+`~O+�BO�9>��b�AY!���%ڼ���o��Ǚ�Ĉ��!1	����`����F�Ġd�p-��]c5-2�
9�5��LF�{�(|����/(�ų /0��W|�����D� �;��9�BW��P������b�^D�Bp�q�
��bl >�3�w1\x��Sh���C���1�Nh�7�Pd�Q�k lY}�L�On�\�k�"۶Ժ�|�c��[���G��g�* 4��V�n�T� ,@�ތK��:%%���a�9��z@�e�(�Ǘ �h��7P�n��it36ͻz��:��p�./y�q��]i�|2���A�r��ݾ���j��@�F�	 h�'�1g9)8XҖƼ���Gy�38d:� a��Fȃ�s�9�K�=:��L�e���|�rH�vV����DM+Y�)�_j6�,��v�U� Ɍ���%|(��Z���F��N���Da��ٍ[��꾑hk�g�Y�[;Xj�wv�c��ǬR��}�Z�M0�3�&XP���V�+)5ۚ�4�斄�>�����]��n�&#�p"����*�*Cb1��3ѭ��)�g�ޔ=���O�Q�1O�l*�,	ħ���\�
�*1�%t��Qj(�^	
R�Gg����W�:ל�^���6NH�p�H�ט���P�S-8���擕�IPn��H	��?'�f `3��m�<|�) �ڶe�d �4����	���*.��͵�;r���ϥhE;����L�9��.6��Pi ��]	l�J�	�����?�����ձ� 6[[i���5��ŗ��93��y�����v�N����c��*����_	�s�����44 ��������i�䁅 ,�,��{8��5������o�D��U������8	N�Nfn���o0����Ǯ*��3|K5p�1��sd�D��z�֊�C�s-��fόor�Gh@j?���^�O����kתe���k�8h���جq�� L3��	o1�M�A�9�X�SƎMj�'�7�3U44'�|�f���Z���k\�݄�����	��в�C�K�2\V�v�@9����o5��`�]����	�vB�d�r /)u,Y/l�˒{�|;�\��3����6���h�li�g��}�c�%������%Z��P��ȝ	&���%�Qe,]��Q����/�nY�����u	�G?@�	�3|X�E� ���>;Z'J��FwÎ���Eh�L�lt���M��Hk ���"���L~mV��z,�H��|V;������`�U��<>���h�q�M�kEA@�%�E��N�F7K�r��-�ö���fG�E��ۍJ��L�_Gk��%G��u��(���'Z��K���!�ax�Y3M%f��c:�&��3Ԙ��D��)#�n��5'�u.
�Ş�碛��]��K��^ڲ\����'�&���(���d��uI��/��%i]�*G�u]��̥p�O�:�Gh��څ�ä-=��z�V���,��Iq���v4pP��E���:|�˛����x'���,���]\�K&T�U9�4($��4y7JKƉ$�H,8�1��z���'�P����Al��g
$Vs,�*�LUx�	��Jv`�pFu���f��ϬRc���r�0�P���T�g����+6*��0Sc���(}�üg~�D�!�� ���&)|rR\M�~G� �s�P��ʜf�Z�>2)���C���i��0]׈�~�\�l_)�u�9F��?���:�G6,e�O0��k,����v@+c���wY��'Ҽ-G_C� ��e�{��ǠuS7d�(�;�A���:�v�yoP�AZ@m��|������N� !:�h��،���;ַv��.� 4x�dJV�J?z��I{�{�ڥЍ��� ��,@u�i��|��3�֕�9�#�)Yƚ����gu��r�{�*N8�*d�g��b�f[�*�X��Z���٬�r�����u虰^���/?zQ��͓Ð������ �H���� ��]�����7�!RTފη�v�+��+�j���"��O��p�X�9�xkC`�O���*%ˬ1�Ȼ9G����fo��R@�]O��A��X7s&�ى���g�Z��D�xr��Xe���&I��Y�� ��j'#k%1s�6��3u������C��n%VT�Ȼ��*�^a�����
�J��I�>��d�*i�L�@��	!�����i�,�=߬뙃Asm��)�!����ea���+�MG);r���q���AW]��֏/���Rf������
p�#i�@��n���'�����׿zF�����g;;�������m}���آ� �4����,|*�?sa$�e� ;��#��
`� ����\%-w`��l7Ǩ��-���6�_ӺH����^�T�X*l��<��G&1��=OB�ѲǱZt��Le�=���]l��a��7l��V]��՛I����00�Hրf��� D�i�Q���1�Ȯb��sJΠ��#��6㖽�b,U\�1>h�c������u ���ۏ�>��� <�IR����D^���Iʘ�uwF����wK���� k���}��hd���}���oDm�_%�v��1�N���C<G����6$���+3�6|a0�&��␁f
�jV�U����>f�Ӕ�JN2)luv����^�^�ڮh$��5�9�����^��}Ԑ6�V�{!S�\;������8��*��V%�h� ,�[? �>#q�9w����0{�$/�� ��N��Կ~ӤY�� DQ�[���w?� �2q])�n��޿�;�_�u��d�ɲ����=`�8��9�}�]cSIƼ\��+���f&���֤g�Chqs}�kL�{���
 ����C�9�Nz�4缩���i�3�q`p�"Cz�Mvv�|/K�Cp'�S�4��E�/UY�|%N�#��i�A��e�rRv�D��Ϩ�(�L��W݃؃R��E�*��D.�i�Y��c�X����X��s� Ru{�4b�,�R\��&/�n�)�9%k�#��^v��&<��ѯFA��d��Y�(M������#j��>���F�^���z� v��E��	4���|[�S �l��W���q�2�==2�x\�Lv0�(�RB�S�<�ً���aY}.�����=1�ǭ;���	F���8ט��ǎ���q���NM���j	cڔ�m	��a0���u9�f�A���,)@��C-�چ�u��N�U8[�䋖]ҫ�O�{(`ͽ��{��]7s�̃	S����19�0�OL����5�|�@�c�<� �4��'�'"�{jY!bsL��d27;)�Ҩ ���D�-����./�l}�,�S�R�~�Ď�'ў�i�@6WXF̱������w�b�1�F����OK��^�#�;����mՖ��p�SA�9s�n����A���FL��Nz�p�n>�Ti�Ę,����r-�ٟ��|p0������pa�A�x@�%�j� ,{d��:V#��*���Ս��l"7���u�p|�YS�/u?�Ο=�TF��Iwi���Gz�-���=�<7�+JH�D8S�<u��龂�
���`� t{&�/�M1O�����Cr�D�z�a��y�Q�'I]a�hQ�\�!�W}L{��]�F���8�8��8
��� ��
k�k:��;��x�i��5 W4H���p�ξ�Y6��J�����|s=�������(��{sǍ.��������,��70��-68����^I{K��_04j����b��i'��Z�t�sg�i뺡K:{�Puib���BHnx�,U���B#�;�5�·�T�v�&����8��~09e4;g�m�S���9*7�����"-U~EL�΂��5����vsk�|�|ލ�}�qQ��Z��/1���������)u���!�l0�[<��.��0օ���5��y0�Z�C�ެn��[���FM�[4�����}��h�󜷒-@2Un��KQ��Lҝ?c�|�uP^�ĄJ�x}\�� }7M�-{C��3u볮aE"Vc��#̱y}�X�Jl=�M��Ҧ�����|Lt@k!a���nT	�L�jQNrY��jgG�7H�U���;��'��.;�1:���1���*��1��乢g�`5S�ί%\T�|Q����e��կ�Z����r#ǘd�� K�J-����8>iZ� 3���U_-bi���(QV���]�U�4�C��'������,�3�ɍ �ּ�лy����Z��'A:�Ǭ��בg�Ņ��/FĥUg� �^�ӳf����g�j�� ��y��H�_-������K	w����z���Ah��jf��iǵ��M1��K�7�6ЍZ��M�,�(!�~�����,@�>+��u�Ԗ�+鋦ru�Ƅ��QL�֫�X�!�IF����<�v�DcH/C��1f��>Vj��/	N��z��v�b 3"5���57V�9��Sn��i<?�ݝյ���g_/:�hhB+���z+@۷��G��u�����j��B��>a������ķ�x��#�-�XS�nuV�.�B�2d{��������z#�����+K�O��*��(�ZZ�ʴD���ӨF,�ˌ�|k�_�I^M*�X��� @�$��
�%�ɘ���D��$P/^������|�^�Fn6�)����-���Ɲ�뵽}��~z�3G+��l���0�y�4}Vb�����E��--tmݶd;����.Cl��qǨ�x�(�0�{\� $9�B�N��[�ܮw�>�˗��ݻOv|t*��YRi)͟�F�5�}�<AX��/'�eK�O0��3O��ʆz�X�p�XW�w�X��q��N
0��L��A�� _%N��qr���c���};^�g2��s94p`��7OZ�޺���E|�����'�~��!t�k|�� �J��cK�H�g�����d�Z������	�b���V�f�����3R��Y�	�Y���Q��}��,��qhv�Xe��
��#�m��e9�E	FK�G��I�Qю�-���58՜��h���"<��sٔ��3��Ƭ�Ţ�s�RI���t�NQ溗�m�І�"�r���9�����:��7$��A��4ל�@�E�7UR�)ܘ=����w�~f:(� ����L�������O�+�w˴+�o�>է���!*��A���Yft��U�T�x@�6ٝĞKY���k�r���L���͂!4�Y�u�P�'�xm��-Ӝ�ĶY�"_G����I�5���
b�J���l�������b��{4�+�L� .Ӊ��;M�%�:̕���H����g�����Q�Z�Q��>T�Z5�4-[�Gc����9q�ee6��&m�@�$����o�[�ǂn��8w*/Ž��m)m0�)L����ח)|���_�;�a�>l���+/����lOD�fܩj�f�]c����(��g��6,�N�vW���z���$�˥�v�����Q�7�qh�G��J4�ɶ��\u��d��>�6U$[��Y}�H�$�"4j��HdVԴ�8gYҋY{�b�:�u�������v��`���I��Fn�p���;��F̗��7|���<�������������ޞ�x�=,�C�4�ź�*�*�رs�$ށqt-���Pcy�J��U��!��ӡ������ì��a�	��k����͐оy��$H/�'/�5>�G��с���Н��7tw�����}c� y�A,�q��w����[��l`��M��o?�y�ݹ��@}�C�4:�oY�6Щ!����pa��s��/�睳S:0YXh}?�������=}�Ȯ.5����HR�v�C�S����G��:`����p����*k�G�4 �����W%��Ja��40�{x�!f��˱��v�%f:ے!�^m9H٭��Y� E���E.,� �"�D��b��U��Ȭ��,[��j�y��H-ӫk�KJ�=8+2�;q�쎴�X�h�rS
 |�\4��Z�-���{�zgg��8E-�	&Nw�����.�nx0F��Y*b۱w���V�|�l�P0�����.>_Ӹ��#��~�Ka����Ŧ���c�\��@/�����į�y^�����`��k�z9�\�?����Å}(�7O�S{�l���n!�Zj%a�b��ޜ����ϸ���������\'�� �H.8{-�����f�u���s!�'׬h��',�ϛ�+셏�i�����qv�FǨ85X�y���R5T�*2�`'�T8�����]���F�dXVD�������RK5��8�؀Ȫ��I�85�����Ed��?�u���X�Z.�"{�X���(3������{��0�^܃`�u��˺��l/���j+���/5c1KO�������n��P�� ����~;��sZ��S���驗�[����\�iX�N^OQ�����믆�&L����ϵ�+�f�*&K,<����^(���=|������v~z���8�;iO��Dop[��qM9�ʆ���>�?��G��%N��g"X��5���{�%�9lV���f1�E9��[RG]C-�@v{/���&��N�-=��QnvQ|h���&�|��Xts�����R���{��
���&�;)��-��P��������ŕ]��+ObA����\l�?�:ⶲY�z�C�Yj���׶(�xt�I)''�vZ>�O�y���z�Ў�]��!"f'�<{���=;�6�g�G��q2���m�Z��>K�%����z1Лl���+����	�#�gw�P����K�]������u&g�'���8������L�.�k�%:UV/m�X�Г������+@k������ƥؙLd���m��M���$��p�[u�]f��M��g�w�ޓ&����6n��ېC)缥X�,��p�	à�/+"ܧ��,!�����<��Ƒ�`���f�7MTd�/r~�,?��5݃V��(�ùH����w����xqE �<�m@b�А0W����5��f_@^��Cs_�_���9ڞ�y'�2�h�`�ܔ�A�F\hn�1���~��;9>�o�>*��N�hKV�cZp<�H����F��-]71�ލ�`7��(~z����_�`�����ׂ�?�GY\���M*`Oc�<\����@�n^��>;=)��,�`V$Ə0L�K%q�\�Ur��� 1r41���Jys�� MI ����,Ldrf8�h\Ph�²�]�ay��!���/���ݡgr˱Laa���gyߙ<����M�V '�^!�R=7tbz�P��{�\�^g@��� 'f[����iøt�M{��Vjl3.�G,@^���,��`�[>ԃ������r̕{�9�g�-)O��??z/$�Q~�SxX6���Sc���0V���7���g��&�_3{73KG�\���Ț�l�`(���v�����*���!��ȳ�����o�h�%����?���Wvz��.&$�'4�F��k�]���~��?ٛ�mM�b���K� 0_�E! ��O*�t�x&s�C�zO?���h�j�&��ʷ��Ǹx��R���*����@�s}����?�M9_L�~��G(ו��Œ�h����h�A����7e�z��k���W���;�9`� ��9�ڰ<�v߱~�`�u�`��36���f�����f#�J����޹=~tϾz�� y����$	'�%\���mZ�)p�-v�|�y��QW���J�\��u,f�QW��i��1�dx_Tp�xߒ��{6��

�"�$7�G�B1U`"Z{s� �{�p8��i`�N�c��h����U�U���M7w�d�4:@�8�� ��#۬�����@�	gf��/>}�oJ�V���Ks��G�1V�������T̆�k3�kPsޮKvVP�jc�|̍zX,k���ॶ�A����a�g#+S�7o?ؽӃ�yD���]�l�_�z�5�����O/^����s�&��T��b�|�5����g���'�{�4�ׁ-�}��ʏi<Dg�k���KGL�. 4'c����)��6`f��{�x�_������6"Բp�x杨��$�L���j��?p,X08�O6Z��L���*��֬�2Q_���Zo�\��8><�{w��Ǐ˟w���}sj�/>�IڊM������T��o��� ����D�N����3tM�VQ$}��g�C���F���w��hǬ����(Ճ���sfYk��h"90cD)�i��������F%�"�|�y�Rkc����� T��E0 e�ͦi������������_���w`h/ӛݮ��U%>>�)f�U��Do��S�P�1��yt` f�`��ݻ�F ���<��� Ø�;w�ګ����\6h�����'J��w�뜂9�sM;�I��q��U�e�b��cv�q��+�|Y����k��ay�f�KL=Xy��ksk}�!j��e9����ۏ?�(	ۥ���l5&S��� �gS�o0È!�9���i˪U�?�dު�H]!�6_w�gj��8��Ki��)�a���v+MQ��N���ve���޿�`|��̶$6��������Q�]�` �+�c|���v��.�e�������/�^���5�4@+U��Ϫ/vf/�2�[IC����v�J��~V��ûg����=}|ߞ ���y��W�JZ��8����_�WȪ�h8�u��s8�/f�����=�Ƃ�c�漹n�(lZ�]����(�au��%���;�ʾ0S
�1�<��Y�܉^ j��C�{�=��7偼k��r�7��#�׼9��N�m��:G
�k�w@R.�AɮV�$�P:�'���F�z��^^�*����ˏ�wo�3�Hߤ�l3tPl�lPli�����\Y�<�M����v���m��\��%��3��7�O�P}X_���\ ±T���k�~B�BLZ��g�uc�H�/tS������_������s��BeC+e�~h궩E�ݗ���������Å�Q7�s�ͅn9�B{�r!2�jj�%���L�݆,؄Y���_���9;���n�M�YAw�3Ձ�f�Ο�/����_���� �/8��Ʃ�Ns���@���J°ٹ�[Z�6+.LD"@��0nȚ��s�}�Ⱦ���ꗿ(��]���Օ�~u�ø?~xO�|8��7��&����=#���!�B
m�~gNP�����2=(����=ﻳC���~QdV�q[�J�w�Q.�"��f[Q��o3�SJζA�T6ϡl�rݰ4g�������e�m�s�V N�(/(���K����Z�j=��۰����\ ��������6�Y`�R�J������1�w0����%	���|�UWj%o��s ����W��W_�ӯ�" #�P6������?���~��~��?��&}}�U��A�W���1f�1nJn"��VeW��!�QV�^ ��e��%�5 0���������o����w�jg'��Y�Q6����cn��w�)	A|���-���r��l�ϨȀͅ�h%崐^��`��hk�1�|����F��"o�e�/a��u�O��r��q�E��> �u9@VVI_�ò�"��O?ڛׯJrxf�>{j�����=��<W�ѝ]�w7��P����&�o�^��*�p�r0��&=s�#'��3�%��ΜK�w����־{�ؾ����_>�o�~b���uH_8zP�z��#��Js}*K��U�wQb�:k2��o�k�I��O�<�pе�6m�Շ�<s�zagdy��N���P���et��#j��m]xq����l�Q�q���g�QyѭJx!5 �,�A��Bs'c	������3����d�*	\U����"y����ٽ�MC��ӹ��p����T!)���$��3p��>4%�
 ��<�[teb�n�2��f�+^�N�{�(��f�ǿ�lH�@�o���@���.������xV+Q��,�g{����/��Q�����7٭'�L�fɏя%�zj&� ��<�`Q���hʴ�i�XLw�`��6!T�z�U�,��ӣIUs5:��|�tU ����w������帞���|��`.��]�.Y�?��d���2&M����UL�C#�@��g��1�zd�1TF���㒡��_=�_~��}�������ٝ�3�!����8/�����s�6刽�4��u�9O��+�*��Kd�����()�U�S ���g������v>�%���^)5����b��_�Ko�6ekN���Ɇ�q.*8
͍����g��z0�'�����`���Y���/�w �b8u�T�zV���R{ƭ�d�k��;�fF , �.�/ٴ� �a�2O{��S� (1�_}�Gw��ɩF�8 ;;;#�p�<\w��+�>c
�zs��͟>���,9]ˈz�ƫ��2E+Rh�tg��J��2֜��:��x����������ȱd���ڭ�UC��h3I��9;u%�=-�e�mQR����sv�����h�\�a�3,,C�F���(���j�$��r9�s��Ȏ�W�;O�P�������1�$$�H.p~,�Sr1I+˒�@���%���>r���ܿﹳ��(�Ӻh�����g{�ᓽ}���h�b��7��经W�b�T?yR�_f������~��~�Α�⻯KL��~��3���=;-��p5к�H����S
��a��m�M��Ε�>B�8&�s}~�̵��������N(��Hw�f��b�y�к{�A�;�;>=����=�r�7��ӻe�O7ܙB|0`���Z�ҍ�B�6�4���ЄԸ	� r\�up"-I��l�a�����!��.(ՙ�M�n
yv��.�J^Ki�y]�`8����-7h��-���s[~ �*Sy�w��5ʑ�Rr���Xo�9�������:��=6r��~����o��y{V�=���,�[����I��?9��S�d"������C�x�oA�{�cv��8�юu�a�� ��� Dw>�ppެ5��"S�����<�?�����-8S�z�3�p�ET���f�v��������$�t���f�2����Ah�daq]���?���_��,���k�ba������B[��)ཏ�=e����34��j�ѕ�i��������_��-�%D��,�,pq�1��q^��XKG�kS��΃i1~�d2W������ *ƄѼ�ڻ4�[-Ta���;	 ��a�S��*�ZT9�	����:�b�9|a����	�a�H��) �X���W0��e�/AX���_j���zQ�F0q����B����F������(����{��~�\}�it�N~�b�3ׇOI���M�t� �ǲ�B��|�޻C�����F݆��`�3��NlyxZ�e�^�5c�.���A¨�A��Q'�t��$���|�u��$�C݋ۛɇs�������FV�E*=��:h�1�d�%�b�����g��� �6w�.��n]˧�K�8.��senl�-�?�]��j� ,*�=�d5�qaE���;�4ƈ9���C@?����1~<��+�s�,}a"������+�65���h~��]>�x�#Qz�G��F�˄D���D-ȝMYO(e��[�����L K�4�X0D�ox�z�e5��8
��m9�۫�����Gw�W?<����������OJ�L�/��@���>_]��@yG���L�<ԐT�Z��vQ�
�%�̥?����'{m��`l�12-�&Ь%�옝�Y�*I�ݻX�g%�9��_��ztr�|�̼������A�Qg�2��7��R��ѧQ́͝O�<\f�|�"YP�~Ȗc
�-��_�stj��MuV6�v��3;??%낓ƃ�uo ��4�}]���˂ܯ��"���q]��<=w��`�VV�.m&`W��-�_y����&S�jI�~���ᘈ�?_������^��f�Cr ����f�ׂ���»�����d$��,�	�{��k�,�]'L��#k�z���v�[����
��ŒR���?��hpɃ��H���95�"~q�Ep�Q��ߗ����g{����~� 0,wt�>��$(@F�����-[����d/_��x|h=��Z�]�h��\)X�^{�Rl�{`+�B[�H;;9=�Ǐ���o�|Ax�,k��`C��c�.��Ff����\��Y����D
):�\wt��g&Ӻ��)��w{v�~?ӗ�Q���Y���ʱRplP���X�a�FM�=w����M��Su��=���[�c�Y�F#ta��Ρ��{� Gc���.��^��b����{�E��݀\ �a��Z}&���_�|}��~f�J�N��D�����åc���Q
p>��+Zע15��v�5�}�x�����w��8���?.�	�b.pt:v��$���rtWzy����˻�Y�ڒ��$i��B/-��!�4uv���*��Q� ����;��Ai\$*�\�5����%���'�U۔����k��v2�ɷ�Sa��8rvz$�����]~�`�^�,��=c����;c��!�]3<!7��I�:&��ׅ.�n�����K^'�y  �b�g5_H��3���9iXy�#���v������6��<ٸ.�Ji���_�*m�^9�_<{l��g��o���w{a�q��[i��LA�p}}Ko8Ȟ�ɏ7��-a�ґ����MY��ǻ���٨�]�`����-~���l-��9^q2��#��rAn��c�긜52����N�}��J�w�?���Ѧ����0.Ey�݂@�Sv������%�������T�0HG����0/=���b}�13Y9����G�-��׏�}�0Pc�)�\p#��/ ����c�,��������7,���AN�/�<�2S��9�m�%���<D���d��'�f(ޗG�Cwl{6ww6�ت�7	h�%��\��������ŧ��uӕ�p[[f��1�\.<0`9�O��0�9�-�ځd��$f�2 �݇J�(ʎ��onJQ>׷�<1Keju�OuT�9���ߍ��(y�j�n���ð�:����	<l�{�>����/l�ӫ�\K���x��p�-�Z��v�]2���h���r]�@]�tsW�n$�O�<3�\?��s�e>�*��^Y��>Њِ�����?��޾yC!����J2p��Ya�12��G��� {���q��4�Gf�2;��ѝ��(}�f#:͒w��z�Ɣ�6WZ��f��
����0mS���yyǧ���c����-7�'BxŃ�Cn(�50�j��&����g׉�85���#��Uư���h�ճd=�J�������kӗ#S}���k��unF����d���@�d�և�7}=��kʤ|��P��{���z|����#�\]]��x]��{݋�#{Tb/b%���p��^`Tޖ���k������KlC�ɸ����;\�a��:Z7���m�ph�=���-�@F�%c]��Q	��%�ML�9��[g�ǺN���U%_2�#Fӵ|�F4裶dZ6���1�⣗TC���Ý��%���d���~�����<7G���P�T���܏7/��5P����UO�<��ŉ��}���&�������&v���H>Ky(ק /�1-�X"������/%o k;�;�����٣�N�kl�Y���8+�;	|��Kr��\��;?[�_?���w?د~��N��$'���Q5B2�X�R'T jN���&e�1�2��A�Ɖ�F�*��ܳ�r�V�'1�T��;C
۬y��,h�䤃X�L����$����r���E�- � } ��yQ����r�X��;��@e2xid1r:z��ql�jb�A�f���w���(��w��V�Ƚ�1X�X����Օ<�w��A-^�rZ<2e�BԀ<�g'GgB� �����# �E�F���G[���Y	\4�Th�|�`��ۍ��(ABM�J�D�x"1�Iu��"h:�)Sr� G�
�d��Q����b^Rϵ��8�<9`�!�L2'��r�2,�Q�m�jx�F�ΞqN
�ʘ�~�J;Q� �[_��w�qrq�}\C�c<c�2273��;S���p��a=��������[�2���,���[gD�"�x��K��V�4i�Hv�Ϻ?��V�f����^O�?���>�
����S�,��2l}����_�,�{koN4W����l���� �x�\_qMo�!��b�r��FF|	5  ��IDAT��fd�"4F�������������3{*�C�#"�˹z�Nȹ� �? �u�NV�eS$Y��K1���N �|j�SҰ2����� �>#�M)5��)FӄF-�>�dg�\����S\�Ơ��c\n�]i�g���v�ڲ��y�_������=J��+� ~�f�N	b�|���vq��(7�0�;j��z� �����a	�l��xf��&�$77[�fܖg����>���7#!� ��3	lN��,4�C�'V �ٵ��Z�h���k��jF�PA�9�w�I���ͭg��܌:�
B6��`� K$�ۍ�PИ��<O�p7y~Tנ�0�1J�K�<Vk=���Or=�&/H��(���4�;�so	8Y�._�����(ѡr��5������r�NH$UTzv�lV�4�.��Įʞ7�J�=]JJ}�'h�7�9�c���2LǴ��|���<�ӣ�~x���ݯ��_<���?����x!�B��-�B�K�s�^�T��;;?Wy����kg��%�ؕ���")�<x�Ò�«w�ĭ?��wj���#�w$�Y��<�����xtLBI�'l�X���u`�[�٠��+SN :��|L:'� �.F��P�g[�W��&��LQ���@����޽{o��G���K���=���dbO�<����v��qI� ;:��}�;iqkSi��..>ٲ����3�������.�x�wo�ٟ��g��t�k�YY�ao�F��XB�Ndˑ�Kv�@?���Bfn���av��fd�8Y~��@�!9M,,J�,U�E0>������h�g<�ԫ��#};x&	T��x�UV�����QgˠCÑ��2a�����g�%i��4DV琬�xP����f@�|�d6�جA���7Fm(3�v�9�=h�Q�7���O�Q+�Ңܣ����J��7t&(GFT}�f��vb���y�夰�}^�����dE�(��ѱ��J�ؒ}�h��a�r��n�p�$�<G����Fɶ��=1^>����U��:RY>�bt0:I�b�gw���hI��0�����N��ņ��K<�J�@Ҁ��@� /��5�+(}����ٺ�*tg�e>/��)���������k(p��Ȃ!�%{�{��؝S?�;�.�9���}���ʝ��P�9�s6���� �\w�ّ��ɨ�����i ��S����V�n�#����x��5�2��J�(k}���$�i���ZҰsGv���1�%����sa���2�*�u�=�<'!�[Cd��m0�L�sl�>�V�:��'��4/^R3�VIk4�3��H6C,F��	�[M�S����e�`��Y�k�����:�u�=g1$�6�M��`ҡE.kq� �4<��x�������\�zP�� �r$��F|q~�,cuj�xٓL�灂�)X~�u�K^�ƍaT+V�{���Z-��Ӗ��I"+u��h�s������o����v�^9�af���T
�^�t�޽;vt|��	�NL�<5Qs��
��Ņ]�k Fb�W�хʄ����&���pgk4�s#��8�u'�}��x�|��X���z�Ł��X���f�f�ʌ;ߘ����h�ԎY�\�1�r f���rt�V����-�x:"ږ@�֊5����L|qY?߼yg/�?���?ڦ<t�].�6��<��Ǽ?�K�k������ѱ�� �\�O�>��@����׼y/~z^��SY�>�;������l̧�)�])�x��̃JU;x@��K�b��B� 11)��`�T~ZE{�NY�X#�����3>�|1ZD]&�Q�
��A�f~���%+-iP&�F��6~ϨMc`V�G�0���X���ݠ�:˄`|�u7ʎ�R�	�X��d*j�q�aw3^��l%<M(c�!1	G��D'�~S?���)�������`&�t��e����ԑ��8$yra�C{S�ɫ�K���V�|�,���غD֭�@`�S���9_��rn�+X��j�m�k�ā��H$P.y�`"w��ה�X�Eg��<ɿf�4ܚ9^��q����p��H�R,@[�0�i	��lȈ��Z�E]�1<|�s���E�Q�~f9��74�� w=�j%šv�5}�U{�h6����T���G�l�C�㚚	tH"�҂q����<� t��>�P�Aˈ�d�M7L��KC�VnFǅ{�ڬ�1i���L��k��Ό˴�]�S�ԒW	F�Ȇ��u`����-�׋��.��!5 ��sRą�|le3�a��ㅴ����L\�Zz���S�k�b����	2�Yc�� p:�jf�r�'��H�^s��ڑ>;Pq�!�g��	`������S�X7�{��7��A3��u���u��4��f[��K��^�4w*�ީ:�+ѴL:<�=����xr㋸~�(�q��*$���ĵݭ��;w��g_��Ky��� [&� ^F�xpp\@�I`��=��ZS
"�DGplE���7�ԯ�eW�a辷��i�iɛ"�of�΀_�1M0� ��DQ�^�#����[��"�p���Zv��bG�fG_	�G�g����q6ir��BI�Z��Ã�\,*�'>���f�g(a.�b�]_|�����1��Kjz�i7�_��{���=?+��vv~����n󎷍�ц�A%Kd��`#�f���~eBz^~�ww�����ӛ��By�����$>�e�E� ����C�l�ߟ�u5ʜ�.�vCZtM`AF	z
κ�I����@��Y+7��|��r19�0K�8js?>ĸ}.x� \��&>#Ԕ ����J�CK��(�:N��� �*�tto�N�YIJ:�\�pG��rXQʙE��.��P�'��í� �3�ݬ����%E���|��:�l.g����ַkQ�%5^��o���M�YĬ2��Z��N�I,�wߠ�An��v�n��5�\�a�W���y��1!m�l̘�e����+�J.�[�������#������ \�u�8f}jƙ�U!���'��U
)?{�a���h9l�K���F(a�I�5��G��Lu���D�u�J�i��X�X� +^���r���\� Cҗ�n�\���뙶����>�`�0�;%�����?~f������a��N�W��Ȭ�<KZǩvD��X�9`�{"q|v�|{oݗ�ɳ��n'I
�$��^`��G��4�P�:��$m}��u�!M50���=�*Fs��f`REvl�,�8�{�ޱH|����
��C3���2|�Y�q��zk�չ�d�X�������Ov�*�F#g���cӬi	�,v@ݱ�1�`�b`��Gs���"�]o(�CBsprdc��7y��w�ޱ��;��k��$ɍEh ��ġ/\S���PWޒՇa�R$����/��9����I�|1fp رD�y%g%�Ȑx(��쑿�����|gw���=��hB1������g�'��n<��%��N��kH, En������|^_.����,� �~�8�a�������9d��]D� A�H?;45�4k	,�=L��)���{}��?�d��=�j%�,���"_ҔE��2�oM#���PR{��n//m�6�H��$�������?�~�v���{��7��낌���<z�3�eZ���͡i͊�Mw�rR����k)�
n �<�)�;^��������b�ޫ���~b���ݨ%$P�\� j��jӞܻcg���؃Q��a*�g���H���C�77b��� �:��Z� 5a�,��O�#�������N����u|��؋�%��#��'Yf��4'm���-}9���6�Z��+>R�	
?ү�+�!�^&M�4E��+��Y��'��->�����vt�JǠ�FY����U�.�����<�\�;ϵ^�t4i�HӘqZTN��U#D���G��n'M_  ���30؊�w�n�UF�9t�q�v�,��9��y�D����!�DtcV������L��PdCn�VW���̓�ˆ�1�%��`C�?+@���y�[Y�w�X�@*KLδ�.�����إl�G��ٳO}i���m����vnQf�g8�#X�/}�t��o_��� U�3�Er��E?������s�.���ĐJ[��MbA�Mx5z.�ԤO_=*�-h�@F|�<W�')�&A�'|��b�fs�X�E�s��ɶ�H�fk��������,��*VA���3�:���o^��Z�A4���q1jͩkY�"M���&ߔ�l8�D�{� =���\mZ��<��5i��L4���.� �5��^uv���[߈�)�r��;�w�q��'$�ٵG�\�NB0�e�*T��d���,  A��̮�����8ı�7d��Q�����-��E7�����B��w�ڷ�>���A%I�&�
x:/ �.%�w���%>Ck��Ƽ:8�1��Ě���5��X�)d19�k��~B�����h�_�I�/�.h�����~�qV�[�sO��w���8Sȼ�,�Je`ƍ���6z7]\13������D�(��b�}����|��]Tz��{��3������ٳoi��!�ٝm���v���d�p8E����f1r��:G��&;-����s��x�����Jw�C��Y�c>)ٛ:u���|������?؝r��z������^ۺd!�做A�6���<Fo�	�<9�5/���M�wa������e��p��C��P���lO�>�g�ܱǏ�5zD�Q��U��±&�G����u�wx�����|���/����wM�����H_;�ܼ5 X)�΀%�|����v��A�a�N*���VG8es=���MS,�n\����*A|1�� ��bR� ���5�u�%Ƽ C���M4��Om� C��CX�+u���{���J�%7��C�[?b!����k�+X|LSlF�L��;����+7��CR?�G%�^�$��������Bz-78�gnX.& �a�υ�b`�d���.[g!L�����X؜�kwB�� ]��5��m�g��l��k���(3JGX�#�?���r�Q�֎�5b�ky\�g��n;FP�,��BiTI�';&�`9�9Z#����[s៶���ݞ��6�4�n��!�Z�ԁt�ZU*�>����~*�s@&��e1���t^��e� ����Y'��OE�Ai쨩b�����9h�͌��Ce�g�>�0+S&���)o��ȟa�M�v�n�Yluv��<5&)y7:�2��9��ؼ���4��futb_}������)A�(�\���L�J�s��!�(��c5���P͂�1���Pf ���
l�{�<F�"�g �yۭ��1e:�:�bя,�*��޽s���S{T�*4�]�M��r,3�N)^?,X�<1�xT�C}���w�[��r��I���/�+'&Ni�Z����6����1�0�z���eRMs�$���$�ai�K�J��̰u�#碏Y�$N��V>����^g��� R�9��0/�M�+QN����D�p�������_��~��_�ciE���P8�l��n�-�}uC{�B�5iZ=��3|#:ʔh������z��=Fr�I�lQ^�ک����q�5��9)7����ݵ� �K��|kן����Cy*.�s�N����*���e���K���mB���G���i����Z�\Ї{xo�'w{|���1X����=���cP�+�T��ؘ7��p����.6v�hg�N�{0��H���=H�͙���<��NA�g*9�E��3N�ٙ�ӊ4:Gw�C��D�M�/j2�>k��i\�Mx��t�5���k�k
�P'�Sf�C��6�
���k����=mHe+�jlP�Cՙ����,�M�ˮ8��Z����g ���a�"ZiR	��.f�)tm����Z�d���G���6z(J�,�Rl�e"6�;g�48x���J�)3�sئ3j��]�j�v$�X>X�^;�3L��LQ���P���,����k���+J��g�� ]�K��4��o��/����+�p�ޢ�a��=�D���Y�}�C��}Gg�V�#{�� &Gs���WsP23#!�� ����y]���AeP(ϲ�C�k�fy�=��:�8y��r}��k�[�7�C��C)ܮ1c��Ts�s�-Ě�B�@-�C�hP�����X���3g�kx���ޔ3�$�v�-	ʆ�����sz��'�Hxf#;�n�i���F�o\�L� �R���2���Dt����w�Ǩ�Z�d�7x~_C�<��~i>�Q��1�5Y)�e�<(�� ���r~.�./6괥t	�W������OJ&I���[ͬE�rk��N�%���+5Ќ�sž.��:dA���17�"��d�X�Tbi��� _��Z��7����94�ƈ��owY����3���F8l$uy|r�@{s�k���V~n	�����϶�|a�����ㅝأ�����o��_���߿KO��#j�=ԍ��C�xk�}�����CF���l���W1�o�)�T���޼���4&�o�]]���Տ�P��;?�������/���??���~&�¾��À[���'����af �����˗�����ƃ�F��j�HtN��gW�J��,�kg�2_�n_���?]�|)ڕM�T�|��q{@���	�o],μQ٨O�7���C{x���\�B{_�/so��Xsn��~���^7r��H�
�D*��lU ު�o�7����Q'P"BñF'","*�o
�9ޣi�`3x����7�1�C}(��&-�qV7�3��O���������M�����a-����aMPl��F�r�Qڍ`��E�q
���'��߼�1GCM��Rj�����Iӳ�ɋ�fn}^$�'6�Df>}����-?<ce��;p�D(2a|�	zB�jZSίT�ς�A���?�v�/����^������-�X�>;�KS�8cgx����l\��ó�I���?���������1JT��*1��Ϡ,�㛧V��g�,7@�Y�.�O�T5?22>]�^�1S_��	�%��PH��"�#C>P��nh�I��	~_Kű�;bC�8x�ʁ���fo�ٹUϮVkB��-��bs�����T_�j�a�DW˥�h�����k�/7~	�.vx0v��{��òŷ��7�!���FM4�`��n�-���H�/P�g�����ڔ�Ø{�CS�e�f�uC��B����֚٬n��o�C��3z>?�zF�R��H�a�	��ɻ��vऽC�|�,xp�\F��螋��O���r4����r"�[���L���Y�n!���ɻ���2���H��X���E�&�Oc؜�by�]퉄Ԃ�T��}P�y�)�3jID��Ⱥ���+{��u�P��3Ϥ�ۗo���	�=j�(%�{<���sv9�5�'�	�F����k���\���X1�6#�V�^^��q�YC G	�￳��{������0.��ݥ3������ڬ��J9?=�������Ջ������O����dɺ��\+T>xpV �]���C.�;'��;]���]_�X,F  Mzv̱6+9��q, iU��V�;D���� �L|8�ѝy�^�D'ӈ�iI�����p=�	N.���j��=2�{r,��1h�-�(�&��eV�.�ih�b��I{�G�$Y�#��jݣw���{G~���|$�V�L���
�3w��D�ܻ����Q@"32�����<�=#����J���������Znn�2�� ���VwiX��&��[%�(�B�	�H'F@�q�j�K��2w-J
��	��0ڦ�H���h��Ea�� � �u�)P~d�N��eag��n�*T���6�Q���j�ٮ�vZ��D�|�U)�D8`$:�N!e� �1	�7�P�]7�٠�6m/i��s��k�+� �(=+��ԋ9���5-�C5�/�>-���c9 �z���4��
�h��"~���F�ãiMW�Ϋ�_W���~���M����s@
���{J���u�Т�m�P��Oig~��սT����6�Di���e��1-��{�	DK��FZuND�9�s������R��@wJ��4���o�X���6;�ج�b����Bɥ�ӊ��	�6y�{�8���^��ЁN���^{+��@� 0
�כ#�i,��>�i����:(�L��A�E&���r�'~ǔ]?,�[�A�	EU�r&�a�|Z!�L�.hcq�!nJ� 1e���ٸ�Բ)�Ѯ�Y��U��n�A�dG�Yks�א�I���@�Aq
��L�N��0�����] ��9T
���=��Kr4�
ly�Y�P��}6�jG�M�m�}���N����Y�ףˑF��F&��`��F�MD
���q/��H���Q� :�gR��͋�Q!�`yO�ɩ�)@��Mh�+�An����29�ڕ����ɅP֧����]���_7�Q��LGȍy|8f3D���z3���e�o߾% ��傀�������[-P��kj��^���2N���	w�)M��p&8l@J�P���wX�2y;cTP�����:lH�,����pÇ��L��*��Uh��Tz���t�͆�@��e����Z�
�~�鑎�r<p� ���:g�H�����[hJt�K�}3!�-��mY�y�����������>��HW�=y\@����K�~�L�	L�Z��d LMo)�hF��"^���-:P��͂��m}b�P����0~(�X�*ϿW�d�
JJ��G$V�%kӀ*i>�p�����]"#�(�&oQ@��W��n�X
x���j6�M����RQ��K��5qcH m6gsV�F[�����h�05��$v�\���mU�yT�);����I^ݨ�d��E�N��mF�z/Ba5�+�����{�|���t�GK:Y+G'ʯ��(<zU���X�G�C�c�O�����6
#Hn����.@��R6I��xx�8��X�3�>��S6�nU�
�{a�°�(�GY�o�/�fWSm>Z����+H.t�-�[���2R�	�%,:\���R�?;V�}�5SUi�2O�@N��Tuqߖ� ��޶��jK>6�fU5޵6�?�u�(�2��t\s`�H�X�Ks� u�}�"��&�N�{�Sݪ7��RnoG�~�G�H��˰W��Y��.q	�H��#Y�x)]�fC�5�&sp)/%��"�u�#�T�U&sc9�R���G��;���L���Ч}��h� ,;C!��?!�Xyw*��x�C):�f�4��64fp���|�:�V�@��1��m�j�����ŵ1Q��Y��}o����Ρ��K97!W/��X�����q��TS�(��'P,6�t�<F�{Ed"-ܭ�9:>����@�5]	��[k�l����X1��{m��*j�#w��J��!{{K���"�M�����<��ՆX�ГZ��vz��e�P�o�J���������h�" 4�Զkv�_/f��
�<H��i��GE�������4��2@��VwJ�].�S�7�F���
�b|�1i#\Ѵ����(ٌC� �1.���Q�w��ɞm�{�օ~�-p`����8�\R��S��� ���"���B�Y<�m���¬��jM�0���7k'� 覅H+�R��
����O���ӂ��q��b��<�4�&�� �$�{B�4�����Kk�h���ށ�Fb�Y'7g��##_EĪ�K� .����Z��$x�q��0G����j���ѱ��HDO�?�W1Oa8��TR,8����-��{*������"d50)�nrN���C���WE�wX�X>��VW<�2/&���/��L�m�䜻TC_guQ�G�&Y)tp@�[�/?��{�u���Z%�e�&`4R�
����Ux_9�*�!��_�wF�&�
�5�}
TƟ={F���}N� ��a�g�97W�4]������h&���!i2�Y�Vz-#P<�l��W#E�b�*��Z[ʨ���~R)�������[���Ƕ�;/N�1][�>�ߑ��ML?P7}�q��\A�qLm<pIA��N���P��Ո��]��#�U$,����<"��i� 5L��#1���/P
kK�����L\��_�naT���^%!��6*���W$:��Z��6r�c���xi�m6Z�'H�y3#��;���� ��*tmQ::�r�Mn֙�������<��-��O�'��FU<~�5��V.��]-�H�6-䛨$
�[O����C��9�
�������A�$��hW)Y.��|y3ETi���z>blW��r��p'�2�/��钪�kd8���1�0�k���j����U�F�bw{�z/��,��Ao��j�0��{y|����C���֘-�(�y�w Ǉ�i�����M���H c%�U\��,H�'Ѕ��܎h����h�������J�t,��i-ݛ<��O�;b����V��oU*��.Ѫ�D=m�����x�\��Vfά�>���z�6r;<�h�T�泧W���:a�oN�$���6�#�Zc�&�8�&i9:��z��?ȼ�$sH����gЖ
�.=v��&��Ȅ\8��8nV�I@F�h-��H.la�QQ�ݻ�I��C�:4���j�#5\�p�n��{`+���C�NG趰%�G��:���8�,���bK�ˋ��=K�hZ�q�#�6����C�s1�ѡ�S �;��9"Acr������8�Q�R�+��b���vmM�D��i$uj�-��c���m��-�9���!6���|�4�*W��r������ '݌�Iu�	�>?�o���Ә��8_8�<w��i��LX�~�Xr���HzK�W�����k$L�ym�:�X�۠}`��.tb��e�/�,�~\,հM��U���t�!���N^�����ɏE׀����}Z'������L!�L���E6N��:�] �Q��2]��$}b3�&�� H��{�3��Uy��re�^�qҗJR�����ɉ������m�}8�Lt�!���H߹�l��v��-�G���C�����Y ��gG������-����Q[�E��T������=���O�wqy->}"��&R�:UW�#�Ժ�\�;S6H��Uc�U��h�~����,�����1ݟ� �-���an.m.��XD���V�_��j�E��͞X�! �u��Y��`�)��R�z�����]RD�y��M�3���T���jU*�@QI�s��� �5��N��Y�`���XT�%�,R��=S��M�C��l�
�˶L��J\n}m��6_���F\��[*�"B��GGY�!�c�QIQ�4��s��F��s�E���=���W<gZI���&6	 o:�ZgT���N	�b��	�C�t3Z��cU��(τ�������J�[ V�# �(��6t�P�'�K����%&����2 ��	W[��an>8�kT<\��B�4��y�0��Ss�x,����MH��T���sB�@�6�&e�g�¤lu��m�@���q�SJ{;���*��3 DA��{�͖�8���Q<J`�ĄwY�0U�5e����O���FK` ��͒����\����-%S��kհ��6GB j@�=�?�ý-�J�k�u�3�H�Y���޿�fK���N�uQ�g�?ݛ�H�U�@C��hUb
�����T�X҉���Z�="a��]�xeo���ϻP���Y�����z���kk�NI�59ꬽ#��˰�t���:K���Du��ˎ�&xr�
�9`~�:];%��9���Z��t������ѯѲ(LU<1������K
����1��^��i]��>�(�H]�*Ȍ���4�!� ���K������^ۊ����.��kڧ���8>#rjq��v�)#��c�
�:V/�5uLʆ��6�FK������L��uW���O1r��D�N�p���I!M A p���<�dL��7�{�t���p���dv�����'������|�����a�]��4ԃbT��s�/���0�n���{�iJ�����/�`�V��2�؂�~L�
jUpV��,��u*��(��2�SB6v�n�l$C�(�����^|Y��R��Ս{腾�C�w�S� ��:� �q�z�þ7��3�}{�n-
fr,f1��jq����}D
��Z}� ^kL��$�ذ�-tW��]�x��"� ڷ#���}w��=}ھ��Օ��t��^�~��^�h��K�y˖#%K31f�Q�]���h��;�]ݾ-�Յ��l�ޅ���w�"��I�r�NQ(���������P��ȓ�jޟ��z���c���~|n�"`¹?���,0H�,-���x�,7Ftdw�O�݈(�T�y�Z��sZ����Y��#�R�hQ�^�F�z��w�h���Z=+�	V�Fn�J�#5�^�
��6�{l,�_T��8�Y��oZk֞~B���'lJKz[��a>�^���=2ztx�Ǵ��/��ų�4����6P ��B��WL����o޼���N~����ٳ�Lc_N�k��l��b��j��XI�H٠����^>�~��y/��%�����E$is�u:I���I^>?`$�o_�"�c�����/NOO?��幥�:3�o�j��e���3�q}������4�L�ʅD	�����c���"� �'t9v�_�n�ݨ=�����*���"|ϣ�f��կ�E���%2���_uJ�(����bgQ�!誁�{���G�>�?�`�+�gb/���<}L=�V_#�؀{&������ք�:uYҼ:_T�Ģ�!f~t�b4�c�h[97H�����u���� 1��ԗF% �N(�U]��������J��������r�2�*�kk��M`�k��6"JɆ��/���|�x�H)ljN��R�" v+��/O�_��w��7��wOI�@K0�a���`3S`@�a�xB:j|�����s�Lv�G�`Kv�a{"}Z�/ C����Ǭlal �R���is�@i���M���5Ӑ�s�g���9���lMZy����_�E^�~�(<"{�?(�M���A^�i'Q܀=��=���\Nϯ�����m��<��52V����T����gG�"-T��u����Tև�n:�ؿ�9�춹�RVbvJTrʩ�P�bɼ)����B�ڊ��/�1�G�p��%����z->�}S/R j\kU:C,�T ����l����.�-,o��u ��pZ��z����>���X�j�4_�x��g4���bWB璣!�p$�*�'_*f~uf���������bF�}��!�Q��9 ��d��
:j�nV֡b�i����O�vmTK��^9?{{�[[iC^û0�O,��]凍Y���T���c��b��ڄP�.jy74'�Xˁc�~����c_6L�P�����Y=�����E|z�lPI�>j4�d�O�}ʢ�d�l�X�8R�0v`���H)��\"5ʶ�7>�����D��n�'$��kM��%��ųg���ɏ?���?��ɑ=���b�Hk�D㛎q׌7D!Ш��ww2��E돻��b�t�Uo~5��Y�@���	t=K�fF�޷�~���#Fpg����ѩ���hr�ם�*���k�p��j �*��y���S���ȴx����k3��8��#�c�Pz��G��&��)�0 �+��t�����9��h]֍�6T��Ч}%���Ћ�#eC����������������"�eU�rt X����+E�G
��I����\��{�҂���&4T���=1�hk����^�}GN��dp0�kC!�I�����;���_ț7/���Wrr|L���P*����X�+B�s�{Nm��%���3]����D��]c 'R��� 9c߼��������K9<����d�zEG�e\����V�Ŕ=%Tl����ե�\����T��zMq��n�}@����]�� �f�( �,���?'��z�G��'��̇ǹ�Q��� �:� ����.�:
�k����;�a�/TH8ȴA���ǳK������̖�B�1e:��ڄjT{mݕ�������'���
ě�J�<cfc��,�3�~����ң�e:����ۇ?2p�~b����C1�ڧ=�LE і[��k��ѵC-O����Oۻ�K���ٸD����zD2�8�ފ��%F�D	�U��\�'�Pˤ��a�k����*�d�c�ź�����<��22��!��G�������VXa⧍g�jõ��}�1r�@E���}u�J���b��ū�r��Y2j3�1r�"�0PƸ���鍶*<KWq1i
 �Z�Co�.ݢF6Xl%hk�H]�.�W6!%ۣ��C��diʼP��0>����`MeM�?j�o��D�h�u�r��*s@%[�[%0;of����M^���X���Kٙj�ph����w��& ��o������`�����[j��n�RJ�W�1���ʨ5�owo[^&O���w,�@q ��+��JJ��esrr� �u��c��T��/6��d�/.�����6`�=!;����W���}��C��3��+ �򫔜��ɴ��T2���U.��Go:��o�T�Q� Bk�)�QxEFٖV-E>���sȎ1H��5��s)6V��`fd}!���#������U�[G��q�h��{#�HM�ה�~�&�����5�H��u�����5D}�pt�z�\u���#]oQ&�<�t�(�0
�Y:�i��}hs�(
�NO?3���ky��yz��� ��*�~�+���K:�x��M&ON�r	�Ӝ�쀈�ehe�� X���!Cdub�1$j�8N�mM�7o���߿�Wo��pJB?b���F���D��d�M���f:
h���x��t�.��{to��H��|8��q�G����*���W�@!���h�B]G� ��:�XM�6*��=�"����aU;�3��Z��ʱ��*Ͳ�E[��F�=Cvx|~�\���,���;�G-l��"�<�Kݮ��3�UJ���dL|��׹�X���I#E�Ŋ6$�7=��b��T�μ��)����d��O;ˑ*�7��wBN����Y/�Ʊ�x���6�B�6pT�����Ci�I�0�0D�F/Y��g��p��y�4�b�Ѽ6�Ȃ���,RF-��|��21��<�6V�'\�_����a��g��5�?���Qř�o��m�g�%��E��V4""���E��RAԔ!|���v��4���p���^k��&5v	�d�C��/HǑ-}l�W�6>��J�u77��TH>�J4@�Z֊ �My��W �[Ӏl�N^�a{�tu�{�V�,NXC*!��)�{ZB�l��+�t��=N����w��e�NN�x�ܢ��<y�7w�r~y.���a�^�2�{f��)�y��w��Bb+c�34l��8<8�~u}�6��d��IDEQ�����9�4-g�'p[�[�?���u�g����g���S�a?��ģ�>�JH�_/��z�+Y-U��9%ɳ��������hTRZ]וI$���S-B�:$; 2l2�*�鸧�P%W~>��A�~�0m�9[G�<� ��M���Q��rz�/�X�R]�w���f��ϻ��9h�+0�թd��B�͌��άr�9�E���r��\ �/fsV�ȁ�uxxhN���⃃�f�\]��>�(>y��N����erz�̤M��.�v$�� �P�qil�5+��A[J���Y�J$�^�<�He5�H;�)���*?������O9{
Y7T�I�?9<��ݡ|I���Vm8
Z,������}�[&�I�׺�U��x�cd"�
�z�!��Կ�����u���@��vw�"X�E���\m�E�6����q��<�_ڛ��v�{m�[�����\^�k�O6�Ɲ��V���wǣ�ḬR2Bȸ��Ȑdv$6�3�T�K���uzSʴ�Ѻ��7y�Q�o9���*���
���&8��`p饲��C���������@>��"���J~��%���K�G;J�,Vq `�ĵ�Ԃݼ���1����"
������SZXK�SK����׸ms3rLz�!�ad�?a4�8y���H�x'a�(� @�G�ɃJ�[Դ���,>^�\ ���G�މ��zjH�X�5��wm��2	 � �X��8Lf����ʓ�۩��p��ue�l=L�ѓ�A��� ���1E��ň � `#𺠄��e#�Z+Y��)ǌ�����������T~�)�W����A�_;����;M���O������_���=I�lH�x똖s�#�4^�~��o���R? ��+��>~�$w7W��?$���HS���<��dL�u�_?�Xy��|��I��n���j��25���
y�WS���f�f�تHg��޵+�(�u��*$��)����P%���Gr�J�l��ĹM~}~��k���P��r���������<����7��S=6Sj6:H��w�s��R��~�Gs"wU��=U��2�J�N�U�=���q��EPW�õ�
@�Ys#�ٞ+V��3���UB�����kf$Pi��ç�N�ᇹ����MrtίhOY���%;iM�8_ճZ�� e	�u:�d NaY��]��y�����]Z;�i��p-5�-ɘ&<��`ha��l�-����d������_�_��}u���3G�ªͱF����@�<N�-�~<L�]<�����Ң#����1����Z[e{g��F4��nQ�w���A>~�"�>����\�u�QM3��GJ���VN?�����/��G���t�ymYd�Z�&��żg�~���a[���/^���K�}������C�o+-������Ɂ�&d������E��@�p��f��,������`�z@B��|�<�����J��ng��W�����
^�au���Y�B_��9`����B`�K�I� V���S#b���._���J����6)�-��	8��[���~Z����G.r�����갤�P=1�bF��H:�S�3�ygka�w�|�t���V�e%C�h5�zu�Y����i_�X�I����u�*�1(G��m�?���sr�+`���au�XE���+^���"$�����J 5��	�M.W�*JC�k#�#MGC��W/N������OZ���o���R���/���G����
Y7΀/�i��N����>�G����^3��Ro��ߞ�v�(O������A+-�hL~@2�(�@cvTA�\��|��n)�D`zO�Q�╅�ސ�J^
y����¤Y[�H�m�+)ݘ�\�)T�x���p�V�*�AV� �L�) ��_����V}ޛ�g4��Щ�B���e)j:r�i�͈��d-Q��<������5{
���m�:���G-���@�*�󜪀�]#}#���j�}>C;OS?����&� ����ɜT���X<&@��` %j=���ݢR�������:�����\'�t{sǹ2F�k��Z �	�FQ�'��j̭��������^��}rviǥ0� '��̵�3�Whk3Kv�!�A���A�QX��S{��� ]���[�,Bx��M�#vi#�?�������4�G�4$k \ѯpo�:��A�i�	����=�����w39O6@�\]��Z.�R;�� ޏ�0ju��ͼW�}�b˵��#�7P�����+M�?>y&{��ܦN�DF�j�L~������/���}�`��:D
>���T��`�!�J[��s��9��l#b��s"E��k+�N�<�k�v��A�@���װ��"���#z��z]�����r�����o=2
��g
.�,o�d6}����#��<���[�^s�Dyg���}�MZTwrq~ƨ	��sp�v���@�������gh�y�M��
���!;z?�M��>W�=�cB�
m���i��� �����^����N��u�FYd:��Zj�=��O�'͕�2m��k��=�`�d��wb�A��R����F�$z���f��$��b���]h�=J`l�˥����06��� �$`��lb��N������˻�����/	�A�s��"A��<�S�9��9;���ە|z.?\���ܖ���`0^���I�t(ȹ��?H�h����R>�B�2�K5Ȧ�\P����T%�R���E:6��|=�k��^��6�-W���M�kU̒�{xZ4"1�e�jч��zJ$�%:�M��8]=r_��Sj�� �_�/�M����Go�i-��9zT�ݫ;K4ik �j����0�v b���d��{j�KY�
�~,���u���V��<���(Ҝ�)?v0���|M����0�%��౱�����-��vR �:?��B#�C�{�8�찗'��T��#��.x��u��/��	�����c`���UC���/���� �b��0)Z��� ݪ%l�|��z����c���t)�{����d�)J�ڹZ�Vt���U���9{��|�1T~�˿�������'W�w	����˯���:�d#Ќ�� 'h+�Y6%��x�Uz@w��5Bc�g����!�o-�Up� P���J�|n�߳�to��b����|b�¢� `o�y+������?�~�Fܷ�������~[�p?3&�~�9AE��m�W�p���֕G�<�-����' �g�9e�F��@LS���x���뛶�������q��Q��Ye�!������8�w�����U
�	��_���B!:w�\�T��J�:�'�b7�j���@}P7��	o ܞ��N��T��O���s��(8_W�3Y�K.�$�}:kp�4��c2XaE��$M��5
�� ��htA�"2�FT�@�Q=
�F��F��Jqb�����"Z�O���˞�h��z����t~N��ʙ�J�N����w��ai���z�D�k��0բ*�XZ�� 6�X㘑&V1�U�Q�O���_�ɻ�����3�5����j:ML6À�%�[�Du���O�,�W	PA�̀*�_��ƕ�A�I��!�	�7a���ٽ�W�gL,��)3�:��/�jYT�L�Ͱ�;���]��j0��m���7��ΏHYټ��u/<�c�2~=�D�tg�m�z^�bk>Ư�s��}<�Y<�R9�`ȁT!���>O��U�sC޼ij����.���YG�~례��Ez��%_�_i�}���P�ԟ=��گ#u6��`���tA�f���"����[�C������p�F�Q���t���3
�*F��5��k� ����5�}}��l}�8��m ����Qg��J�֣tɵ���L�L�9V���Z�hVށ|��)/�)����o�}#{b��4Z%��t��~��l͹|A˺�+��m���:u�JI0ʣ.���
���1�wU��+��������@��B��1ʷT��Fh0Ɛ��)6� ��5 Cd��ۗ�{p��,
�n��ewkʮ�4��>�5�k���>��u�����u���1�SDVQԴ�Fʢ�h!`����X���lcꎚ�� �"�	���;*��?�";�����#��.��Ѻδ!=J'y�1n������O{x9��G�~:8��m�)�Kn �	��N����"�	����(~�V���K
��Ԁ�����)y;�[[LO�1k��.�˞9qhiE�	�tab#|ws��p��oo�`��������8o��Z���T�G ��q��76&�=�����az��l�T�7�F'��o��*��I�i�/V�����J����S�D/"Π.�S�ӥ��@ݒ�E�p�}W*S�J�NL�SK���9OF�o�Y>|�,�7�?>.y|��qF�����Ek����YPZ�Mfv/�%t0�;5�l��M2�x�Kre��+�-b����:��jDc�9��!�jW��ܐ2���󛛵G�6͏ϣ͟��"P����騆�k3 ���S�u��Vp��k،�T0�~�{s�NJ9�G�
8,�u���x��$�ݣc~�Z����)����z��S�O��6�� �n�h����Y5��J�4��GU~��F�8{c�~_�9�wCMsv���VVn<c�R;�4!���!�?X�k�F��竛;9�r���ӊ,�7Z��IܞlK7�Vm��rHKP�@D�q�k��́}V��\(U]�}�)��TRlM�Y�&��a��V�*��w_\\���ό��R�A��X���Ćx��݃��>P��og80
�]˝oܾwy�/�5��P���wEKysr�$�ɅU��[o�iq�c�b�r��/�f�8���AF	�k��xYU�rȶБ =�v��
�iM4��k��ږxv%�w�n�M�׉����'���ۚ}�0�|���(d\P.�&�!�9z�&&�M��+w���*[��9�ǜ��N��aL��z{>B��:s�4P��_�k�XNP�kg��6vP�I�с�5֌��h��h6�C9=����1��̐X�$��
 ����I�9��Q|����P��a�|�-�k�.���l4V�m�X�j��)�v8�j˳��3�<es�Bݘj�CXB�0.ₒ"*)�7�	3\��1�^zj�=�
����[��t!=̃C�/�u^���R<��<��Š3����habB��玖ڢ���)���|��҇��z���G��1
ˮ-�����q��x3lD�I�ST�z���z�Fr=����{��������/QQ����F/�_Ȫ��F��O,s�A��X@I�'|v^���Wr�jb���1(kMϥ���z.|U%���ae�$J-�6�_�������m���.�k�1���uV���-�+/0����c)�
�=���\�	FުT���#q~l��aI��lg��z�L�v�>����;붣׎Z�c��(��ͽ�i
�)���Q�,�BF'd���Ǆw"���fK��ը��lն�'{;ی�!� �{�����-�n�<c��^AJ���G7T=�>�?��/Q�H����69�H�ˈ|��8Mgg_��p���܅��U���*�{�͢.TТ$ޏ�u1ݿH��_��~�7�ӥ4�"�|�|�2�0[����#���ɽ6�>�^/Y9��$q����4'.��z��o׷"g�g���G��ݒ��c��v � ��{�B�j�u��E��f��[qXo� ޶SF� ����x��$}�D9��>X6:�{~�^��W����|NC�Q�7��䚁�����s��uic��X��Q�l=m����8�F�|�0�s�4�ü|dٯ�W�7�	�֯�$DJoM@Q%�83�Æm�9������)_�;�I�M��.���_�����b���錇 �B�l���2]������/�?�qX�uX�Τ�N���Yk�8*�GTG�S��e��]����c����S��o�:��op�V@\US�E�E&�����F����x�����y�'�d*�]KU�̩�sVM�h�*��iz۴�GG��n��ޛ�y�l�,�j��fZmc��E4���][�d�f�#j�E���Oic\��-x3�K@<<�U2�)
T>�ԐxCn�p-��X4fmN�S�y.W��FY�xv��5�C\o���բ�7�` ���U���}	�o���ܲ����m"uo��ီ.,�cd�p������n��ܪ�(��k�X����߇5L��7h�rn�Ś`_<�~�9:�d3�V_�s�4�1p�� H;����4�5O��w��5yI�qi�xq}MU3m�x�Vz��-
`���"��r)�wC�],�����^�K:,���h�5��?����M��� �j��^&@����M~���|��9��y��b�hK/"��9��Ѽ�>}�i�
��V��
�2z�u�1�#~���&�-��a�-���drDnWNI�4��ήL��+Z��'t�4MlO��O��/���^%۵E �����=Θ��V��k���`�ПE�L.WK�弾�"�y:y������R�6��~�5��{��9�&����/��)��N��_�U����&���nR���P��g����r����{)� �79w��,-C#�����̓\^�0 ��^u����s�t�0Ӓ�_�P�l_�Ŀ�>�Y�*��SP�^R?��;8�F�kb��h!�j�
ը���e�V�]~��0z*��_zԶ3'}�����a��in��K�!��.v�rdr�$�_U�N�����*@f�(�4;���ٚ*����0��
q��r-�O�I�uo��
l���XF4V�{2i��ؖ)K��J��Yy�F �IԪnK4�'*�tR�b�u�_3��ח��(�\W�f$${2���T�ᢓ�9:�7S���ʑ9�x���d��`��i}�z���4`�<K�KS����(R��«T�7AU5=�" �1&Y�a�_3�����zkF�q�iɝ����[[�MA�>��5��觶Λx���W(��������̎6�R�nNA�3:���^��~)s�ap�1`ĸ���~;�Gԋ�$���37���kh֏�k	O���! ��x`]�w�Q+�YZ�?�j�P���(���C�}�����N�׺�����>�x�V��������iUo�����W߱־>&.l�=�#���ڑ�y{�����Y�'}縳=��P��������;�O��&_ 7r�Z�7���o����'*��|�tl:^�� `5�]Z�EG��к1��SCb�lc���v�֟Eߐ��ճeZ��x�����#�TCo%w�'�i��nSAo (��ȸ=%����D%^ @�����￑���E`�i�Q�������A;P�����S������� ���͠5x���4�f]v�۴�M��=��-V�n�l���T������lɷ߽���]��t:J{�3?7��'Z:44�'���(��XJ>�#���d��l��{��|� �yY���(@Ph�5�v�?��AMd3X[�P��m��͐'|Ѱ�V���ϴ#�6�C3t�	'����nYi&F���(#]Q�S�������C���󥇍n@����$#>/� ���($g�M�',�op��䎋���;Հ�9�������䝠����D�ί�nnn��F�!��j�=������-�:��	��k�ЄU���
����k$��(g��s�6���Ə�q6�%4D�fI�8?%��c��e�B�0y!:������!+q7�;�'M�%�PRY��ط�9�m�ak��A����
9��S"%H�h����j@�Y�������j�
oE#
O�U�#���mT-!]����V��9$�=��g�C��7pԆ������5�,��Ӏ_(h���gY�e��7��
�\_��?�*2htUD���;�Y��\5 ��6������_�@� �u�R���d�.%Q�������k��Ӌ\T�n�S������m���>V�ju~U�_���f���C�����`��s��i�E��^b��X�W�U��=��*��� :�6�֪�Vc�U�I{o��Z����9%'�=7	P@�6f�Erj��������C������"��L���9}�2�3Y�g��5�1����?S���3-�Y��W�=c�ׅ�f*�\/�4m����B#{l[�k�u��=���;Fd4E��2#�m0���
]4`K4��3�Z����oS=2�R�4����������Jߞ졎)וE���M���ӱT>"�����v�iL�m�|����X�Y�:&�fk{��C[V$�C��C"�?����Vk�0^���������YD4���J��s8��
��vh���
���� ̨2��C/��#����ߧ%�W�ӱ_(}�Vm�&�}� �&u5��|�HZ̄33u�~���Jɶ2�V�G#��-Q�1�u��FxO�/�kL���HG1��Q�5�@5:��u4z��G�9O�ސ5r��,�w핒�Q��2�
N����$���/�T(�֯���(�|?J�bxi�� �]��U���a��:¿�#��e<U��L�q���9z&^Z�C1��D�
`�>���D����xxt��a�#�v�(�����AA�KbxJ0������5�þ3���9Y�9y������v���ă��\�/����R���5 f�?�Zm�SUXP3�-*X߾}˔���0�4�՘�3�(p� r�#5��+6��-de�eZ��d�Q%EI��	�m�)��i�������S��g4�^�Eʲ��e���)ᑦ�ԍ9Z�C�7�G7�Q�'�3!��A����^Gv�;
�n��$���;~����'�򨁄~��x���:J��B����o^c͗��36����8���__G���~��9�+|�b��G*9���m���+�����˼����6IFOG��i�u��1ޡ)\��b�=�����VH՞� /�n>.���6+�'�|�����'�����`���M�R�������1�)W��_�V�,�X[��5��Gl�|����v�5h?_<�JSԌd�������,�'�\�lv�߃���wC�{�j�س�`��RE�x` x�Y����־��U�"� 8LGf�����j�r>"i����-<����?蜭�zL�%��kd��}�?�L�'-"uH���>7��B��m�?+�����
����+*�s��=(�C�(Z�d�`eb5��ϣy�i�<�cߥ9���K�Ѡ��~]���K�MS�]QP(�@��U���פTP��/�W�.�~�~�G�����/߳�Ѻ�5M�%2����Q,�'D<��]��)�����SHӀ��qF���:L��U0�kF���X�kl
&�/e^re�so��<���A�k��6~6I��j�V�aq�o����� P���0w����E�ǃ��x����*���l��!wh払��oKP�]gh��n��h3%zD)��R���h��PR~�F�����A�O�^�ko�x,)"W@W%�B��fKb|_MP���!/м�7�X�fV�@�m�iZ�>�ѯ�`�⩍Ѕ�aec��>P 2���W�@"b�����?�QN�O����Da"c BlE��6��y����O���	����h}�<ͻ�n�r�5��Y�f��?99�&@Q^z�����͵|��?�E��E�7�>�f�;�Sl.4`��9���C���ҟ�rc@�A�N�D�����?��WU)�EG��r��ߊo�9��7�N! ������CNcK�YE�ks��fOL'��S���[� y̏��Q�߫.�p�G�]8ց6���0l
�"R�Y P��
�{�hl��P�'6�s�A�^���5�]��B������[�t)�: � �x{��SY���n�z�-��Z���B[сה�(H�-�
�n����^~�9L�J(��'Gi]�6C����6l�K�Sa2b�)Bȿh;�ƺ�l1�jt��+�M\#"��ǰ�6��?~���>�bNEa�	��1�Ħ�9��NQ��8����O�y }��x�v�C볝�=y��B������^Z� R͕��`}д#�"���[i�Vv�hu��*?>�yuw�QV\/[��q���+�Y��+��pl��4p�1�Kcu�����4�,�F(>�f�xR뫋�s��im͎�:U� ͈5�H�<Bc�\�v����a:��N/
J�	9J�2�>�9��Z�*��S�B�����$	�,��RG���Vt<�Ҧ���
�2%�6����+��'�І�F��0����1�(_�oy��͛��Ѣ+*9a�󜸓{��}�5���aO�G.����W��N���˅w�L��3ϻ�U`2]�$P�)(��szz���q΅�q�Qj��	�cm��,C�隡ƚ�&�R�AIm���V��gJ����4m�)��b�S4v��4�e�^�_i=���vedF� �}��m顔h�#G���Z=�Eb���>�ύ��qB�[��y��68��:�k���-��(a�%�������Ǝ�Rl���l�b�#q�Ϩ>@�8�op��<M�~��R�W��H������Gc�����#y���|��[�5��$�K����4�u��7���Uu�8�F�D�[Ш�/�A���6/����W��tW�O��xĨ�/"���ޯx^>�cy�N�?em~ۤJ6fbQ?r8�C2}[Iz
�ɼ$IK���:�W?6#a��ysQBu�%E[�^�|r���u|�n �y��b��8���qC�k��ő���E�;�u�q��ш���q�駟���gLy�Q�� `���	x�1u���L.�o�s��c��^�t�bU��n��dKo..�� �W�rw})��ѽ��&8] ���C�y��=����e�-���
��ۢ2MM��n7����ۡ#4����o���m� F�
�c��^���/mI����%	�v��յ�^35e��8��`sK���N����]:���Æ�� [��I��n��{k��_���p͔�,x�����Hũ��"F.�ހ�H�U[vv�d�ޢ�����!(Gv{2��>$wh�=R.��=փy�)��S��V �ݍf>}>�ݭQ�]6S���ۑ4�G+�7�q���D(���� ���	��̛��h:hP�#�(�:���ٙK���K��1c�����]0��W����7R�_�����`��	��_D�+M�D#�E[��C�+6^Vo٦|hr(��,��s!ˠ0#�K5<j�ܒ��.�yT/:���)M݌��TVP �|������X@T�x�@��i��/���#O3e�U�\�i��e���g��w �א��͐2�Cf K�k]�h��Ҕxd��Z������=bO*�K���1g�Ta�ϕ��DD��-!j���ͣc8?-Z��_�>t#F�Ab"���3/�?1ϖ+#qb5H�h|��������fDrm4-�Z�����������_�|I5jL�M���j<&ɓ<<>�
>�	�q�j�C�w��Q��T�*9(��{Ƶ�j	7�T��;�>��D�
����b5��US��c��S l@������?��D��8`F`l��J�O��S�`-�Pw�r:���;�3f�6���>7!���\F���#�nm9�`�u�6Ǣ�0�56����u`�״�%sy��?�ډ6��7A��m���l9�z��	_�I ��cgb�XzEi�b�{�'x���������C����{:�|�����C����>��d&���b���WN/R]����e����7��yH�9g���P���k��ɳ��;wh;���$��=y��OF����� ��Hk���`�Ѓ���&9�wr}uE���`k����-k����7o^3	 ���i|W�N����T��Aŵb��ӹ�y�R�����Er�V��Y�U�ˢ:ʈ�J�^�� KW濭+�KH��F����uAq���@��RшB��QG�`:ڝۥ�y�j�T�`�|��R(�N��c��*�^�VTF�c����(��8E�	��x+m����b-�>��q�����	>нO��d��	,���m�~�F���+� u�Iy[�'���4�슠�b��@ܲ���� �o�+���+Ri�� [o<�&sc˾hU�U!�([�*�T�XF6#�bB_lx�Pd�Z�V�&+�m�e��"|~�޷NW"�d�mi��ْ�f����H�-^]}�y+���а���X� ���~$_�jA�<-��/�rqu� X��d�1�g<�a�q\�%�Ϟ��$-ʛn�MtM�&�x�O��h��r2���EkzOj2��}k�"e�ſ������H�5�����H�`ʟ�͜5m7��Xe5�0�9��;B�࣏���;�Z�-2��C5*�y.���$��˛�ҳ����!�^��s�e����eeӭgӜG�>�wx�8-VL"�4ʀ��*�t�Q����K^&R��{��|.��n�"4��a���f9J�>/��ZK��I=T�$��x}!���7���m�/˳&�(�b��2�p�V�9� ��r
L4Z���K�!�4���P��:��E��g7�Fե���&`��x�{j�T!�Ʊ��e���k����h�O�^p���@����~�6��ij)�QNbk S� ���Av0�W:���9`��DC8%�;{\'� �f_h�c(����g'��z�q���am����H��IZ�,�B�fw_��Y-��gc)^ �yZǏ��zS��'�B����cy�*��=ޮ��� �$x�����V��p���i��5�Mδ 
�b�ށ�����P׈z&;�����g��t�i�ONX�nD�9�Qr�,�X�;�v�{��`E��YF��3�FH��������p{�y�$p薔��=��tXC�Z�tl�d�{4�;�A�!�=�R��,�ި*N�g��7@�p�9�(�)�s5�����|:�"�=؛2u��t}�Yi�������*S��v*'J�^l�O��L߹�k��ɨ����m�<R�����xͤ�(�ݳA�tI�H��5(l̂0aZg���f����4b�P�{1}�����w�7���3!fp�H�(.�w�X��xx�L�Ң�E04��=��J�G���b�	�e��r�5o�J�(T�ņ���~s'��5���~�ҏ��^ڠw� �X�|v��l�r����Z�@P���W��%�&�ڦ�G�����)�h�h�r�*�:[d����Z�r�ɵ$�[� ���5h��+=+f�}���y��NRw��}���
�Q$��#LO,1�,�lQ6��~ �Л����v�P����>� �ɋ�#b���?�,�1 :���D
���|����r}{�mD&S6�=<Q���CC��;1��2R7f�d�Ff �d��)R"��1���x�pp*�Ye�kQ%�h9���Q�|P~�a�'Ȑ>:��b45�$�Wsij�QZ.?�{��>k��ע��5r�l�7��eQNr3|�9	y�L�ѹj��_k��@ʣHA��s�j���4��(��I_RwE��5A�̫����4�O�+��|�Zt�1<\�߫����%=2�H�e-�E�=�6R����P,��k(1��x*q ��x!
����B���(N�������������SL�����+����@�û_���-+���-�:r<a��f��9z"�U?��U���¨�a��qe�u�`�#R��V�ۻr�~�lmS3�|�H��s	 �����c�@>b4�zZ���m͢*���[1�Ϙ��8.���,�zkMw��AB�ޡL���� E�7u����!�S��p�7��(P�
=��[ ��}������tI�/������kyX�d�c��7c5�"�u�X�"�� #i��hH-�߉����
�	�X��V�������(��հg�Z�t��w�����t��ۙ�ʵ�����f� ��!��B+�d/�5���l<e�X��RޤJ���,��� \j�Ϟ�7mF*����[*�.�v��-��{�V)�If��ִ7t����p�4b}�Q�_s�|��tn;A�1��G�I	�'<$��qA˹���j�o�R�U@J�ӌv��p�`P�UIv8��U�H�6������>1,z�6���MZn-ɐm�0�5�l�*�HT�4,'#��^���$hH�ú�*̃RP�^p���Ѐo�u��&G9����xT*�aM���P��Y�߭/�(J��Y$�+]T}\t��o����+�[4�e&���A���[hب���'��ߓ4��@�Ԡ!8��a�xm퉬1�I ���QFVC���v� ���%����6�-9yԶ R}_ξ�� ��C���%P�%u���e��w3*���*:�c�*�����������+�d���2�Q��=���[j�#�Qyt��Dq�;�ё:�UG�Ꟶ��s�l�u4�+o�`e~J1���*u�R�_�n�T�:�N��Z�|��W�����#\��?V#'�%k�}Z��`ˁ�_k}ݛ��ڲ���vʸ�N�k�eG�֮��ޜ�U^���i]���BhJ���s:C7�36�h�5P�����kV_^N���S% �i����j�dA�k<2�.2�
�! +Nc/��D�78���f%�R�#��mF��z��&a	����]�O��H����t���&���݌k��ܤm�c+�Q���<}�B~}�+O�=�;���ɖ�e�4ٱ��GF�q�β Od^�7Ftʃx4��e�f��bA[�@R#�����}�j�@�h2cO��d/w!���"���l���F�Z��k�?D��\$�|vu�� �  ���N���B� �
�h�Ć��N�c��[3�ٲ���., x�k#�{ ֭h�U0�<3"H��3j����b��5����cm���$�]�E1��,}�γ=��,��\�z�74��kXP�t����N�J��IKN|Ǔ*��^]�`�j;�#���=���m�F$&Κ��U�'�V�2��2V���8�oQ�]7O����o�M15'	M��tHl�wg|3�$>���15ʌ�U=2��(]OԌ���gr~~!���^�}<K�Z�s�x����bn�5w����ࠠ����*�$��1�.�q�:�C�:疼��Q"��=0���3pse��"��|�h����Y!�����-gݖ�t�u_z���j�u��]�;�N��}ǜzm�8���QA����Z��e�Xl��ݑ�{x|"?��'y��~�k���%j�G�_����bᡃ�q��T���/���?b��m�+�;�����a������iZ��s���8��
�H���u�@ݗϟ��������Ü|��^�:#���ܾG��d��`���{ۉ���ѕ��Sq�|�8��^m�9aQS�B�� e � �#O������ٿ�&G�
X�����1�ކUTI׍~�u����|�*���uy[����S���C�ڣq 9�S�o �1�pb>���a��ϱ�4��mF�r$S�~��'fz��f�����^��7oy��	� � ��'��iM�������e��c�p"����d����mc��msK6����%�����ͅka�C���x\ek�Xǝ;:L����'
Q"�	$|܋�ӳ�V���������Fd�`�0;�ynK�~0�5-�D��/��|گ���Lcy~vFG����<4����Qo{&;z8�a�@�ܡ��d��o�� ��r�>��u� j�5�u^���}T`&�{�K�Ţu~��ś����39�����}�(���(��f-P͊ԶO������s�5��s��x����;	<���\�=�����#��Ջ#9:ڑq�)W�o�-����g|q�m}�4TY�ŋ
�3FS�
�T�YU	�s0��L��vl�h�N�M�ֺ��,������`�=p�XS�z@i=><��>h3V~]VD��Y�W�� � ��w��kt3��;M���D]�d��F*��Ȑ(â���cT����@��DTa�0"�8i��B�c�F����^qo���#�b��?����H���|���w�?˗�k��L�r"}��e�E*i�� %�k�\ۨ�� Y-��3Da(:F�X�f�r4���
dj�-�	7��-{AU�3j
���Y�>܈�a!;ɍo���aoZ���g��t
g@p��7"�_\�apzu̓��YW+�+��[sV�^__'c3�W�f�~�k7@�9"c ޽E������=$0���҃�& m#x�0H�7"b����:+Fy���d��VJ��i�V�'�k��E����p���*��nV4����`@${h�Ջ�4=�6Z�����W@*G��M��5�h}>��ڔ~ȳ�{u���;_˞n7�q��G�k�/Ѵ��k�=*��k��`ɫ��q`\7Ϝ���U�I��p'+��m&�VE����+���s��ː�&l� ��v����#���#��*�z��ԳZ����8��=!�]7|�^F�l���Ԇ��=�% ��̺fb�i��jAS�,3�:�q��I6��{H��ޱ�l���:����ڑ_~�U~��/�����[n��	|��nۑ	q*�R�ҋ���D���ca��A��6٪�d�({bcS��:����ӹ>��l�v��_���)�)��*]�\�#�W_�?�% w�&������������d:R�~��h㶽��ƈ��5��H�E�WW�JS^�p?�J�R�09��!�"� @�na�R����&a�
t�~�5����ʯ�HGx��P�Z���i������Z{��2��=�zhǚ���HoT�3cKI����+)�;��g��R����O���Eq��d���!�98>����%�I(�bMs��o���	�fT7D�f��iD�$X���\�ik��	iy���ĘN4m�|4��-�g.x@DŘ�l�И��nz���x�)�9{1݌Ɉ� _	t������t.�0�fJqA���$����ѳtN{�34�}�"�yn�S�Δ��E��*Y�+��f��g�e�&���9�1
Y��|��Mk��y�~�	�|?�f�2��d{V�Bj�5�_��v��d<��<�^��F���>���FD�(�x����2MhmWT���%1�Ol�B�4ߌ���,m,�L������y2FM��	�ݧ{��t#_/��b&��|��ƍJ�yC�%K����س�&��(!�S*��
o+�]�j���^�e�`��=�>���}�=������j���n������4OFy|ï�RK
��[k:G�)?'�; e��Tz
ҁ�����$�2nOE�r�����7M��KNd��Y�Κ�V�V���:�#|z�@�7e-�`j����W�qw��ϩ���9�ۃ�|Dd(�{n�2ww�i�f����C��zy�+��>������N0�ƨVTm%�TK-^WZO�Eǔ&$! ���vL�^m;��HӉ�؈�!+�q��k[�t�>|������w�k����B������/�kV�����Ȣ�֪�E�LQ;e�΄��k�j���R�������^�v5�w����t�_�(�/����ޝ\\\�gZ��O�\ự�nM�Z͸�+�u�^]���5���ZĖ��(�ȯ�wڞ)���-2Jk������K��o��W����gt	�GTK��ˈ�3^V=T9w=%i�p:�,Y_���((��������~jȋE����E�����0C�1�M ��X,&xf�������J�ުL%Eyedo�v̭�2��}�}Qm�����Y)i��W�7�,�(k��i�K���u�����J�� ���4��I�B	X*Y�����S1=/(�MA����\F�7��\!��,ѯ������K��d�fŞ| %W�%DŐ��@����_:dM�wc�<�h�^N��OrX�ӟN���_����>��խ� _(7R;Z_4 �M��E�d(I����$ѱxӒ=�2澩5&C!���gVH�C�QJ�#(����׆5�6�v�b���'/C�N=������������f�����/A��SZ�6[LHrڙ�wH�\ȗ�ό�q���GB!Q��{�+A5t��<�.*1�����	R�ggWr��K 2V�.{�2{����$'f���V��jD,Z�����s��\�\��o�p���PE��>ћ!kj�FY�9�^[x�su4�粨.]�[3O��$����ܞ�_�x��Je�J3�U�]c*�s��S�d��fd�#Z���<o��e��6T�����5��y�R��O��T!��Ħ�>_��J��{\ۀ�����e�~oV�jT��Y�֗+��R�U¡�P��M]�w++$
dw�b'rs}LP2���G�d����HN�uZo?|�������ś�J��?��_�1媣���'�B��.����l�H������������("*������D�J��'��EIj�A����	+-5}�N!6v��,������р�l�@�l� o�|�����5tN@Rn�]i��ֳ5�'*6������R�*M�BD``��� �Jq ;XfHO̩<����dF@������׺V%��)C�L�D�L��hu���`�xB��J�B6��p�-y➂tePD�"*P�1	������G�~��Nd� ��.0f�Ǌ���*�W�L�b��E���>�5�s�}����ކ��*���X��'��0:��ˏ�E�m��ߦ�r���"ͫ��x�RF�I5#�	�J!0�����@�� p�u��4��s�'и�7�lf}��tU��*C�Y�hP0�O����n~�Z�Z;QT�l����U�M���L���n:B���>|�,�ϟ�"��t�%m��Jf�I�͊G /L�E�H�|�l�'�`�aŝV'a+N����p���P�E
��-yA���.d�,�_~O_k�X�HWYǷ�Y�~�J��j�W��z!zǁaw��@�曔�k�̼�6M{
�W���5y�f��f�i��(b�2޳�I��/��<#c����77n\chx��({'���R�8�ǅz�����2�����#S� ��\"=����1�&����A,�e@0_{I�:��I3.�������o�*��4�eY�=5��m����{57���kW�{���1�!4Rlt�s���uڲ��*=�}�{�5��v�Yr�`��J}�:2��]���������)K�|9h�y����1{6z_,r�c�] �����\��IiB��+��=��u[9#���)6���͕6�II�͐����`gl�m灖;?�s�����ո�P��ގ#V�@{N��O��d����1U����׈B���!�Զ���*.Ԁ��3� �`��.�@���J7���q�>�M�'����~� �O���˛���ӭ)+���b0n��`
w�� �N*l���`����S��M�¯#?�`�q �@�DJ�F�����#v @J8�o�*&ު�"���z����������	���ճtm��?���&o��V��v�+�,8'���{��ujcq�\^�W��4+U�k���R���9v��<?��X�%Q ��dl&i���	[��I����3�wo_����ҽ�t�bŨ��h8K�]�Xx�&ςP�O����jg��1�V�m�_�ppi%�5��[��7��Hr�+�s�@���9����'�0�O޻�E���(�Y3�	����P'�H�&JLO,f���Atޏm
|���~m֪�G����b{���ϯ���bӭL��a�daE��0n�
i�#g����'��/����U���oՊ�5��B�(�M���@80,	�B�o1��N��(������%���Y5nn�{��WCy������؛vGn,ע� ���ԳԒ�ѱ��]���}����k[SO��Lk�����(��]Z�d��!bǴÑ��s9��^���,m-�ͅ:88S�������I�׺���{�������oQ��`p�e!�seP��׮�,�a�.�ϪGļc����bF�6��D�u�#H�e l��a���&��b�h�Z�¹]>$�#Y�4��L��P2T�<AZҭb8�����g�����Qo����<[[�H?;�5�͟���>������[�=�E��Y �<Cς��^P�ߧ�z�~={}�G|}a��d��:���"�ڰ�������� 5�6����?��u��A�cY�X{+�d��s����,g�Ρ�gLa����&f�����'*_뇇��ҳ���Ȼwo4_r�$[<R> w�{9!�SK rw7�®�� \(�A�1"�Dҿ�������)���k��suxx�i!6�?��g�󬚓|fA� ��g��O?�۷�����(��{+�\E����7x�IP;�re��P�����Ng�4�1W�6��.x�
'[��;&��-����X�ك�O�=hЍGi,תa���\��p�h��Z��䧟�_����G99;�Uz�G�g\�X����h�9S~N��n5J�ei�"¨�Z=���.��N�8������OcJ}��.T�.W䉻����!ԅܜ��8�Žݎ΢ o{GKAP��|��1)ft0BFz�4�^��rٛ>�u��^�&����$à�/���f�_��J?2Ag�� �]P^����/�?$t|�6���|CºG����k9M_��3�����,���çB7�\��k�fk^m��߀��\W,\�a0�c�( ��m��&@�N�4Ṹ��O��W���\>|>��®nQf�r�� 7h�Io��.������mo������X� \NU�L����~�ز`�N�2t��r�xΓ�!M���j�JQ��	^h�\���R���hq{1F��PP���"+M^����WIr�PU���c���jJr�����'J_h�kƫN���=�0f��A6]�j}9����( -���a .���}��W��XJ���|?I{e	�s�R�����F4�$��# �t�\��}�>��D�A�����T���8C3���N�S��ߒ��?}�x=��?π��I�������կ�}�;� �B`�핪����j�tMR������*�m{�j���[�߭�X6yJ��)�����^,��:������Ľ{�9-a֘y�8�ƀ^���<y�̽+�ͮ��	;X����7Q9�h���Z����96�7a������r{�m��`ca$AA3e���	j�g�B���ZV0�Ty#"ه.$��PMJz6��k�����h�P�����`�<��^+�;Ðә���y��02�ؑ��ac�nx���} @���ruqAY��Fڍ �s�y��_��<���o��_2���)��S�&��  ��ᡜ�8���}`���J<JU�ϥ����0Z7���Lks����7�7�)�>~�\Ĝ�W����{%A�n`�mp9��DM��Ku�`.�
p4�ޜ)K�����'t m�n=��{����Q����y89ڗ�/O����!Ȱ'�0�U�!�u`�X��G� �z`�G��^��ڰѺd=���br�N{,y�<G����O�m�A<�,+#?|�e�ʥ�g$�p��U����ײZޥ.�T���5�dC�����]�5&���YqP5����t�b
�Ds�r��2"j9�ǔ۠��\)�{�Ak�Y?L���M��x�+lER����\^ަ�~�6׹|:����n����nҭi�'��<�zəN�߄,�H�_�z�y��e1��{T�|�����o�ib�`�g,ؘ��m�מ)�E�~�xig��� W�#�\a�@�L��m�fРU���
!)I�eC�y���_��}��WH�ֆ�\r���&LL�z�����Ҥ�=�bks+#�o��{�02�B�Tu��]���m݇$aE2oLV�
!�e>���)���X�A��=��_�q���I���:oǬ9-;5"���T{;�������G�=;y���;�.�5���������W�{��޾���5J~J5`�>'�{<?�@͕imH���f���lO��z��B����I�/SO��M4�O���ږ���E�����-y�n�m_<,N�أ1e\����z��F��"!����j`z���y¿��s'��}���ٿ2��4.�F%I[A�Qc�ã�޾��o�0�^�D}�3�P� A�:ue �3�����f�z**!�b��AAWq� ͋�)�<��H&�쁗��7�.��?���|[P���hpW���k7�Ҙ��	��ƌƿ�e�X�&'2�Q!� F�E��=�Ցi��Zsqs+��Q>|�� ���K"ΐo�v&�\O2��1@�Y��L���e�T�k���槏&��Kے��_�KÞB���t���;r+�\���*=���O�ٺD��ٔ<k=�D	�7y�2_1�����yJ���_m:N��!�s��_��qCg @��J��C2�'�ք��\�kxXM���Á{N�Re�.�9�md�U7$]र�^IM־�ů��676,;lL���Ԭl�:�YKaeX��?SK����]Dt�~�7I�h� �fx7>��/�0XR`]����l�D ��M�d��G=O�����ņ	�88���y[2�Q>��e5����{��Oev�c1&k���^�ӎߋuj�-�[a^-,k%W~nl^�=E��"F	�b:���]�u�`i0*	W�/`˅���������D�{�i�%�\���8�P�D�ig�/U���\�8�����:���C������`L�\9e���fgToE��y�B�`:zFn$C�P�j�	ys,��|�&+��سCE"<�/���E�D�ޞ�ٗ���@_c $"2V��敏O�����^?��W?;T��L��y:���?�T��WT��?S����)p��p����yu���9�Ǵ�t￯Cb۞��z�������yN����cfoj�\ḑ�j��-�gc��ޚ�{�E�
H%��A�5����
����q��Qs�����������W*�~��(au�C�V%�����tm ��iD#|���&aü��m����W����_��6��!���}�8�F�H�su�0���HZ��<R(k�pEn4ܸx@Z�z�^��@�W�	%O��/_����]����C�܅w(8��������_����vrt$΃�N�]�SA��4q�5ه��t�YZ��5:�HB������e	���O�oB��k%Į|�U���zYcT
�M�Tʷ٠Q�F�5��/+s������<<eeX���bMz�.������\�>�������b:t3 ����0���g~�=Վ����*Q$/:Ԩ��[�� g|͵!��f�{���B�A�q��O!�=�;մt��Z���.m ���Dh�H��Xǔ��P�ȷ�_��+`��ݎ 	��fUB��S]�i�26ZoH����O��zmܙ�������v�C���&m2��x[0�t�r�mw���MV��7�2.�<���xĘ-� Z
0����A��si�����Nߡ��$NTZ��ث;��P񀅐�M��L�I��G����gKί�"��\���"�fȞ�����Y��d!ϭ=<��˧��Ȟ9�M+�q����Ҫ��o�T @�{�tNEkz��9��[��h2��։��7�P8��J8ڕ���,��
���"Y9�GY���J���Ëe����99!�[Ys�|��\���1`�;a��	�+�=���������|��ρ�<�^t�«�Ί�d��u�i͘غO}���;�j�ISY�m҃
��z��(����U[�ո=��[�~�t'�X�w4��_�=?gF�(MN����'u����G
�*F1ē�գ��;77wr��B�>�� E;���15l	�9��r��N</n!n�+
�)��{�z=��'dGgz���^&��u��up|��1�Y�P%=a�� �\�*f��y� �����l��nl�hv/���l��3���7p^����3�d��0s G-�$G��	0a�wɹ��O�c�.@(�yx��Hc�yx`��ݫW�w�b(O����d�����Kh'ܟz�1&M�q:%�&����F�^����*�����t����D��Q|1�ŝ���Ӝ)�^'ؤ�����;�U:T����0z~cõ��z
q	�oʆ�Y��a�_Q�Z�������ҵ�UЪaє5�ƪ(m|�=5�����d�(�[�������$�k=��/�m���t��A���>o�?�Mu��,��u������q`vl^$J�"�`H�/.OT�V<`�:o%����V �0�/��?h�Rf���a�4��H�'�������O�� �l��՘q�$d�GaC3՞\<T� �.��]�ju5����!!�]4����e3�����{�ez�R�uoM-��{�Q��ufB�D]���S��ʝ��q����U!8��E��)Pl
�y(�_%`�;C^Q��)`��8��I�LYv��?z|~�.�������{�1��	���M�׷2I{��(	�i`GX�әz��5ۛ���_���L����\�2��NA����6�mY�>��x;�*0�z�IV� ���T�qa����d���p�4yG�w#��J=mς��{]>.��RK����k���߷=`5�XV��	 �Î����8��۶��X]��n� |\؟>���,c����/]/ pﴂ;_$Fө�T)jhMC?���-n`D���1���6�.�R����:\�r ��o�wp��_���ߢ�k���s��a�k��>���;��*�Ne�
��;�����hCk(B퓷�5w��x���Z>������X2�6�jӖ ��]��F)3G���V
s���!�#�5�}aa��s��\������?���+�;�l�����X޾|M�yV���ʊ��f�d���̿L_��U�~8g��7]�9`J��^�\�Z
a�ъU�?��^���5�*`�g��X�m��m�� m��P/��An��Ǉol���&ާN�{+>"4hr���#{��φs��{�~ƍ�_�ҿ��^�A06�'�D8:0&Ɥr���$���3�f�F�s�}�.�.ڎj�P�΢���w*
z��Vƞ�qnEt��1��F�׉V���gL�"�_;y�}�~m������X���hJ�V�h=����e��|!�wجm�P0k�46��*^Tѻ�K�ø����C���H���ƒe�Հl��:���|L�6:�l�${ _ٔ!E�J����U!�&��$�����v�N��J�{n>-
��x�ʃ錩���G�_ҼK���5��)�G�N-+/G�k�]?��e;���-��=��y��;׫
�d\�h��<w�U��@bf}sO~fw��9(�>.�,H[��|���]!7��Ф��|o�K�3i5_�Ϟ�F=aHu�6�_v ӵ�s�*�w�Nӄ���z'�o^����1��I(�G�bA����b���JӋ�u�J6>)Oh�g���<z.{�#��Jk��,�ۀ��,�}�ۺ��z���;���ly���w�#��(<P�ٕ�?w���ǟ�U������|��ն�����~�lyׂ���i+Z����0,�]s�4����P������ܨ��k?)t 7�8�~aH�� C����-+�ၿ'�0�YIW|�(�,��&�R����*Bk̏C�	z�&y���0p��j���ϟ��i �����5�mx�����Q6_���o�Nn�Yf�''�$1Źm��r�Z�e���i5^pΠ������.��>ȷ��0���BQAg{�2�(��d1�gLW	���1�)�d*=�~���nn^�F��	=�"B�Lm����2
}lQ}9�P)Y���� �ML{@:�T��������n���+��N�iإ�L�;L�Tz���/��:l5�'2YE��������"*�����J�$�s�����;3:��h�Z�j�F���#7�l[�/��/��7Y����8�ڏaM���h�uV%+�}���!Ʀ1o�;�2���R�S���Ү	d�K�&��5%�HČ9.̋���$�U�2��?���V	���>o��Xf�� ,�S�8���1ګ�\`�+�B���ӿ� ��~i�B�%��F��>�t G(`���a�X��� � ��%��L,���5�a+̒ȹ�E���ry�;S����KL�|�*�mъ�ױ$rS��Xa㥤�ţ5��?�y��3��]�R��缾g`g7�+.�'%���W�;Q���E�o������\5hm�j�8ԹS����NΪ`g
�_8�m��Zm��K�ݺo�ܶ%�A.7
�vfrzz"o߾&w����n֛�� u����?�o���6(
.[5HDrN�{����	_�F{khɼ�U�nt���6�K�¦�eՀ�쓸���C۞�z�{�|�kUZ�@�9~/���߿4�W��8�]�l�������v������ ���*���v�e-!�1���z�fLè��}��k-����[o4�\#��Y���V�:侩����i����ū���?��db�v Vy����Oٮ�� �aK�qu3����\\�3���J�+����&x���i H�гo�M |(���˷$�%��(}�� WW_��?�J_�%P��������{>S��BASFy�M�3h$���Y7ԃí��#{"��h��붐ˋ+��?'��B�ͷ���º�d�̉Kנ�B|���7DG��p8��I�r��� ���@�NA�� �ӧ�4���{�W�r?���qPJ���1������k�����Q�-QÍl��i����q?����t�dh0�N�M絈Dz^�wgbFtG�.� �ך���ѻ&�h�U`�7t��<=�^����S�b�c*
��Y�W���,5E|$ؤ��9�n���C�0��̔WO��͒�]���tz�#X��c��1Ļ c�a��C���~a	,H>�wx��})Q��4�6�v�5�+{��d��q%��-A�`���%͔��ī4��Jp��,q1�����x�f�����Jo �5'chm�F���2r�Q+V>���R-�9@)N��P�>�'�e_�:�d�ZA�{�d�?����h�]K̼h�=!J3Q�<+���$g�w�ǥ��a����|�Am��$_� �5^/
�.'M�c)`�a�@SJ��T*
�s�k�/=��(�F�F���8�L������I
!)+x�z=��vI�	��Z1$��An��y��ռC���<�@�*.����
1Z����
��]�pW��e�l�隔=V�3W^��I�q��ρ��J�}(^;�?��Y��g���M;���Ό��g��g�o5�W�>��T���%޳����_��g���=q^A��R��~yKS��%��@�K �T^�~M������B_)g���1�!H�F1~̨A6	�,��֚> *��)i#��c׼�`-�:��0@�Q���� .�h�1Og������0��A6_7	�!Q�V`%��M���!�9��;m	��KX��p)�X/�a{��l,��*l쳩h���I���ǖ�TX~����<9���S�Vg�6�5u��,Cq���k��ْ�b�H�z�Hy��$d��B� �Ms���p����W��|���;��������DR.�= �O܄Γ͠�6�ߡ1ǈ��z���ծ�T�&��y�>yAa@Z�j�R�VD�:��ް��@�2YeK�5h �|h�f0�5�Xr�7�C1�TՕ�����`�˦ǥ�xD������C~1S���'gLJi� ֦�(6A��T�x/͌�� `� w��o���1ܧ��(Zb_	)�{t�1q�U�W>��Z�:.\������hg��W�Y��7��$n0�M�3ǐ<J@} �>����ChA�ٰ�F�Ʊ���b �N���t��)x82в�gŢԜ?�@��8!�K	M�	��·%�76z��y)-]��UR��&ŷ�����	4�����U���PX���
Z�������wOl˥s&�ZyF��/��Q�P�!�Vs83x�}Q������dP��J��j�h�eP^ZS��G����IX�����3��ν��D���e�ڝ���;vy-�t�����d�_*����ش����N�B�=�9m(�vw���K����3+����h�� �*T�[����ڨ��s��/�����,#Oj�� �{�Y�z��';���
�G����읡�]y�^�d�m�Ba�k�TS،���V�}�>�p��"�z �b�.��u?I/:�wa�u����nx2���-�c�N�Tcw���R��H.0�(��`����L�w���CU��͎U��X5��%���b~�}a���9�Ll�f@-�#/0�����kwJO4Ș��*S}g}$�Ypn]�\Qijr{�������M_ `���bp*�W��ĺ-LH���X�iK�݀\�A�:ÄQ�����X ��o�ͭ����7x����d��#z!w�3M ,��e��3�{�N/�i}��\���p)!ȟC�s�h�|T�NӜIv���D��/� ��aI7�u��c�,�U+5+jj�Q�]�I~0�PR����y]��~�y3)EK�3Cog����[��Mo��s�3)��b[?<7�zt�}�$����T;�>��/Xs�(v]	��0�������"7�9̴���܋������/���[SR|`
��:�؇���41[ �5���%�)eë4�rl�\�8��'�<`M���3/5��EFեԞ"��&?���®O��U
��qe��uwsv�	�ˬ�|��4y�s��"�a�x,l�+x�]T�]Z�4�Ai����)*E��h{����s���	���Bt��A]�}?�,q�8�U�z�:��B~y>y�u����N�����%�m��~�h��Q5?���I�3� aX��I��G2�R����Q�����C1����H��G�C� ܳ�C����C�to��D;x��=C��'�hU,l������j�`K(L(:$񦣣��l���%�<�+�8��r�A1��qRQ��;�g��ÿj�6����!��|O�����{�����=m%g�y`7>CO��\�3?������B��{���Ʒ�A��W&��ë���y� 9�3�7�=�>��85'�ck8����$b��58�B�8@��K��=Mg�5�~/���^�e��A����1��X�k�L��4^�B_��.��� �ɯH��L�Z�� 𶡯�Z�b��f�+$$�V�6(����>���"�G <+�'C3 �6\��aZ���b͞|(@�Y��;]TJ<�h��o7@�Iw�,�	�3�0�A�9��|5�H��SF�4� yِ�&�("K2TOh\ޡ8h?=�n/�2m��O;�j���д��R�r�Fb�A���A�s����#���N1�y�f�g����_�F��?��Е^
�vg�C�1r�<u�69����uļ��G;��hq�1����U�95Eχʱmm\��zN����RI�]|Lvf�Zc��a�z�4֥�c><, ���`1O5��ze�&��0��-�*KY����e�
w���Hb����c�%5-�~kE�A�z'�AX&��7E�mIb�d���lx��:_�zt؎�4��%�m�q7U\Yߡ�N<ܐ�,����:%�s0�X������>�Il�����#w(��QL�*�!k���{�i~�\��Jn(�3 �Yě�������V;7a�OS�H��\�吟�:���{���9��=�	�sx������*����]^��1Ǥ�G��V��\*�H0?��EZ�����{����F�YϹ�O�|��L~z�C��~��|��I�9���C"���$��<��|�Tf�Ї����(��י���Eɽk�d���'ī��ɽa����=<�#���+x_�R �g�tk�{��/Uy�D���oϽ�UkՓ��_��H[�H���m��߻^_����Ӷ�Gx=���^J�sN���8�!w�7�9x)p)��63ܓo���{o_s1�!虅�;M�X�R7�\~f0hJ����h��� M��O��?�/�(���7oH���AV��|Y��"2�2��W7�S��NS<���6od�����Jgf�^2|�t	ج��$�{Ғ&(���D��zyzD���b���)\?�i���D��p�WJ��9�4<i�y��q
ɶΙ�����5i��a<e�Ga͇��ގȅ�x���Vr+��+cR������-�{ȡ�})A�LA��M�9M �����Ok����r��)mN�)��Z� ���I���u6Aס�~��ws�(Pܨ6���l�sP�1���CX�	�g_�E�F��g+hω����T�D��P�~�su�Y�I����ʾ//ߞmu�g��J���	uEF��?k4,�E�)P(D�t�G�ZC����"ND. g��x������I����TO��+y���b��������aG#k>�aKѻ'�c�
Fz�`i_�&���/���*����?��g'��ʢ��$(�����%_��Z�����C�UB^�
���V�)fW���-�e(#f���Ɗ�7[q�YecՖv'�V݄:��
�A�����x��ޮ�?�x�6`���B�+�:T
$�4���y��e�z�<����\�~PTU`��V�<&a��2NL�G��yg��J���?8f����[&�S!L��h�PIsv�9�����;z�non�˧�����0$/�?�Q1�k_��R�N��]�|8X(VK�]����\�;���
D���
��j�;1^�1�r �}p5�f���F�����20ʀ,�> ���^1L��]�O [�+����I��סr��u��q��A����P��ߴ�g9Vm���<��d����|{�m�>nC�z�{�������j%	��5�ǋt���
��
���<./T6NvX��2d�����e!�W�1[�|��&�[��ƴ��� �����y���&$���L�l_m�� Ds�� ���G�t��]O:����B�S��WO/6 �~2��NO��o��˗�����T�&Ո0�z���l�<�B=K�Kc��(b:!zS��jj����~x����r���s���x/��ᙧCAs�@ҽA�y�ܴ��kָ�<]�d��*���î��qc�x��Ȓ�S�M��N�|u5��=/ W3��q��l��#�I�g?*|4ߚ�c� �o�<��(V�r�=��Pz�@����Ds����쪌�h���He{�鐣�tS"tǪ@ � �W:@q���Q��'�n`Q"���"��F5�����qҿ»R��:�`�O^v�>OA\��p�3V��2i��Z�y��:�7�`U�ނy=��[���s�F��%�= ��K������@�bu�s�TgP�*��wS��z&o��\����y���۶6k��)�]A�Z��D�aT�Hu��F�a���G�Tݱ1"#;#X��}ُm����:*��Zek]��-�az��?�,E�����=�KK��J��
�Q�xx�/��a�`�롅��w���i��I@����K ������u�����yek2X�$��Un�⺿���~\��{̟ͭ�"|�YRn53�� Ƒ��C׈�s� �P�)��m
H)`�0��b���ptF� ��=Ͻ�A�s��[
�t�nW�U�ec#�@���.��k���>��P�T9�޽fue�s���|��l�No�$�n�={ل�tT�*i�D�h@ݻ]���F�P�׫�k�~}��$�;���N��7̉��]T��BQ����?HgpGs]`�[zJ���UBnV�@��|����1��&􌾰��+
O^'����O�_����'��F��c'��5��#:S����'��G��1�V�����T��E�'N_��C�{�SX�������y���*��~)��'�pj�yB0����q}d�F#6��[�I2
䗟�_}��e�W�W	��1�댊U 0����-�ʳ�g�%����L�N�4��؍ �����A�a��m&^%�=�����c�<T�<f�]�^��Z�JVX��Vr��p�l��& l2ɺ�%�~+N��d�v��H�YEd��t(�,�\1�hƭ�%Ön*�r��;���ƀ��F���H����._��:u�6� ?e�j�����	�گ躝E�M���`�y��r�j�Et�n���uUf�,A�)�z�8�N
���=</롻&���.ͫL�y�g��8l-f�j뜑��
��M�ZWx�����zHe�am�����Ѕ2m���Un�!V��Ayl�ޓU�9-�+y*�S%���h�+�!o1�ec=��s[�geN�-��z�⛰L����KJ6Y�(Ç@R��ŷK���?X��$�C�n$O��+Bp�O�qj��zVQ�د�<�۱�|q��2W�z�`?)��=�,����:?���9%����|�(w�7�+
���[�,�u���6���<�q(a�1)��^ZS�������x�F�k,\7�V��aeߏM�|�_�ާc\#O�*Ͻ�1�}�p�����sT����G�Gr|n���]�E�q�=Y��!^B���	�5hۦ���On��:Uz�(R�*̘+�bɏ�hM�ap:a<��2��;���A9Nwfrv�����F���MD��'�vSe�G����&�\�6����J���K�u*3�j��t�`� �iN�R����:=9��t��f�v���g	��K��^&�ܦs�����1��+x}��!��,4��֜>��+�L��	�+�����!�P`��)� @�� ��ى�{�Z~��'>�{k�φ��jB�0�ގ����"��[w�;=="�C-���Մ)G� ��w���=R4�3�M��k=��j�6��EA\>g���E'�����9|��=gt�C�u�U6��xD#,�b/I��`������-�4WW񗍣�2=+崺9�e��;pj}^�۞��w�=�B;����g�.bѵ�+*GZ��-��;���$%LI�v�i6��%�t	��X%����j�5���`8��Sf��S$�Y/vٌ>�^K	A`I%`C�&y9J�]'%	��B���]_-�H�4G���%�����V:����{d�Uy6����)��]����$���}o����o(�W��z M�C`�3�j�Wo
ïA?]�3�ಷg!�{V�ڼ������skT�U;a��r�k^���P6�&Y�����zuCA�M��kG 4�����!_I��!��0�Y�ɧO L��}��6m�*􆡙�٦5'���D�rE�2�Ͽ|Nc�g�@$��J낭ړ΁6� �b��PXo�W��3(EG�9�%	9�e����0ƴ��z�)�K�O]������� ����_Te�6���[{��Y�o�V��\�7�M\����g��g�~ey���j�����3������?���{���Ɠn4����R,ˁ�� W��x�lz���� 3@�	�W�?<ʗ�o�:VܱW*�x4�#�NшM��{�1�U�y`�����8�����"���i �r$��%�����ҹ�����-��������z�B>�as�9��0�h'=���IxO���f�:��Aj����^�=>��3{	P�swyy���P&z �{�� �"�#��c���c���v��t6��Lk��h�:!8Qq���k�%a�Yĳ^iL��������L�����EEZ[�/�xcY����)s��� m�W��xd+��)��|�����M��H J2�G�o�f.�����Z܄�$��]�4���Ґ��4�0���{�
��aE=S�ӝ�oZ�?�D�d,b���.�W�1�
5&|F���VӋ]ܭ/J0ja�][����\�g��@�?��g	�К��Kt+Jj���ա��7fT�`�yB5�t�V��2!u5e>Ɇ��o�
�W`/�o[������p��s ֭>ŋ�u%傒3�5`�\�Ds�x��<QŃ�sB9(������G�(��/�/��=g�֍�� �C��*�OZ��oG�­��V 1#�t)rTo��z�d����@�d�C�\�@�h�a	N�/�	�G��T!1�__X/<Y�wXZQ�)l١�#0��
���*��yXЂG������2L0������pf��}M2��G'�KU~mse�Ɓ�y]��L�眀W��r�/�x��P�e_�z�����ʶ�[߇����)>����j��j�mV���QJ�u����=���c��m�)}��Y��S����<��n7/�<��@���V�33���v���G�l�+���{ϗ%Γ�;��M#�� �&�L����A84�EżlQJ���A��z�W,�b�z0���	�P����鱼8;�<z�>�j�dNӌc���%��#��w��W��';rpqE ʅ���H=@o�U2�6��'H�͎����ׯ^&��+�&��(��1Ɋ oT�L����{3�g�O��(�s��[���t�G-&�H�7'@�JJ�N`Ŷ��lH��HOf^t�>���t���]7�b��c�{wB�D�֪�j���R�S�1�HI0ߊ�Tp?E/@�b�
&��~QUn��F\���	�Ux��}��<m�f��i��qNU8#�cTG�B�NK���Q��( ��`��������W��l�刘�ite`�zY6�ݕj�
�{�A��2��ǭ�T=`�GOŕ���j	����$*oG��~H#Ik��`��֛!lo�Pͥo�0��8���;����Xw�GkHJ�m�:'��pA���/^+��3��������3�)�+�y��T��>��6'<��66D�����r[�FBB(��s��Wo@�f���fqy�w�(J߁�Z~��?��Ã�$�v����aǎ%�=�#ջw�$6�I��	�������@�m:>ܫ��yu������+��esJ�;�0A��&�PY��ƪR[+�p��5��=,�"��+k�Yz�\�ѹ��h�]���8u�5ĸ���*|��魚UJ��6&�%��>�nhT�? ���=��b�4��￶��s��9��6@��]��L��:�2N���d���׭�S}���9_���ޚ?���=�S/����A�J[��6D��kee7RyaaK�g{o���z���nn��I��]k�Z�\n���F�cN憴E��c���h�<:��^<Ȱ~L�v�	�Xϰ��t�I��;�A������M���Aq�"�z�L����O�J�Wrys�Έ�{~���1}�Wس
&:\ڼ�c��i�;iL	t��� ��9�D$�',�N �W	��t�g����w���Z������r���ڗP�5X���R�9�A��/i@�#2����/$c��� `>#P���ce����k�∛d��ʢGað!|�#��"I6K/D���V�5��c�XQ�S�x#��sV}����D��T���>@��^9>�ʻ+&�bgՑ����
!Z4�}����ňt<����X�W?W�o49���Ob5Ѳ�ݸ	ռz�"��c���G+/�
��"�eg�,V�_a��������<G���ccop���E1�׈�{4��R�P�2䍐'*���u��]�I�����D��
�
+�'Ⱥ@��
�*�����ms��b��<=�#$�.T���ś�	܅��(k�X�'�7�T��)Wm�}��_���-w�V��K��[��r� D�\�V�ʆ�����(�~q�Bک��<�t}���#��� &���+�^L�jgT6b��"�AY��Z��Z�?͏aȔ%G�n������?==d�����<�.���):�(��A�XA���{X��=�c�4TFE�{1�O'*����V�b�������o�=�g�-Og=�����Y5����Ws��=Sa����{~�O�k5Z)k��:۞��ð�_��={��>	e�3^M�c�d�����k���}6�Fb7*��0��2\2���U���C���;��*9hhO������$�^3�,< ]Spx�����`�����]�I��KL�P��x�q.� X&`r����4}�����к��K !��Hm ��c��Q�����8P����X;8%WU$A'��V��(�a>����;l��7L��	��c0c`��:Cf@����������r>n]e�Eh�-}������W���gY�57��3$^�_�:6C�	f����XI�b�,]�����񼟍��*�>���5C�AJ�?�Xk�y]���PAY�{ΕH)�h����3�D�j챜��C���΅`�����V�#U.�F`yun��J�Ƭ)� |��BQ=��/�T+�v+�G��K�s�AB�I3@"�Pz��ɿ+(� <]���6~g��������ߞ*f`�v�R�^ �83$��l#�kK[^��Pࡖ���jh.VYe�>�{�rY�)S�ָ����$n�Ȣ�Л<�M��R����<A9�D"����Uk��t���j�FJ��c�����kY?�������)����cg�؝sf���{��#c�&�wN�jՠ��N�u���c�w�}�4�=	��kϩK���Ga�a����������:� 	pQ�}=�,��;�"����xVj�5�2�bj�V�WE��gáV��CTwk(gf��Vv�wW4�18+`m˸x��۟+�������{L~���=����dR⦱���̼�k<1������j��ݓ�׳���ss��w����ak]��_�r��r�1�Xȱ��޾{'/_����������/_���5A�.R���6�H��g45VT��L���(�zǆ�$� x�� �b� ߼<�#�z�3��c�����oO�����<���{���
��Ym�����#��q�c�O��ۧ=�2�(��{���=n�jz={��*$-�"�$غ��������_������Ԩx��2�k�1^��&�膊q�Ө#L�wL��As[;�c���h������������y��k>X��&�)�4gXcJ�qE�� �<l�ЭD��jE�rn��tt^tp˓�LS;B���^���rGD�����B�n�U�Lñ�H�����
@UN�9����]޸���+V���M1SLd��-��r���p�g�]?����V�%�>��Cƣ���u߲z���H�3g�w��`�TV���T�����R�ߐ����*h�h��_�DO1�-��U�]�t�4�:ǋ��p�W�Ur������x��S �%�^�V�&�h��x������T�j�������Ge���x�B�p�8?<,{G�Ҡ!
ψ��(��m^����(*Q�:�����ᒮa���f�����JR�¦�i�h����'NR�U������R��#`�|:���vQ�>��P��֏��N�_�!���_d6kXR}}���v����	pY,����k}�����(�J�wC���@^ߌ�G���G���{��b�5y��������?{�8��Ûρ�2�m�5���<I��5��$3u����=��r���&����4d/��j��3�J-/�wy<n�͗R��]Q
��U&K]�1꟦���`��������\>~�&�H,��PZ7�Г��@4秵
�����YgyI�n^0�x1 j�]�l'���~y���{�!7La���y���(�͚����Wc_`��z)W�7$`E�áoyn����{��L��!�����) ;�PG�!Z�F6}�X�a��7�����N��n���]=�4渇{�\��QӾ ��YE�2t@���]?o�W��a�����\�_���hN�hU������m��A�y��>����.�[=D�y��r���3�P�SD����2:^+��Z��`�ѰPǢ�]���ݱ#����{}�L�s��|�2�Q=��i
�pP�aΕ�����Qu~:*v�xn,�GDs��d��L�}b�L�����.��e�n���I}�|�*ԥ��J�r�0xr�N��h��ZI2���ƽ�H��eP�¦?�ӭ�*Q�HY�r�\��+%�E�RQ�MoOd����o$�����B|��)�M��XU��[e\����_c��������w�����큒���&�2�P<sYq�u~���hΔ�+���u�A�ﻻ{	���/�kڟ�B��m��Wh��@KUG����*�>��^?��[E�Y7KND[N�:=D����ih\`������%�`�2�R�E���$��p�7>'���=�ź��Fg��	�d:�g��Y����?U/����������j���թ�Զ�����J_��Q�T�Y���]m��4�6�/@���<]��d!�c�2N��X���#��U7f��8
f<{�2o�H�+5]�(݌/��&�E��{g�K970T��V=+���^���t�J����"#���i�n���N�3މD+��
�N�3$xq���iG鼾}�V��� ��<Z.�G#l�%��r�l�wȟ��M�������d�\�r���d�nG�&�=n���v<wx߿��^~~�C�y�,��a�A�,��� (!�i�+po�4um�B!a��}E��%�ꃹ��O2�ŉ�{�Z~�����ö�2���3�ZQٍ�Fv'��|�����˗km�4h���|0Ӂl�<_f��?���*����q�6������Ұe_4�g������5�b
����{�1:X�#;���~�G�O۷�e�t1c
?P��k����S���*#x"n��t�	��;͜��B���̨��C*���v8ɇ����ؘ�q��\�,���\H�)a
��/��I��2��B�N~�=������
<�P3�&�h.��f6��tmeܥ��d`)���&
e!�ߧ�n��t`��!�^٦5ǂ�L�MR��-@MQ�Vz.�w:p��#+!�_���m���^�ɹ��Y���]����fu &R7H>�J�<U-վp��D�7�w�Ha;��$F�X�����m$�(1.��������%���w?���	C��_�2���Ǐ.˳���N�'��e��ʜ����)C�h7f���]�F��銴<����~��g-*R�m0�է-�$��4�R�>�
�*�*��WJ6L�7V��W�sυ���c�\�ƕ�ޙ�-�H܋X���Aa����KN�S������2�G�תa����{������󺗮�;E>z���4<2��J��Y�I�x�@ �w�0[���=�t�A�8F���P�NmT�Y�V��!,t+R�����)Ð�=E%w��%;�e��A���J.�� �����۟���s�����D6ٰt.����ՎH�?;9N��*^6��:)�j��C0Ȁ$�5CoJ���>�r����>r���h����O����y�����j��t$����p��)N���zD�(����6V��av(@Jc�a�����k�|�R���KmA2�5;�p���;(Q7��{�P�ch؁���,RЪ�З�/���;5��O��+�|��=�>��X�Y�E����x<�wx*A��d�jO2���T1�Uo��s��u� �mX,z	��[16���M����UT��T��Э�J�8
�
��`@��P�[9`��m����=^�=u����*��-�B7��`�	���筏<�}{�7��.��uS�I)�K+Fc.3��H4X�ٸked���!R�J�r�zE{Br8}��o)D�>�T�.�����������աj�q�k��m� �5j�
�v�B�s��[�^�% ��NO�����~�iAt��ZM`vpp"�ۿț��e>`����D揲����ĭV`1��&�v&�ɢ~����ߙE3PP���h	v�$(������ ���ʻF��%���3J�����M���<!�X�Q�I��X�����>S�W�W�9�4��p;�؈�����`�G��U��!�g��+���(��d�� !�䠆�˛���Z Z=GꙓѸ5�Cå�~���k��I�����C�.�
in��!��`v6-�`z)��iL�{%o�jzCc�&X	����6�BDr�z�!����+�͸ǹh:P�\��k�^����=�����T�/|�]��n�sT�8^�h����/>|����V޳Q�>�mr=���ET��P�������w�p�@Y������҉m~��F��M���gޒ�?�C���F��<v�B�ުJ�D^̑ D�)7�\('C��F����� �\�L��'@t�@@���.����)�ސ�s�yrys'_..�a�.���SBJ�ʌ~��eN�`�s�d�ie#��S��P�Q���D�j;��-���~�ߺ�:K)^���:�>��'�����-�h@Q���8li�uV�Z%z��,1�H�|��*C,��@�d,�����2N�b�>1O���}�$v�V��6cȳ��t]@pU@�Ye�k�%
M�)�5RM�tF~�(�1����=,^D7�P�ﭢV�@Z���4��<^œ/��#%�ڽݚ�5n���7@���hI�y������o���Åt���r�Q�p�BX�k�9}�����Mcd�Vͤi�VѴ�)�ku���54F�i˦��V��Ą�P������d��xi��3K lg� }�zX���Ra����r7���uXӢĲw]IB��Nw/V����P�%�{k��Л�C�&�*��z�r�n��k��&��J���"�c�5)�N2 p� �=i�T���\�2��jkj�1���*Py��{�艖��kxh.0?P��+Ʀ<����q�x8We`!>�~����Y�{�|6�M.=���7Me�pl#n����EG4D�A$C���Y��
&��f���?�e�ͦ,���'Ŭ�,?_As�l�Pd��5��z�+��Bv�[�ٍ�șg�c�-����I�
�����%2��=��X�߰p��No}e	�M�}i����F��Q��W���`�V�$o����k埕z.1]F��ͻ�s�<�0�qM�<kIϡ�C�yC)�����Ez�N����婼89���=~�
<�$�E�㊼j���ie�|`!�`�P��Zb���!�51��9?�k�x@�m�<��m�\~��QT�\�{���K�6G��|)�I�ZP�I������B���m�a!&C�~t���E�,���8�:*���Ib쏊����^�2�XXKQYi��0}[Vu��~�AX�W��'L�U%��a��`��@8�ٍ�j�4�ᐘm�E�����r,b��ƺ[��l��ak�M?a{&�s���G-�`I�z�4'I��Ѽ�������py�� i�Ϗ�ϓ[����UgR=\�!z��Y��b�MX~�Fߜw� FGh�c�Ѳr��+�S�����nN�@O�r�`%�����Z�MY�I�y�m��s ��!�2q��Gr��BVm�������s������+���B�O�p����V�sbv	�@<�LĢ^ԜI-�I�k�P�H�X�$D�Ǹ�zM�0�4f5+0�y6@ ���!5�F�§��VV�5���yؔ�� <hK#���J:09��j!s�"o�=��~�c�{���r!�r���P��*�>�5C�Z�Xr��̽�����=]��V^��\0q�����uV�[~d�m"%Ͱ#���Y�4&ơT�>�>iv1�#�W����'G��)]�)�Lc���h��y�^%��I[�3݀�KL�t�錡��b��M.�WԒo�S��c�i`z�)�(Z��M ����fU���/��\/�;�m�U����6�;Y���Yb���l��,j��6ކ.C^�nz�u�6^��Z>�p0��8�&���s�]��54W�h���_R2��0�9`��gTo��G�^L%�M$d٨��Ak�y꥟�[���A�ʄ��d�8��D�\�{#�m����pW���?�(~ 
&]޳X���T��;��g���+٬�.E�M����P��1�fWpb������T@I.�olq�V��s�}�c� �(�1�)���^7>��Md�v�${kC�5n�(�}=�>s��|2���Ɣ{Y�u/�0s��Xܡ�Ij�(�a�vY\�*���5�3�
I��^�&�2�]�%',�h�&�^�Ȳ����6�P�*1�QU��{��7�VȐ�}N��y@֣�8p�YZ��,1�y���5Z���E�}i�)#�D]��"��\���[�T��r�'u�$ؓ�Ԟ�"���0��*C� �*q3�&.�;�<�&[��#��� ذ�E�i�Lɧ���j�|�j�蘄�Kj�ɣ�a陯�>i��@`а��������M�$��$���z�ꕼy�ZNO�)����_�@0�I���>���������,T�����$<[�=(~�$`���0ѥm��+�����r��t�6����rn�	q�N,��A����;%�$)��k�dp���ϗb�ګ&�y�$��`	�qL$f.���@��t@�}m�;1q��y�치H>d��6�V�����U�7��ek���8����.}p�GЖLTT[����Q$�P��+~s�s�RGA_���Y���:���M4�F�֔�1� �����a�|�t��?>2%`�8Wn����\�f�ëI[�b� ��(S������wv��y^e��!�"�
�VFN�4c̃˶�o��}3lH���~��U�QN��LєGH����{r_!�t7k��z�=����ߍ������8_��T�(�v���8?=ؓ�g���Չ�{q�-�xe�y��m���7C^+��^s_��&Q�L��[Wc�5�wf�������h*�`!L�חq���Ɉ�)N���ۼ=�|w���i)���+`�J&�-G��'�8��Ve6��y,�h��9d0��g��B�{0�\U�U�g������b]�!͊'OY0>� %?�]���8�u�y��\�P�q�r-0�yf�ߕ���KE�^��!G-���sV8��	�b����pBM���r�ɮ~^�+��N�ɏ���JNMFV˼�+����ry��qd���,q֒Gs�RTX���%{ot&�h �ah���!�F���1PJA��i4���I��`P�3��.�7�F�X���g��L���^n��X�aL������ƿڐw�������S��������ݏ?Ȼwo����{j���k��Ġ�@t� O�X%"����i�9^'��KT�Ů�o�Sqn�s�rU�*i^�-�@��j3�!�cߣ�%9���B*��܄�J�8�B�'@��TLvF�K#"
>��Ri�s������\���:G5|JN�QD�c�+[�@J���)Ʉ�XfQ���Aif8.+�)���5��
ـPS2�~
&��[�j��9(�aT0��e��c0�9<����k9-@>��\G�O�Ǥ���Uo�H�fd4.w�5n S����;j쨛�D99��kϊV��a0� �\^I��nV�E��{�M�jH�1qqp�^�MzrL^�L������oߴ�u:��ֻ|��g��#��Oq����h*�c�w�{K���
���&�c}����1�:���@�ٮ���nJa�
�V��|����kAe =+Ea�V��T��m{������5e��	��p��ڟ�W�# :�\_]���u���$��,���5��d�1��х`�@޽~)�߽�ÝV�� ��i�Y��	+�y��Z���i��?�N�"�eԾ���g�J*�������[�j�3x7���h<�pL�=J��y7�\lk�F�:V�}�%�Ԍ�+s�6���y`�k�K<4��5}�F�-TƓ}u��9���Q��������lѹ�/�XLzL:G)��6T��Y��'��ddn��Q�k�?��*K�d�����P�nd�fL2���g�4���;4/�B�6��Ѳi�&�ޣK�9�.�'�V��9=%V��M����"]�a�M���6�?��Kx"F���o���	��Ğ_���kĲ���Y�G��lm%��4���jXw��h,)���Kځe�p-O[mrMbDsRxՕz�Txn ���!y�d*'gQ~�?���!��eB_//� ��G���2�k������ʦe���T^�~%?��.})���g/�Xa�Nc���'�3Gsճ��~�W�8��z��vX�$�;X��p�;�vt����WO��연�wzS�*sM��0X~�����[]9�G\o��}�A�nR�C'*�},O"v�ۛI9_�Ϋ�g���q�HYH)�9�nU�t6�D��4������b);����Z) �K���dP��f��p�q���=����YNg��i]6�--�<����q��旄M� (��S�&@�V+��x��.A|P�p(D�e��x�����V4���$��D���:�����a���F�E�) QVɈ]<���{x��ŷo�� �Ջ���#s�H[F���f������u2ή�6�f���}�!U�Z=S��2s���+A�@&���_>'�5�p�<�Hys}u��w!˃��'f���s��%��Ț�-��
 ,�̜?h�cn��zm;�����U�{/O�>hQ!��|�'�1����L[yyz̾������B�T��zű"��*�Nʘ!(����2����\��P�8�� T`'�{�d`�URݼW��)>&)�V}�P%A��-]�`F�;/�h&��[H��0���qvpe�i�;1����4��y���<oœ�g9o�0�P��ṔDN#�����1��.K�ʩ�]��=|�����0]p�)SX�P&(j᩸���*D���ZBnK��H����+�@	����jU�M;a�COK~l��������}�=�\��������QF������T?T8�ѵih����j��k38�Z�t�{�zK�A����5-n�̬e�		���Ps24�ؙ���)�b5�b���t�n<KBc�`O����9w�I�_^ȧ/��ׇ�r�����k%2�f�)|N��o��M������~L����D�%*� �}�I�]]��y�{�?a�)+�����I���dQv���v��
ógX�i$��F�g!�\�#������"�*Bg��J�jv�ɢ	�ҵ������$W��赵�x[�'��AK��Y��Z�?3�Z�9fm�g(4��ܛ�S=�����d(_��>s�S�恅�bi�m�_�F��"�3�w4aȾ�R�,x�+��HV��{�TB��Q�L��MmW�8+o��K�{˳�yh�yJ��2��T�K<��Ӕ��E��'���x�K�<��s�A)��8����̀א`�T��;Sz$<G�x�u���9P Ž�3m!�v��Ū�'*����]>\�EV�S�C���OS �4nn[.�2�߱@���EN�ښlhH�
���8�����R�6�1h�����~���h�9>��G�s���S&���G��kK��dMm�	 -pƓ�����!175��3^;�P'�)� ��������MQp �EHm^T�>@�]\&��*�9����͞={�� ������[y����G��l�|�k��W�(S�&�(G�Qlf�m�@� /+��^`�w�@�+��3�����C�y��R�z��H���8 �Ғ�=���zJAot&%�l�S��ט�L�p�z�U^kx�ɞq^���Ļs�j��E߁^ ���9�0�:hJylK$F�5�6m�0'�rSjt+�Ale e�w%���=��r/ƌ�j@�=r�G��y臲��$���K.�l���������汁���͗��{�Y���T��j�;A٬�IА��0��3C�t_�'�[D��8�-�=H����6H9ɻX0ި������<�,U��n�X3�M�ɉ�jBn�a�����9x�����ق �Y3E*D�n����%�	��=��q4�]���͗r}7���G�?L�xo�����=
1�o�Z�����T���G���L���SZ���S����&������k
�������������鳜���˅��T>�j�i�`�<�t�P��������B0_�%�GS��w��[7]Z?��j$%
�&4-���s��Vc$HI�7a(!4���ڃ��ޔ�m�� U��l��yj�n(�<]A?7�UiB�=Xjd��ˮA@���ks����h�TLL��
]F�Ћ��L��90�3O��Y�X�D�W߬�7v�P�'�½	N�m��)b��7��kēxk��z�ۋ;T�ڬ.A��Cm���A�5N%���/&ֶK�h"�Z��˫;u��
Q�je�s��5�J�k�	�@���OF���9�VD��	xO右��0�M`g��vyu�<P�#=s�TV7�?�ۤk�ޯ-�Jv
����F.w�I�/8�f�S��\� �A. ��^���%ǽb�S&"J-0(�A��w�;K�$��q�p⥀���nG��h2��@=��ZiMI.���i,����n�+�
��ӓy��$��Y����5��h����.ɸ�܌Ð�Oh+'J��������k4N��t{l��h��w��N��R8����X�zky,�Az% o4�X�W͜'���,E���H�!���
I��Ï^q���F�p��$�EԱs����eԐ$��X",�"B\��Zk%A������ ���4��^)(��c��1�ͩ+~�xCY����Zt�/�;��e����a�His$�D��EN��W�xHr��<M��}+w{����� ��ĕ,�|�ך+=(kqwC~|\�� ����\B��ki^�W���ş����6s�m��<�C�t��2�:	_�2Q%ɜ�^[K0G����Wj�l* �^"�a#��3y����`����X�Zq���|�6�ͽL���{��s�ӻW���5�/ �ݗ/����?�:G�p�K9u �w���}$ǧ'܏d/FNG�ߒ@��O�;���"��	�E�t5{���h9��֖��k)؝(�O ��<"����I�B|���}{U���b�����coC2tg�`ʓ��=@�R��8���q_�n���5��[<�~u�$6��| R�tY�{h�T��!�܆��5��q�!̴)��/��^�H�N�=1	1	 ��dF����ߌ�`�[��x���* �3�}����z��"fc��)��U����\��G�9@���
@V�C~���VO5�`�qc=��,/XOG^�l���|l��^�N�s��f��� �;��5���on������2&ϲ��;�B����TL��Wӓ����R`]�)�o B�(��j[4�+�:PPdzS= ����k��kcF��/�
WΒ+@[����� �{�'虰�����x�=�	!��;�za_���W��)���+�=����I�q��{��]z��{��L���u�͔|:��Z�OR�0�<Q�_V�n(���cQ�M]ogОЭ�C��t�k�i�"�Twv�r|r(GWI>>�˰\���W�
�h@��1��ֆ�愷AF�ϟQ����M�q�5!G��ў2���G=��Ωv6D��R^n�6Ve_�ju���� ֍���a	�\��Z&L�� �XM@���Z��
%�n��cR���߫y��G	�*�:ugz?&?fZJ��?����@��ٚ%�2�'K�/	�i
���q���G�5;hS�ߵ:J-i��ѭN�⋫ ��t���$I���$X���U�{v��������;�w�ⰻ3�ӤXr���TDUͣjqٓ�UY�N�MEEEE�߼<�.;VP�p��M�V���Z�D��M�;jd�� l�ʽ�r�Z�mW�E�v���ʑII�o�<�:�,�2Ec��Ec�dXh-��_��}SB��Kfo_9.��ɰ_��V�O���9L��e���7hk�-2���m+^K ���{�t~+w�O
�:��Y*�KN��M\�Y2�Jt��e7���"���7c?<�-�����O<�G�Pa2�ǧs�����p݋�{��p�gd̻�k�g["0�A|��V��y,t�^�)�\�5I��Y��]c�R�6���f�a��������ܡ�:�k�d:���Bȋ2�#��V��й��ݙ�;�ks#�s��y�͚�����n+ �^
s� ��i��63m�ob8o��ã�!���+`?:�E/S98������<:B �l	�;cL�Q����{65}���	x�����G2�������˰�O?����!�@1#L0$k�|�u��Y�������}E���inڶfW��da�w�5yt.�1��9Fʹ2���X���x��~Wz.k|8��8�Y����c�8�R+��nK\�h��!�� L�YJr�]JmCm�{!�.ɲ'���%���pz�Y:��ϣw�R��x��t4b�] yQ����9�U�鯶�7�b�B�2���h��mO�R-�V�f�?^��R�F ���;&a;A�-?MJ�Dv��Rz��Ľ���@a�;����-`�{��y��[:՝�>ޘ� K�[�/MՃ�z/�6ƁgZ�ß���#(�/�<b���AU�B3�4�N(L��H�$+��I�e7�צ��	ɳ<��1� ��y!q�M�^��l�A�|�X`6-����gdVb�K^��(�ɂ�N�@�*��
�uB��ӎ&�|�+���I������P9;qBK�<��l��dM�lD���|�	=���֐�찋��4�W*���n��U.�k��k�����{eg���'��(����'g��ڬ ����
�Qov��x��	���Sl���C�<5>�  ��IDAT��̓�5�Mr<����������87����՚/5����u&�//2�j��J����U�j�7��z�k�v��տ�Ŭ.�͸i�ō�5�� @�Qr�T�U�S�X�n�dG*��nͮA�[����<oit���Leo��&�tb|�
z>}��ϗ��P�M�Vo6��{�w�B�!�vL�f�� 5������&LPMkƌK���4�Xb��Hr˵f����Q��|!.��) H�;��E���VVڰ�yc�D@�ǎ�����H�������`_Ξ��tˀ�kg�i;%�J��M��t�]ҟ���5D�����iY��f3L8���������r}s-��M��ښ����ܑIH�7��P�������8�����W�7d?��X�X.��_{;5��>
���&Ԓ�)���K��noo�/�E.ί�E
�4%6;d�ɞ�9�ƂC�����8��󹜟��Bz�/ ���K]'(;���[7�Dy�c>�t��O@з`#^��<��&���G��ּ��������;���?�!����uy/O�,5�7ȝދպ+�Xf /_�c�{����A� u�`��R�@�R�t�n}.�=��7L3����X޾}�ǱW�i�\_^���h�����P2 *u��� f����������<N���]�	��ĲE �;�����0�k���G��7�/S�Gx>[�i���`|Xx�U\��S����|$�����z/���v@�����b�W��X,Z$�O����_�c�W$�`��b�$m��(<��(R���!M��-a����rx0��lޑ�X�A
��W˺��k�fو0�+ �~H�yr�k��	��	��^�����H��1倌+n��<��(/z�aRF��A�L�c�Іb!go�d�ݴ�G�X��-wd��V�ܮtM�rv���$�S�jH�no���lW�׭lN0��'�Du'�R�d쬹V��5�%�d'nh�J�����-O���+ӝ����_�]��q�����'��0���f�	�<��C��AJ7����U�	|�%���T�q��y!��\���.6����f;�{�
�z�/D��KC)��	������FL��e��S���H'DR�-�ҫ����&�`M@w+]�+8��0Q��	j�P�C1s�� ��eS�:$����;DC�&�F3R�h���l�Κ��6�G2]��x�a(��vK�7T;�~6�5H~�x����b{i��,� \����eC�^��ʦ���_�=��y�(���S��kj���`����v�`�Z�f���(t+�C��jmX���K�`Q� �

�k�Lx�b��{_��o��aI�*_�~0�v�6=�D	+���Xe �j&
����Y�����߾{K�����脌J]oe[h�Sp���ݜW��rO��`���K�&�g
�޼z#�޾�I�z|LL�r)}�~k�F�Y�Km�'��?��ى|��@���eɲ���ug�g̼��+O���[j� �&���Vuyy#w���:3���H3�����υ��>S���)�kh�a�I09 o}�{��s1��=��F� �l�[+��5�<(W� HR+��&0�"Vtp.ϟ��o��V�4��\�絞õ�����`��ѻ�#�qK��f�u@�z��^�~G��%�cclg��2%+�Nt#o�* {����X
�[��4�k�]�gz������LHZ�q�.����m��9*����~�^����850h0ۺ�LW�w�e�%��"!� �je���a��lt~�>	?���^|�O�=��5<S]�e�-�L'�1��յ�q�,W����bE1 �*�A@��B^������K�V.M�U�e+����^tw��cA)�$�Cʴ}����ұ��l�'� �xa��%�Y�T�d�Nk������X�fsԳa ��X$L吭Y��`״n77s�~��7�gq��*�UW���8c�,��;�*�]���SB���}=��s���S�� �1M�~7llʘ<B/ŎR}2 �L�y�|O^�|.�������>$��������,�ƸUב�a�+;��\Ia�Tr��rQ��� ���D�VDɪP��8۠�z?�4a[鳥�j�sk���ʿ�I�o��<.�<>�ƍ �;�	���Q�-A7:�:��=ndO��F��mHQa��\��.�-�P\�rr* ����Pm�SK�2���8`V�Z�|`j��j��y�O){&'���0 �S��`׵�k����B���k��e�6{�2� �V1��D3��l�� Jf�#s<\����KnΗƮ/JC��:���k���ڭX���ڃӗ�6�9��&:��پ
�e�C�b�^_=��\Ϲ��>)�z�{�>) zx�u�����lRVYc�v;ȡ�~��Ka�b3xxT�r� �F���7߼����Ba����,�}�����p}�@I�#غ��frۭ��x�A#��5��pCm���[���r�MI�ں��w�䧟��/�+�{$�&��ټ@�>!�8p ���]���}�^>|:��,���%�i��=���C{7���l��-�g06`��ϦmfdZ����X�ر>�r1�����U01]m���DA��yrz*�}��<h��Y1���b~��ݱ$KMOgY5x[1������1Kn(�b�����P���|�F�,Wg/����OIf�H��ƺ8a�r,�*|���b�����9h�Pd0A�ł�c�T�j&� �`,=�t,F�uy&��q���+c�����*��7J�&1Q�!+xx|$/_��cج\_��[ǁ��c0���^���3y�浂�c�ꚸS<��k��|��=�E���6�=��ٞ>�{�o�>�KF�j��=���~9�Q�d'K��H��\���1��?���%K�t�I��������}�z���A�{�}�4����:����|��	��xZmɩic|^���ַc̀��;o��}��w��v?�C���k��O�Gݰ��d��&�7`̍B�ež�8I�;{{s2�?���Ĥ =�����h����{X�xN�Nr:�Y���^�D����O��`�M6��{�7#�޺�[��#J����zl77�,�_��խ=�ٯ9�HU��Qdl�!���X1�������<��T�!���O�g�%$Q�2�}�7g򧟿�����p���~�or{�!	�����V��Dǚٲ�yc���{�~ǭ�\�5��#�4���A��,A�`R�SPT�ZY- �x����'W�Q\S�κbT������G��p�M�JFqjh�h�M111j�i�J3��]e�U��"(�j���a��?fA�J8ţ������2�� ]dIQ�K�P�ciRvк�1�cƿ�YI
����-X%�=��P�R�GбM J�v,��C�E �����������?CoZ���E�f��6�������ت,,��v��Yq\�l�#��\q��|�Wݖ��{m�o+�u>7M�nr��RC�dz��ةÌ~�P��@��*�K˝�݈0r%�����ݝ��;���Qn./4�SP1�G�FO4��ꃉ+~�����7dd�d:�;���a���b��s��e�.��}"p���y�V�2$��p�p��o���~%�ִi�FS�gg��Ἷv�ol�a�9�} ��fPfv�X�58��r8b�koal͋�/�� ��������z;J=����]�`�1^	�����}9��;{vf������=Jw;y��˞}��SY��X����/������ȱ\nȮ���hƭA*��-�m�1�@� ~� �M������#?���u��0^(�G�!���5:���C�iH��Scc]wC��:������C�rPf��Q+ۀ3HF��4�g��L޼{�NAݬ����3�`mK��}t�hBº��'Lex�� ��pOs�AvJf���/���͝�hįj�����t-/������d��!3 ����=��X�3}{���!���lވg;I��͟k�b`�i��/�"�6A��8 C��=�'
q����em{���s��k�w�c}��П.�&S'�=!����Ru�V�4e�8��l+��A�<u�̛Cҗ ̌����5����G�U�֪_Dqe�aLj�ر�{����=^�3�+������ T`���u���N�I��d �Y��A+^���#�[Zx�d>A�f�{sG)R�S��`���\⾽]�s�d�i��������!�Y��Ef�+y�_�f��[��aMl"��4L���s[Q�>�:9>����}]?{d��qw���������єB;��G���_��o��i�#d4������X��	�ѓRfF���	\�ÛCMkͨ�> �u�.ڤ�}�&6v�hl���ҹ�$�^V��n,}��܉G�9�IU�������nY�TKX]YP�O���[~J�؍Ðg|��FU��gq���EX�/��Nçmٜ�j�Ggݨ��Q�{�d�}ڰS���k���3��Aw�y8��2�r���y�1^�h����Y��!l�� �^����S�CW���ϸ���k��:��[��_�� 2ԽT�Q:ﱕ����`дq��6����g�U��Aq�(7�=�5|�6~0�څ�(�L l_�I�p{%��7�˯����� ���̝~��� a���	s�5��2Aϲ�`��i��xF��aԡY�6q�P��:x�e,��6oa���ty�@b��y��b+�/ �$�_��s���|bz�<�skJ>�ج;j�,"�L�=D7 ����ə�Wo���9 �k cs�_{���"�� ��TP.���5��*�9�~�S��͛7�׿�M��������[R�G��p'7�hn��=2i {�3+f���ѕ|�t�uR<V\M��Z4�A�P
C� �������7�0fw����澧 ���'G�\��:�y��ugz>}���G�@�1��d9���(��� ��ΎY��/�����7���������������~�����F��?}b�s�����Z~�uyys�ϒ�k+��y��J�[�~�A����N^�|�@p�ǵ����6���Of�r�@��gq�o��޴С��!7�r���fT˦ ئh21��,�兦�2|���G��uGc��	��r=P�9j�S?&�5��Z@űA'�{^sڅYB�wl��� Dw�$�>���S�����O���~Rn0ͮr�qqCG�����Ne�C&�q���NDh�֜[;�MP��9��`v*�moE�����X�!.hŕ�ɳ��*�/�H��5��Z���c�#��ފ}�ݜ�g������������`�	��f��3��2��l1i� ����(�g2���)��d���H���l?�!�O0� �
�D�E�uQ+�҈�τϬߓ�b��>��4 �Z[�"fIU%�z����bJ���"{�46G҅��.��ߟ��TU�������4�M;����'�={�M�m�#���<�U,c�:�Y aev�]�܃.���ȩƒ�w��fKva�Pz_0�?�l>
���6��z��IE�W	���n "y���b
��[a� �e0E�5L��nlXkb9
Ae�������X���s�0q�#K�5G�<��M�aBi�e��� ���6��b�b�2-3i\x�m�ٱDp9(��<D��B#gdGԯX���:.gˠ��͒%��X'���ez˃������O+�A�d�qV4�?TTLs�Z����[�#fZ˼����d6[ ��OĢ��E�6(�zK�N��%?�L��"���Q�كM�����D�A����4^J� �tK�)��� �@<�]2� `�2e�>������tq��)2�9��K�`���F�۴�[2Zߞs�G� D�OhXo9�Y�U$�%�L� ��zb�I`V�N���{��o�a܉w%-t5�
6�qc�n���C=�c>W���Y7��v7�is�X�{�
��\��@0H�eƞ�M�'�ON�ڿw���Ɔ��Tc ���G�qN4@H����Ãz��2+4J�8_<G����o��N��L��\K�����i�!}IQ��=P��?�g�>�+��>��z�[d蝕��AK��k���[��1��9���/_�" �z]�K���x�� ��q���m��Y���ǖ�-X>4,� ��x,9�a+hhy;��\�'t&c��vC�����������5�����?���5A�;�(����?��~���O��/	�&�j�z���p���^�����r F�#��'z�%��ڝ�%�������%:�����ݓLl�}6�(�;���K�-��0|����eȻY�l�#�K�H�6������bp[��6H^s�0���c��ޅ�%��dܭ����@���
{��2����P$�}71F
@�I0��0�Y�/�����.�%��;_+k�X"I�_����|8�fcT?X��boT�%Sr��# O��� ��Y��e����䊀��t�Ը=mt�BG��T�kRt��ɄR��)��|R˻7/��n��x�n�Tgj�Ѐ��ώ�4��(4I�3�q�7 �N/f=�n#`c��m�2�d���f��$��ny]P�t>%6�t��,��>Q��I�E&�{&��b��c����L׀(AD�rp��sT�KK��-�dUV���
��6.A�� nRvz8�rdCKrL�YG{˴D�M&{'�S�~x|��oМ�s8�M����?�O?|��`���d0��[^�������r6����dKgݓ��m�[k�X�_�y*ZL�!Ji�f.J���j)���
����]^�S���f�Mj�#W��j���&\�|��;1��l��Y��t{��M&v28�Pۆ���l�\7�)�WېJ�w��9�}A��Bd�4S��@�BX����*���bk�������O�xKi�� ����y��>7w���sK��#I-D�(M�uc���h��jDR��XW��n�43=���=��}fa�r7=���MC���|��I�����k�.�Q�6Y��U��� ](�`���(�������v��������C����ke�T��,hD �����M�k���	�щ7��_خ'����1Q��{���3�������o���H��ٶ���=#���_%3�����d�v(�-;�cDR�P�eD�.@Z7,�lغ���3u��1upl6� k�ݷ�ʥ�t��c�,J��'��3�1����}���o�6���IL;W�1A� ������M0��S}��f��L0-�6�O��������P�M&�d�G!~��H^&�g:�Ƌ�$����[�ȅa�20��W��÷,�n���^M   f���{M�ݝ��".�>�� ��
W�x)����� ���"����Ç��?���,1	m'��m��SwH�����Ʊ���i}�.< 0���o�5A���g���_�Ң+�C��%����U|�>~�(�>~"p[� ��Vڢ,�C����)��monx=fO�9�s�6��a9��R�r�y}���I%(Xш'�Y��V��R���=R�/ ��L� �4�|M4V���D�p_^�>�5�|��zGaX��uE�����߳������ P� k���b�9�4�uqo[7:7���mx��Q�}�[�YI1�79Pcldk��v<x���ִ߸��98���1��:)����S�x��9�o ̶�Q�C��
��G�Ƃ�&,��AF�kȮ_��pK
���S�����	��e�{�t&�e��<5��\kP�g쮨�X� ��1ddAj+_�p�1"�P,0�oأ޴���cc!���K �tq|����f���C���2b�at��9ű��nK0�׋o�@���|���Ŵa�y[m�:,��'z.�@���}&M�*w�6W��&���8�wX��Vv-6�k6l0DS2n
�^Ǻ�g�ـ��x����l�dD݌���4����k�d?�ǢધC�����A�U�>D6��E�2lZH��k�+��Y<v0V�C\����lI���6)�<k-�كf��w�uy�����+��-��dڒP���m{��]\^˧�+�ίu�\o�Zrʮ����6��"��_$d|�n��|A�j"�ΌI�� �Y���؄���7�i����a�9 [�'n|���65�ay\.e>o=Ӵ�n�'��gc�Ul����t��ap���5r�1ѵ{qa�� ,3ˉ[��@�l�o�ȥ��j6�/��5�Nٔ*!=�R�0X��y��'s�fY�)@�b�7Şg�a9c���x�m��\?.um�sO- ?F�5S~V�i|�f྅�⇏��Cp�<���d��,E�1�2_�5��9l��ܚ&
�v�4� 6���}�?`�%�NH�z���-l"�P4Z"e�0ضI_{?h�Z����^˕X&�=��������d[���H�Ͳ���1|E@�1@W���{����*���~d��A���2x7�=�t���U����o?~( ��*�z��bq=#�~���� �Ei赆� �x��r����6W�+���������	�{ހ���.魒 
����z_������ޘ�����!��ǹ�m�=�Y �Ã���<d���&`W�|���d�?���o0K����R���O�Y;�Z��X%t�w��$$]�)��+M|Z9ܟʑ��ӣcyvr&�_�$��u��T�}�����F4� A���OL�)Ǘ�l�涔$�M&n`풝(5�%��^�2���S /4\���4���Ʋ��v�����އ�.PKǃ��[�2�ޔA�O��p��?����3�uZ)WU4I�y�`AE�3ѬO0��鶪ʂƆ�l�cz�6̜�L���<h�C@�W�dOq��}���9` b`�rmT;�RK�8�q���L�z�T���<ɫg��w����3Z!��z�˛;��_���!>XJi���� �#��rؤ�=���7���+9�l�16WflU\�A3���w͊�AƵ��D����A��7�f;X���1l^��g�],tWrx|*'�^��W�ҫ�o��W�m!�F�`�Y�����`<2��;�j�F�I�u�a�n������v�V�&���@r���qO��Yn��`�ez�����3vB6����+46���C�`Q�D��s����ܻn�[Փ�!���i�\S`E��y���)hs���~#���|b2p����{�T�r?�b����'K������&98M�ڌk����A��,��_]2#�2�к�7�̨s���2j&��	s5����R��nT�;��\�5^����Q���oN�gN�9�ݢ?��]���ʃ7������_+г�>��x/��w�_�5ŬOf�ؓ*c���J��Kf��
Z-�5wy$��D��ۯ�sO�u ����]hΰwX��ේ4�hp����>r.h�2��H�Z�k�#�|?}��g� �6��+ �}v>��`	��� ��y�i�<A�6c
�	��=N|�#���K�Ϛ�a�ahsk�ɞ.HD��c�0�gi#��q��{r�qgrr�����9�Q�T,M"�c��t���DR� �e(n�BkvòC�����G�s������0����Wv)��&��a���,%<�ue��HV�p�k�q���qW!��ѣ* �:�k<+ �̙%P ��n���������1�����<y3���=�t�R؉0�ŷ������i0y��O�"��r׽  �����ޯ6�K��X�����TILN����%��?c�.i{]G� �6��2Y`�*�5x�jot�H�l ���{� ���� )�a��j���\޽y.�^�h<=���#�t0}��b}��r]���7���)�r��
��qn��q�XStsd\�+_��(�Y���w�Xk�Y�}�M�щ��-:e���|���6�����Fhz��k]rFg���3�k� �MP�,�c;����4��\�ML�.;���|Yj?��������Jc7F�y�	���v�B ���:���=<�����𑵁	�~C��43τ�Z��a��n����2��� �.�E��z.�z�_��ɟ�%߿{!����Z�u����gE��_���Kf ���Q�@���{A-5pl5�A�7.֓��Svʠ���w(�fSJ�ذo������~'�O�ʍ?�^���ۭ��e#�5\�M�:���P�dj��#�?|&��P��z��^iS�������e3&h���)(�(���1���nZ�@���tRi@��!86���5Z�ϵ���ɡ3E��.�Z�����;S�%��Щ�e�ǩ�c�u�z�X��y0]�,�����1'�ˈ(�l�!��~^�s��Cc��~��}��f���`�1�ޓ�@~� �\�΂k��̒��Z��p����?a���+zO+s��5���«��CS��<,��b|����S�"ig�be :��F_�V�����`��,���趃�������?��q~	`a�|����*��d�v=Jp �XI��<���|�ߛ�*e�.�TU[�i4�P� gu�L��$��fzwc������ꆆ�(���YC&/b�Ko�1���I
�!_C��g_Wr	�[i�{��G$��e�g��k&+
¡�B�`{#t^���M�U��K���Eo�0<�P),9�6�1���Fw`��vUv F��D���O 0��� ����_�J�3��އsk�<c�o�7�A���rQ������WIe.o%�H>�6����,{�H��\$$�`�`p�wޫ�c�=�0}�3M�j�	�<�-������1�(���$ 0;�q�ha!�p�Wt�#T�a1�ٚ����c���d�un�Owh���u}U�M�̑$S�\�㉏��٧U�� �~m�u�g� Zl�g1"M�C���Q���`���Lל������W�rzz �{d� �7_@��m}�G����;&�M��q��X.�^�W�#���, [�Ȓ�O�;K3��=̂!-�-��T��<��un�t�OC�� �Zk���b�A���������֨����fe����DM5F��� 욳�������n��Q�ci�;��Eq�uepdDg�w�,ۃ�����A��(���X��'dbpiW�z(xby�G�jJ�)�������ټ��G�d���Y����.�g�?}'o_�`�6͕ߧ���_������7�1��E&�' ���B0k�">AJ���f%+P�+o[M�yߒ�Hl9_��6�	�,��/�ȿ���~�?���T�.�D��@�7Q����a�����ō��p����Sщ�<� Cn���o5���S��O=����� �j��F)	l��|����J�YP���"�'2ۃ�\�NΤ���ׯ�r3C�wxĲԚN��Y@p��Lo��s	�vhw��3�<=��ܾ$ 8��Cb��vk�y��� `53>�
�Rt&�G�$#ꁃmѵ��B��"=>\ɱfn�{�9�<Z���k��KE3 ���@�N�����G�8cq��Dդ�`qtL?.�kh���[]w�O̚��>㷼<VkO�Wh6y����{f�6O����G�',_�>�D����+]ם�{K�{�?��=\���h� ��u�l�C>��Z�k-4&��i%��Z 8�[󖃠����ָ�n{��$�[ݚ����y 8�����IX�9����4eKڨMd[��W�dP繖�w�˯��Ȁ��T d.�$"�ƬP�����n�8�{=O�O�M>���2�H��c�✪	� ���\V*(eU[�V��܇���Sh�����.�{��7�LfEϛM��pnf�G=��.y}���XV����s���,W¬��{�O��! ��?��=�	�)1}���ˢiu4md*���N�����]�cq-����q*\�#�Ua�ăͯ��k�b�\U�z��ټ�8;9�:�AExm�>GT*g(c���K��Ur_�8�Hp����y��݉Უ���R�"��v9ώi ���V����a�]�3����'߼{!/^�*�Ys|u�Y�Xg�%�W��q �/m4�u��M~`���o���Ƶ8&e=��}�j�y�Q�GPV;.A�M��jEb��o�e|��Zx��@2�A���n��e�-����>�G�ƣ��x��EVu�(���ux�I��/�n�d������^yf�<���C�[���jdE ��X;C�l�^��푼�9�g�������%�ӻG������m�0ޤ�.�.ҭ�M���dF�.Ǵ~sG=����N�`N�Ȁl�\�������n�}o��tf�x��ڻ�4=��d�K3+�(��6���00(+U&�y��Y�P����AjO�N�Q�`�&&]B���ypl?�T��g'�,͐�N؋[8���� ��vqn� �BU`Ֆd�k!E����������Z {sUM��
� b�+�^�s��a�y"iqdS���e%����;��������`�Z�g_���tOB�Z�X���ډ��B�@&�z2L�G�k�}g%����f���n���_(X���.̿*��. \0����|y� �,͂9�Ȝ�[j:�7���H��m����c�0� ����s}痢ٍ ��yO�o�>([����={��6x�+/�����|����@��(�� ���b�>�Xj[|uu�5��	�=��M�~��9$��)�&Zu,��ق�˟�,-��c8��l�f�i��ʑht�|~���Q�Ꭰ��	�����u�1Q��hΙ(`���:�O�7zNk/���b-�n�3���cؚ2���SG&zM���M��b��Y�A�� ���$�[-Ct�Õ��j	�)JE^��`d�̒	���ɦ�M>�2�OA��ߍ�ܒcꂮ9��se350m ��
��S�/�L�~{�r�G�� ��.�ą�w�gn4��^JN;o,I2�W0ާ�e^<�;�Ϲ�Y#��/�!#�2�^��m��Z%�J㈜��w&����šAz��-3H�M���@R��=/>]&�&JG{򷫼4]Jś��z�uk~BX{c�H&�Z���������߾��4	=��-G^Sβ��1	���g��z��ޓfs�?;[m`9f�V����r�e��h*1ۉX{1S9tz�l��l1�T`���	"�jV�?Vk��zv��Xn�G�����2�fx^�]�k�� w�x��%GUC���p�;���h\vv�1'�/<��QP��"7]'1{�X���o���:d����M}��T���-5-�)�>��>ȍn������h(߮�;����6L�ǂ���N���c�Q�P�B͸�O�eӘ�m����t~r$������q��t�Uc�� tO�Ol��!w��:�Z<��;�ezv�`l��1L�ݑ�Q���QJ���;x� �w�u��Y��'S���^6��4f�10�bf�[S_�6p���6�m��oب�n�	 n�7������Ť��kf����]]ޑ8��;����15^��|��\t����Z�J}�^��Q�\�yWҖ]C�� �C�vgJ�8?[�Q<U�YL�P���N�)��ٶ�oϓ�<yp{<#5K��޾���'����F:��� <]Ȟ�翰�����B|�6�t'�w ׃�-U��mp������B������~e���c�ݫ�S�< K��k`6ݓ��S9}�R^k֊�f:��M�F0��f	6�9��X/�h�Ƶ��׿���
�k+��а�s&��o��]���@p����l\�]b�j���X�QY�j3���by�����\t��Kj�(�g�o�Mz�9�)�+m=�W'b]��7r�n���l*By�7��2Cܚ�K0ԛމ���g����cVsʾƐ#ـ]���I���Mo���w��ˮ�������M��J�;��5=�lH6��:��d%*�2���;^��4�x�kb�-�(3j\�t��Hv�pb�rAN#KQ�O��� '�.9 �. K��?v~>7�|Ubu�n��¬TR� ��d����JQ	�+x-.$�5_/������j��^oܽ_|\]軂��������!����j���>���������n��.�{սݯ���IG�I%��N��������o޼b�-�:X�-�h��g�>�Q~нq�Qw�'h`��N���5c�� ��W��i�86�8������ݫ��'�g#�����k�waj������,[M&���5��Ï?Qz ���n�N�[�d�3ĳ�W
j�������`pxg�/�Fb�*���3 �et�u2�Ψ�O�L��VQ��A��q�Rdǎ"���RS7J�����D�aVZ	�0������=�0�����O�r�����ʴo�Cc��`���J�:L4�b�,�Dc�������̽��p9��	zZ����)�]�%�����	-�0�ԗ���՟���l,6?X���v��W�?o�8�<*+� �|��������]u>������{���e#q��V�\���g�p�6W��O��^�I��H,�[6(����}�����n��9����nŒ�����] _t/�;����A�NÆ�Jaa�rvޞ�/4�`��#����g���l��/'$��$�Զن[ŶdM���um�QވR��;�t~���h�L�g��lژ2������ �N�|�p�!%X� B���RO���@���Z��6~���_cW���EO�g���t�A���s�0#s� ��a%׏�X�ty/��O
dz27(������P�q��n��y�� n>�r�۴V�٘b:�1�6�Cj/o4��o��h<@i�qi����:ms65�EAxc0�|� ���ȣ�%H$"�#�)���8��
g�-�����rlp��e�q���� �ҡ$��)]�^�׿�S�Dbv@�?�ևl(�O�\�w�z��3ۅ�w�94���ڪ%�e���5ۛ��S��ȸcc��M�}�l�)��;�^�If���Z�	.)>"Е�`�-_D���|�s��<��/^���'����U�R�l�����@�O�}O��`���B��QJY���u�_ǈ���T� {��v��O�야T�Ǘ s)�a���d����?	FTX�b3@��� �����u�� ��w���������/�1N�����ƈq(�i!{g�L$o��Vɨ	95ac�� 7��7���߬lҌ�����Sk�Hо0~�$�g�Y7[딄��Y���8�Ǫm*������28ӂ2���17��{+�Yi���F���(y/��t����K.�U,��t�}����X�f�F�vȪ����{����W���h�q�C��~� H���o޾�oD�����_���es~�+���̻���|1�$!+�G�/<x�6Gcҽ$��9J��b�Ǻ/kׇi�u� |}��������3Y�������=���A������ѕ�m]����+?����Sf ���D��J�
x��>r��cW�sl�)�	ݗQ��E�&b�]��?�ަ��o�7����5�`��40���z��j�V�`&��d��^��IC�W'}���o0;&��uFC�"�`�0���\V��CIMY�g�a��g_��L�|��Y���[�ToH��1����l輱�5c�ll��	���]͹�b�U�jQv���qi#��{i�a���tJ{��\9�%� �]_������"�Yr�ύP�Z2�/5I�E9m�	&I�뚄/�o�������� -J�`{��<-����ߡ��Cl��]��ڞ��o8��J�02lɎp*Bc�1Cd���9(^����k?�I(���@�/�\<Р|�����!��H��v����&�p�E�h[姥� �3ާ��nod�t�ʃP�e5X�$�v��Y���	'�dz����h"耭�I���!1AXo}&�wC��_�����>O�+:�}h��w�k� 	@���yg��!*ށxT���2-�ao�ц;;0(�-K���2BY
!���1��(�~p3��~� ������tu��/*��w�a;�*�y�F�����μ�YʿG�R����]#W�a۷�9j��{Ɛ��U哮 M�m���ِkq@}�X���WG��H���#���Y#o_=������� l:�e�`+;����,�t6�%���	�&a�Y�`��I�ĉ�p��ʁ0X2��L\�+��%��\�ܻ�w�mQ,��W��]�{Z����=�4T��w�MUcFꍁi����Ɛ|yp���vM���H!�%������₞CT���]�T,6ۃI���OnuѳL�c��d�k^(��.��m&�����b����LA��p���43x=d��	��R�P���ӵ����=6Y=9+n:j�|��^�����9V,��c��� 3�泆Ǘ�3�Q`6h&��mz3���UWc6B_& R��u�,��fr||�)o^��xo��ל�1.���k�R�R��pF�41C˴R���=�Tl�_�M���M���(
<�s�/�IIv*�� %�=�~��X{v;���&���xllǔe>����G�+f�g�����Eև�M*��Y�3�k��^P�9�A-xq�V A4ĮM4�x@���"���y�5zXҞp��z!k��+����=^o:���}�Ҕ'JS��k�p�M��o��~��f�r���> ���ߦ'x2_6�9J�{5<��2�H{��n���nQvnh�`W�ٞ�W8���G�]��17([�(�2�$��'MdjطaL!6��3ǈ�3�5ơ���ƃH��h©���Ѷ��5?�`�m7����:�a0{�G�m{x��f'EI��}v_E�9wd�	���e�F��RlX�G9Ն�oM/���A� .��D�����9z����>f.�n�bJ����G&v�wQy���Aی��<f���対ƭ�yϴ��]f)IyF�1�$d\�Ï«�W�?�G<~�{IaPv��˟ߢ܊<��a�	�� j;{Q�3)��g���P�+/{R�c|A�<i�r���߉;���D/��ǆc�$;헍�Zk���7o_��?��o�+�T��I	$�3���ԂN��F�U6�9� F�+����(Y�M�1�Í�B�zpZ�
�j������n/�z��MI���xa��Ԍ�gL�MgL��,���g�4 �R�tfVC�Νqi����0H�`�fYc#�X�ݖR��#i����ƙ��N�t�M���[?n��<-�����8Ql2���C?�0�n�޼i6�{�j�c괱?Ɛ�e�С����4�=Y��R�z����M��-����-���̑-i�\Ă,]�������K�m)��SX,�� ��Cy�옝���*?����9�IE�߼{KT~wy-O���<4�i!&�ʁ�Gǜ��N2\���ֳ�S9;=V�����\^^����+�,ph�a�.���b̂��:t_N�M=p���������?�ih�jo�P��س�ڻiń�^m���Z0ΪÈ"h�H����6z�lh�6�����D]���G#��AE�X�X�N(5a�*��4"W��s�vK�T٦��eݑ��x���.̺��̭��I���q�Jʭ~�]���|���@�c�lYjB��l�=]e&�5�ۘT�6��Z��Rk����5`��JA�F�e���o�SS&),��0�ƳV�`oyD��2��'z�mh���!F՜�������t���md`�9��C�g��On0�2��0���>�+�5��|�ǐ�l>E[�^tZ�Ϡi �!sXK7i=�&��agh}�L�ibj�B�C���s}7�y,s��??6	��ǲ%�%�mM2І�Jf��q� &�G[��]�h�wo�O����^����䕉�%��s�f��f#�,\�H��[�m��{�d��l�d�=� "��#�K�V���JR ���  �`�|�ټ{��v@f�^�.�s�E�c�4�l��<��v�$|Gfn�gP���6� ����;Eb����������J|�ݧ��-�.K�<2��`S�yc�������0^�ף&����#� % �Q3����w�������O���o'W�-%h�it�~���rpt�j�h�{�ͭ�C]ݗt�L��� l���jI�H���Qߗ,P��5�%�^,�0��9���Up@a��KѴZ�6�xU�%��7��W�ݽ�#��Df�)��4"�3�f���\3P�����l�r��l�I�vR�e@"spQd���{��6bPv�+����f[:/W03C���7�;u�fq�И�	 h�7����!���+�	)6@0Om��� [�+Ya{�x��|��]x������i4�s�r��a�yb�����$���?�7k&���=<���o��˗
���>Cٰ^<̐�z7[vЁ״�^�;0�=��P�8<n.�����p{�!,��J�Ŝ�YϡJ>���2���g��a�^w����;�l7ۧ�MX�?O[3�.%�)
��W��x�*˺�8�Jfb@ݗ;�,ջ��i��Gf[�	̅��:mn�-XG�i˒fJ� �����~�g8�v��t��.!;6	�J,x�$���I�k|�Aز�$�[���?�-%�30D��`gD�mK_��|��Im��֍�c3 8�n�J8�L���k�W'����μ� �9r�~��Kg��r�����/�K��vs�lQ�����%��5	:��',0V�źq �Y�<rg�0��֝��YT1��	l�q�<�_ƲQd�*g�i��B�3���D;����~H�j��O8C�>=�,�Y��׌���$SY�k�ց`�@��ń�����ٔ��8���ز�e�(�����@૤���K���b(W-���L#0����PD��`��v( wȯt`;�y&�e�9��c����_��>�?�v?� a;`��K���f"1�k>B��X���_}_�Z(�Y��Q�:
��W�wC�:�����&������@Zr E����&_��3��f@�&��zf�j��>?;��}-o_?��ә`�8
�m`���̼x�N�#����rs\3�.�X�+}O0¾6D]jc^�O��ިfl�ÖS�S���<j�\�M����oدf���ܙ���M�a�VG�i[,Jnz� ��pZ��$F+3O�Rlٱ�j�$�^krN��m�����ab�QKAO����f����`{��� S��5�Wgd��xp|jo�G��;ol��6Ks^~��� C�@�11G��fɮ��6D�@��7����M��������;z��u@���{���ჷ�oҁB�[������� ߲�|���-�}�����������o���?�����#���cS�|�3�ܙ�y��� 䃞A��cp�XM��׿����/!�E���E= �f�����rj�����g�7�}E�w+&ێ�����%�)tY��W�� @���ak#ZX~���Gc@Kl���+�N��ф��Y��6��B�����t݀kk�;���X�EYa��vB�Y+�͜�����-A�ϲ��sGI��кL���m�*l8�I�W�E؞,�<'�Vs��l�O>?e�l ����`
�&�a��-(`�ƌN*��K�(;e�Q:�P��M"&�6p������ ("�묜�u���7=,A��B��\+p�5GR�-B�~D���MĿ�Q���w-1�H�R��{F�`�h�s�}��
l��0i!�U�����6ޖf�����
�|�!B
QKLA��C>o���6N�;�$;;�B�9����=�"��|=�q=���؞�یF�Y��K��$��d̼�Lb��Ԇ�7�	�q.�л���]��z�d!�f�)��^��)p ��������-��㕝��Z����o�[��hO�r � �Hz��u�8C��Ư>�3f��cd�F6�Aÿ}����l}U�d��w�S���6�Kv���_���0�R�۽�9���:�G�aJE�T�#�h����F#Ƥ���<g���K�!���s��N�X��/�#b�,vb������MaGr|4�������}�悂M�{���k9>=��ޜIG*�n�B�R+�s���Bݢ�6,�v��,d��˚�&{�n
1�Han��#�,�l[�Wx'B3?_t�Zi25W�䈯Hг��`��k�Ǜx������l�"fv���[c�R�Zj.�Q����*9��0fL����&����LV�^�M���ɱ�grx�� `"Cq����g���`�/��$�@�lgmkǜ�BoA�)�o��]	{����\��r�m��6|��g:�@`+n��Ƒ.�8�i�.Nf�h�E��X��nl� �G���$U=ˣ @��׃?\�-9�C�G���?�`�,���cv�<����Ņ�ܸ�ۻ[+\��b5���B<X�eXk�3H`����V��X��M-��gh=�\{��Xn�uA�6��g_6�lڰ���|�C�Q��yʆ1�����G9�c�՞U3*�¬��LX����F�A�X��e���p>QЅNA#`��ph�ߓ���Rt�z�_��>�>n���^�	ڪ5�Rw'�1���ZկWw���Vno�,}B�S5�>TyTO|ll&-L�ϱ>}*o����;6+)�kH�a3&q.]66nR��_�l?l �:�)�&�Ed��g��ϻ�'\t{�T	Z	�O�3�*���_��|������B�4n�C��1o��R�qx�l�M�1�6�5�P`�M�,pdE�̓3��`�3pݎ�O+���I�,\0��EI3�77y�&J���W�[,q�\MhI0��Wm,x�qN]a�(w���R�%�����H��N�,�J9�y�=k�w�,���R�<ޯ<��ʟ�*���;�<6V��q��#��6��_vB��$S�X����w__�������R ��# ���#�e�x�ੂ��7��ીT��<��T;�5�C�D��D�7���t�~��3�b"��'����2���0�?�E������8�`�{o-o߾�wo��^ܲ��a����N_����s98>����{a�Y�f�kU�x
� 73`r���=@��uc"zȟP��a�9�XVޅ�q��7�	������H�P�}(E�v����m�Ӥ�-�=���7v�BS0�6�P��`�)(5Q ��'�`���������왗����z 1_Ϟ��;�B%�-�!��k�ԑu��"�osndN��9�f������<�nK�U�Ik��,&�LA߻�/�W��p�٣	i�iזE �,(���g��2�d٨Tv����3�MSfс� ā?}��>���''g<$���=��ї	����^`�`��ga|� � �АP����i|oj��3*5{�X����{SJ����'e�.��L�1V�5����Ѥ�5]�+����]���l�9Ӳ!�4U������(`�=���8��Mk�%�2+,=��Da���h���YG�qjJ��U�L:�)�Ëk!{�/�U<>�ȇ?�����d��@���;y�Y���3ٟa\�J׍>��*�{�[)�F̒\[RٳB�+|��>;v��?��ǇK�Ory1��é��3i�� x/16���1|����C���^�e�P`8?b�l� 9�%q�����#23��p�o6<�hxQW�9�3�U6����v�i5a������=��|��H_��3Ƃ4l%��6Nr��w�Y���aO�2�4��D����zH�AMe̒8HB#�yg���"�X��n�f ���cfli�󋯓��L�)ƍ1�2a�l\Q�;�,:�I$«��\H�e���)��A��)!�0?'��sc�0e�[o<�X�h��a�b�A��1(z�ѥn�U3��NlZ����5`_��s��ZR�3dB��t<��2*���a�� ���4���~��%�o�K���hX=�����h|���,�4yd��v��"v ����;Iė��%�+eޔ}-��X�� 7#�I�)޶!J�_]�<�H�Ʋ���� �L�5�1� #B��N�֞���Z���?������7����v�R�5���lc�8rM���pdV�il+�D$��J�G�����1�Щ²��B��(�/�uـ�W�4ٽQ��4�ޗ��	1�xB�FӨ�:�3ЮE��� �(�Z��;�,#F��7 �]	���ٌl����}�S��#Š���6f��A������d&E��g��P�J-F�G��wa|����s�j�)8cq<hM�0����K����I�5����Q��50�0Ǫ����cR��:�[��:�S�?-�@��tГ����Uc���sn�4��+>����!��e�5��9�j�RdGقo׻_�u<ڬ�8#�B���6Q����g"�b��7v%���������@�7o8p�c�t+��@}��������lA'
�QF%{����k�r�c^����Α��� ��m��h��f`���f*s��Vp�^+й�(��3yX>��C����s��JA)5� ��G��v�6�d[���X�u�^v��]Row{[ɡ^�ýVf �>?���N�����
���<��K���3Ŏt3:�FO���Z�uI1�:�z�!�	;H�m	��%ܘx9k��C����uL����fOr6`�z���!X��e�S��p#�4�Id�c�H���)�+I��H�����Z��b�S�����&�zi�K��U�m;��l�9�Z��3`L�+兖���d�Ò�}�,��=�rjfƲ�1�2l�A��|���8xّ��`�M�p]���P����$e��KG��q�� �wk�ސc�T���Y wR*"��'w9�����"����-�7R��.��߀A���j�}��;��)�����,����H!���K;��{�dؿ}�4�u-Ǔ,�*}um�ُE��+XR}q�񜙾.ʾ��S�c��Ȁ�����8ě2�{�AM������y���K��Yr_� q1YD�Hf2��`WDN�e�]�s�nX�^)m)�Gy=����/ �����`���(��,�(3^��{#glo�rM�j��6��i�@g&f� 	'x�S�M\����]���=Ql�wu�TF�</ZK���t���:�����h��|���/�����|Bz,S�ҡS�7t����i���̄�3�}�V���_�˛{z}x%+����1�r�pb���pk����@�
��[vu5�&�֛�=��]���+�E	��F�����PW�)��ˊn��%�()�u��z����{R��D��7��~S�fP��s4�
vfm��,S7��7>L�=[`0�� ���Z>�]��?�V��^<{%�^��Wo��}�ם4kͪA9�>���BSh��$@�y��[kǟͧcF�4�R-�Ӄ}�q��cls)���ۓ��5շ���)�zd�o�A��{��ۗ�˕�]�98F�8����q y��7o���T�l*A"����k����+�"��5���J �@���nl�������4�}����N��eSә+t�R ���w���%�k����7Y�1����aYp>��YF�L�6v�]Oz��`�X<s���eX!I����	c�!�wY�2i�&��{����c��!��}�g�<��y�q���W���>�L�iͺR���.��8$ݜ�*%<�'a�Zwl*aI�5mR[�k�zg���u4�5�ɮ��֞GN��y�z�;�V�w �eMg6����=�5}נ�D6��ĵ@ l+s�g�s��]��X��ܞD���5��p�7�AB��fk��R��|?z��P�cg�Jt����8 _�]�����?VׂMډ�e��RM�ٮ@��_,�"��Ұ�)�y$ʇǕ)D��6L_0[~�ž#l�wU��]���R��b��jU��+�G�����_�u,Ar�(1�G� ai|��������4p�]32�f�C�"l��%)�I=�WHqP�8>:b������ř�m�<ْ��b.��y�"�:����jw]|�$�L�������7a��#l[S��K��3}i�2�BT����;��9q���@��V�p��ݡ��>�����,���Je�|�.�6W��H�KB��ƚ�ҽ�c9:}���X�Ɍ,�5�k��&���8�'Pv�X��M��ņ�N�_?����m���#y��DNO���Սl&9�{���U"��#�x�bI���hd@gf�:7�L1^��x�;1(�(���iMe��p�Mb���R �OX\�!��9�n9�-��F�_��[2�X��D,#��-rxxȇeL8�cS^�MS2�S%ޜ�\=�l�!�@9_L��1����~(�0[ˣ�>:`0�{��h9���\�l���&�)�x<du�d�ʛ@���e�άi#�&�5�뮉�t�p�a�^ق\OpΡ�����ꁁ���m�ق�6�KF��AL�P�]G<b�������7Q���X�Y�3�rh��Ҧdk����}��BO���k�/o�< _(ABK�[0�����86a!;�]�X����k�6Ɗ٠�g�zOPZ�D�	�=�Ъ���X�6������l�Ɩy7q��Q�rf�zC�`��A�� #�~f(]�m����� ���])�ÃH�e2�(-�t!��H$mv��gӇ��(v����1@��a{������۲?���'Qhv�q����OB@� ��Zs�1�H��zAb�o:�� ��nJMvZ���|9k�R�P98����5��4��5;+7ވ����1y=}�L��2�m� �b�_j���� �Ї�ź���$LI,Z��W�q�P�����c��y��j��b�`���롪�8����x�t�����Og���BcC�.l��Pg��`���'P�C��$G�
�#��<"ڍ����ʭ,� >����<#{;>#��s���1��6@(�c^�'F�KLnԐ�i�-+2V-�ȼ�^���uq���='�Ę �Q�$x[�G��_��>�b�#�B�1�$�������X��������R���G��z����`��P��m��ղ�NJD���I,w��wp�OxՓ��/�0Cd_ى��Tb3�B��q�Id���)0zsQ��z��n�3�F���_�8���;�t�(��J&s�G����ĺ)iL	q�-5��1r��뜐h ��+>����/00�ñ,fa�[�{g�@����r�_�-YΣ��9w�Ն��W�y���'�R�_:A��ռ�~3��B&cW�y[�%��Cb7?���ZZ��s�_�	�����H��YF\3xn�2F7�M3��!���M��H��_lݭc�C���x���6�s<E�Ɍr%[v��� ��?����5�y�S���n�1��FA��Y�M3Г�����#��L�j� 3�(��@�A�7�Z� =wh���A�4����|�ؗF�	�W�kj� �K��k�e ��P��i���Q=��J	�=���ޟOy|�sc^i+wNd�8���s\�V)�;��E�����b��R�3V�����&J�cI��= ~{����u�1ݽ͞%)��/X�,��9z�]UY�W�~;�GS5{ ��3�v���q�q�CMMM������N
I��B�$��L���(��4i�Sg{>ƢۺR�s�M{UGۄ�/����]َ�ܩX.�W��K��z�Ӎ3q�h٦_�Y��D��k6���[��,ͤ�����'����dJ?! 0��j�3�˪�� ��`�k2���,�R�x���	l{�g�,un��=j�`mRF+�A��i�`�4lx�F΅�~U�W�Ǵ�@�r��$��BI��;ۗ$��� ;C^��ao�vLf����̌��$wJ��gO�e�b�Ơ�l���u X�I��6�.�aB��T��u6��Z����Ek啹!wc6���Q���|����ձ�)�/^�$�w���[&D�6�R*1s/M��X7G7җҟ�y��A�:��4}�>À�2ى�zz�=��\O;,yV����������W�@���������۴x0p���03zu+"��D������Q�����+v��?E�(�A��n��i  K����}�2J�=�Ill�9l�v�`&�c�>g��;W�랜�����`��m�f�g&��ӏ#Fi�rm�GC�_�=~&����a!��F�]�Sd����.DZ���#E����z��|Ŧ�f�f,���BZ*#��dD7_�w�fk�ܐ_� ��8����<<=��.j��y�c�^�.pوZm�����M�[�m_�U�S8�����k,�������k9�I7cr��py��������p7�P�b06����'���� .ߤg��w�����KwD��u�=[0�hF{��d�NL���}B� �Ck����S��GR�����6�����;6�yr���!x��Lkm!�)ۏZdvj?K����z.܅i����69@q���� SS�A/X;�j�Qh��R�9�"Z~_��1�?,�r�x��e�1b|-��#����c��ؿd�pO����L?�6^�ɐ�?�V�x����a��Qy�?��2�j���Q�ƺ	���c�8�ʙ��'m��umDl�M���@/��U�6v�"�ƙ#[<[o[q�>uх��L�8�ckA�BȖ>��e!Ho4еьiF�i\Ph��]/Y���2o�=P�$�`�W^��P?7F�EFIM,+Ƣ�N���������=7֚�>h���� �X�����g�� >�;����j*��sk؊�����y��;ۯU�Z���a���]Ve'z���^b�BKk�qۀ(�W�{�4ה5���{5�vi����s4�,�iY?��ΡBg,���̊�l�'����[o��v��� /�iL��I
p�g$�oYAJm���c���~P��A�;��d�/�i��
B�I袬4Z,J��?�9��l�l�qh)6�x�knMm��ҍ��t�i��UMa-�r�mm�P��U�� b!��
����dNhBv�l��z�e=ma�{�7��K��:���L������[�K�ď��o����s�؋P79]�l�N�4���)�_�t%O˵JT/�VU��&r/��IAZ�����yu�Ȇ�p����)�,�(�.��.�`-�d� ʐ�*�N����|d�˛�&�pJ�1��qE����A~��=O�!�J��z�k����xb�Y� �/�p4!(A
~l�Tg���~�V�ᄎ����ۇ'� Jȭ�
��Q����+����o�F>C�cYr=�������"u��l-�M2ٍ�u����T���_CV���!~L�&�B`LvMǇ��Pi{,��L���ć�jzr�v?�T��c�����]�Ѳa��N|�`�r�;Y�>7C�,�"H�M�A#��~��yG���f���ڴ�[}� `��d&h�Im�֭�<E�nH�x>�:�	n��R_��{*�A����ǁgb�h��a^���wj7��f�	��X+��-F0;�@f�ש�[G7 $g��h6�zH��(H,(d�T<�ʻ?��S�pPK�3�V��\Y�n)��m���V��\%
eh�Qi}D{�6u������|�� l�g��b�2��Ѯ%i�*th}��e�����g��A:�`O`٣fr� ��1�1u�4�d��5ܣͺ� o.���c7����Gz�k�2��-�ʍ����4��v��,նAv�R��k� Ҙ�\�u�o��Wb��c�#�\�Զ�M�m�%4�/�fݴa$v�W҃�^J��������a�`�Ր
���R��,K�OҜ�)g`�]0�61�\?���L�{v\c�i䐠[ݼo��Y��<���5��db�K遐�w+����h)xv����ͺ��1�<S���x�-h�d7���^h�<g�R�[{���J����g}���W��w�@���ϧ8��w/�3�����=ڀ8MO.��Z�^)R����>�j<��X�#�=�ؾ30���{y���G��y�c[�Iu�՟�h�\(��R~vO�d�Z\[(J
��L�z�����7�»���E��A>�y#oޢ�qKğ�whK�GS��`��GVMϵ5D���fK��5B_��������.��.��6�n��Oo��aFk����{�?����c��1o�����ܳ���{�6z��9����� �d���Q�&��ehVQ�3� ������G�����5RN�,�M�*	�Wl���*M�(-��v���1�q�N����q~`�R�5R���TN�}��������=��y)e�)�iƺaK)a��d��s�С�-2w��S���[+A UX���i+�Lư�[��W���X�2��?M�Tn6	�ZY���c��[���>��t0�T��1F�� �Z�a*Ԇ�&�+���Ӕ��EF�WW%����74\oi}7��j��e�қҩ�ĺlǄoҡ�`�@L�FW|��0݋������)�͞�iI�\���[��!ȼ�Y�`�k�,`������}5��:LoyD@�(�C� ة�@�������&k����^�7Ԋ6��v�d*87���O� �� �.���{���-{�M�4(�VF���k�u	��s3��Hc�" ��w��*���G�l�;������Wˈ5��R� ;�@ZR�r�tٯTA���}��߷L�>�J 0}�љ��|v�W+��m�޷���E�?S�14��`$-Z�PL��Yi0H���R�c���3R�A<@�y�N�U�1��/������\b�*cqF�l+���xe�l�����.c��'���r&���+�X��~�2�ۃ4Dϧ4������ud�P0�Ki��=���p�����p�_�+j���\6�0cՓF{\ 0�~�2����{-�m�6et;������ˁ|�ث�=��k.�h�|v� ���l��uj)��?-M��O���7��4��7o~�>�ĺ4C��p/��Y.�����AN�����%݀aL�%u%�ī)��D�oS��=��9�Xuus�(�������_Pp5�ă��r���l��(PY��h���K��?�N��To=K2���t�dzʮ��
�V�t+Xe��ݍ�����͙�W�:�b��>C4I�}�L`��B���/[�<qok[S��sf��=Zk��/t�9�-�;��d��hT���<��-�����9�b����AN/_�f�$ヶ��T�����w��؇�XZ3��%DڨJ��t޵%�o �^ e�1=O�q\�ؙ;=ꠠ�@K�ʹVf�QW��z�(CA:=���ef@�Y3�d� s�*U�Uh�����:�wi��P��{��]D�`7Y���:�����Ʀ2!p�Z�8�/��3]X���,23d4M��!�0�;���Ɣ�B��S���!��b� �<'X ��lrA@�3a��n��-yo�U2��U���їܤ�^��i������qCFUؐ���%g?Z��sv� Sa�r����y�8ޟ�^{�� �q @�3L�扽Vw_\��1���Gs��z�����=}ɎON4H{!�|������a��w��X�
��L���Z����6 �"���@��!+��MN�0w ���á���$6��]�-�0R<�v��|>���Iy�0�_��ƽ�����s �	`�e�>	�>>��W��g٧-H� !cfs��4�13PηL-E��q��``��>ˤ�\Ki�-3[@�}+��"�m�P�j9���yd��FGS��$k���0���-L���+|��I?t���A�J�5V�n}���LY�L����O<�_ɀ}|J�W��:��V�`ѿ��@�]@��o��`=��%A�@��&��B��Wm�ԭH�s�l[:�seiٛ���f�M�g�1R;hB;,��qO#�)X�U=-�c�m
��e �8[l�&��f��Z#̭n��(�u��ܛ�-i�����@wI�[z�EӢ�t�6�$�]C%�V�=�:%{X�
�Y����O��Ne<�|yo����B��lT��BA߂�R�WA�#Q��M0��n0�|��8�����Q��[��HFG[nz�� 5�$]##���EMv��R[�Oa(��g���w���f��-h�1�9fY L�&���a3�љ�#�m�<$�e8�ϖ5�#�+���2����o��&���GZl�b�D:-�6��ߣ���܍��S����ހ��^�PP�Q�f���V��W�x�q_�!Zph-A����rv��c@8^9H��f�����V��[	iNI{�>��3��Nx��`�s�fV���.[�FE�zyF�6�^��`� %;�X�Tb������5<Ps���  ce���f�[T�ff5��u$��Z����q�,�XM�H���g�	!��g�Yn@c<m	��&��c����}�����bE/L��lѢ���pk�����JYV����R� Q�Q����k��Y	��<@�t��N�x���rA6���^	��1X�����@k�����L���C-�YE���}MkywK透�7�i��M
���yJ7氡m3����Ͻ�ԡ�b�����9�v��{��Y�z�uQIi�2&>��L���%Ϳ�:n��_���>펃@cIq��G�d�sg��6��*5�Hw��ka��sdf�=g�����Ҭ�����J��w@��ߐ�(#��U�8;�\��y6��­z����E�A���C�_Ѐ}j@�"ȐnV�<4�J�G��f�+��@А57Y|Ѭ;b������zi6��矛7 �ѯE���ѳ�ښ���ȼ:nH fq����vH)�,g�����i��$6�U�J�~0K	h�6���^p� �����wt�͝Fd�u~����~NM���*���k|@�*�#����I��j�
�ۻy�E�b���#4w��_hD|����)x���
�z j�T˭3�g�@A�T�
�n�P�'���)��`:����}sh�63Y)�\nL���2�v�H��ȷ�{�/��K��ߍL��|�����$�J���D�)��V[
�k�_�Uy�B�c�~�4���/�[��C��Ƙ/+FȘr���W4A'TPW�cM��-��v4���X4CE�zm �,��Z��U� �xG��{�ч�0�&��UP��vL����q�b-�(z��/͒�O:_��K�,x��
��@��W�%��4ZUiZ0���e�V�͟�������Ҁ��ʨg��J3!��vdD/���Vݕ��NƐb��,XJ��lM0����X�&����)`%�님��H�8zpe\#*����n��Ƅ6χinBy�tA�)l]zOx�5J^Pm^�d;�e1_�z��Q0��i����v
>aR��Ohܺ���-��ﯸ���B6�G)���69�:�xz2�  �H�\GЌQw���X��7_����W/���^ʿ�}~G��'�Ә4K)Nf�����X�͗_y�>�I��I�H�&�v-Xb�~��������7\�@־>�׀@?�o�I�ٮ����Ǧ�ڨ|~y!��_t>����L~��g[���u�g�z�N+�gd�E��=��3`��>��������f�W���,m�幤^�LE���.�Ǘ�Y�k����S�j�@��b��)o�m�!t�(?�Ap�~�~��4x9�t���0�F$��-MSu��Aʷ|k<R�M6�ʎ�wh��ةx�W����	�6BH���,2������b� ҹy�Q@l�] '�Y;]j���O�*���kj��jP�{R0v��G��{aɡ�Y�ϑ��#ʭ+���<�l�Z��ƈ�6 f�`[}���+��r����� ����x�de���Zf�%�yA��m��/h)��M2���y�Ыh6�f�Q�>]�YX�� \����~��4�?��r	f���l���1؂���Dc,}lԉ�&����1�m�Ho�L�g���R�)���dj���nJ��*���!(��g`:���f�>\9�����;,5@�҆Q�5	X58�SSV���s�����P���f&
�c��>_QE�x�,Ɏ�D��tU�ِ�*S��E���  @߿�-��%4Za����:T��A��U2����~����\d�ڡ�� =d:���l�QX��}S�^�f��]���W,x�F�[�3;%e����;�E�&�&�ͳ�Y�ۘ[��
��|� x�e�=Gd�d3V{� X/d�b��b�Q�W'  �{,`ꓥO�Z������b���ɬ�Ї�z2ς�iz�f ���d��4��o	�j��� ��,e���@����}���Y% 0~�M�ŌKMߖVZt��|v&߼zI6�=ʇ7?��u!l<�6�cg֊K�u}wjAPô~b���.�9Ă탞���1[��.���>�w��ݯ�4����R���5����φ�p�\�O����l�w�0�����bU��Or�T{�+�A�sJ�I��J'dC�?���N��3�<�`�r2N�%=��_�����lG'D��k�	����;��Ӫ	�8�k�*w�G�����<��'��&^!�ߏ�� %����R�o��-���#v�G��m�?��8-�ޏ��E��y�4��g�GO�E�6�-*��=x�Ul`�<X���E�7Z���m�@nܬa�j閞LGG���Ԉ,�[
�VL��h��*�D��i�\=+\��8��ݝ�~�w���Z�'VS,��k$�Ejs�)��- _����͠Eʐ΅�Bۀ�6D3��)��9bʢ�;q5��<�Jc무���I�O��<t �3\���&·���DkE���¨�`}k"]�cyc����v�uI`j�v����ځM��J��v��ZC�֔��G�
(��}�>�0��e�9-'j�����稜��� 4R�"ͦ���B7p�_9��H�JB�h���	�UJ9�_&f��]���T�C덂-���FL}a��At����?��l��=�//��#M
a.�E�F�t8�~�QƏ#2uS��1L���F&����q�6�-�I\O�|��^c|��GQ 3����ѿ4�Ɔ1���R{_��+Ǣ�u4ۓ�޿��+=w���F�ޒ��o%�*�����	u_�Uzt<R ����h@4{��2�{�+L\b�d#^F�<�Y�U��P|�n � y�}XT�ď VM�O�9Z:ƖY?=�&7�ҏp)�Y"�:��Z���|�~_0瀏��ɑO5�����/�Wbg�-�2����vV���.�lUW_���l+�9p�9���}��9Fm�������HZZ��dlki��Z2��TX�<���d����dN�'r���x2�1�c5>S�$Jh�ofh$-���[eWR�Gl�S��~�q�dд]�t� iI�`�96Ū[C��������]ab�v����[�y~�l�֭� 0>ҴmH��H:�,$��ћ��/�P|�w���Q��k)��V7�N5�tu��d�`l����w^�Z$�������#�a ���Ǳ�Aɇ'v��dq���3/	Q�&����+!r' q�<�� �
��Wy��XU�WNډ���C3�ޥ����H�Q/[��������9B΢�`���)ɭ���ۧ�t�A0}�f���Y�ZV��:�+d�hVYe�y;y�I�,(�$��F:�Ϫ��c��8K�Օ��˘�4�b��"ƤUb��Y���oBWscV�x�}`x�=�$(�#�"�Ե	�!^�)*��Rv��)��*Ѻ	b��S��nS$�]��S��}��."5�y,%�2B���D��B��#�1�0�������g����
z�� TF S���f`ӣ���l\�=<7g,h�%s��X����1�5{24�)�&������OG]$�-l,�����J��������]wR{�Σ6z���.��nB=��V\�����У��q��%��(pLj�lL�9y�i��6��5�u)5��A_���Y��@4g�9O�rr4��v�t�.�d~ˎ2��x<�}SF����	E<��`��כ�Wj��|��Gz�g��V�K�a���E�{�Nߓ�Յ��YS5��?��M��l{2��dH����ǴW�<���U�f�G�>�f'u �I`�1��a]�f�՞��,(���׾��k��sK����бbZ������r'0��a�X����
0| U�L�(Wp?` 0f���f����^fQz"ƭ�H7��)v�*�1W[t$�7ik�S!xĸ�nG��`�J���g4hI�x�|�}��O�ĂI�i,M�܋��>���������s���:��1R;tI�~e!}��h�j�XY�f;u�B���ug�b8|#�յ���/t~����j���\�\�P�Lɡ�}L+�eV����\��P�5d���%biL�WUza�	�|[Z	;��>\���V'�ç�3��"�}� #���C��&���F9;;�>�&�r�3fF�:8���U�繂?�(���,#������G�4a�Ĵ��"lT������3wƶ{hN�A������ )Z��Tr�r	�Hc�� ��h>�I}V�؂Ք�2f=A,;�>L��V�ڧI h�݈Uf�q��Ap�^[k��龰qYAE ��W�=����i��k�v�S�n���}��{�<Ӓ�7�����@�t��uY*t�3cQ��Ӎ�G�S�(��i8���	To�
՚��������Vt�Ƿ��$҆�Zi�7�f0�3���Hm��O5��f�e�HA�T�K]�6A� �������6q �7����U�q��L���B�O�<����䄽���VQV`�0]1ֽ@��E<4����6�7Y��Y{ ���2�a��d�'q��r~<f �m�`o���+������F����|���r|rf@7X:,��q��heU�����b���c&#��ޫѠ'/.��9^xK˛�H�S����vG˵,�s��_�c���[�e��yf���ѰO�sdۣ�,��f܇��f�Y�"��vi�n�VI�۪�鵺�(�������~���+��pۯ�<��� l��R*�[)�sW܃J*o��B(_�l�7Ǧ/]a��1fL�0b����آAD���!vw쁼��+�%�Q�˵e�P��ϵ�3�Ǥ��[�gO�Y��e�b^��+��lS��dG���'�����؎����+bi|����3�J����C��3�/_�>	�^��Ӹ�n0ؚԵ��Z�J�!��}�%���mwҗ����{e�K��f����h��߼������Qe#�4J�j�Ķ|�U9�8+E[_@[��גqcD:0y���F�\,*?��6�[?lryb/9�G�����eHo@��~��\����I�7��d�G&�2m��Hoi�4p'm����i��W���Fl�~`�G�&���ҹ�����Sٴ=�n�ugl���"=��#����M/�&Lܼ3�����=���ڻ4��ր�� �װ���V#�j�"c��ZT�f���:`ȁG���=��& ܌��p@> u�4W��.��m���8�|M�vL��Ls{�!K[{W�hc0UV��5bH�A[���K�Y���B�5��Cu�V���
4�d�X�� Csh���|6��ٓ�`륒�<�=g��t?���V�k���z1�uJf���h��H����}�#�*#5��:DW�Rz�5�[UR�>��W.�GC� �|���+���"X[��j �R�aG���zX� N� �0�yi�э���D�Ǥ't�pva��g�3�OU��O'�����f�%��d� c�'��6K���9G ��m)0BЇ>����<,3��i�u���27\.ٶh&�n��@{�/^<�����tH�v2>�g����W�N���[s���= ��u��ߺ�.�fV�y
24�{4|-�ۆ5f6߰f5Nf��|��+�@�M�}j��]�}�w�������d;���.��b����X�O�������������gub
l-�ڛ:���t�Y���$�F*z#�WL�!��pDI���L�&:6��_��FP �XU�D
�6�>�;�ٜ��l�۞�����Iؽ���3ưW��E��"4$Xn�����vǱwIF�F�8	P��X�x ��l:L�-�w���^���i����P!�@+INMO6���L���7�[b��u�q쀯��U����W�ܝ~�����)�9�I#�T�ic[%ѣ���N�TP���C�nU?0J+wb��~ѳ��#��U�X��CW�QHl�ޚz����'���V�H$X�Z���Փ1�ɞp�hD����=K���ژ��F�j�u�C�Ǽ��uh���2q�;Ӌ���Q%����d��|m�Y�LZ�������yg��P���V��D��?O�w�.05MC��\��
��f�n*��43n�l`T^��E�zh"����)ڛ�]�L'}�4��.�ct{GiE�	�e��`:sc������16n|�-2��+XqG#�X�Yb�*�:�!Ŵz���,G+��kY���z>�Q`�6����|4��O���TN��u��ʡ��-K��������߿_;Z�[ �bLaC�Xِ��W`t-�7LiLzd��Fp2�Y9����!+r�ۨ a+��>>�����k�#ax�L4���+[<m��?���M�߿'�;;=�R7��鑜g�e���<�ײD��7d�+ث
dDNO����L^<����4�l��X�i���le�)�r��N?n�������[ts��k�[���;��z�t�?`A@�Lotl�=/s�7�.m�V��'�)pM�������R׫���4� k�cu�5�Z�Y TzTR���ɻ�W���7���d�Z�ʠ�<�z�`��jg��3�I�'�.)�KD�$��f�v@L���/�X�f�? �DZ���R��{��C���@X���G�����K��Qj4�����$@g�3��Nxdޙմ0ߝ�tN�tL�iS��]^t�Z/�,@�}|4����F���Ky��RǺ�����ǰBT����t��fk�p}#?��������6�:LtWy`˼��`��L~�n1��o%���}(��b>7{���l�֧��k�I�Z�y`�C[T�3�Cv+�w7��WH)���+mv�B$�L��4�v9��i=�Ԥ��~'|�L-Wսi��{�r�e�|�RʸEg��L&�3᱕��8u�� ��Uԏ�����M��=Em)6�����J�j�)��a{sT�3��u"n"��vej������S_3|�h�Ɨ>����k��	(�j#�1�K  
��AkY�Bv��5�b�o��U ���{���mũ� :O��3`i�'�����!6��X�&]�IՒ�NS��}l�������7��<�y���˼�����'�l�b��M�w�)X�]���V!��,c��\���褎O=Ҫ������ؘ�~�ژй2pK��:<0_���`feE�V�[��h�����fi+9:���]VmF�z?�:��Grr4�W�.�˗�
��ɳ�3`'��݀�f.�)Ѕ�݇��r�v�=ث��TY�¯��AT��( ���b��ê)/���7_����/��G�D�`S	�SI05�<�=����@AX_��pt:���cn*݌���潬g�,(���yR�5W��2�1�[+gL�H�t:��}y�\�P�uy~��t�����L�@v3�)at�_�����=���kG��`�̞@y��7�K��1S��>����@���=͘~�-�c��'��S����r4�P�@ �����:�g��g��ܗ�#nH��YA������#�=��^�k��Ҵ��X�!	i����g����o0��@T]��;�i�}�סWb���}�o?���?�C��4�h��{�7#6�r����.h+k���ox� I`n��F�}�X_Ο=����z�J.u���CG0������=j����J�~�b6�`m��Z��g�����AEq�"1H1�vmPGg�:w��7��w�ϼ>��]z&1�|a����iQ���iqE��=�KK�J�O�
i��X����8�9B�j�8vx+�6}���?[y�{��N����-���.t�O���^�ȭ�� ���Y�'F3.tp�������t��D}�͉���|4��N7��=#Q����&؅U��s���aa��a鯥d��!X�DY"���?4-KN����'Y΍"g�@�{�-uC��zt�G�i����Z&�w�� ��ـ�"5Z0C���z��0���b�|H�:ah��GN:�W��.,�n�M�S�N�T�g �[hd֤�:�&1|�Z�?����3��>7`����MHR0��)'�L�	k|��6�� Hz��+������z��4�RF%#�hE�t�SLz7�wp��]���~>rx�"�VE�=sc��a7�+J� S�nK�F��b�ۀQ�ecHI�����D�Aϳ���J�	øF�"�g���ͫ/����|�*!�o�7Ҧr ��b)�c�/���c����
�9� ��K��,�w� Ṿ׷_>�9"����K���I��w�`hov|T���X�_�*;W��^Aߜ׊E��@b3�������V˛�p9{�9�(����W�����Fr�Ꙟ߹|��rv|,�ހ�x���֌��.�1���p�G���u+(�gzw�tkW�u"ۍ�):i ���Y�k R����;�1��w��4�u,����ϋ9�{z~z�Jţ1�׀��UNڽ4�cI�5˭"U�Ѐ�ȓ��>\Ƀ>C�Q��Ctς�Hٷr��<K?2��LZ��H����
�1XJ��׈�������k������k_/�9��^- ����eɧ0x{3��ܧ/��0����Bpn��J.t,��N�>�I<��s�LF$8>K�3�b�`�v1gE�T�E3���ul<>>*�[p���MVg������܊����~��;b��I�(v���_G��`?�j��T�f�J��\Ϡ A`��P���J����]�h�H*v}�I:��;�N�#U]�ͤ�q�f�e��"z����>nVp�F��)m¡}{'1�S�Rk��B���5u"*��U�U��X�E����K?���r���z��ئ�4���=p��G}TV��
�����㓂�9�-�����Z�A;t�@�U�0��*-u�A(t E,�G���LF�)-#08�������@m��}�ⷦ~H��r"�}��w}l�}=R �H��ƣ�\�&{������)��(WW3yZx��uTI�����{&k�����^�1�(%���B� �����.:�$��ڕ4�BѦ1u����i�	�鰐c��!D�����U��r��f���8���sM���m$���Va����s�Uĭ��6ǆ�.J��Z��r?���:(�?*X�[����`��CD�$[O��>�R��
vX�d%�>l�f.O_S�K"�"��!�`,�Ntv,_<?W �B~��Wr~vҸ��1-�����
^R���7����	�
y|x��"����L��/.N	�c̿�(��hBAp���Y:�a��`=�(����h��cfL����-����ʌb3k�jVΒ��%AE����!�?��٩\^����1�-�]�U�2� 4���!]���7.��t�������!�ϗt͹l��-Xw�R�Ŷ�3�x+K�pm4����:;9#}��B��t,G�~���L�}����R�f�c^�	�.w`�Pxas/�=��2����S>c�:��"X�u|`��p{�qw~�c�P%⾏��D�����&��;���S�OUR�4W����ixuӕ�R�	�8\m$簤��3S���H#U����{���ӽ���U��;��;/2<y�����(E��$R��3�-�μ�7�Z��:v���j��4�tM�8NvV�wta������=�հ�	��|)��$�������f3�&ޘ� �X,���t��t>i�u�`�j�0�!����C�8v!���h�C�R�GQ{'�oN%�x�=�6�   �����P�y��ڹ��}<�S� ����q�(�}����#ոZ>�G�Mds��u}{#7�wL!�!�^�@@x�4�	��fzv6����as:�Ǜ�������������FK0 �W�c���iD�����,3?�hb��d��������'���?�"jztL���ޚq�ۿ���B��[Rt��&�.����5��tzL p��!�ԍ��t*���?ɷ��FNt�O���Fz_������ӛ;yXV�!�c~���ݘ}̤4X������� "ֱ��C�8g�ٳt<���B(>a ���^Ǐ�XT��( ������/hL��+�Uñ!J�|b�����LƯ�f�J=0�d=\�g"Nی�ъ��2>'�����������e=�*�r�A�
���Ӈ��+��� �m�\x+�|&P�F�B��5@s�-��F
B������x&���|���d�g����i�خ<\�D��(���B��BA�D�諗�)��=B�����"@99=��^Bsrj�~L�QP���!]R�R_j��`� 4gR�O�<�"��x��StW��4v�y��0?1�
(��G2�~�
�� �(=/���5��YD�|V����	{�*���*�E�F��������暕a[�4hr൤�]?��y&ձ+cLQ�FMXn���3=������|�J�]q�aׅ�Ll9vJ�J��eF&��x�M�f)*�?��>k��wb�J9�Ֆ���C���CH_��X�6}(;M���{��Zp���?k߾��7]Ʃ�':�f_���R�KuH,����n4i��L��4�X�W�u��-���� �QYyZ6��P��H�,�A�Hb�R�\���+ ��1F�|*g�4B�r\n����{-��3y�i �2Õ,r?'� l�{Ƈ�{9;{�a�heE3tO5�$<8�c��]p��i�X��<t~��t)X�qF+�zK[ �r�"S���($�yKf��wz�|��7~�wى:�U���e�>A�}Ą9��=����ى�kE��J)v107Ԩ.c���r�`a��5)�4Ԥàu� :Xl�X��}��!=111uL
T�W��}�ԍ���psê'c�z�֣����X�f_�g�e,_������nZgt�~����Tl��|-�EdE"y�%�N�gC���clW}>\�i�驥�Py�}ۧ`�D7��y%�������8q��(~z��<�Y�βx���nHF����2=W6��m-��@+r������* ;;?��F�h�:�ʛ�Pg2_W���u��FN�ҙ�����}�H���6 ؍xv�[���mO:��ck'�"���樖�e�~�(�h �|q��|Nݵ5@�r���W���ƞD�~���ml���Ѹ�/��u�1z;+S�!������Ɉ����w�qʬ�L�q�	��Ę����Su� ^Tѹ~#=
L�4���ՀX�P��F�O��\�M��߾Ԡ�9uW�b�l�WhH�!���x~}�7��p��>��U�g}
gOs2ZO���NNLO� �UʬN���\.V�<1���F���lvV���^1�3@Zt����sj\ ��x����1�[ ��cT��\s.a+�h� �'7��xnM����o۫y�A�x�.��#�����!��Z/d�s�A���[�3?� U��h
�1���h���8�w*�y�=� �w�}-����7_}��@Z��5K3v^��d�uBꪑ`؉c�`cn�3 D\Ҽ$��Y�ZO� ����e�&{l��v)(�����h���&������*�}J�u���2i�&�xu��Ӎ����K_w�n�|���㧶H���L��4����7TS�ؽ�H�/w�뇌�h����@ώ(��l-�8��f��+<��@�Kh��#�:Z��\��Zq]CZۖ���t�x��Z��T.u����i��Y!�
����Zvv����?���x�>��Ke���W6+c�K�'c�-IZ���]��8=~��7EϠWa�,�Df;�6�؜����k��iF�4Mue��~�ZZy�@EK?�U[�BlҀt�3��[Cc��h�Qaf	���|��:�և�h�B�.�i��� ��[Υ^���$��� f~~�V�_]�9I> ���˚w�����~L�`�E�H볣���ǅ٢��h?��, z�J����م\>;՟��-��.	d �&
��n�I3�[s8}����
)'����t�����_`��$�X���y��%���>,����EO��<>=0���}��BZN��Y��YY��jRi��7�L0�Q1�,�v:���R���v*b}S��,� ����5U�h ��[A�2��.k��!`��#�^� ���8���!�V�Ɩ���͹��<u��Y��liSu]-CJ��Vg:��Mx)?�pδ�r�쐞��{��}'���fɉ��5���P�+1wU<;q��j�Q�=��_<���������t�_ɻ��:nf�0�C����5�5�C{���)���hO�qsvzB!��-����s�S����ͧ�i6c	���j��Ȓ��q�L�)�� &�`����s�����3}���Ĝ�|��9��?��OG���#��p�Ṯ�l=�GG�O����M�������fs2h˥KԼ�d���@����5r�0�Ϧ�1��zy)��_���~{/^<�[�F��R5=����~���lA;����?͘Q0)DN�����G��ﾕώ�e��������>)h�[꽜C�����n��UZs{��΀�����	CX�
Ú@?g-ثd�h@u�vu����&��6�*{j�}��@�/�}F�{��C ���]�.�I�U�H�p�bɺ��7�! iǶ .m�dcj���g�i�2߼m�k�3v4�v|k��3c0�����V^��I�,@�QbO!��[$�^����d���_�,u~Fy|�Ql�ke��]&
�(����]g���߱*��7�5�c���ڊ��d��%>�������O[d 
)�?P�Vz�ш#�6�8)ݳ4"�r߼<W��r-�{7�I���x�i:���ޚ;#�������{������-�/�l>��"��B6I:��SJ�q1U)f�Fs�"�����*"�f1H���f#o"�=����KKQW�`�� ��jZ	���Q����Jnu -�%j�>��sȦ�R�Z;�ښ��C#8t�� Zo9�ۍ`���!=����grk���UJF˭g��/^,x�"�)7���g�c2����@� �ՠo�n�P�?q�L�X8g�"��b�����H�������mC��̪�Ě��o���"$O�֛L h��yR]`d/��U���8�W�)5_
�9y|���Ĩ��$��8��P�z����}2gt�sٵ$�&���=$f��aO��M�WJr�A�"���c����`0�ˋ#y��L7��\��ٴ��3ołEZ�ab�;Z`��dƦ��NR� �d:Q�����l*������/�����G���Ç����Q=E��&h�þ^l0P�ޥ�Y!�'�o9��:_(��n��@L�p���t�+�OOsZW�?<�+�������J3ť�����c��r4�	�?;�����<�hͬ� A��/_Q�R�C"z�Gc��-E����{ �<�~��g����rusG� su����ghR+恆ֶn�������5p�V0�sn�%c�{���V�̠ˁxY�(�洳@E% )M/ �H�����J���%��Y���`���|����鉞^+�����Bp����Z�7p�è��Tף�d"�g�D>��/	���:����87 �?|5J�z�V��3�;����%�^�Ғb������>M����K����?�|a~�B�u�O�é�1=��0g"�����P�66o�5�����5I�%�M.LJ�	{)���؆U�S�`T��>��P̗�ց��I�9Z_i�Ö�)Q�.�E�s�:�+���+�SA���v���9�w�W8��Re�ִ�h�dm��==K�R�v�3�?XG7��@"�u��L�u�"I�R��܏ DX��2`��v�؆b��F��?r����[:�A�	|�r�upQ�'Pl*�xV�YZڂ�j�r�Y�0Y'�_�%������y��D�\l�#�C�ܰ�v.�z+?��N֨������y� �t�x��7i��	ݵ\ad�(�*i���p���U"���ۨ �fۥ��HX��lױ����H����>�[�%L����:"�0�i���Q~�y�BX�zgO��Փ�UY�e@2���pvrB�1��;Ȇ� �dܗ��Zzے:&��FB���]X[�_��t�������}��N�:���Eń������%_+J}b�M�_./N���X�m�-U��d�����g���:ٮ$���Ú�)#;��_ؠ9E�-�niNۗ��9�'��/�n�s��D�9�x޳άR�Ңn���&兓���Ab�*��Hm�ܴ\��_����D������_�_��|��9]���%5%�œ|���!_3%
�rtr��X�L��Ρ����شX��C��׍�CVT����(��IǴW��庺���z-��?���v���Bd�����a�5:�� Z��O�~��F�2H������8P01R�3�.d�>�z3Y�f�����OT/��<ȿ��������<�"u��% �5�W����`����o�&l-O��cZPo����-"�M��6(}���m��T(`�e�@HyӛP	����U�ޫ��� �ǇG=�����^(�7W{0���]l����jS�ʸ��3(K��?��~��9+2�\ceX��1IS۵9$#��>��������!�j��W����b+��{큯�k�������`��1������a������6��"������בޑ�c�7h��,��3����A��¼F_a:���C�r�ә�C�[c�o#��ګ�Y�A���'���ދ�Ã�߽�%9S��-��FZF�(����h(�T_��Z�@R+��%�jb�:o�� t�2�K��z���qS���{�����޾�Y?�Rۮ��E��|Q��TJ�����(�x����ש�M;S٦�F���U�|QSU�ߩP���\^�t-�s��^���w{z���@v{�7�4��Yg�ҵ���Q��]��e�#�>J��lZ����B^�y'?��ш����%,ָ�#��"i^a�N�⚹�N�4u�;��4����uk�1V˭o�K�.�"
��8qc�\��ŉ�4Fb�*� �^5�yk��L.]��Br���&��Y(�����۠���~�,�e��,����ȼL"�#{>��9�z0�G������m!8Y�t
3��ʴ��P���4W����8�����'*;$Ƭ��<s~O�L��M�-،��e��櫵���4Ax���l$� �1�Q1�{ t�F�`\NN�>�H��f?/���g�@�(�{��)�/MT�X��]���͵�~�����i��9W;(���%�_2ewz4e�B�[��6[�����3�ф��`�a��b�`��/�� ���(tE;��F7 �o�gSn �bV��ooi��Ï?3=}��+ÀǶ�nXI�J��Y�3�[�o�k�Tp@��!{G-Gf��`�1�3�4-������\Y�bq�ޯ���+��}���'�!D�=�{:�M[����)7�������H��=S��GC� DHq�ok�m�
��(������������C���x�3s�޾�ׯ��N�$���A�U�om�&�n�c8gg���^}iZXGN�b�S4��Rt��t��;��^ӂ��Hf�@i����R��:t����~����/�_�~?�1p������c�3M��z*J)B#éiԺV��d��1� ����|(@�y��%����,T��۵��Kc���tЂ�z�歎�\�q*S�IԜ�+�^��UٓDO���w�2%�^�c����"р.%(� �5ւ����I����aQ�1���ּhZ�'�����{�s��ƈI�Z�"� ��xVM%�?��S0Rw�#�p[�H�\��R�h��+K�ʻ�m���Gb嚶x�xR֬�:�o&rtvN#K8 7�4����Ԟ"�>�D�g�v|��'��
BV�ׁ� �q��7����7��A7�2(h)��\��lt����[�XCmR���yy�%�����ȸ���܄�p�*᯴���W~Y�PW|�5�5��6�5����zRш�f�\<
����P�Q�����~|r��&̼�֮a�SkG���6I[�(��)b�}���[�c,%� �]e�(7����W�^��퀯�W���T�kȬz�g�pU҂ӯF�Ubj�Adz�#�x5�����߿��׷a��\=׌͵�� �K��(f@��̘�m����i������~���$;�nzu~`.�ӡ���1��K�߁ئ���j�G<��D�0x-=�0��X�AfՂ `�+��Cm�M �����]p,e��e�Jl�S?Y��=]gi�ϚUۈ�i���rg)]`�a��ݽ~<Ăy.��o(������9.��zyZ�� ����gK���+^���!�E�i8�T��(��O�.�뜩P�`��Vv_���8�K#z�zՔ��2v�Ґ��-�%�	��x��y v��>�1k����t����@�a�����p_�*�bE����_T�bl.W�[2�- 4���4�I�&�g�]�X���7O�������?O�>���&�c��z�뾃YJ#�4FP�.�XѺj���L�!`�>�a�����!����:�>�>WAy���h�j{ٞ�:�$0�ڸIp�}�JIL�J�QֱyN�	��=���-F&���{�c�\ż�t��l���sNm�J�4�t�Ρ����O��_����<�����2[�X�v%�-H�`����f$MO�<z"���Z�mh\� �֘�V�SFf��J[ն�+�k�C���c��H쒊Umbt�L�m֭o#��g�tMÛ/�>�ѣVW9�H6Qt�l^"�^2�uMQ�_����A�M�E�lQ�Y?E�$�\Ϣ7�QLED�B���T�;�ǫ���B>�����7˄�4�E~�1\��~��凟���|'�w����b` :����}�Z�5+M�N�.ܟ%�MpQ�>�4P���h�$�k�*7y�nft4<��q�kk]��}���i(l � �`��	гH�.�D;�0L8V����燴%&��.X
m�����ca�Aϲ�X��TWG�G0�[��"������C������Z;���m#a~��u��mt����vG��\���Pb��LA՜��`G� l��T��
�N\'�
o޼��zG��D�.w�����3�h��R7u�Q܁1K�Tx̡U���A?�1(Z|@�]tdN�r�M�_��q�%ǝE]����Iw�xx�(z�9�E�)4d�*�i0M�tX�*�\�������5��8b�2��3R0yҳ
��4C*#7�:��d���"�d�R���Y3x�M���s��7V�G}_f�D�i<T~rt߳-��Z�?���9�:���m�1eX���`)�mI����?6�a���ζ6�
L;8ܡ?C�'��+���%���]�@p��d�Ц�p���EE�2�|��@Զ��\v`��u�Mu�����~�ػ�p7��R���Kl�2u�[L�^�l��	q�{\s�M/Y�-sW��4#�Xv�CM����I`���I��>���,�!�j��^�q�~�װ\���_�7��s@`�N:)i��t7���I���Ys\<w����9n1VйbM-p�ӳS9ӏ�x��}0`�g��L�®*�n������N�:���c����x2��c���x�Eo+���!�sc��_\H@��x*�ф�Q	��Eb{n�j�A����~d�@@P_ν6z�kщ8�4�sb��~J�w���V��7g�@"�j�1p�� ad�K΋^��[���/ "���&�yE椶���`lʍ)b�3�pn=�(�A�Ҧ}2� *K��h`%�0�2�n��$�RhM�cm�X���>q�B`S����@C�=�X��f�$e|SNa���G���7�ۏo�i�ש�I(�z�c���:�ɄA����Z�9o�.p��\��y�� #@ܿ� ��A�ɪQnZݾ͸��W�(I��upG�K�^7h������|T[ �)K�BY�1�BщR?�l��f���H^�s�0y�l~[��``"�T�c<7wY�&�\3c4(�������h-8���#�j�]N��Zg�k�k�(Pw�:�h6(˚h��HyFv/�pN�়�-��B?*�߱) /���c����|U���S�PF?��M&=173����ez� ��Q����\3B���+4�E��,!�k�Hܲ�3Z��X�%�GO���6���U^��	���"Xf�1��2����:��|�W��5��zc������?n��������|��o��Oɮ���3Ʋrs}%�٭�g�0n X�Ig�N�+��6��cu`ύ�7kL�xFkT^��"_ަsi`1��)+\n#]�����8�k�5��И|b���h8�4�3���+������~���5v)E�y�Vw��*�u��h̛sh6
�rn��h��F�	�c�2��`���:P�_�p��=D� +4@�l��5��kR�W׷rssOF�X��:e@�*IL�J����}n�Q�/��T��
�+m*�=�5o1�S��7l��*F_��ZR�^zG����^<Ѭ1�Ҳ_{|}N������|�X�b��A�!�׏��æ}JWv���55�YZ���z�/���D{%=ؗ�f�O�밂�ڏ������o��ﾑ)�O��$z�n�i��>�1\�Z��4�G?��ݭl�%] `��?���H?��7y��'ZUP������;m�ȸ}�5�����!�źEY����eű��!�l����/H��c���k2K#�j��6 X$x�@l���\vC�Q�/^��T9��0� ^�Z*�(�n1��6#U�`6�\��eyCf��U�7f�|�9XT��X���Kc2������f�'�3m���j4v%�*���>bV!�^-��]<͑�1��47f�����.�ְб
�"����i%?�������凟o�Z��z�* �@sNi�&
VAqn�&�Bo�'�4��K��n��ײXΉ�=6��P�>��ܫ�)ٌ�bVq��&e��J�n���B2|�D�ٷ�8�"Pl�,�o����7}g���C�f��L�3F��K��a`\��0�q�u�hag�>�MHo^^v찷�4C��|u�6]W^c3��2��+w�&l���N_:V(Fg�<�q�`I1�mfV	miW�{�TT���T�>�L�����m�h[ɓn��͖�
����l�x��W�ZM3�6+���g�L���gHKCl�h�M}����>Z_h����ġ#����Uy�Z�ta�q�湾(a��9����s�櫗r|tn�?^��Xe�W�s{,�ŝ<T���;#mJ%�EN���y8@aBV;(6q��G��(g�D6)@0�^�6' "�U�7 ����##`CvK�V�㡋̓�*ۺ-7d�r��ܫذ�(X��hЧ�F�ͥLȚ'F��8����딦�ڞ������ߓ���x� $�Իm�gV�A  �v�6�\w�LZ�۬L#T0�ȼX�ұ� ��0&f���N��z�����#���Z��ǐ��,->�C���H80��LM���@��W����?��R���Jk�G_�f����Yf~��+��l��ƚ�l�䕹:�����(Zp%������]�^Z�*�'G4�'�V[V�4h��[�Y��䛯_�r?�Z�򌙮�+�M�|й�=h4��~	5�}�8NBY�6+��T3��
Y�Mk2$e��Bd���1k�>�$p�f�e�[��w����!d�[ڱ��)3��?�J�W�q�^ڱ�:=:���b�*��K(К#�@���A�g m��Mq�F����$$���m;�2�ظ���33V�D$h�|�t��t=.��3E�6�up�-�\���i�,n2{8�Ji��������?���W0&�Dr\`��lH 6��=�� _XLR�n�ۈ�F�`���eT�*�;[5�Yy��42]s�!��$ӣz�<�ߙ�73�8� �E���� ��h�R��aԠE�n{`}5-*�U֕/�� <q��՚)~@�1/hgD�Eɨ�@�9@�ɍ-3�5�(8-%Gt�����òQ��a1z4���)*�<���/W_��oS	�9�D�}�ʁ�V����8�9��pO�W'>ؠm@)}n��93��+��X���n�9��#��V���c���]�N��9�|0nouCDsw릷3�AI#�-L�v �m6�׺�Uݹ9E��fɈ�PP�j�zk˩�<6��d@�	��N�z �.��pn�>颊��2u���ݧ����mN`�0�����2��= <���^���uNnhb:� ��m��[�cHi ����e0��,�؟��`��0%�Up�1�A�x�1U�n�`}5ǰy��Cի�W>dLu�n..��K�(RU�~)��ާk
��XM�6?��<.t����(XeE�z�X�]]���������8a���! -�=�c!�ϑ̭Mp�=8��2S��k'�SD�`�,��k�X6�Px�M8VGk�4Esn8���>���<��}`pFmKH ��U�K������}/�7�ƚ8��1���;lN
 $��n4��eƮ��Sb�C�O�ާ�\��������)�j���g����c;3XG�mf��E]���~9�?9>�:O?0}!����� b�޽�8c���-�z��d
u�x?T�[�-	dz���L������{Tp�^b�"�����oo����򕮥z g�k<2���,���)��0��`�}����ڎ6��w���e�Rp�T�6vX]+�(��X��7�6m�J�Xద�
�yaB�%��Р ��Ԡ	��#k�6��}��Z�^�FG������$�n~O�R��`�����LT��֏j�R ���g�l�>�
�Q�&ɹ�63�p0�R��֊��^i ��{�՛w��׿�(�፼�~�:I�GzL ��G�`��L7�MU�[�Q��HSY
o8a��:��Hs����x�s�����6���s2���͗���i,�)~��+9^���w�X������|��'g�6[~��.02�8҉F@�5�>Q�Pyj�}�E��VӰ�~��q�Jl��<cXbAgO'6?I`�YN[z&��5Գ�1H#o�^�o�Ф��:N�4�����c��h����j] 董�>��h�go2`L��ٚ6����x�,��Eʀ����2]�H��!L;9��c$S��#�I�LU}�'6P�CWs.���4�*�=�.vև������SЫ��|=?o|_�=n5�/�QL����y�� l(�⽶,�ؖH�>��݈��K��c���L;�y�������;�WR�QG2G�7�L��{�}c�Q_e��+��I�x��`�,=W��&�G>�X�K}f���y*>R���u	�a��k�\�)�0�&�]��G�T�����tv�m�o�,��
��@@hcNώ^�͇���O�{��|�v&�'�d�!�/k(Q��e�Ҏ���+�w���\82k��[���� �<�#��EFݫ�T<�V=K�, ��z�B�SL������} ��u�����fh�Mߝ��|�MZ/�������J7�cӟz�e�Z� ��v�[���� ��{�_��b���J?~��)�ءs邸�hţe	d�kn�3`�����[���w��B�=q��'W��t��{ ®���^\n��>��б^��bVV�c��`�������=#��B���>�|����u�����6�-�n��h08֯�\(h;B��^�L"*�+(X�6k��:Y|7�jĭ�-�3]ݴ�ݼ�b��:/�g*�w�MK�`Ȯ�ʊt�
�@t��ߌ:̻�G�K��gR���d���V����g�$��.�Ck��d����	i 4��p�����ˢ�/D�3���""��W�V_�F�b��I��l7����6k�́:UG�2�Vo?������*��\��|ôc��K��F����|��`�#g�;�K�{l�vb��)�>�`P( 8:;���F��mz`d��13ɑ��j'�_���iʯ�>������.�+�o����7�h/i�&۬0�h�)G0��%�
vp�ɋg���7��~������������00 �B�R��b�M
3�����ф��֙��,�F�!؆dƣF�g�
ΫS[��6�X���΢��؄���)H�rK���M,�
��E#y�����?Q�W� �w�����N�*Y�+S�h����u)��A���C�|%�
���� ϟ�^#�s9��F�����1޷8aԇVz�����j�������1ǰ��#�P��$���lsݬ�����GY�8�|���(�#0R�DFc��\M'hw�gza]<�Pn�8�^�2���H�?�޴9�$����߼g�ut��֊�~؝���?`E�{����ʬ�8��M:��f��� �#�{d7JXI:���T�����]�	����ޡ�|��C����%�Qv�t���Vz�%�]���Vϣ>��{v [V]����eA�H9�н�8�'�������Ȫo��M�իSfhVI��4���'���B~~�A~ֳ�y踾 ������4��9[���_�)X��؏)Y�"�3h���V�ľ@'$-Nt����a�(�/2cw7���[�9pZ*t��>k�=����C��x~9v�&>G�m�AHP���&�E��
�V����ֈ)�<N}�9'����$��`�L;��9������S�Sk5X���\�5M������7��� ��ݖV66ӓ�b�{4�ܾ\��C}�@f���������w&��;�1�iu��);�ɀ�{�/�)�R��������;#k�F��Ȝ���(������B\�k�m-ߓ�S��c�'�[�#�./.�??�ȳ����p|�|q,{�����a�Y�=;��F�)*�1��37ﯺ����������t�R��v���I����ʻw���������ՑTG+&g�:�n���tnmZF�M{�Ԝ�'�D׾ӓj�}�{���%�e�,@�&�l�N{�]<��[kBR,�&����KJ�<�3�(ͭ	�Qץ��6BQ�>�u>�Դ-�4UtM�:v�R�VJ!N���H.����%��n-�Xb��H�J�L��*"B�օ�Ǒ�xk]����խ|8�����A~��\ܪ���+Wt;'�'�\q�4~L+�c��e��x_�v-�o��M�lsp0�p�H�r6 u�Z�s@Riv�K̼@��C{�>��:�Z����H��߳�18����3[�dXIrG�i�+:
S'��FЄM,��iY�a�N�"��k��
�6.��(٬�s�J˵wC�Ͳ1�]��o�1tRZ�#�(��q2٦�eO%S��"���M�O������Y�:���L4��n=���2&��.��IE`ղ��R��S��b�2(�m��z�>����9��~w����0nB���?p/.�B~Po�$�X6N�çKV1��a}��.m���^�����lcz��Z�0xD��E�ٗ(�^�\��85]��y��P8q��ް������������͍�ݎ���OS0��P��a�ǵd�k�P�~
 ��aD��AY��0�k�BTy�����=aOràh����z���j%�z��ܤH����f3m8s�s�Q�"Y H`O�F�2��"�ɑ�b�,��Sc_�������'�wǬ�5(�l]��Y">�F: �R#0�3ܢ�X5gW6���E�9�Q&୳mğ!���]0�m/���&��@8]6`�&��J�v%P򾺑����B	���s0;#���(���4�������+d��@�x�R����`����dүd��<�b��C~^���b|y�����[�ɡ`�Kl|���x�b��r��7v��I�=9a���Kt�Oc��	{`�w[��hA�B���&,^[����\r���l>����ѭ�tOA�7�?h@����#��5�2�{�������)���[�=�WYm�)Zs���t�\KI�*���E��4ϺACL���w.�q��|�T�:d����g�r�|�t���L�,��_k���D��ř�h�󴾧�*EU�*��u@Q3�0B�+'���������7WG����?��,�_)�p�І����6tjgTU�{&E��U���md�Mk�ǃw�ǉ��g�/姿���ߟ��Ory��!Ҝ�6�%#�x\�t�Oͯz���f>�5�yd �/2h��!�%AHmZ9 4���L-�2`��h_o,�mF�r�א��\�x?��^�|E����)���$������c�.x#��2W��..|���g�_\���\������@f7�ө��b3Z��'�b�RB	ød;�C��A�bb~��ljc ��/��w�v�k!����iREY:2��׍�Gz�p�_�'�$��y����Vv�]����nV�*І���W�����]��Ɯ\��G��EWQ]��.T׽\]|��͖�>t�^]^Pc���L�U��ҳ���o\� ����]��lfA�r�Pۦ��&�ֽ颋C���%�h���*�CZ:�c�����QV��(�a����Z�x/7Z�kZ͠�RNO_���-��0��C����H��
_Wj8��A��AY6�o����C(Vruu�n�f=�b'�7Jp�\�����%SĿȴ�=��(_����dCAϴ��}��������?78F��C���Z4��{�M-�;�n�2�}^��3�l٭Ͼ�1a� �www\��]O������%�C�?�}��z{�0����ۗJ��SW˶��|��W{��0��̎4���l|�W��m'���Q�b�&@*��T�n�����!�����?��7ݯ�smѥ��g{���A�+ų�\�* ̾��á�?���yy� l���\�ɗ&�� [��9\ϊ�~��Q����-��}�s�7���_�$�D�����tsM�1c��o�|u�l� Ӵ�~�3���y����	����})�^�b@��#��-�c2�4�Ԝ��� I��>J���N���@�^�#SX���@�_3��Q>~�$G{39=��������B�z>w<a���芮��l6��$��P2�/ɢ�_�{	1�_��"E�J�dW2��g�X?QBg�ϛ/[�HIA�_t6��6h�ި�z��1�2���m�tf�� Ktʦ�G�I��D�r�`�r�îT���K�C#�ñ��p�+X�U��݀ړG��R{����lG�h2<������ry� �
�r��Ԅ ����Ժ��B�s��]�{V.��AC|��!��1!�n%����� #q�!��p8�>�� �Ĵ%�\�	�tv��|���6"����V$u����"���yD8NjF���?��=<2k��z2�1Q⼼����k�-�����:�=c9덵�G��5� 3�ED:�s�";p(��*Xw֦�!�)uaTܐ:�p �]#WȄ|a�3n>�X�E�[��5K>���	KK���h�{};`��lQ��Ǐ,��8� �5A�I��ނj��_�b�IF��jҎ�hz7�8B���є��*O!�f�������L������<m�FV�'3�����y%���Ɓ�$&*Xc�F��2=�hM��3L��~8��e�+����hc�;J�W7��pwK�|�0 J���}��~�x�i/3�C����O����8��YZ�>���v��.n�:��O�5fJ6~.��W3�?�`����l�刮Y�`�Z9 0i�ֳ�/f]d��E�0��vq����;��c�-��ڶ4����#�V{4�ؿ�5�x�=�pKE�FR��!�fe��ݕ8PE�bR>��C��mdC���u;����*2��+��u�|ڞ�8	��Ec��
{'2�8��$�|P����$;��<:Ҽ.��?���g"�jLa��pK1I#��5N� ���u�q?ջ�,���"R���b��JL�z�y8��N㦁�o9˨e�_�gU��d3mj��*�Ũ�������4��b�F4P��@or�(X	�1_6�4�P�e��|8����#�GlHe���O��w��޸8�u����y��6Q[�|�����G�Yo��nRO��5g%S�N�r�-HJϞ�=��t��Z���^>�3~Z�Ӓ0��QZ��'�Gm����h���	(��A����p^���<���Н�"��=���4%)�ƽ��Ew���&��,��,(��^�❛�Z�rR{�1JB}6�}�EU{���Z}�����Y�T�����;}pP�V��[�g�\9M��bJeG �����h���~x(i0���>m{?�3@��Yh蔚( ���Y0T���/Z}���S:��|1�w��Ã�i���V�Ł0�ŧK�ޟ����]4�a����׷alj�g��<(en7&��_��b�:�5f��.��Iؐ����K���b��D����ϱ ��JN���	��ۼa�3�H
��P������Gg(�.L7%����1C�j�
�jyITf�����w�r;�E��S�A�M�f�n�*�7�B%�;��Z.���7o�p���į�_s_�Hf�i��r�{��R���=�'4�P`X������6I�F�bڸc�Yj���I�쐋�G	/���C�Jw���u� WA2��g�5t��+�V}�X#tv�Ė|O�ؽ�0��=n�����iK�(���?P�F�d����u��6H����0��(л��3����U�;+���(����|Hc�,����I�͆ F�W��r�ױ"�2���-m+���g��;�	�g�IX�O�Yk~��y|lY�@V�/p4Ƞ�*|+���X���+��K!���A���e�x�v����H\�W�:P��d�~6]�s�P��u"����Q}c����]�,Ye�m)3[|j�q�Y`���z_�z-Vs�7�.>��۰s����|\
ff{Od\`$����O*c����2�[`�f������_�0��Up�$[uC7VN-�U	��J�@�3��Adg5�sY�~ �����V�9�O6�9��n5�@*�0*�u2�9�J'v<�Γ�d�Zf��r���q�M�Ѿ"�Ğ0`+3G�A�Mi��+�	��빂�1��D����P7 �>��Y�bT�6�sE�}F���?�4'*cW��}�E�{�j�){b���\4z �"΁-�b�2�l�<���Lc��Wb��6=�D�=mF-����,â�'ц�d
{�m�`���Р\�`T���o�4����L/�5z|�L&�,��h�K��7md�:�،��G��h]nK����4r'�ۈ'zf+�< �;6	P22@7�䮮��^���u�/a0r�<DU1K��k��Y% S�U)0A��ZY}DƋꍃ��䀚�eJ彾{P�z$��ו�X�j�����c�zqʲ"���Xk�>Q��LW�;.�6 7�/���9&#%�qww�����:��sQx�՝�=>���[[;�L�<Q�cv|�'�S�t@�����t��&9<>b֠ser�y��3/u}��R�%-5� Ѓ�J _���+<��C9R�2o��`�?!0�b����l.[z�y��\�5���|*�DU^Idks������ze���D1._]R�ɻ^b_'
�z��)
���L����[p-�5J%����B���K� E�]�i�,���2~��yS+q^�D,�gnXRd�9��?���(��\UR$�¹�r���}L{����rA�`<��B�� ��SE�8$.�0@�	�����Xd����:�Ѵ��`���l�u�t s��R���{J��y���g��n�O3) d��]�V�1�@V�-����~�⡭�r�z���6.���ͦm]��
�����}]���SCN&��ѐ�ܵE��ߟ���Z�#�)(�QS	��ʉj,�Wb9���W������B	c�z_[�!\ݘ���9�<GPtI�=&�ףy����*~�X&� ˷Y3��`�4W�dUS��t~_سp�U�g ?�����.�M;6[�w|�2@eȓ$o�3�e�2�X�ShN9:�B����o���w��|�g�����8��h=
�J��?y �_ˮ23%��+��u/��>�a�sSY%g�<O�?����u�!���L<@ܜY/K�`o�:�um;ʦ�� 4�h-h� � �-Xg>��{d缿����֒6ȞB�)�xi��q�j��	J%�a�q��_�U�͚���ΐ�5 V�<y�3��K�g)#p�Pρ;�LYIȅ;l���	&�ؘ�X�C@���.����O�uo��X�Z�u����=�
�v�����Z���L��?7`mj��(�`���=�ͅ;�Q����+���պnXdK�5kF�v�o(�RcU��E�k�o��+֚����5�3�U��@����7u���8ܨ�1ː������|:���o^�����Vx�;�����~�h��Z�g�7�����/�<�C�1���gF��~t�_ɇ��3�R�>���; ��Ս�z�F^�yKeuf����iG�_U�JG����͑	`vYs����/XJ@v��~-���䧏r���ig]�(��	����������?���s��S�̿��{9z�V�å<��|b�n&����(o�!��W&�/�%y9��CY9����ZD׺֐Z��@{�d�\��S��x4�[lk�O�N?��� s=���ތ�;�.F,6�7#��}.�j����xf>��s¦sFy��d�-Q��zsK��_dW�X�R���ceoe�ˤ`J�ƿ���\\�%tt���͖���V޼xA��������'�q8v0h;'4e�܊���Ą�6�g����棕��At~8� �[�6�
R����{u6ۓ��Cyyz��`���V0�a!�ۆkC����3�����x���о�5������{^ʚ���*Ŏٞ^\i���{�W+y�V�ro^��o�{-G�{��*��t��ٶ��Y>|:���I>�_0�j  	�S�mR�Ӧ#ײw���نi�b�x�Y��^o��h��]��Vm��͝:Í�ksn̾ѹ&��昤	�zs�B�HA�����{�5T��gtu}-�
�+ځ"K����h ��k�7۸,�}O63˹�E�vw��z��3���>X7r�"��M�%�����;aF��`ƙ�Di�?4_�,;d(C�6%*�]���P�V#��R�gR��"��/�}�"�1D�E� .>�@�:d����XXM��f��A��U�>��YIE�;�6#��ȴ�Y|H���֟��joDr��T\ s���^����-9��*Ҏ-�F���� >%��Y06�d�@-�/��� ��L�S:�Zڪ�����a� ��������B�wv{��gU�l��b�p����]�7�ȷ��+�+V�T4���P�VQ�a��+�0�h�����B�����l���v��lQ��;�}^��� �Gڟ�7���"6 f$��y��:pKe������1�l�YYl��#���У��&s��:6?�4Z�|��n�+��c�0�����n-���T	��7�R�e��}�w �}�[Y,��޲� ����C��@�䣂HfoL�c�$��\�����T3���:ɯ��%;���{y��a�U�{f�v �u*�7S��l�#�Х�X�1k��ù�]\��̓|��'�܀A�D [����\(����^�u���g�O_����R�{-SdU�bώ[+�0Q��gcH!�&����	���)�
CZ��o�$B&�>x�[/���wQ¶��FQ3��[��[,OoFF�N�O��1�i�Hh�X���b��ui+4����������	e�4�A���G�(��yA�}h|�q�7�A�E|ٗ��-d����y��F��p�����y����߄��Y��P�3UM ��pK
W�m��8��1mA�)��s1��2a�=�cF��+�mY2dM�Y��+nW�:�~�tآλl�	��Vi>�9y�{�"#v�����h%ݛ�J��UV����!�A��A���}s���[�7ֻ�G����X^�<a�wp��g8<\f�]�~��;rZP���R�į�|�$"��g���~��<) i��%�N��Y+0ZSF��s�g��8L�'g@$��e/��8ՠ!�r�@k����{���?R��t����х��Ρ�\@QGv~A�F�>��pceD�h`S�M��$�e;C�e���|�3�4���I���#%�i�������u��Pmp�DLw׍��ʥ��4㛺:�Ձbi8��%G���GCYL�L���3_�{����w�'�~Qc~��Z%)�-9I�}̚?Zt������hPCW�N}ޥ�ip��+��ۣ��Wo^�k��U\{�A�uV$X��rd��8c�Vf~���o���̖\x�? �?�~�rJELy��.9��H�����##�3�u��/�Cqr�X��1�J� �O H��Yֵ�,��̽�鶀�\�4��	���M���Wj�k��ᐞԐQ3���m��OO�F�B��r�@=�l��L��k�i��[Ě��i�J��΢7�uh��n{��䒪��_f�d��#���֜s�N?d��=����ˑ��B'7s�T��1��� �z"�p�48�>����|>{���W�3W�~מ���;9}��Y��w-��x,�zK0�bCM3;t6*Fj)�J?�!\��l��^��D;����rr|hF4[DVG�tL6�Cھ46����N���O�_�ۿ�GtR�[�` 5�|
@�bT��Q�:X��k��hO��R��ե�N�e����L�	6 ���,&G2uǓ�"�O�E-�	�Ȣ1 ׃�	�ˋ�Cy�շ��?Pg�熦���#=Sr��4e�Jπ�#~�CĞ�<m-��ܫ�����&�P�	/�Yp/�@10HL�[%+�"K�I�����͐4,Uܯ7>:9�m�@�}��w�\��ߨ�bc�_z�w3�0Ϻ�R~7��u��-�����V
��ܰF��LXzĿ�5�轁��z@\1yWKd^ʾ>g�eف�X��cKy�F�������#Jh-�0��Z��/�,��Z+%Z��x���gyr|�_{�ʅOʖ��߱~�����sN⻈B�t�/�3���N�z���g�tq�{�徲��ׂg���Y���C��o�>�3;' G��]_�u�A�)t�1+����6����V�!a�����M|:���qN$���Q��m~mN��]�=KM[}w�����W�{�|�tE���#m<�J�U����7j/~���rzth</�c��B��?�$�����{���󕕳����̠Q��qM^0�A/�"�� �xC�ǭ��2��I�t���SG��Zj�j{p���\P�WdPЭُ�|�geY	i���c��?�Ӗ	���!���l��:@�]v�z�.;�k��^%�`�@�2=�`�O��EA��(���t�ӷ\��D�<8�����e�����rd�Ý��K �vͬ#�#8��Y�޸�'i�i���Zm��<��	o����$�뺽~�J���?�����k����܅�D�I�E��Q؈�5h*��U`}���/�I�[o���//�l]ܐ�&2e�)�CP���2���~=$�f�o�1:!^.�?�� g��&K��Vm��70?��=��+f�A3�&�H�E�e��t�XMb�kH�2�VP��{Bv���e�4��(]��:JAPr��d�4)%=�uéA���� L�[�oP. �r�p �s�(�M�ly�Xՠ��9t���"�)	����b%���罗%j	�����SΟ�]8s50�w�\���XVP�� ��9�Bgr��&ƌXs.��{����j����������3	��k�m�d�%�s���&�a�n�q�w+����Vrtn!3s����j-?����?�(�w2Y��Z*;=pB���m�lz*�rȸ<�Y�CIL��w��h�l6`��- o�%�����g ﲗO�2!��^�N��i��ғ��8�5ӿ/n��\�`�)�vO�/�o���K5*;w򦟶se�����-�a>����@!���'>0��N'�N�l%:��
 �i��. ������꺟�qB&�8���,|׍��[�X�0Iɻ�|$F��?x9Y�/���qc�C9�i�Y�X7H8WdJQ��@���4�]�� ���D^���M�1
���*g�a�����)�0"=:�&
�~ 'j�4\|����-'C��I��wC��v}���w�<��][�$:=Sr���m���\��O��3�tqɬ�g�4��
�v>~$��\�f������٧sF� �W�r���_h�9���}>n��s� �أu��ڐpd����YS(��2����G�I���[��<�
qNz��*�(+b$x����f��T�.d0_�3�����Cva��q��S
p����?�E��mE�����fZ���1���c>7� :�l��.��l8�J�_}�V�����&���F����{ v�D��Z��N���.��iڴ�̄A�)P���G�ܬ�3�k�<��m�UE.��}�Kܟ1�r,2����qѷ�yŦf��������?��#�`l�e�z'Ʒ>��:�����=G�
�!��{ c����X���7P�E<Qi�P���g�&u [�I{��|��W��w���K��;�z��v��,J�,�dZ������߫O��r��ʒ��w�1�,�!���]9]P�A��	���`��.�(`j��DF �Y��Y�2|���H)C'�MO	9 zը�%�)�^&�B���ՐW�F�KzP��7h��ŀ��"��/6!��Q��@�F^_�w��
��Ƚ+boR"t)7$��%H���c?c%MO�z
и=N���1��d�Y,|?���N�̈́������=y)���]�(�J|
��@�c'��I��C��������ӿ
{�E����W��?��wj�N��!E;��.�ͺ�;S�ǵ�v����_�;��!��I#���7H��b k='�q���e23��贫��>�zb��\�����՝|�t!?��3�3��?kds~q�r���E���Ȭ��?f<�aУ �v���Q�:P����D���T�e�9C6������c��̮H�=�eI��f����
r6�<덥�1g�%�����|ˬ֭Fk+L^�qE��kk�HV��~Z.��͛��������ZJؼ�����8:y%��!`�A��gѶ���Ϻ�Oz��M�cN��S+
R�Q�왡��
��*ٯ����y�^�e���y[�RȖO��㹮����	2�N�kP.�jo6Orsw-��\Q
���F4��fWfN��tu�#��LC�V�-g�]h����j��/o�L��#���(K��_�C��/./�`_l��s�Ё�o���,��gj�z����끙G<��cȹ��'f5@8�� ����r�������y� �hz���6�q߱��ӧ�ޯ_q�e�l<d�\`72��sTAw8���Y���325�3`j7𽋛{څ�A0J���1���;�[��l��Qk?�� gh E��_��]k�W��:����-aC�1GY٥�vE3 zO�f'4F����}��C���I�ɻ>���xl9��!�I#n��H�|��������q  �G���1�4�[��"� $]G~߻w�������U��U��؇��{�$���ފt���C�<�mu�7�@��U)��-����b��ْ�0{�DJ.��Y06{T������۷o�����Y���Y+�G�A*���>��>����z��}��A��L{r�@�FW�cs� 	��k\�V;S�4  ��IDAT��H.�čS�l8�W�7���rS�c�����|L�g��i�� .8���6�_��r(+ڴ��ĚYhr�s�F��%q�k^|����ʑ>qh����Z����I���,~ϙ��.s��$�B�lk`!�&�I�o�N@~u���Ԁ�pɬ����JWq��4�e0���1��������e�����R @���yf&R����2�/�˒"{-��ߧ��6ݚH4�lElv��j\�U���������� %�e�l6R�(�6���g�U��ԸA�q���`5��I3]����2�*����Hj]"�%��g�h1��F��V�u�̑���L(�-X/�^Ûs�v��a�sC�s�~�)�>[O+8;�<>|���~>ӈ���m(��9TP��� �����-2S���P�����������98>!�F$�Bs��Xl/+Ӿ �\�o��h �(�!���T󇰫��=�m��e1@�_�(�Z�С����Y�Ƹ�]K#��!����08ƉD�1��U�t�,�d�2-ϑ5S+)� ˵��¡�-t� �x֐ݺ���.C��ь���Ip<N�����[c��ҮΒ7�Ig�g\z�o��&o�^��A���Xt�!v��� R �K�O{���<cY؝�j>+s.p��W�)�@��{��ʕ~�v�T��:g�g!��e- �������@����o`(5��hԭ�ussM"?���X�C��A
�������Z�+&�,� PRY�H��
20��"�c�D�.1K���s#w�Y�˚��5A���?2�&O����XU{��Y����ݝe��Qk�*��Tq-%�>^���@�+[f�w4�u�2��tО�i�q+w346혭Y��Q́D��i����II �E�J�<b�rU5�V��
�H��bE�'gn��&����F���� o�z��A�
wl�  ���xd���g�Q^_
���!� ��1��xF�kǆ����z���~J�q��X'p V�����Y�Dd�h���F&�Q3�9�
r�gAѯ�����=�Q�)�\p�2�](���L��W�?_�&�U�b�o��1!F`�����@���ҽQiA�jkõ�!�ӵ�������@6i�H;�c����,���
"?gL�G��A^���Y��b ���T|/����l�s��e����LA�Ϟ#2 _y#S 0V�j��Z�ҡB̲B3v���������!m���eu-ڸ3U�{v-$AD8�K�u˿#��+6���_���!cZ&K�e�|P���Q�eI��G,@�0Ĉh�&H���K��л8\��z�4�9G��E
\,{D���2Ї�޲���ͺ��v-�|ƈ��F��_���{�5�%�Q��(./���3��B�'�ә��ʞ�����`)a�zg�zt~������b5�5�����4��<���/�������Y>k��2�#��ɞ�0��\��ɣB�|�Wi'���5M�Ȏ�^�.p�`D��}���rt��D�v{�&k��$)���Ue����7�%�^I�|ʵ���d�#d"rg<a�;i�HZ�C#���D�C��D~d�66?jJ]V'@�8�|`\�:�������9 |�� ��|���� U�UG�Ӄ.,���}�W6gg�~�'�{T��L��2�'� ��%X�4��d���������.b� �xV F{�)�_K��9~�k������"8fh�-4p��5��/����|��^_�(�LDʽ�Ri����|x��c�z��{�H���C%l�2��ˠ ���,��\�W�6�~�g��\r)R�Y��.����.�u(~�8�`ɃY��]�o���PDӁ�����a�	�(@�K׋��lXr�`��_�I����ąg�jӌj< D��	D���	�6��[� �V���8!s��BZ�ٵK��+��ؙ�<��.ȌAE	����o���>��^�(��a� NЅ�F����33g��������g`�?BCQcY&ȧmY��	�VH�k1o�X���W�����r�⥂�f�p�S�5�R��+�5�����O�>��oR3 �wPj�xÌ�x���ٳ��������½�՛x����d��g��Q���]�;���S=h�Q�޺�w��(@
2J��C5�RL��F<Ѧ��b��5�����k1�d�jo��t>~��c'6?�ְb��b�\��b3�?3���o�i:Pb�ag�$�[AU�g�VG�G�䇿�U>|� ��(�p`|]�UN���$��"�Se����;����y���O�8|��^�\��$���V)��qp�R�|�,���Ff�5F\5dqM���"�n ��2�6vVf=�v�{Km#����<uO����`iP�V���"X�W|��L#�5a!�j�2��s�<��� 0��_%e�u�([�!���v����3�q�Kc��B�I���L���R��R�[���:�-9G'G���2 ָ ���[��{�e[9�-H}�� j��Ŗ<
�*�R+$� ί��M�{vR.�S�Wjt�Ր�h�L 0tI�%����B`� Bh;f�fE�U��YbP�e�H�/�W0.f�<P�����,�~�?~A�p��v�8"pw�ZD��\@y�(�㱪���#��[�G�}�%��ŁM�xY"1�, �32�q.�iA� ��lٞ�� �J=Mgّw�ޫ�������G�BϘ)Bfm�P vt�3s��Q<�;(���6�
f�n�B��1U�)����ڳ��хE�QɃ@ �#1���0����M�ٳ��]��ߣ<�k��S�Ĳ�ô�<�[2pB�@�Mh����;F������`�sc#�_\\�1��j4똤��οF6T�GL>G�����b]Q��1���kkX�X)�fd�BH��E���.�V�r�����hH�^�v���4�zv��CF.##j)$N��0b,3 "�2Y��A�${�Jܸwɍ��������]Mo���1��eV�-�}�O)�j)�Tbc�Lg� ��V%�w�S:�Ghw7Y�/?K���(�{;!� \�$1 vL�ު	t��� 3�g�C�瓣m"���G�aN.�	:��#��������%)���@�zK		�F�~r����L�7.8�ם��a�U����� r��f�{��*G
2N�SPv\ɝ﫟��RFB�� C��^����(��&{��pϳ�q?��BpD��}L�����󿼼� 2�*�v`S�,�V�Ha�~@�����҂8�ـ��T6� ��f.���)����Q�L�0���5�pWlZӞЎȚO�&�x�A^�#��\W~n�|0� �4a�+G� )�<p�y/��s@6�3g^��i���vh��m��&2;%�M@1����<��'*�7S���Z��	�[���v��Y[����HF��;���TY+t*�V6�e���n/WVΝ�J%S&nȫ�-Æ��GR��9�<,X
�W�Lʵ�i�ѿ��^�fg�GKVΥq�f��'	K���N�ν�J�X�:E�pk���i�>�A�6�ۋ!����q6��bT��3�9�Cd�(�f��&����uZp�0�hK&(�SΩ���L�6PO��ъ9h���r_�Y��b_�s] �Rʃ�#��9t�����TlĈm���6��:`��jt��#�\\��Y��gewt��` ��Q�Ӭ1���8ܼe�:��M�<7ſ����#��[+�nצ��Q55� H��k�Z�t��Z���#i�b	�l��:���/�R9�=���)�]�xWT��Yv2{��ДG28Dv�S�%��� �uZ���N��K9�_��F�b�2�dwX��y~�*�"�pO��!f�:�n :e�����(�>lk����EVn���;�Z�f�z�)[�];��D��\����Oȁz��qJK�6���k��ml����vq�Q�+U�i���s���~�&����9�EF'{@�K|�nY�����`���Δ�:�I��XU�泪�-h��$���]|B1�G��gg���t�P2��]%Hv�o׼^�i8��2�QO%#d�� ;A�ω���q^ٚ��71n�up�,]]^]�[���"���n�La�)q}��4 »������0����g^RzH<V٨�zb�+9�3 t.�K��8���<��N��83yk��_3��ӵBG5��a]|������&g�~��G�C�������ÿ��AD���|�Ohk23�����7��8ss0]mu�'�[�M�*������L�n��NX�`����H��=���Y6���ؔ�m)Y��͝�{R��Ͽ��o��w��ٖ2亢X-^�(����QC��w�W��#C1���G��$��O�{fy�+�9	I��04�D�E���Jzl��Er!�c�p�H��`XI�͍G�>�A%���M�B�傖 Sg_82��U�e�Ȱ���La�d�b�	s���|Qh�k��H>�9�2�� ��3��6�"��w��G@��p��^s�`X�$�uL�?�z�H*�D����h{��ȡ8 ,�@[gN�6
s��6>��|�6\�Sk���$ȂmzN/�m���*���0��Q��'�6�?��`�]���E����2,��ڝ{����� p*��L�b����.y�q�����es��L�x����+A��?�f�m�G������M���UMG�x~M�^�F��\hiz4G�И�Vc�����=v���z_߃�#�`�M�dB	��l�u��dC:�^f��C��$%*".?�_��������V�[f9JG^����}bG#���*�kV>7�����h��=ۆYD+��e͋z4�*vo	{�GO5�Z�+Oˇċ�Z�1�� �Y&�M�k��-�ܔJT�����`���>P� 1p��\j@0#�g��0��i��ng��pPu1佟�΄"�I�y�xhޔĉ�i���i��M��Ujs���2���x|�c��y�!�ë��-��Q;4��)������5+��Z����v̦�T\������'Q���LX�Χ�\1G�Xf � ����u��`��g���u V��v}yC�d�����qY�� ��d:`�s�$6��N��=`3ǖ����`�dj@f��Y0�s�P�E�w�D�l��/�����r����cc��i<k�{SJ�؏���e+�Ṡ��؏�dÇ1 �rt�S>�S0����'%��Ӡ=�R�ֺ�	�=pI4�����N�习+�|>/����f�1=�l�lg_2��.��b�<�Q����=��ٰ��G�;�������4%�mvG� ��e���;����@·d� ��g�8p_ˤb�+�}���6�	��%��S;�C�ㆇ�g��2�Sok�$q|�b[�D�ɋw$�w��#����q�d��<���/P.1�M������,@��(%黺�.�� �����I͋�3"s8zC����wE�@���S$�erZ��?�Q�=c(���i�,�[�(0�,6��siP��V�٢�?�0��7q�\B��S� h����T�\�:��j�nl-����G��1��{sF��%�ɉD�Wg�r�8���n�`P��e��F�⨳�� ؖ�lD׏��w�z=g�ݦ n,/v6��.`��X��|aDb��;[Rߕ�Q^W�3�~2��T�Q:�2�,"LJ,`�Cf>�zQ ��0&�(��mIp#��
�I?Cܙ}h%/�ۯR��'>�g�ؘ�� YN���<M\he�?p-�Qc��y6�x7�>���=11`ξ5s�� >���<����Im{��iphV�g�����_R�b�()��C�x���R�v�X������{{r|x ��G�laZ�m���=pВ���9;�	l��0qQ��X<��sg{�3�֟��'?'_���C橞z0N�WB2� �a͑��⾯}ZDo�*-��
*'�F���c3� ��X:��MGG��2���#��#{�6a"����Z�!�AS<��x<�ΞT��4X���b9�ݻ�2C�l-p6�j��g������	�=[U{g!�ݧV����5g��L29�٪��W�W��&�'/���u{�� 5��Z�<1�^��+h
[4T$�v֡K��@0d0;�p�lA9��I� ����¡�.f<w����0%�`����%_��_M�7k�����L�H_f�Z��s�l�H8�'��7ad�Ud&�����s�A�w>U�3>8�L�TU9��%��ٴ��Xj�=	#v�	���;�dd��C�@Rz�S��p�`E%mdJ��`/;E�G�w�J�$a3��yI�g_�*�tڤd�00`�4����:���k?Ս���:!#�)��`��d�ߒ��\��3`�7;���R�n2�á��ID��C�7�E�X�"G�2_�ʃ�71�׶B��Y����#o<��ۃ0ğ
�G�K��^�e̉���� �#HW�^owS�2�R�q1+@�7XKP\%3������l�*2U��M 3�C� �W첏m�r��dZ�l-��l��}X�M2F���M+q*��g�q������L8�p4��h���@TbLV��؛.*s,���w6�/��Uٟ�"s�|&<�i�q.Nv�H��_���Q�/Y�a��P�Q�6�� fv/��"�T�ll��r���?���}����ذb�J6��5�4R����|��������%<������ƳQ����~�C�z��V���g�}�z��`T&c�������e��d}w�λ��[���ܞ`�%�4j*��̵�O-�<ʶ�����G��H�g�m��ǜ*�a��FZ%\%��S
�>���!��_�o�I|	s�Ƞ�@7�Ss�%E�n���c㨩�
X���v6�R~g7��M�d�n_�\� ��a�Y�R@�
x�\����k+�c�w�Z��p�F��ʫ1�gyךt�y̦f_)�\�s7�7�+h@V��%u��z�Ɯ�FI�Z~
�Wu^p/��
��E >�i�d�o�.���d���%>�VLS�t2SЇ�oK	���b���ne��h���T)�u��#����@0M�M�,ڶaC���*��t�9A�6��O�Dy���e5?f�0�]x[�}�HK�2��8�6�Pd���8�~Y(2�Wkd������#I]"`��.I�g�c�'��y�����'r*n�r�V�����MA"I(5��d��N:t�kz^]����*�-�B�.5�d���������S�(5����Pj���b_��ߨF�>vX2l���9�w͌���e(�c`�P����̂xg�`ݑ̊���/4�W�J�JW�v�*_�E�8j�:R�I���S_�rt��*M���~h���,R�������ޭ�)ILr�n&�QG�q��k+G�T��!�>3��Ǣ'Z���t�@���D�ë��W28��I����ڜ��G/����,���1�37�A��h��w�:S�a)Yr��vݰ�9i��3p~�z����N6���q@h��������(ˌ�~0�s��Ǆ'��4�IJ>��]l��l���dRu^z�s̀�.�:g�4Tޒ]��]�6�	!��2m�e��f�t
�,��3�����
�4���fQ��k��ܖ�4	ұz)8���:=х'Mݒӈ�c��I�������H��N|���ͬ�lG6 �b����2��2,UgːZֵ�(ctM�)��YD 0�BH��� �q}2u㥴̛�,��|���+sz�a�ʈ,%c��^��e���=1Bl�@�Y��@���f�wVѰ̝xi�;�[�]p"�h��?d��rE��7d�&�cĹG5��c��f����;���t5�N8Ѹ��� Z���T)�N ��L'��%�W�ސ-�&^u�ω��r�7^�hAf\�c1_��ފ2+(�Vl:�P��&y��9�����
2���{;��ǭ��r�<�	��ߍ����0qھ�P�g����b�ٹcٵ�`w�h���W�C������,�iy�~'9���5�̏� u�O)�a�����\�|�mT�*���>����ss���_�O�K����?c��r������í/^���<�6���R^�ܞ9�ʆv'�m��\
ʲyM�B�#߸�T�u�HA|}����(~�Nԝj!�X�����[��D7�xd?��zrqA��` �X�T��?/w8�<<��f��cN�����帄�a)KX1��\�d�O_�sjW����J~�F�d���� ����%�����8'Q����w��g "f�<Nʱƣ�� 5"��%J�d�0�{
�<�m��Rc�Os�#��ϱ�����V�T~<�BB� h��A�+ױ������^��X&,!�#?��܊���F��A�B�&�;Nl0�$~m�K0Hݷ��(�Ȼ�B8��f�X��*��3X9���+����PN��+�$�3g�y8.�2h�����x���`0���_�_Bj2*	�w�ƞ7טΔ9X��6�ns('�3֑%M�#HC�9��2m��8hvϽ�ރ�d��qs�f�� N�3���:�9�O���
�v�����<��Ֆ 
c���}�[�%#[�Q'��y%<4V���)<=0���8��/�jˉ�ӆg�`β	������V#;�C�ڹsłxc��<�P��{WF�^�|���lw<��w�3�B�jM?tK�ɂ�%���$�������,�d��<��jA�$h��M�Cd<H_�r�Π%)W�Ĳ���ۚd�����m�uò��c|Al@�`�dX8&�1>�%�5�[��6 V���g����ga\���8���YY���l*�� '��  xr� ^�hxt�zuæ��ً�w�d��� �Qq[�8�3+}�H�I��6�A����++�]�G3HΧJ�- ��h]�	��RY����-׭b��]�~C��X
�#+�(����.��o��b�wb��R/e�/��<�FyQr�-��_����Y�LMp(*��\��[�g��=�Py5�ї6!>'Dv\�B��0�o���m�M����8����O����;E�"� H���F�F�CEr y��U���;�tehH���峪Q���0�m5z�9�%^�.88}
6�Pj�̑C@3Fbh�2I�>ϑS�ka�e�y�}� C��fo�?��A��$J�n� "�~�*^F! 
r}��0�Fq��R��|�_`�@#s�H+�;�WQ' ��IwԹ ��ΙC��3N���VP�T�7�Ü|�v'��K� '��M��	������ls9е2�WG�w�mEi�^%:�H�B��Rf�+�EA��%Y`��D����#$���DQ{$W�=��{��S�h@�rk.h�D�P���{@恃��4��r
�x�A�<I>�T|g��k�A�h>�	�L��Vt��V�[� :FH�A��-	��em��VP�v�����^R#�p{��i�h�>�DW ��Ȍ�#��I��ހj����A��Ӄ����*h�͛�|��TO�e۵A޶���HH9F&w�b��vS�[������W�}X3�&ئlPU�����ס�<�ꔐ�ϝ�1�sr����n��Oe��//߼��b�"�mv7�5*�=�T�Z��Z��)�,ֵG���Pů�̬J�<���/J��28����g���e�}�/A��f��D���N�����2���X�@Dm:7>>���-��o��>4� �i`���_�?va��5E��A�D����ԵiT�g J���r_)��x�	�Iݐ���Te�ʦ���uU&�����Y�.���R�,��<B�r�t�N6z��jK&DG��n�y8y�'6[���З�s�u�JF�t㎯�Q���6�$kseCbU�b���e��(q�8��D��Y�,��8ѕ�Q�J�%�r�0�����Iy�w�&�y�O4;|@���(cRF
u�������_�΀jSd5|�㿣u-π���4^�A��<U_�q��Վ�|�'�
���,�,\���M��]�� u]ߗ���g/�u�w�âtp�a3��J������3q,8�ρh��S�LE��ؘ����sόi4�$�!I���yː��{��A���-�YlV��/r,���y�u�����^���F�2~EGPǕcΡ��m�ԡ�9ޫ5���ֲz���d RY�H���V�]��8�W���E�/q {���5��oX������k��Xc�K2aJ�X��4-F��QPcY����n\fD�y�5m:�b��jo)���rt|��e&{Os:��!�7���;I��~��Ā���*�Y(���j��{wv~E1ш�Ax�����������(�7֤��:�)0F)�mV����ٛ7v|�'+�kh#������Bp�_j��"Ƈz��Ǉ̂��`~�u��%HQC�A��?X���uLk/�d��M&[�e@�`%J�,i�-KS����>9��~-��^ʓ^�+��5_4��*��V�#��)���k�py��p��
�UJ^+�Ff�O�	�f(hG�q��n����������y��a�!�!����RnÕ�n-1x�	 �r.���N�L=߷���.�L��y��;s��.y&	�D�Y�bc�\K�E1�1QTf$Q�G��v���5�&�h��T��2�LNf�\��J!>��}p� \3��.����j<��ڬ^0�
V��ғx�3�R���Π?�C"���w���Y)4IQ�������8�aTA�|讀��1�eo9�H7��7�� N�d/�9�y�PfL癨4t���:`��!;8X���S����5G&�?<r�E���/��J�U�����YhE#�:����k8f�+?�g�z҂��3<�x:K$u������Xg��Y���~�喔�J�w�Ɓ3��(;e'�҆_���.*l�4n�7�</Ydgdq�JyX�!�7vX��/ �sx�G?��5y��������\�ڗ��^-�SVA
x�n�|S��#_|b�Ty�;@Ud��C��־0<��ڔ��K�Z�4@��f�/k���e;�~����~ b����� 0�|>[��:]K'�5���Jju2�x3���Y����;����If�X�P�"x��0V;��ސ�"��c�ym����'vC�V��4�C�n˒�{������F�m�R d��u�Ա==��J��ˣy��H���(��Z\^]�_~|'?��蘹����t��F~���	f����g�[̓TC������t��)�\b6�[�_��Gy��K?w�u���L���Y.>_|ͼ�ut|��>��S82Q0w�.aӓ���Vίn�͂(+F�@��͛S�曷��W���u�Q�>��O���a�_��D���뾑��߼~��oA@��^�,����bO��ɉ�|�J��ʄ-�z
�pnS͌DxO��?}<���+�����[�����~�е/n�Zʧ�K��?VNȶ���޲�tx��˿8ޗ?����.�o�����?�u�w6B�6�:A���7����#�>�N�ۋ�ͻ�����[�o�}�Z���7����5�W��ܣ���EFS�)96��]�ݨ�V���9 /7����K�-K��W^ZO ��N_7�ͼ��-�k���2@�T�H�;VҬ@����sV��[rÚ�`�� �V�� Y������>A׮����@<d�TYC�	w�	�ad1��Y1}�)tzrD�u��Y7�4E����LX�(��22�f�mN/�'P��iD��y���D�z�J^�:����_�E.�%�<��@��	v=zV��H:���Ԅ3g:�i2�L�a_�<����
�O	���o�_����I..oe�h2l���q�A�Ro�Q�aӞۯ�W����e��D�#�=�����ǀl��ê�\��{K ��I �~�)i5D
}U�X�>dy(�!􈺜���<��%����4 3��9�-��(�ϭ����<hI��j>���l�<��h�_���r��
�~<~������4���W��8@�(�9�T�����3��; ���eq����Ҟo���<@�_���g�Ϣt� ��gk��E��ˡ�.�+@X�_�Q�3f��������@3%o�C�|b��B�)���S0�/AF����ۛ�b���;`�:Q�0±��&h��a\�2i�;��`�������m��F`Ӱ�y���n(_?{���I�%�f�����������}#G��Og�j$�4~#��jJ��r||�n����f$��͗
�.�w����ĚS��h_~�o�o�2��[w)��?�$w��F�����ߓ#{ `��mi�Y��8�X꥞[�y�Y�.�y_��M0�@�W
n�����~q�r�D����R������
�~�Z���kuR����	�1E��zA���J��pO�2�b4����V�.(�� ���+h=��YP9�{_�����^�z������w8�]�a�[{J�s^"�+�~��'O���߽���)�1kz�˿��s���#�V 9s�ߥ*�=}���
캬,DG�O� z��cI~Ҏ��G��_ɫW/)��A��ٝ:�')e�8��� �&	e���B����������ưFcĭ<ޯe�l����,?����9A�=n�g�l�I�l��K��ȁ����&�)��(���T�������AWMy�;IM���ӄ@b���?3����Z��(�P�!���H��,�V��}0��5�o��>�������R�����l�.�+K���V�"��{�gᛯ߲���O�K���@u:����?T�~l]�]O]a��h8u�H�˕>�k���2֧'��ׯd��l�r�?��uc�'4�P�V�N�Ԛ�Axx�0��Yp���?|�k�C��b�]��`��gE�@����Gc.�nU�lɗ��ڌ�����8bE�\S��3��kS���c�}q�2B��V��eF9�e����-�Nq��h����x��â?� �����/����\r��p��{�57����.|�覞�-m�����>E������|�Q�6��\�W ��\�˭���k�d�r!� ĩ�r1B�(d'�\�w�e��8#l|�~]�2��e�\	s�D��� )���?3�]�� �z�x��W�2��	�
�6���Ջ'ꀎ�cR;��7���L�>�� ��?���+��;}?5��NY�������3�������,Eh����,n��(M?ګeM��!-)1�5�sA��[5�_+�88P�4�(g�R��с�#���f�C�?NX��H��8����̸�sp��}�\0C��[����L�`�y��P��EB��;�s�v�� ք��Zj]s�>��b���ƌCt��}� �(ϵ����7/_*x�q] LN_�ț�/�	;8X�Ȥ���x-��FZQ�|A���"�ں���Z�}2�2�w�:& �!���ބa�=����:7%[���FƤ�hK�4�f(��r�����\^�\��^�d�?�T&-�(H[.y_�Ԣ��N���NF<sU�Xv��	�u�g�g��3��Yة�>(���{S���b��K�ԇM����'DN_����G��>g� ������LnP?(C�:H^`�*���A@��)i� ��T �Op* Jd�9���;�q]@��9���=C�e���B�1� N�%��	VSw�';����}��6:��b|�{5�[�6����}p ���~��J(����+0��{dh�olmTZ�����KygQ_�착�W�f@�[6�p�V0@b�@����%�b�lc� @9�J��j����������˰\�,q�@�25�������{�>^�3���Y�h��"�X�E�c��0���j��c�����KC�I���=�s �����Si���~>pp�\l�)���Q�Bݱs$63��y�̒�8 �fF ��X�&S���X��g������%��Z���E�����Mҳ7~����3#/S>;2�A]�ׄ�R�/)}�Ld�]C9,�/Tv���K �<��R~L彞i����<�_�Ry_�İNc�]�k�;��Y��g�EĐ~��)����������ت>~)}�y��˗�Q��G�5���Gy0_2\�u9�ua} �"0�f�����g�ՉY���l��ŕ���(t�����7b훯�w��ZN���a`Lʚ��Ƥ�( X���Z~����7��l�\��/�������=�rs���͚�c���h�b�f��̌�׳9Z� a���_��`O�VB��d�  �������tY���Z~zgC�'N2���٘��)B���H�{ )��Q
F�L� �ι��B.3��B�� 1�&����m��eR����2TȢA�	��C�z�@����9F�4�Ig�G�O��l����5O�~?���P7����󥗖L=����M�\(������D��t�)�@R���UڿKV������&Kް�}3(���[N�'��3c���@�><���X��į�+ 
�thM5�!gâ���x #|Z��@�N�H�� ���i�LZ�M��,�S��{m�e���{��|�ݷ��j�̲^=�Y)X]p�(�YG̚]��}�,?��R���� *�=t;0ˆUE4��x�6���s'K�:�A�u�phb����N�f�E�l�-�oTQc0y2
�Œ���
�O_���|�J��5�2D3�U��~�8��xm��X��E��-6�:�3U�y���QFE��"��1�o�<��� �P������fm*����!&J4<��[rB�t_�.o����%X���	/��r8�7.����F���Y����P�z�C6�x_����%ϬߐHz��#O���ͧD /�,���U$r�ۮu�.M�ᚓ��^flS�r�t6���
c�F@e�)>!�C%K�?c��ؙ��E{2M�*�������q\�M�s�ן�僌��Z�������~����A* ��O*��H-A�'�!p�c�g�h��_���X��fF69�	ْ*6� ����7����"��4�k��]�Y>1�@��R��̉�!?A�O5�K����|�ա�o�J^��c�ѽ���[����<(�x��a����j8���������?����wZǤ�a�Sqw,�k�����UЅN�Wo_����7�������#*�#}��b���R�_հ��8G��*ࣛ	��� =��|�쏷��f����d�)�#��	�@\+$@@~X+��k���A>���+ �O*�i�=���P��F�4�y�L�Qp�αL�o �/
F6�� <!���X�O5Ҟ�S�hZF�v�':tN�L�X?=2�S�cO�\��%4���T��Ӆ� &�
Jp�
Pz��T�{ �O��G'���賽yA�V�~^��������֦�,
"| �w?���:,-�9vSf�l� ��8���6�؉p7V
jY��By�|/����W���GHSy�����3������T`m*��qF��4��
'���޾���I�Ċ�	�z���P�'��mFnc�Ls���p�<`�%=\W�
�s�-6+�_|J��a����)�(P@�(@�BAE�g֚��%Hf��uJe�@����7m�$ˑ��̏���<*����Wd��"��_wegg/�KNWwUe��q~���*�g�Y�FOLdE��]�
@���h�e�y$s�7!��⪸���}����!S�Ɓ{o]���(5�s|,�>f��M+9;ڕ�ߡ����|�I؟�M(�ֆ��D�)�{�'A��p}�?�^,Yzd0��<�/�2�@p2���0����H'�ߏ��n�ʏ���Vά<���M9�N[v볜:�'�m|��⧍5Ĺ��ml��Y5��ɹo-�+�~d��2Q��@X;���eŲϘ�g���JA�?��6�ǻ�S���h�w�R�s�ҽ��H^�|J��Ƌx�LJ���+d�.�!^J[��e�9 R�pY�I��p��\90����(m�ַm���Q�W3���lX����k.G�?f��	���������1#�+�9��U��v%C��6 �C(g�Ӹ/RR�E�X�a.#�_d����x���3��{���7yw[_��|p!v�yإ*�oͶ	
�^�1T������P�{{����OKٛ�ʓ(��(O�3�c9j�ɏ8�ٍ|�#�����g�1�ӣ=��\^�:�x���F�ޒ���~�y\���ry&�v���JR�jJJ6�S,�b5�V��3¶�� @�Z�zm�	�"�1����>�h׫��k�F5Ʉwq�T�{C�a䧧g<o4B�"�N�;�4�*�*E�\F��R	W7��;����≃�m�J;�D�I\�\����gY*p@�M��:(}�G�	�:��1�kB�0�u���8gf��D-	2����r-w�6=��b!3t�Q���V�7J� a�R��6Ҫ�e\�u�鹶�~��4>~�sp�> <�D
���Q�2��U8֡������V��A���#A��d�2S��ˠ�gd�Й7a&e� NzԶ<'$�

g׋�Vf��MS����I'�Y�	��D�5x�)3q )̖j�%�0[���]2�Q6)�x2�V*�V�U#]%e�Pt���ftrt����,�u[W�<�U�L�x52��h0������zpr��5\�k�Y��/v���=<<⚼���ۻ[���3A�%K:��\!�#(��[���L(2��]ԖmG������m��.���R���$�=<Pj�����M�n�R���Ŵ����=��['���9o��N�)�+v1o�H���S�9a%�I�7J: �뉐��f�*������Ov[�MK`���
h����I9�2�n�{�x�!�˳�p�F8Jm��I|}�Rne �^/+�u���u�������rX����������%J9� �G&�*\�\^����x7�s�R�J� ʙ������<��J^�y	��r��5����O\�0���;5x&C@=|l2 �e��-�5���\�H��C:<�r����;�A@<	�k�Yf07FyCYm�sp ��p���u�lV����x�D�X���!4��||���.I:Ei�X����+��v�qM)I�����m4�ì-e_'�WYq\�]_�D���J(4W�f�*$"CqCCW�������5�g�t�(T��n�����]���4��,f3\m�����5:=9��o��n|����]t��qଘɪ,�����7������R�!�.���?�*0��hdߦ`����G7���h@��l��!���:N̯o�LA�zK����v%E�B�@j�2_vB`c�Z s��1]%:!d����d� �55 ��4�窈Ӻ������Y30�<���ѵ1
*�º5��d�����k����<;���.[)�JTp��İí��Ad�(�{����0�
L�G]l��.aN%@@P�|:���lײ���%�ZFg�Rin�ϯ���K0fG6	3Q�N����ԛ���]vE[��\����0m��h.��Er3�;��D����[�J�5;7+ޯ�^��T�S4�O�y)k
���cf�j�X�F!�&_ǮDj�A�C�ӌ�c�h̬�6�7���_\^K���7ک���C�W�Z���Ϲ�V�G�����k�^��;�ځx�,h���J�V��g��4��N3�|�*4!�y�����;&���#r�:���x���R��X�d)�Ҫ���$U9�~K�Z��;���|��)��y�Q�H�r��@�7��lÃEw��b��WɼXh-1�:�t�=�S�0�G�o��{��ð-���WOڎ��ϲ�@��_��o�	�|����� @�^���
��:\�ɧ���T���+G���]���/�|~~v�=�+�2���6�:��7���I�q�������XE��o��U��!�̚��5�2��LB̜ð�rkQF�
p4�e�p�a-��/����:���B���" �kC��{�����fE������쀿2�|:@�]:@8�CϮ��,2����e�>گ<KY3{�6Pܮ�pЮ��*F��D\ J��j��+ƈ8���	>���Ȥm|�@�rqf)f�URhч�k%rg9���yR��\,��&#u<�h�#���4^�T�% i���p�ᘜ�N1گ� .��)��Ƈ�Gk�f��Z�qX]­� ������)S ���D1��<�p��W6�ѡ�(�ݙ����]u.^�U4o���Bp]h)�HnSK6�h}dRr`�YRE��p��}�c���18����dB %f�,�k��c35�T�2QJ��c�8-!�\���S��yW�A+��3F(��n֞%������~����TD��D��(��z��ސ&����H!��qq�i�6�#9��D8]lS?N�K��g�������.8ϳ9��h�����6!��m<�F����ݵ>Fx�>�;��
��h\��9B�:f�Ak �;������K=>:V�'���A��7�<��k�7
���g��7va����3Y3j�`n��D���OB"�lBw���t�x���]��m�Aؚ�/45�>��i.e9�
a���^r�-�� S�ppF�O|�����\��R�H9� �$)������zY�PXJd+|E�As�Lc�١*.%@����}ֳ�2��noʸ�m`�n��-c_Z�*xJp
�Ɔ��)�j�pg�(<�aơ~�ֲيĆWj��xD	�h)����M ��u�����T�/R*k�W��|j���m�i�1�x�������B�8�5����F�{
(S�o��Of�WbU Z`ٜ2��x��O]P���·K�.Lw9O���od��c�@>���lMC!�]�+�!ȫżA�~sU���_������ޯ����Q0W�e�|U��!���A�ef
��l����Nh���0�؇���L�2{x��8/ϡ���/�Ut^�x����pu�E���{�N�rm��f�R&�R���&�s��L�)�:oM�	`6��-8�|���`�������d%�)	�8O8v��k� )���9q�*T��T^�
� �� C9���a�C�g���%�I�����L��?����_�?�����X�_j�9�k���.������< ͸���*��>�A�Պ|������$%��Z�!i`Y��tӎ��fd�v�ۖw�����g|L�ㄚ��=N��i�Y�������u�c�0�>{pD�Pjt5v�����9-yjk~sP�;NV�$��4�(슌�O�e"[5������%u�R��=f�{�L���X#(j��LT5�\EL=�/�1μ2��G4\^Z`��c�>�ߩ�yfv�����
�K���Ý���_�ݻ���*�H�ZVm�uN�^�9<�9r�������]2����.�]��_7��{Y���AI�� KL� �R��3� FU��Gy���׈�5f��z\�@��`�g.�s'݅�3�Ҡ��������_� _T
=��?�~�~�%�a��\B�ʲ�A�W����!(dh6+� 6�r� 3ep�M�Ȁv՚cA�G��n����������@\�]]�!�.�@ϴ�*j�Qj�6c�%=�������=BݯrY����^�U;k�Q17~��_!�<�u�B����f�؃�_��/�A��R��w$���סo���`��r.�����<21yޯ�;��-�WN��I��_���"�㟂p��΁G���;<��I#�\�\� @<�e�l�H��{��F#whT��g7*��H�	��2�=�[��&�7��{@���c���99Hp4ˡ>�' "G�D�K#Ao""˙������Ĭ f���t��c��q��Oz@�e&|é�u���ŋs��1�����'�4�F�ޥL��
���=yz��r�0��0c�'�1)�(M$Tԧ��$��':�j�L���$��+B	e���9u��ps{K�<�V&zۘ~O�16�%+��(������2�lFϝ8� ?����5���}�`�[���)��2��> ��Q{~VЯ�c[bp4�b�8�򿪒���$1w4t��i"+���5b����P�dA�.�5shl�9���;!��d�\R&�,���`(%0��_�l'ݙ�.A��\^) �A�� o2��`��Y��l��qͱO8���.���^���5+�i���U�lB��mv���6s`�D�����0��Z2��:3��zm�Y��8H�X%��T.R+�zr�W������+�ٰ�>���3��� ����{�����A./.��,���I��g�Rr���(&R��~o��8 \��
�P���®��Rj��������|�+�x�]�ވbM?���8���L�R�ހ�U�)A�H20�h�^Խ T��2( ���w�f����#�2R�����ﲿٴ�	�&�(o݊�"�e�������i�e��E�����@�;fƔ����ߋ��a�O|�He�&��\�.��3�D�ӒX5�S�R9�/�uC�`i�y寁V`�4�)�,8\������������	�o�<Hso�� �����PP)��`� � �d���'�����M�!)>aH��wr���ZN"���U������5=x��i�,�J%�V�W�2�(�`3X$��m�A�Ue��BV#E�� �Ú�D��pZ߼���xf�_��b�K��pri]�n���Ӄ\_]�|�익b��k{�XU<~�.��!�2��?M*��"}��`_����M����Q�?���a㜤T�1��	PF`FN�9OH|��[y}�BV�؇���ӧO�L.�Y�lgwB���~�,����gG֢r�������	��3�ob�;��3���ug;,)B#l��O��!��G;{SfW����� &U�Y�ʩ����n�g��cd�r#���8~�	ch��	t��e�FuD�
�V�8��9�s�]}�p��7�
��1X�%.*Z�||�d�3
}�U�1�4��$Z�g����G�L��e$Xn[��?�=I����.��f
�?}��;�B�?�E�>�t���y�f�- Y1d�B�|-v��6�z}�z�e�9�t$s�����|����;e�ޮ��}�燓}��u]�~!���w�rqq�`� <�A���!�su�Sf�����.s�Go[�Y�af�Y�؏�'�s����K�H������r����#�����<��P�����g���A�����ã\]_���>����m&��^�f+�#�[y&���G��� a��i uzu#?~6/�j�+��-:a��S�D���}A1����Mz��a�[����`i~eYN*y0b��d`�*�ݧm�̓���G�gQ�X�r3�������@��2�"|�;=��-}�r���:ګd�[�F��!�$P��*&���T�ecB�^�C��#��!F	e�: �x�.�ކ�9�m�뀨�].�t����<-�����~q��.��+@"p��D�>V�uRs�*9Y�R%����Ή�玠*6MyYO�+��3y�Y��T!���e�`&>k������!���_��4̹���}��0ǝ���qɩw����x��1��S�������|��������FX}���P�N��D��;��Ucf�M�����gĽ�qGɵo4rX�x��T����T@�~x�SW����Kh��`o����a-^��a���\��(�sڎ��5]`����j�����.�]���������:���х>�7�����v�P[v���Ƥ! ����r$ �
9��Ȍ֏��5�Z���сYս�v��QF ��$@�����J�3����+M� [h��>{� }(9@g�"�����zf@%�X�=�L��������1SR�:0�q?����"@4s�-m7;�6�m�~?-Q[\=�K�,�Eݳ�8aMmrs�� �Ѓ���x�d����}#���S7ƣC6@s�ex:��4�:���i��q���C��G� �5�F܏ �ϛ���s�>���F��s���f��a_6����Ȱ��2y�0�[����lS�|�����8�m&�<�d�QD��M���.a�&n p[/���JO��6���wЂ��r�Ә  M���a�!��R�uU�\�)+���sF�~n��ɉ��p�a���X�Ϝ���ɦ+�֐u�|xg�;um��>}Ӻ�l��Ÿ����Iml�v��(D|�e){�)�qG5~���ip�� �<�pοp	;i5��1�@;mhg��@��a�0������Yܚ��d��-�r'F� ����6�Nښ�V�"5 �@}PȀQ��uP�$�a�(ҶE�[��Э��{ �e0�
������N�x��|֗}���Щy#2�\��}��x�òc���H	����x%
�_�2�m~!BA]�ז�T�Z�s�t�0N2܀G�=���X�q]#���Wϰ7�[%����@s�v��iD܊m�� L+8��[�b�3���W+�X~�� �����a'�W��a���rN�
k?�  �ɮ �?c#P�P��j,0
�	-	ľΒ���i�z��g�Z螚�À�`�,7j/mx�Ʌ�6]��[[G,#媌����=0Nu��y�n��k���T���yy%'{�LΥ�1� dA�Y��p� ·-�#�ch]����}y��l�cy9b(%2���!�$����>prSJ�M���n2! S��s��߾U�wn���tU>?�볽3nSem��\˟/�>9��`Ӽ���3�&��0Je�ܯ1\w�QaV.�ۍ��u�7�����l���%�9d�3���}wO��N1K҆y�y�+ �� �]lLv���VL8<�D˒����|�`WvN��s�(:/p��=ܙ�������ͭ�Y�k>ߣ�	�!2���_r�%�����\�˺�r��͚%+�g��Ig%mQ�Q��{�i����#]7�@����
�٭�n��'�� ܫ��7�9������l�! ����y�ѕfb�бZgd�9s�$Ƈ-������[n�n���6���Fd/���=�W�m�K�gL^5&�|Xd�0��Q''��n���;�#{�\�8���������m�����w?˳�i �5+J�=KM%�=X��T,�Է;��l��BU �*���*�N沝	�4�*�d��7��h/:ʣld}� �G���ll:�qIPS�Bڂn��K>ŚaZ��(�,��&��Y&���,��$<r��ZL2��l��s@�A�M��� �(�'�HrUV̒b��I/�vX~GatL�Wu,����A>+ {֍���X���f⋶�������7d�)و�&��Gj��a�fQd�W��8 c��RNm���ξ�o:��ߜ�ZC�]{dz��Z�����o�aB!�C+�"�ђ,�V	�'՗6�����)������/�\�9��|R��#~)��:<�RQv��gT��%6lo�y8��W� ����Ӹw���9Q@�;��ת}�0!��
���V�{��~��p�W圙�a4g�8��ՐղWc�)�r�0dJ��;�.׌�`|8�v���N�稱�;˒g���beI� L��wa���C����F)�3��^Yd����H+s]t��l��k��q&�/ײQÌ� �]��r�E[�5��!n����+Q�xtdb�(�҉9��F�
D&� J����G� ��Qm�e+HC@m���I�Ō�yxpDb|�<�f����RY����&.=�6���f���m� ����r ��=N h!rQX���D��JHl�z>�@�gI�R�`�G*�K�M�mY+�Ô��:��E��ASr�äu�����Q�˒2)�.�u=k ��xef�����ށ�J�ox�,���X�,��$dY�SR��*��q�����h�`���r-`���W�嵂xL#��~|���G������N�3=�1��v�7�˹^?	���ă�`U��\/�qE��v�\,���I��:%���°��}d��c��2�w��p�� ��x�/_����ڱ^Q�BL���>	"[	_��O_0�|yqI����K��+)�F�>L�5�𪞚����#��3p��wٙr}IL�6�Pg�X��� $�`U6��u��2��$�<K�3]{3�C�@W
^0@%����;�k��5F?[�J��U�C���&�{��e�DQ��$),�y;{c��t׭��7v���*W5���1`�נ((.i'��vK�Q�Q��hk���A՟�P7K��+��Xf��"+��iy6����ʌ���5Gꛁ����L�V�h�=�*�%*��p�b�&���AK�U��	:4����X8�����`�Y,�H���Z~d�JP�J��ϫ��Z$���9a�w�[��\_Q�/�u���C,_�O�eڂ�l��SYH= ��;\^7Xlzk��T�:+#�ft�G��LI�L6p��n(�f1���[Y8ǆ��:ȶE��$T��o�C�vk~
3��Q��t���8WL�8�-�	����6�k'a'��I�n��#����y��J
�nn����L7��B��*��G ���{� d�*k�K�]�Fⱓ=v�MF�n<��I�)r�[[��Á���av�EB�=�@bɮ�c����aӄ���_oU�D�q3�����ZF�P���B�.���˕�{����|�Ϟ�8?��cd;f�.>�ںe_F$�RA�
k��]�k�p�!{|j哾�����|��}}f�I8& ��J��ӽ���>��;rt`|���1[\�	J��\\���NP��0p#�Z�9@~��~C'o%�LN��1�ƞ�kY��s�������J:�.�)�0�P�i:�Ryh"�-Ud	��SX�Ԇj,#��_�w�3Xq���&,�m�s2)��|w{(�w�,?A��T�i_~��C���3�c6�;���JP�x��A� ��V��(4�A����ɕދ�&���)�?lbL��s�e�N��I�8;�W�dg_����Z�FXm̹��6�)�8bizUK]_�y�s�ޡ[I��]b�ןt[I����:�Ⱥ�^?�¬�ya�;���Zf�<�`��G�^�=ci�G�A�w�|��7���o�R����u�������G�x��X�<-W׏ry���o�`��qL}6�Ȅ��EBG3J�)�������G����=��\ ��&t��#�0�d6A\��!^���v~�ĉ͑ެ3����W�{��s=a�@JN:Tk�>xژA�aC��<t�F��j7A�ͧ��!��BD�4����X���nP��	���z`\�t?C��{ER'�·�
���D?)��f���;`#���������4�i��Z�$�q�a��1�:a3��7��&fH���}޽(I��V�X�\�uTI�&җ<	��Ȑ J�9��c�A�ip,
�ǌ-��F̈yM�D�A��r�">�(�+�{:���OC�e���_H!��E���t�o�)���2c���ץ������<.�����l��s�������/��A�cs���3�Eu.��9�54�Z#\�3��Al�Eq�3f���2�VWc�c|7(�A�aM�r�n�)b�d���ُ�u�8`�5�|s��-Y��d��Q�	�*2@��3Y7�dL��	�"g��j>��ƹ�4���qP�C���씗MKtM&q�n<o��� ��47è6� (��u@u���9�h��ӹ �$�ɮ�&yԎ�@��M@�����v�ԙCM�s#�繻�L����L�0�&�n��%9VcqT+_��f�:�H����6��02�)���'�[S3��o��L��U4��wԹ���cF��GCĎ���>2aJjj!����G�s31be�t�@�"�Ub��bI2�q�V|��e͌�IRd�=���S:����eg"���8w�ZX.�
�;[U���K�vG����{
��g'�pD��r>�X,l&l���r)�:Ws�k�����3�HНݰ�����k=�5�����[x2QP��X�QK�eC�9=�3�A
21�"�G��r�ˆb_���g�h� ���ϫ�_tm����V��g&�]�neK`� ��ƛh���L6�૪�������+$��1ު�qAf�.������3�Ӊ��>;�Y����0�� @(W�����q�M���-nW�^��z?'���߾y���^���}&�f+/#r�xJ�"ǵ����y��	z�����͜��i�xF��|ձ#�ld��&y2H̷�R"k6pTGd��̮�ٺ��YHP�Ew�u���5�Fߔ��=��y����S��0*�WF�j*�e2����H�m@�y��� ��3|�eU�� YXS-�D�y�rzԨ���ǔ)b8���TcN־s灴�.��	�FJ��,"qu���S|�$O���x�,�i��Ԑ�3[��̌\ň�]7mE&he��R��&����wdXP+��ŝ3SM/6�)�>u��%�[�g�5�m.��f1d��F
�pQd����� ���W '�����(��8-����vf�t.���):�j�@ �C-�6�p�3=8pr�m�i	�+�l[\Bd~r�ڷ�N^�k��s����7��7Ku�/�,�b��H�{��b���i!�i��ʥ L�	r�Y���c2���:����l�O�e�!�uSڿ33�R2���D�2�����8PԺ�i�V׭�@�S��H�k�{G�(�`sC,�a��R�!q;�\ �Dv^�Z��EJ�q7*\ˮ�,��Tq��*������F�տ�gsf�+�v3��%��Ũ�=Ź�X�_���8e6���Οsk�d�0+��'���>���l`��1{6b�|&� �}��Mh�j� �O�XR�-m� л�7������N�MwLc�u�,8]�S98�Sg�d�k�`Im$8(��.��Y����,	F�żÓ�#��w��7߼aC�+u�B��P� ��:��a�q?	�6��*���^�ŀ���F�:������3f-��|!�Y0t=������ �p�6�� qy�L��ၼ<;�?��w��7��f�c/��K~�}x�7Օ<��s ko2��^�����v�����&ϑ�l���^M�;*����}F������\�>��Ò{3���8ԕ7_t��8lm��Vr�0ˉ�wf�ہ���t�Ob��ܙ?�9���ӈ��\�R���.!�@��@<N�)ɺh����}��q{�Y�etp�u 2Y��v�3�f�j�r-�)3ۉl�Ja=r,�ݵ�?���	U����������������E�Ѧp_ò�q���0��<H��
���&݂�.h�%�0�c�k�c2{�.�k{&|������\��7Z���*�;��i+�����Sc�e)1 ����gQ&�t�5�Z1�1V�1C&L�M�A���+uR�Z愭��&�&�F6^�/�G�`צ�d�l9c���{����|�/xq���n�񷈄�|�	[PL�2��Vͨ��覮Xs�h��bL�/A�{ʬ�}j�K�P��1�6�s=�ͯ>�#}w`�����3Sl�Aؖ��6��[����R�����v�W�.�0�"�E�H 0�}�\� %��5�Y�;��h�ĺB
lM�#��Ze%*�N���\S��|��C�u��[����<��0�g�����v�`O���7H�u��ֈb�Tk4a򿳍�;��A�PR*��1g�%��#��,/QAݯFY�s����11=)�yy�kӚ dd]���r�u��ՆeO4�3Ƴ�h��y�h�P�"H ������|"��"G��ʞ�AZ�0��F�pg/^ȣQ�SM��"C7�aW���Ax�4�P�D���Cf�H����7���f�#7fڲ|; K�)���y��u88, �I��@��xo_�y%'gg���G��%���zT �1Qأ���l�u�<<?���95��΅�@?���Ń��%� ���l���w���݉�M'�gz޾�FN�'�8�1�'s���H����5 �&�����P��X k��$�4��ٞ:u�;=��q�nFP�3S{�׸3n�p�+�w��9�8=�s~#o4�е ��r�Z���ý����3�޿)��>u�RS�e	|�͵�� �C��ɼ T��H3l��ݩuâ�bkw�b�=�����MOv�l~��ɀ��<{Mh��ĭ_���䛈OB��h�Iò�����,y�"�'奶��Q.Ld=6�E:���g�q���(�!��08��j_K)�f)I���]��'��hm�;��N�W�_�]���'
�rݍw8�����Q/N� T���͋��x��D��w��dr sqq->\���̤.:K4�#�Y-p��ײ�`v�L���34�j�&Њ�8>)]��b"+H[T*t^���y�Df�^b�a欂���R߈:��䠷�h0�W�A�ڈ�����,PZ��ms��3q�V���w��"�n� Fc���h�<�(8��@
J���r�A�5i���ʹp�
8+�w�X�m<�~��4H+��˞U�E)�!��]Y��lQ�ST��d׍����ʺ�89���;�aSc�2 3��E� FK(��R"�����f@��2 _�����;�7^��s�+��,Zp����q�� l~�V9�����\2gP�J�j�({L\a3�P�~�ɽn.<���9:>V�y �C��̖�AKN�����+���|=��s7Cb"��;v!����ӆ��V7��\�H��4`����v$C�R7����5�N�����̀�u+�i�w�,eO/�x_���f��Fq�������񣔟IGP2�wM���F)��|%8D�n��0 �JW8F�e(W'u&v�%�Ί�}���ZP&f�`�h�7���*tD-�*�b �����N����X���=�g�o�
�N�����{px$��?���r}+�n��LdUF`6e"�ȒR�kg��>9F9���	+ ���
t���	`0����P;M�����.�/�^�#�Dǝ\�J�2�
�N�NN�i�����ܓ���Օ~�����׀�}N�
����>W������w�}Kǆ���V h��ԍs[��q_�j���9p#��S�v�%�R�gb�˭��ܰl;r_��ޔ��?=?=0c��N�����hp��_��(��\H�k  �������><ڽ./�4�\��O�,8�ѝ@͔�� P�>8���,�r{s-�Y>��Q.�ܰ1������Hﻮqr-�^�y�2L���H@�vJf�����^�h.�ƹx�^��l�%�򊍢�=��Fu銌K���1{���>c�.Ǔ��eM�{���S��U(E ��m|rL�{���wݹJ~�J&,�ȴU��qRXGXOt觰�j*���A��<sfD�8d��)�l|��z�&�5x�fkQ>Q�-���C����<��|����'|�v���L�O�t͌���!�$�<�;^�����^m���8�1[ؑX��_ˎK�G�
�:�`l�{�!�2�9���fƥ��\_�.�y֕K[ٳ�]҃�6��1z��XC��X,��Y���8�hF������)$cTӞ��/�L0������a�!S+k� �0���%���hC<��G��^�&��n_��󽺞�˿�p���G��*���M[��l8i\z��#qU?e�Aߚ{��4l��a���ףa4�v�(K���D����#2����y }z���(@X�>�W���5_}	Ϙ���SI��a�	��Hn������_`��&�B�h������Db;2A�7���A�oo�I��8��N����F5��~R��6k���np
4��y�HYGZ��jT� <&0l���vG� �0�`7��"[�a;|��p!��lMGg.V��aԗ(���a�Թ��������\���y�b�	_����yy�BNO�l�Om��ΐ?+�9��3��;���B-w���pC���+;� �A��ϼCg�:D����B*{�~�F���V�&r~�ϒ2"cw� 4�^��h���ip6�ޮ�������QD C\7
lP^�� s2�H`�R�|#�Ŋ�Rȸ�8�gG""|p�w"b�5Z�a#�.mXt��#`D��؁(��'H��|���ÅF�7r��h�9����>+�����謗3���#���7�oy�ߛ��7�	��'��y8��� ����/s=��k5�چ�`(�p{/����_�s�q��eFPj'�]<���� T�����$��â0�c��Z�u�t����H��q�.`|7��;�=��#�0��-�@W>��Zf>|�g����N������^�>�����=�3'23wJ�P2����{� 1�p�����!@\4��@��-�}�f�����@�d�D��4���<$Vs�)��b�ȵ��.�ċop���
���)�� �(v�� �������b�cd��А!�a762Z�`�JG�W9Ήb����S>e�������t�X��	���D��k�/.6k+�Y��(
٥}Lw�S2�NV�µ�g�Ɖ�&?_��}'?��^.��)ݒx���wb�1+�_2�\�Yk���krx���ɾ�lX�k(�p���l�۔,O��<_˜�M��x�k[�x0�^; ��D�	�CX���=�^���Q����>�g�A�$U��X�~��r���M��m>��V�w/ҘL8�7�*�-�r�����E�d�R���*�ǌ��cǘU�{Ԍ�o�����at�1.M�rph��I��'B'�5��OO�n��s�8��^{��@���G��k�xm��05��=퀇1��r���Uq�N����ȀJ?`�_}�_|��5Pg�4��:�l�)/?J䌆�dx�j����H�ٛ��G%���1��깕/�7r���k>�g���1�+���]5���.A5 �Ƴ:A^���y\s�Ԟ<�<�t�7��qbl�+�{�^���:S�k��Θ�C ��)��Cpl�S2�}�$�^�r+��/_�H?��70�����u�,mm��<W���:�Pd�ȩ���1{��{N��H��;��;ӆ��� �~�^.>}�\ ��Ý|����o~���?/V�FoU���y+��� F}ݭF�/�������g>�(q�<Uc�*��{�w�]�lMӏk��f��/��'u�P�������������#}N�������O�0�=���gdT����Ay�Zb
��uB�Ɛ����3�����a(ǈ���NtD�?kp������<���;!
0������Kg����0��;��</�ά'���	��O_���w�?���⑆Y�)2�(U����m���8�O�Y�Ae HlF$�	"�:L3�=�0�`��Zţ٭\��J���,��~d�L��L��������?/�߿�B;x�;�XN_�r���
l�m������\e<�~@�ji®�:�X�OS�0��45��؈��!R'�-��kL��f-��&wd+mw+Gy�$���G@L���~Z�� �N]o�<��K��l.x��M���X�����ݽ�{�;cVq���ऑqǑ,����R_>k0�I�������_��*�`3Y��\�=˿���>�N����:��Fm��u/�����2߱ZQ��)�%[� ���r\��<?.���[_?ˏ
�n�\/�2�ɛnZ\ `c��Vz�A4�!&L@$���y�ꕜ����������~��L���ܶ�%_���b.g�Ih����:rXS'���֩��M6�\���dc�[u�Z��8����LzNИD#K����ีR���ku��Ռ��f���kΉ"B�w�	�j�pd�U�*^U���T���� 6���L��2$8 J�bC_-�0�{5�� �A�Ǆ6
�.f+�U��p<���6�7�p�G76�)C��tY|�8v���į��ڗ[K�{|�Gi;���xc$�r�8u�ڭ�ۿ���8��g���\��ȌY�����#y�2��Һ�,��w��s�ΆDE�Y�̖+�ц˞@���Ov;SX@��%�U��Z3e{+˥�Of٢�Ȥ��7:UеKn���,�����y�R���FR�7�۱�-�	�<Z����2���
 ���7pe��uc�5yZf�Ѳ��A3L�&X�3*������A"��V�����Ϻ��Qͧ	������ޝ��IQ�N*��s�/�v����9� @�W�q��˛G����h�rv�/�)���(����H,�`Md]f|ɹ31+#����������~/?~���&��!F9R 0o  J> �Zf�&���s�$�V�a���֚�-�vu��ԁ|Ҩ��.���	��2b� ��6�$f�Zf# ��u=�M  ���%��'r��ʱ�	 \~�r�����9߰4���X2%������g�tu��jE��l-��q� %�тEu��u� �3;��m���@	����{����{�3��O����#�bF�E�l�7t��g1�0Yv��W ��l��$76�5a�1�#˨����+V�� g�TVg˽e�b�d!I�ɬ���M�3{�3����|ɺ�< ȹ�a�GٲJ�g��8֕=�SG,*c�Bf)�����2"eswfu)�`/����F5~�/���@B�`~v� >�/��+��IH���~{���������e�R� $l*�2N&���8Gd����I'�|�Ҿ!;,{;$��YM��4C1����u����-gKf�0��y�n��/��.�ٝ�ה��Y�6�c�&��;�Ĺ���S� \�'g�����>3�lʭہ����n���+���턯%���Q	�R�0\f(#W�5��]B������)����3ٸ*}��h <9:�໻G��{.r����}�c"u|�./^|Gm�5����j�e����X�i�s+�ӓ��i)R{q�N�_�F�0�8�Ì�I;��I����B��N!v��E���W\ _��5��1͛1�d&5p5*�F!T��]##�ؖ��a�2�o�kEĿ���o��?�A���Wb~܋����� ,��kʩHDw�o�'����ʜ\�Jڐ{@�#�����[��%q!"K0i��ѨI�F�f���m�&��R������]���Z�A!��������8{R�v/�r� ���I���L�I�H�<4,����©��bM�-o�t�H|����u�̊��U[ Z+�V��g�:�H�����r�MG9�ϟ�P�	�#��@��w�t/��7�.f`aydԙ^���-�(��_t�,;4~�tl��A�Ɠ�P�V�v���d��D���Gyyz�6��Q'��{�܏F<^�gĮ�Y��]H�>��<�	��Ņ��/��~��]�0�;N����3�� ���U)��ٜT2N��NF��F��F�W
*o����I>|R���fY�2�@r���� ��w�g�dάq��a�w��z�AVz�s=h��N�t�6H�d��wy}�@�	�s�b�r�ҟ�}F5�G����SmPK1W�8��e�q���s��f��B�[��z���zv�(?�S�ɱ�Z8�s��/ձ�V�� leJ���vc��>/�@/>_��왷�zu��)Q��(h����C�ާpk=1��]�T=u���=�<[sz�	�&��h h�qp��E�Jw�\����W��� r�Р��Zs]ד�5�/4&��t�(�&G��?�����Z���m�Ql���)6+3&�o/Zxw�e������F��������^�no�ͫs9���������;�\� �أ_n	����м1ed�k�Dmg��6o���lvy#�/�HzG���3��/_����w�o��]+����`M����0�q����@�w�?ȟ���dN�E�Y�)�#-Mnj�l�0`o�3��3��������w�w߽�W�^(9T�3epQ�&M-���	"����jV�f_�AZ��[B����x�aʲ�o�zԺ=�y#ۍ�Ѹ�D�xFէ I4�@�?�`�8$�`#��^tv���ܢJ��P���=�{.�l5^�B阎6�_�=���w`����s��u��R2��Fhڮ��aT��=���|�1�#s�lO�,x�/����P�|R�����~�j4�ԛ��6�<�f���B6Utb�}��kx�_�geJ�k ������W�/o/��~������*��J�}�ᨆ�8�m��g��(��m%$�L���N�8�QC�qR옂8^
�H5��K����r]1F8rr��m ~u[�g�$$&)1d6D5!{�M���c��e�[}J�wJ��,�D��k�CL\�~G�^��έ�B,�5~�	��F��u�œ�޳�X���i���ˍ|Ԡ��枿�]��586�IZ5�¦2!WD���2(���e_�����8@���G�d����J�����O�ۻ��?��۳��o�Dw���j�̆u����qt4` �??=TA���N��GF��� �	���7f���@_9y;Coso9;�Қ����U`���5y._�������Όj����Ҍ��_�k��3E��)����˵~�LF����{RPy 1W7���vl��R�D{�}�Pv� lE�4� �JvR��� ,PF٤{����-���.�s�;]c��+��j��V���o��~��<i`:[��ᐥSӿc7Ym�0��7�L��
`pu��+y��3��X�O�XaV���$a% Z|&J�^>�<��a��F k���?�c��Ջc�c>����n��h�O؜��4��������'�ޙ�<S��@���ءb���C���ܾ��s*P��&-�6���dbб��+���e�G��h�B <���9��B��䐶����Q��4 c��&0��z��0�祄r}v#N��(�C
(瀇>
pCJ�r�HJ�X��L��u���H�9t�Ƶ���B�|�b�z��_?~����,���^���Ȏ����̖��z	�]<�C��o��?����o���R-_Pn]�I�ܞ8�+R�����*)��6��3���1B8�����h��z$�*�*��%�ؙM��!&�*�;�j#�����ѡ>���u�T6��W>vh�D>2�rt������[�P�l��_d�b��_��4 `��r2��'�aQ� �`d/E[(�����`q:ͦ��h��h�;�_��8���^i�t���Z��|)���g��'�.i4��ф�M�'6��g��i� ��/_�`��h��/��F3��'�����Rs�y� �}%r���+Y�˰ ��!$=HrC$U���đ=]p5�^��\���������7���њhorP*�>��[��h�������چ�C �?;����U����J9�����}��A�G�:����U��>��yDT��r4F��ٍ,X`��7{`l���,{�<�����aNE��34�,8{�!`�� �;5b����� � $L��.H$=_p4���aIx_;�V����H����)�6�uQ�g$��1K�(��|F���#�Av�ț�'}�%������ڿ�b�M&&�a��HY�s^ƚz`Oj��ľX̸�K�1���P��;��^������N����8M�{��-A���.[+;^|��?��Nؽ<*"�/���1��2�CB�A�IEq^��l���K?@���AԌ�2W��?;��6���;D��_�8c�`�Q0�j��Cg+����>��(=�ZTX7+ʎ �5�&�R�l����$8���&Xy���K��;=�eO��Qet��Qr+P�t��{T�5��kyF�罼�t)gǇ��8��3^V�x� Q~�M�^d쾨�G�N�foJm�%)�����G��+~��G����2/�Q�O+��CU�Pa\_?�����+E}��?����۷
�����������(�%��>�?����g���p�AZb��SP�y3t�.�1�X�ֺ���Қ�#�#;���)����F�Ys�Ҵ��tʔ��k�R��%�e�Ά�S��l�s� ht�r�A�\���k������M�a��)(9>i0��\v�r���[�'r�X��RbL�������fEP4_'���K��iG�w����g��1;f9�V} ��Ϻ�Dcl2p��Vؐ����Z���,�c:�u��L�I��������?�᭮�C=�OLm#�6��5P�o�1��ƻE�! [ s
v6�>�T�%:e�Yq�L3-�s�����z�\���E4ǔsT0�Z-)Ȟ��=�¤��\��7oޒ6��G������"^������+�@ǂhc�l	�H0�W�<g�
1�J�8M��7��f�z��n(װ�Z����N��F&�F�7 hv[4�:;�.:�
�>]<j���@�O���L���Kݴ�tF��t	�����١���:�l��rG��r� A�K���}�� �5��PY9������B�U������������f��M���¥�,�^�H�#��c]c�w#]�^�l<�����,o&S�(�4pYDo����a����kg���[��4��ݷ6ct��P�f��g��0 =�����=�_=��F�Xw{u&����8�a��a8S�9,h�!�F�g�(|_T�Ś���I�s�L���yޒ���Z��<�9��U=!X X[��@� �
ggz=�q�q�Q��'��TN�O�=��1��R镝GG�(a��2�38��3x�:�s��3���?�Ӛ {4DI���I�ٳ~?j���l'ʭ�F�{
Zv�a��nh�@����L5pzR �Q+�5�x��ۙ�og���p��%KzYn���;����^�"�U[�u��3�
�*�w3�U1��NTܟ���t
�8(fun+4��M ^f:y���}� CI%Wpg��R��AAؽ>�5���"����17��nUp�`�[���o���H�c�Z#��ﱌ�'��s�u�ks�kgU�qsaOfZ���r��R�#S�;4�e����|N�@�φf�y@F�e����M�]mv�o.��1� V��5QXv�Ö�;��]~�7��/�X��;b�⠰^67�D�.$�x��}T0�Y>^^�-��.�r�	,Y���M7"�����a7Ep�Dl*S\G�!�H\w6�2[&����x�6G�f8{�}Hp�G�C��GY=/Y�=�^�h�6��������c��u�TR?����aFE���[ &��e��a��z�wO+�
�B�k:�<B��]@�~����nlx���g��Ǎ���kd���bM�������?~�߿�o߾���Z���K�+b��|Y��I]�l����9�;�,�'K��4�Zڤ��Qgc�LK��; ��fo,4@^;�J�ح+<��i���b�9�0!yH^`ܙ���<���s���a�3��c�= c�G���G�����H��d+% �ۙw��b\Kg>�B-Qf(�Ed���ʋ��\�k�iU���'�F�2b& ۙ��19�8;�hT�G vz�^����ߤ�|%��9-������v� �O���L �y'S�O��~�+���%�����!s)�4x�'��v��;9�rl{_~���1\��V�1���j��쥝��(� �PFa�5�{¡�
~�i�P�g������d�s��<�Y>є��E�)�Vq��xU� �č�qP�XRF�O5�d����yZ�������y�K�\O��^7П�{�'�5i:��6�cd:2j��� ȼ H��$HàkiŬOK�Dg��d���C�e��Gy�9��k�ɨ�-���s�|ը��r��|��?��ى>�%U�_�|%��$���X�C\M��A������@sd��c�{�cM��3�p-y-7���_��_�`c��.�AE���ق�Rfr�!�X�"=���
"�������o~#��^�����ם+�;wHo:fr�ѱ����yF�"}�لU� ��E�Y=�wJ6M)���)�x��gz?�m����h}�,2�m3�YkY��*�^�)���y����[1�hc�> �c�Ք���2c�ܫ��� ,�Y+�@vi�1kȖXpq��[=�3v�"��l����>3:��/-��@M� �b�0�\���Q�Gv7��q �R
���(�ISL9�Q�*�: a(�K����3d0-B����_J����@b�	M{�7Վ����!!	��>�����������ol�_Zѱ��Iㇰ�e6�.��d��n�Ȟ_��i�L"F|���aJ:���7b��"���(m$`��/OLϐ�	r��sM�V30K��W��:˒1p�왐5ƒט��!��ڵ��������?�L=�
S]��9��KXp ��ʏ܍��<vV2��缴&���t4���Klz����79?P4/�\��-�
Y)������k�ir5bB���j��zޯΏ���'��[�"��Z���Y����輣-����[H�� ̲Y��	Y�`�R�U�`�\ٜ\N����)(h5�33�Xu��`6 &�p �� �A�##Ф�������/{���$��)�Wtg7{�'�t��@}���;kU�,f��j�Vn	Q3s���iU��g������H���%��O"]k�#27k��Y��:�:ב����u���ݨ 
یB+�qS��br}Q�� w����5����;ո|�7��N�a>&x�V��_ �A�2 Ud���5x�XGj���c`�B�S���d#��1�9�{�Yޗ������A?`�Ʉ��;{��s��!^ýIy�5xR�y�32�e� A��}��,(Ӏ�uV�ЍS3ZŦ2��ڸ=��ʎY	@�^���&Q�lE\��g���ǗXC<�����&4�Ⱥ�涑B٢l1{�q�&��Ǆ�)�q(���(����gř�yM��T�t1��6R�r��72=���2g�q�p�7� Ci�������w	��N>/�3ʲ}������=�H�<��B�B�/{�:{��-H�7Ԙ�FJ�m�y���M��o�t�Ź�u�j����4#	�:׊�!d+�nP����b���F����^�k2�m뙲&"+!؊�8� FUKPg+���DQ�m�@�Q@�X�Z�(�-0�
Ĺ��p��,�f�B�@pչ� 2ɞ=�:�E�`��ƌ}>�������^#�2�2S	'����6��xͬ�b����#{Z �<ZɃ�r��Ӷ��5Ŵ��c�`O�N�C�@��e�^��'?LwD08Ym�T~&�M�H���ک����W
�>_~V'��c�*�=�/jM2�Շ��껑×|&h�.6�*ٶ�V����F�!���2 I�c��U��R�Ӝ��� �a��)�}6�Y� �4
M
�C��z�{� ���Z@�Ղ�r;x��gk��td�ɝ��W����iGnt]yyޅӳ�� ���2g,��?FK��q�Dl�cm��oc;)[��}��6��0� -�� ;[� A �wGI^���~����w���7g�!� J9���3��$2�~�����ɉ��������$�w.3$x|�ӓ����l��q9%�|�4��ݒ¨l�.3�Uv�`ϡ�!���D�סi��c<8������ڰ7 n��y��j3��XKK-bRsh����;�= W��W�姄Aw>#X�.�4� �HQ35��Qe��((���iƪ�J4`�#�����wv�$�B�׃#���o2�η�^�k���L���������I�®R �s�Q�kբ5r��E�;ytî�H� '��zD�)3�ȿxU����_W��-�Vr�	۵�@�=o���g�H	�2�]Q1�2�	PRs�dB�x;��6�YEr|ܰ ��\]!��G%��a)����w�p�u)�.� �~�Q"�g0Zfy꒽E�{�?��g`�����Jd���ĬQԪ&� �}�
P����wz��<dK����5�j��?e����o qZ��� K��2�o����d ���f4�%�i�������Z�k/;��R��l���ԯX��M�>"�`�Uc��umݳ�Ek���R*�����u+�xx�J�Ը��@��ӧUK������~�eN���5 `)ėS��s�*/Y�� �5�S���uɲ���b>.f�b /�L=ή�Df������i�^3F��uT!S��yW���V~�؍��� �C��kݵE"�Q���%�ߑ��y�Iy\q�"���4���qM^>�YmL����$��;�mP���TB]q/�Df�r��ʜ�!(ɢ�t�kogwl���L��2���R @֬y�Q6�0vm�p��}C�#S��٣�s9D�E�����%��oi�3&�_s�S�ٚ�d��O��V>EŪ]�h��=���k��v[�<ĉ-��Xw��YCUܧ�]O����u}�Q.?~"�	2)g�/巿�3���dMsd��Enl2F�P1��ϴ�l���<�yn��_��pj����%�d��F�-��& ��f="(��]=2^���A�b�nt��B�z�_O>���Z�I��@g�f�K���b,�a#pg�?��Zׂ�r�Or�ֿ�������o���md���(���;ѽw|��8Bx26
�� ~��o]�(s�>�{p$�g6� ,�h��m�	�\)���%�k��5��bh�+�4h��#�
e/C7ӝ}Ya�1d_l�2f��M�������U��K���h�%#D�8f��E��@nW�ǥ��	]�c���;ty���6���]����1��c�����ma�Әu񎃑�t�:�hu�}>�������7�_�q9S�C��a�M��z��es��C���L��uEr)K�)��������3}��Q�;�����@��� ����ʢo,������}���mH�W~(��nWx��i�lps�FΩ�� �tn>�Ò�)���w�э<���2��Q���B��"v6h$+�IW�x{�	&�V���.��Zk������2.���Ά�W�#�D���!_�Ot�V��U��ԑ�Nܲ1�n�X���#ć�;�Rgb��#�,m��>����5�*��4���lD�yk��N��P�0t���$1[���t���r��c ����5�U�^�2rg³e���!�|�x�O��h�d����0Ǟm��lAD�(w��H�A��r��)����#YYD".
y��פ��o�� J���]�,��8 궉55d�蔤)c��c��ʜf�R�)&��Od��Fd��c	3Y�E59bf��)�MP*�ߋ�3���M�4�2����(������I%��%a�vD{�iM��몵��7�	f�,K���e���� !�\?ȊN�����c��V��k̻�4��)K�]� hz�e<�!@
�V�6p��>I �;��2e�����=5[�q?Yg��Z�}	�:@3㏷r���]}f�	�P�������jǙુr�#,��8N:y����!?g�C,5�~�AaV�:��y�~�-$�_���(*��7R�-���4��b�z/H�E� ���`���ώS:�Ŝ������x�Lk�x�X`m�n�������|��+ٝ�ZCиZ0sE%.�(Ggr���I�.j|�z������+"ή�����[���.l���4��ג�4�N�f�+Ol�΃'̠4����ή��Wz�G���
���J"��OG%c�`�3� B�f)~SR,#Eb�H�7+���2t������X���vU����Mv9� ۓOd$m\8ҍ�C	��E��/_r�:y\lm6Ҡ��$뱊BWðb'���z1���h΄�*m��(=������S���E�ot�<�Ti�Z��
R�j���r6}�*;Ȉ&��+,����Z��8O@�!2�q���^1@X�Er�o�<(��Ԕ�w��9]��2n���<�d@��x�ɴ��T[~j�+��A�l�!y��џ3郜_��ˎ/K�t}�0�<6�`5ժ3R�K^��P����ы]4B&2&]�un5Z������ڌQ�s���C;"a�"���xI�K\�ԍ�I�|��O]�j�W�e%t-Q�,��6�RQ�M���ߕϖ۽�}'N���I� ��k2��3�K��Qzή4ιu��d{��g粸���Ǿ;�j���8���[絑�m"�G��4k���!�j�8���\����=�ו�c{�=��g�K�w^�������2E"�G$מqȱʣ�d l�|���!���~���V��T$W�ў�O�ʞ����n���:��0�FF�Ul��O���
��J= �|��rq�b@��H-�k'�@ �BIG3�^�egY�pu_  ���r�G�w��F�;̂^�<�5�CtƁ�ӚD��������ͳ}�s�V]�]��<�eB*f��3���i���Y��}�<���;�sy����F}�,e�|����<�05:W�晠�� )�M�,:�/�W��	�	*�	x;��|���[d|"X�k��5f�&���q�j�T�m��T\�(�{��'��\������M�$7�41s "�:y5��3;O;O������vW��b7��UWf��`�gf�@dUQ� �"2���>���2����O�C�x6۶��-�丳/��B��#d �y{i���������ً't|x� �w"�b���6lK�����J�Y�K��.f��]�_sȤ$߲�)�/�3 �,��|�����rZ�.fY���Xc"���PG��兯�ޚ:������c�k�&?%�3NZ;N�Q뵊጑{pשj4bV�7���Ԡ�,W�</��.*;m��j'=	"hs�r/+�8J2سؚ��۱|ΑoD�Ѡ|�i�`�فU��N�N���v���8����%��r�.�b��9Ib�y�<W�_����@��/t�,�7�gz8�i ��ZD�0���4��<ؔ~�Sw����;�zH$&ZT��� �	Ƥ!8�+H�l���`)���k�����V��x'��sM_E��N�	w�LQ!��8w�����V*��-Jh.V᜕�7¼�6?��TǀA��E�����6�%E2W#r5��' � �<��ժ0_g_���a˼j�jo�Dj`pU�;Ir��#����dD�-���R�C�l�~�~�Aت��4X�����/{qA.��I�e���P��$WS��<��S` ̏TB[��l&0
^��[&e�l���7&	�%m�*(~��؄L
TF�!doӑ���!j�F��>���B]�s1�3���i�Q���%G&���x^�5K2vU��8��v�g:�
��M�N��q@� �ť��x�o��T;,�z�0�{����M�:���w���]<�v��R�t��!(� ud�젪�FC� "��ts����3�� ;V��	���UA�Dg7�o5i���8P�|��ӓ&�aՁX�8}��}6Z����9��@{9��)��QФZ I����T��M��Hh�����p����b�k�=�9p��|����4���j��Lr'��Bx�LK��+G��yL��k�=Ēqn;�ע��zD2e�7�W�5r����g�9�T�Gr$��R}_�槺���nuUPެ�Q��)���x6�i�������/��sN)T鎥P�e"���b8�g�}� �f�7��#6��N{9k�O��J�:�K�������㸢�E�5���ؠW�N��� B��b�ti��ӧ�����:�XZk_|��n�׃-Q؈̶���od�2�O5����ꎓ[�Ya '�|��J
�԰�O�)��N���^r�=����Ex/�ų����0�].
�6�(���;9i])������$9
y�����N��M:Αp��s{=��_�������$�ۿ��޿�_�F@��/'�/�!��� �w{�F�N(���E�R��64# v�-�E�ջFc��'�-�ㄭ�X`;is�v&� $�(%��e�g��uè�i' ��`¨ތH;�Ht� (�'��ɩ�Rt$�Ks)f͠�ZL$m�C`�k���cj�&"�� ��P�I��v�����?<4|h4ox�U�x����%H��A&E}@b@s0b���pj���zT)��H�M��M��La0P8��vG����s5��K��e@&�^�'[WHTaO(��\�1�H���LY@�$�|6��,�kfQ�2� خP!N՘�Jy�3�);[�� ��C���(����tGd%��-D�HNg�j����a�#��¤!E��g3y{�F57(�LX��ǉ/;����`"�e��RǕ|�Ϧ��y�T
�c2���*�O�� sksiL=�"��ޯ9�9;���}r-���&R�^sv�Ö�#KA���&���,U�&U�UQ��`3��&f;ܥ��8m�-m�,��RfIBݏ�1 �/�j`=�����a v�G%@@��<f��i��p_��
�WΦ���A�j�0�(a!��砗̩@۬i�kP�v�Y��	���8&;	��Һ�%9Aw�ɞ�ۆ��Jtd��� �m���`u.�t��	���L���i+��Yx�t��맷�O���G�{窽�8?.�N�<}.�[l�.I�+ҙ����+= ޾{��^5[ۇ	��Jg5����6v��`�#�^������v>�A|J ���]��T���5蟌jG��7�D���^���I>r��E͡�*Ƀ�MJe��D��q3�ȎAYV9���_}-��YD9Z~:���!� �ӿf��0s�ҍ��^щ�s8�q^��,'V.�mx8Z�����"�A���+I]��g9EHZHa+as�߇{��xU#�U"�krW����@������k&���qD�Sռo��9��I%TJ�T5���80+�Ӆ4CMD8��T� ���0 )�`rʭ����7Tz��Q��AH����
"#��`Z��Ò�%\+Z����} #����h��f1���0�xv"�Th�S�����
�XRၘQ��f*Щ�d8&
�<g|~��;x-2��H�̘ʕؠ l��l�Q��k6�Y�^P�Ëہ5�7��,�cY�xg��څ�D��٠ ��@qM�^��C:g����Q���� ����E7t��{�wxC"��:�$e�������ܣ����jfZ&e(�������d�7��!lke̊0��28�)�l����S���ͻ�n��/�)��mV�K�I���x{e��7�B V�iH�����mv��'<�	�eMp��N�ά�&˔�<�#Et��(K{�!/�Рj��Fh���j�B��4���$i^ޟ=J/?{A��� xF˪'C�R�j��#xf�C�]�}8�c�ȼ2��!��X��6�~��[�0����5�����w�O������38�}�B��������:.��(���_�o!����gH�m�g
�,��u�W�����_�W_}&�����NG�C���o�=���N��r�~&2��p�����@��w��[}����8��e�6�l�$w$GQ`;y�`��u�(���&�QW�y�.����,��UL�jn�����R$7��ŧ����B|/�u���&�;s�(ݬ�d��/���^~��}1�d�x�����-t��ۧ�\FE4�(u/�������bc���3���O.3{O��_��\����Ы_�	�a9�����R[`����	n�C��M>ھ�8xBH'Qs0�zv]ģ�76����8K�y�`�����{P�|��[�%���,4W%9�A`�
+�A�Ĩ���$�/�N����Ww�E��w U��+�7.?Tjo,-Sh���@3@�0�Qaj��&����V��h+R�O��S��* �y���S0#ڞYɲ�IR���6G �����bm�󫁇���A���L��0��!��Az����H!��"��j���c -PeR���IR�^�s�В>��"�1 �}��j6��C�d@ Fi�d�3����4�A�!N��L �4������Z��#w C �q*�԰c�=\��V3��f:����}6�ǚ�r�2�NY& Lج���3�b�R?���Hm!g�ET��~_���<���s����Lk�];��&�E�u2k[��nfb&Ru1��J����`����m�x]j�ۑ�ΎS`��Ӊ����o�����߿���^�2?���<������5����Mp�N!�>�t��|��0�T���G]Cc���,��;ݽ�_��~��;z���8N���c~��9=�~j�k2�G� �4� #��Ӊ�I�uد%�DH���.b��Z���~��z��ZV���9iXM`-���kKQHjs���%}��`װ*Pl���s2�5Y|�Q�K9wn�C�p��A���Lߜa�^q���f��M�����V`1}rT�ͤi�xIl���(@Ɇ���H�� ���?y�B�^~��&p�h�.�#�e���a��.[-�YD"��ϖǏc���#�D5%��0>�Q��D�~��}�͗����(����$N�d��;2_�-�	����i�t�]*�fi���#��I=��ݝ�SY���c�p�@��#�Mc�1���f1�(RTET ��ǴI��an�Ül�j��f��3J&��b�su����I�B|�@_�D�7`��������+j�.�`m���x�9!�Um����|j��H`�!��8Ѻ
���g�@Z�Ӝ�B��{[ǉ9F� 3��a�kL�l.kAX8)X�[f�
&?;�`��xY_@	���l^V ���Щ`��;�tq��.����3���k���3)���4������X�yl�3(�I���!�ٳ])�}�գ�	f-�r�z�uhL�T�����ݥd	
R��BZaԩ�r=��B�u)f�)��M�P�p�)kC�aɾ�6(8D{mV��66ּ����Ԡ�c \E'�B�T�[,�
섧j}�)v���G� j�'v��$����?�\m���6	��|A��;2�;Lg���}10<�	N���1V�Rq{h:��1�t>��� )����N4/UVO��8�8�T�A�Ҧ��p.	�%���)�����:M4�5���̦�h�Mf�z�f����K�pX�E��Z@�&��tV�~}/�\�Zb�GC;	�`�[3��jj��o�f6�n��$��adP�·Q�Y�.V�<�ƥ��Ѳ\iX,���k�8p�Z������7�#��wَF�ؕV�h/ ��+օ
��E������^�����>)/6��E�g�_;3��aw{��sd��Aw��b����B΃�r>+���O�ѓgO������/wt���%��zVW9-Id�A�(T:y���W��D����$6/��J�sb�˯��w߉��]��������_�v=�7��E<�X��l N�2��O��W�պ���p�B����kg�.!�/{@Ip?��ɍ�����P�&�$�R�eϰ ��0�/�8��ٿ5Q}�$�c��ɃpB*��UPP$,r ���ߚSʙ�]�#}���S���l��kΧZ#�p��������8�J�jd�0p3�ݓ{-�C����L��䓶�3�5�͓S�<�XT:^� H�t���[�-��g,�<�?Q��0Y*�U#Z`!b5 &�qS��3����l�wPIo���l` Jq�o8i{�� �8�U�*�cS+R��eeY��$>�t���!Q������u�\5W髄%(�c�-�AB7j�A���p�!���}Qu8�4�j5�$�R;���l]������ B�ͬ�T���H�u<�1��*=��3�8%��fhR�B�w_"�bi���Ym��,q,y8J�Q�B�8%,�[�����ś���0��Er��f�[��򮠝A��4H���������3�_�&�,��ܪ�}�RC�p�G6D�3M?�6t_��U(h�����R��d�f��1��@�W~,ɣ8<����e|��VT����r%0�Dex�DT{�p'���b�����
m_�._EU������&IqV>x�ΰŅ6H�WkJ!M�;�4�����C�-�рK���ى��>J^�3'Hf4x��)����-X؞���O���/���K�� 
R.'@�:�DV�ж�\���q����,����eI{yrHNQ��?��~����?Q}��`CQ���T������T�S$ȲhF�Xaq츜�^���~}�=���?���70��.m���h�q��� @��s���we6q;$QkT	�W�#rp�2�� �$DG�[#4S�P���@^.�Т,��ܕ��)p�j�ae�U�S�@UU2��$.F���K���Ōc�h6^�.͹f�H���R�h�91F�p `?aCT	����Ų�X��nAmu 㐯�>&S�2��t�T2�4r@X�����|���I� ��.�`B��f�=��8sG;���,B�4q4I���G�*�XN�� &;	t������5 g£�B͘�!������%J���b�VL:�\���-~�c�`�*�ϖX����zFj0W�)�9�M[W��<���D:9Od9P�>��1�w���l�D�Z��F�1��a3!��<7Cݨ���,H�g+��Y�f�e{�uhL�c����i�W����ܲ�~"9e�i2a;'�(��3�6���0>!�w
����b�c���Sp�T`�AmުB �e��j{NQ�"��28M�'�3(�)Ƌ ��y��y[�Ci4���08�"p4L�0Z��+	�zus%���ő�9{��Xi�t��>x�fRt�Jw�e��R0k^p���t#�E� ������K���[fC2�m��d��2=,[��8��Y���l�d=����� f�9OK���n/�k5nN�Xn���Չ|�Cj��4`�=S��_��
��x�g�̼�g�J��׿���fY��7q<�W�� l���P��q��ޒ�KjUdQ�SN>���������ǿ��^��J)��������������}�=[��cWt��:{'�����?�[%�@�0��4K�Kw��:�D��E��-F��ⴰ+�Q�r)��
U-�[]R��7���-o=�ʬEb0*�����h3�� "�Qԭ�/]� ���l/��,���{})��d�1ԃ�� � �ah�̈}�I�ιF�|L���ݺ�viH��Q0�����ּ�2] k:%���N�����5����>�ִB2.t��K�[Q�( eE/(� ��Q��9j��(}g#�KT��&ݢ��k�9�vem���h�i7�6���n��z[�vWf'�`[��$U�7�8=�I���h9�,��](,�` [,B�+���A�d1�f���m���F ��P��\�� �,h) � Fq�$��BC�<��=g͊A��$��������$t��mia:�Ty¼�����ھҔ9y�8�ä��l�̃�_֎����C�Nt���o�ӻ��$��:3�x�>��H�Y�i�J)k-��i!o��פ����'��M���b�b�1foYp;�%��0�B�+��{1=@c��)GK:�L �ʅ��&�?,	�Z������`�/����Z���T�b/6��aG���;&\5'����+�$�*�h� ����|�bLۤC���hi�$Id��نb-��y,"��!5H0T4����n9��v������U��ò�^>F��|��H��^9 �JÔ�1B�F(G:���$2�h�{��MwD�����[	�!����ǻ;z��O�l/�q�,���^x����D���D�Y��͸�	Z�k�HH�ىr��
��Nqf�Ӽ��M��ߧ����D b�[)�Q���?w'�� ���1#%Hi�(U��i�T"��� �`+V���]$"P1���!��i3�^C�����������[�@r+�[�]�-����5Х���w:��O�b��]��W��� ƙ�u� �2$#�4�c�u�N,���P�����<W���Z��џW�����nM�Z����_�Av�Fos{��Js�?��S�͋�� �rAɉܡ¾�`�Z�p�gU��;�H��Q��=P����I�����t�fsV!;�L��3"��at[�՜^�}qO��(N�����Ьq�$������ǉ�8q�QK�Ց� ]�K�s����{��	������!%`|0O���0(1�T�ű�q�X^'�3)@`U��(Y7���TICs��������F�}�^�)�B�it:D ��l�YU����9Bd0!�+b�m$�xm�ø'n?Ri��ݛ�r���W����S]�����Q�`*G�։�k�Pt�s+������|�t.�q"�=�MՃnW3��-���c ����@�>���7�nr� ���%4~MC#Jߵ�:ٜZI�+��q��v��*���$��#^�$�q�MR�_rgu�H��ԫ�Z�dX����j�Xi�'�,D��ӧTP&�K�޽��גjp}4<�$�j��n��`@�vt��
5%IgA�C�P��b٤����b�'/��_�x�h��@6�	�WBUmI���TsP)%�au�(�]ƺ�)P�!?Ic��%�xs��_ �*j�Y�!�x�S�3^���:H��(�4�M��s�3�P"���qA��B帢
0�5���.�C�郍B��\g�4~���@%�Ayip�X�!�P\͈��X��F��y@�2�1�Mƽ�����5�8A�*��k��W����њ����,a�d;̙��[���j�"� h�C��������W��1)�4��n��'��~��H�Or�v#(���h�l�}�4*����)�sx�`�z��Mb�iKɼ6ٓ�J�xq�:���@�o8�ba�ɣ��Ѥ~�ꖜ�UspJ��A��q�qM%�*���X�@q�����CO���u���o��q,��w߈��~_�[�m��r@���xr�v�z�p�&0]w�r���(;X�:�����r2}¡bo	|�g8H��߂�m���d}����	��)^,U�Iʨ8� ��*}�3�W+++�WWv���f���&��ATz��a��q�Ȣ֏ �z���t����&�����#���Wm�!�pJI�2B̰��^W��0H �YO7��W�Z) Q�E�� ���O�|��@,rm��bjR��̖KSſ���������aI�jAS6dwWV���+N&1���z�(luHI�A�($iu�g 	�#��lQ5� ��"����i{B-�
�`�u�$�7|�� *K4���8��8���X[5��j)|4,t��6 @_�` �5�7֪���R ��d����5��������>b��{	������-∕�e�יp�h�l�IE���7��.���)?G~ Ҿ�1Nx��N3=�+���`/��L��%Hm��o����f�:�(�ҹ��^��|0�kC����R�'�j�������X3z!��o���'��*����rЛ�m�M��eiX�ٌ��+�OS4�c)�=�`r���JǬ�]Hasċ�ЩYS�-%���t�lTϥqf
���I\"�XO�UU�ɪ�!��R�am���l�7�����j7�X( <kb����>����H��Ir ��J�V��C����ǘ�H��x신��/� �+��^ʂ�VK9=; @0 *=ɉ��������䇀v�ǾXm��*���Ԍ��!Q��#�U�XBZq����F%oM5/�G�W��o�cE4K��φ��a�;�O�$01��2���?����$�[n�]�z�(_�4T���؞�Õmd5�(��YS,���x@�A�ެ�����']�TP�
�+�ޕ7�{�I�,��_~Eww���;��u��}F_���B���?Ѽ�-{e+������B��9y�����!���_�[�*t֐�׌�ť�^|j �H,"�{�d2�������.�,���}Yj��AU8���ݗ�F	pU��
c��4�M ���&�%d:㖊� !��k7�P�[**_j�*�ь�\�qPG����A���5�Oû�B-�c	��=��z:$�ddE�5xwj@�bF�8@D˵U����b� ��>e�d���ȁLb2��P�{���,�{$י�j�].��qg�P��U<;]���\[����SnJ��0|L	l�)>h[^[���,,�GJ7g%�n�M5U���<��(�� �������l�T���M��L�*�����D��ż�!�����a�-����i�Y�LT^�8Nq d�-3� 'r%!�X��괁|�mSZ�~"ܘ�Zr�η���Sq|� i,�;���H���'��R7v\Xx�ì1Ύb�V-o)Y:.%_������צ�-k&̄�5IWB�<���\��F����v�+����c�:������U�+ ��k�w\u�[dU9�{F��iɚ)�v�q�T*�Z��[�r4��u�{����1�-�9��+�����6Z@c'�%��8S�܀_;KD���@~2��wa8��KV�lF��dga�u���>�8i�[��'[�I��E�͛�~��������W�{O���D9~���W_���s�s�Bۺ����.�)6��Z��P�h�f�Z��b�!+�yH�Ę,��fBj��Z)q�v��}nN�i�0�\pri�Z{�|�c�,R7���j�R-��%�굚'��7��=r��s:;���+��T���&�a>ze�%${ K
<j�U�!f��x[5~w1�
�Vb<��CE��I$��Ġ˪�\/)�����Zh`~�!���#�6K텽�N(�((!���� ��C�L	;����c����m��Qc��r�;ԍ�KSS� �q���ۧX�e��P��`\�lT[^%�q�2���;;��l�CA�����`�Z�V	 �k&� '[d�[:l�������+H�f��0�`�l��*M+d�ɵ:*�l.���&Ci�����Gt  X+��	lV$���ǉ�9H7��T�4\�ʬ�F�jV��H�T]))�P���$���0P55��&���8�B@7�9j
>V�H���QI�z Xl�g�������+;��U��9�&�B��+�r��PO����]���
j�M���,ɭ��*��a@i���)�
��]O��r�m�8�a!Jմ��{�U� Vܙ7�y`w���N���NiY���ㄉl�3~bL�@��@���]��Y���Z ��3���?�Kn]ƈ��>yrK�����+f5��d.F�&y� �hQ�2�4���`��1�0~��q,�~1��0�"z~�U������R��%=\��*hB��<�FE�1���;���*���eR/W�b����� �f��6#}JX�	IuU�m}Asj�38 �^��-�"�q�!pAF���c;Y\6��AB���o���5T�Z�\���܎���@d4�um�C#� �-�H76��z����jk� �]L�kc������Ђ�-�V#7ه6ѿb���~��f&F�lD�~{����4�����B=L6VM��ZJ��@kX5�JK�~���]�9�$6v��`6����<�tCZQ-�X���<$�j�h�S R�������Ɉ=��*mz�쉔����������5*\��h&$C�� ���)�&Y[���Y:�U$���%�	b�/>��'�����i�[.b�#�xn��~5�U�>�QiQ���]��Җ9��O_� G����u���;��9�"��#W�@��5����(9Ϧ�܄E�����YT�2w���6�XGT�>d궋/ۛ�(����êS h@�D3c����{��AoM-@@q%�˃�$*�ܢ8i���I��+���;yi�+��v<r�բ����k�*1��!WX1��@i�Q��k�\>E��;N����In�Y"���8��RS|8ء��00R��>3�Fy�z�R�/6r�'`�7BC�нRl����T��|��Ԏ�.�i�c�:��`�%�i;�^~�6�tGbr%����}v���`�9��U�U0����8a��t-�R�܋�����ĥظ� �Ьnj7]���/�-��D�MO�(���B����BƷ�Pd╥J-���YZs����SH[J���������`H��W�WVs���ǩ}>�MtTK�L�-�Ǵ�]�eC]�v���Ad�\�4��_���a�?š$3��ޝK7O�I�/�[�Nhk1'#~�Φ6�`8���1kңx���}��6V�`� �.����>CG@�p�Җ�}Ȋ��%d?[�3��ȻY�1Gsc�$�@���I����P��؞j0�~�0/��7�E��� ��;Iْ`{Nա����A�j�WF��ԭ��@D������GI8��_��ŝ���k죿6i��p�=��I�L2)k���6f6� LL<O���L�ֹM��p�.�,Ӿ�d�?�=����%['�����{�h��)���1�D�.�%���L��e��$:Y��Be����H'n������*q�]N9��r/��r���$�f D'm��ռ��p�"t�t���y��l�U�rJdC��tbS�"8ME��l��F1��i�9�4�� �Iަ>� ##�U�&�����ˌ��䀅ܳ/��[�96����$a!��4HUz����z�WfH��!�iYN�k�V��nT�XQ�%'�2�0\nB���ڣ�4��n�1F۝@<$DR����3s~��C����G1�P3&�D�U�Ge	���`�-��7>��$龻Gc�6k5��s�ܼ��5�)C��m��0����~b����c�5@�ǯYuA��Zپ֚�%:)��֕޶qH���7:ť�Ŭ�ǽ�+�Kg�� T����C[|0F��V�G�ZMb����,����9%��>�$�%�sw�q��?pT37�|�	���7�3c��[$�ϕ��%҂�ٲH��l�V5��N�JVp�:MCQ)��x�����ȹ���C�m0�����W��E�V���l����I�Q��s���B���J���ү�����I�s~N$��fN���(�ռ���lbl\i�m���W�0�:I@s�b�	� ���t�u��X�v(m�سk��Zo��4�lß�O=�A��y��s)��ײ���t5���2�,�=���'�/��x*�EQ��o	1x��¬Ķr:��S���Q�!0T��橷���D챚��� ����Ϊ9)��)c�� ��Ĉr� ������D�HSC�1mܒ�u�ާ�4���՗*��a�2Pt"�1�7�X��J�œ�!�B���5�������o�(OE�)����u��!bPQ6%h��QM��~�̍4���7/"C����Z5r�P3u3����K�x�0�PR�n�����[�R����&���Ur/|9� v�J8��N��J��t{���4��1��l�$b~������~��Eo[��*��6fz^�kK@��
�n��cI�zz����ƥ�֭$��pFA��+��XםZ��3�J��ď�����NM��uM�TO�F!X@q
:-`3�F�K��W# �vK�&>�\w0� ������1s�~7qE~�l+	Id!�}��X���Y�K9�/|�p8, �^�ϧ��?O4_E(S�{ʼ"͛����
���^��@S��5K��I
 l2	��N�"�}�@;&���~�7d!�5q���*���ݚט�^�x�L�pĮ���1����V�����G1+��v]�Ӭ��8!(�͒07$ �+���n�i�,��;L��{�I�Ԉ��j�M�����E:t'����7�8i�c ����'�8%ЯJD8�v�����������$	�v0�$;^J�����VqohG�5H0����6d5��U�؆�`/u�I)�u�ޯ�ۃDfh���������'ԣ`�.i,1nD�܂)\`��>Gi|c�F��Ѝ�PK�����4Ot_���m�np���E絕\D�3���1W����+Y�������&A�1��G��~ �|�>��l�|�`�_ZI��Tj�E�c0cL�$u�C�
�ll�Y1�}��恬��������'�C�US;W�jřo���b��K��@����m��aZ�]�e���+J�k��Jy�Y�.]#,���k�?�{C�����j���s����,�a��N�0KO���@��?����Q�tZ>�h��Y8��y��!F��~������4��I�<[=���e�6z�+�jj�I��gIWx�~��l�]M�88y`$�8rG����\���p�ԧ�d�~��/�I��1� ��E�x6���x*r��r�[v琞�mW�Dg��?�����PIԙ�O�J�l�P<�3$�tKb !'� ��|�~*�w��G��cg�a# 5�-�4S�4Ƣ0�o���'�]1Z�����Q֔�mУf��q:���W���\�6���GR/���r�.�	�_;����n�tk�&�b�ۈHl���U�*䌧Z�;�M~2Ds�i#�"�ab싗�*us@ry9T��M�#��ǆ��%>_ ��W��KZ�X7�Sk�\����Gݨ�`��9��K�Y�[�l�C+Mt)Zޓ`����=<�^�\�%�l@_c���e�´�a-e�ݾ_������uss��%ݓ�C�\I�!��3�	_4��sM���%٣{m��l}�w�^?X�6 �Ľ: k���*�.����^c<3 ��NM��o��".1���J$&<*�{8�����'*�D�Áv�{���,p�*���7���bf�$�պ�ڠg#����-���P\� �1�E�N	 L�%�����&ֆ��Ƽe5A�6�v_ԝ�_;�J�˨#�I�W��j�IQP#��M�=��bQH�������2w_JL~�h�6�����O��!�x�ӄD�E��|/���D��I�j�4�ސR���,�Y=z0���s��`��~F"�,G��u��S2&%�L����A��j��٬޸�c>���ڿ}�e�	"ނ����_���~�k��R)�u��������{�H�D�_�5��8��ewCZJ{z��,�^�O�M.����n�a6�/1%�Y]+iD���@ێ���dn�Ӛ%|�����o9�G^;������]hlil	\�1��X�k����@���k��l�/ss��+��h����5��.�1�����,��t��[!i��7ZH�S����bo����&������.Ӹ�g�:��.�=X7ZY8�� �N�3�[% �<��@�Q���4n�ṇ��8gzww���1��L�zb�2�"8����ٺ�K�8�.�������<{��p|�Uǹ��z`��Ý�d�%�B�ɀ���:�%ߦd���$�j�mڈj��(�=�(�U>���պ�D��q�d��Mtig�Y@J���L4��I���E�������1�O餳67E�¨՗��t��F�s�L������vb���Q"����f��X+���-�_+a[~Q�"��9�3^[ꮯ��2�"�����	�:#�	�6�
�Gm26����ݪ��V�6�,��ރ�����`i5���^�\�D	'` �T��U���"%�Y��j���-��<]K�������-�����,�ؾ�����<���\l��I�ق�5�د��j|7�x��k�`۫�mĻqT�t�JS����� kkޢ���]/��~pnе�z�k}��:��/�o����[j��@Ÿ��:�E� 3��L�|y
��.s�Q:�B����=���(���㱲������\���w�뎞ގ���̀������^�I9�����	��#�i'٘��	H����5��  �~� '�W:ivg����	��Q���ql�v�:��;L��f�g������%�+����:[��=�ik(϶!s���'��fh�)�¬~#�&h@h���n�瓢\����8ב~��}�������UR��<�ڠ��#)�^uX�EA8�&��XͷH��p�&HI��G���}����{�QZ��w�����Jo�>(��T�DnHI����������_jC���	�1Q��� Q���y���(�RnG��8�͗��$:��j�-���4�ɍ���;���xf��}��B��������|�-���nշu�����H��l���XJIsp�=[�ؾ�՟���],�z4׻�!��Km�-�_?�F���`��1�k ��s���Z݀�|0O�A�K�Ǭ�[1Ν��{�q�7�Z�o���۲4L�fZ4�ь�Lb���Xe0���ݵx����[������L�zX��R���o�1���Sb�q,_)����Ѹ�hO��K�9��� �{{h>H\0J���Jr7�pv8
O�]�/��PR���9*�e�^��ϟS7k��[b9�4:�$Hr��
�d�!��iW��$�n��Yc����aز��%�y��na�9���-f�A�N�\H�ʶ_�����|G���{QCC$�%E�ΑH�ě�Y#zw����X�TKx<���ڂhª��h�Z�z��H���������0�0�߷ʱG.�ն�]��/�b���G���KlC�۷�$Y�q�x�{Z�2������.����V\�$F�*,QC� լ�m�Y�7�?�u���b8�k����`>x&����2~��F*+���?���)�ڞ~wr��v �X�����)�M��*y�����!�HX���ԅ[�n6�o��#��^�-�[���oT�����үv/��*<k�wSVh�Z�Sw���W�F�wrO�1p�T�|g�s����C�-�)���P�zV���6�%�q
'F:�_�k	���O��������l��'R��;���^�t<Kڧa���u�:s�B���o�j�9+��Tcǒ��%Z�r�O�O
���pb5� ˓�i5[��/}���TKտ"Cڎ�v�J�w1Sf��
J�V�d$��Y: �0@���f�>�be�xZP&�+GNG� ]F�Ot���"��BB�bnZ�Qnl'��f�7��L��ƪY�c�ׯ�����������#�v����r-��&����	,�v󋵗$���w]��#�&r�(����A�3q�m冡���y/�v��=T��Fm�e�e���Z: Ѓ��&0����][R�ͭ��"�4��7W7�7.���O4�]��T�V�K7���ފ�Pk?�f������0�h�����)��&��w}:�!��Xv̱_ݶ��i��W㗹C�ܶ7�
������S�ȏ:lPbJ	����#{�(�^�w��k�,[�æ��x=�ծB�x��|��*º"�i'@��v�Ź�$��8���_�E��JMy�^pد��SJ#r�=��� ��T�	��c]`�]R5�H�HBM�2���7g~>sb���;v����q8�x�3�ގ�/��{��>��O��v\x�J������ۅ����5K�n��g�=�f͂��<&K�L�5�N"���R�k�8C�e���ի�,̅����>.�[��x!��\��- ��i�xGT�~\w���o��+��f�N��I8 C�S�����h<(�s|����OJ���ҁ�p�&�v�6y^5e��1����u��x�8O�~��|>�۷����H��������_,�]P핼�ݵ �3{tL����r�
�P� $�Y�0n�=���"��V�#F��1��P���26	`b6 C	��V`�"I]��6���^�d��n��- {þ/ ��;49�#�� ,�z��R�Z�!�\����Ȓ�f>�d)��f�޷�z�RiΥ��l�lz�������-	�����۰�,��I巒V����L�!�G�έi����Ee��K}Z�!><V���>J2�sMb��v���Jsܽ��ܨ�?|n�tcoo�Mu"։�O��5(%����-����!�/J���'��%��m�2����y�:�������Z�&"A! �4?4�!�N8�~G�~��_��gODj�_^�N��9Yx�����̙�ʋw�{H��4��ܶ�<���j�D 4�d�09�L�E�T�9l�rjb;!2�:�l7c}��Xh�<��-��?��Nq���8�*[�ݼ8_�<���Qn��'��`L���, f�i�j�~v���\K�J�]a|� ���ۣ��fz��qV�9�ԇ���������O�_^����׷�]&�x�4�����:��R@���kA�����~IDޛ��V���=w���1.���w��OMؤ��M�@P�e�M�:����B�llp��i�[��7��w]�;BDv5�I[CU�V��ޘ��?��4�nKS��khNZ|>�a	�0�����͏��%]�ZK{��~3�jϥ�ׯ�~�|z{�ϯ����>T���y<�ZR��V�2j��Զ|��[�I�t�S�h�Wi�[Izi=�J���ƣ�۾���f���O4ચ,��dd�E�w~��M�G�/n��_��pc}�')�0�����NCQL�N��|�ѫ�_Ӌ�����d�93C5��A2����P��|/Ұ��^���'4\])�3�5[�5�b�N\Ɓf�űHc�b[����N���JU{' yS���H��$$�[�ubA�Rް`�q�
W���{$x�hqN�G�2�Y����d�TʼI�^lT����%IC�=��l���IU30�4k�Ӣq��8��R�$��I�k�j 'M����PD�Y�2+@d��ĢF�tx�vVm�=��_�ҟ�������|9���,x�f���8z� ��N'�.Ϲ�$Ő4t �Q�c̒�=K�j>Ɂ���!o+�SAT������pP�|��%qa��t�Ѡ���A�[�{��b]����3�D�;&����~�:�I���i�pBC�oz�R��=�✆�E�I7śP���j��\�	\��h�m�.��~-���Aci��d�es']馡Q��{Zf�q���4������ъ��X��V̓��y�� 9KV+Nk��KG���W_XoJ��0v��;�cj��v�v��{Z�� �܎����n��D'�f�4��>��)
m�}]/��%�{хԀ����6 y�ά�`G2q
�jܓ:g4��]��q�o��#]s(��r`7�[�q.�I!�iq�>5�9��pϠfl��PJ�ޔ9���~<���A�B;�-8<{=J��n�a�}ȱLծ��m���	\`�1&*�シ�q܋�$K�D"��;�FlG>1NN��E0?��AB�%n��҃zZ�w�n��J$i��IP5��R���;�us� ǥ���%�`�Ӭ�g���;U�&1����F��9��r����Y����w���|O?��f�+�y�v�O�A��"��륝���n*�	��|�(��pb��
�R���*�h�D�@{~�j!T\�]16#�)�M3��oh%��	�0T/�ZIfJq�LM��0��{ܟW�fd��rj�H�MuKi,���T{8\X���{�V��)eu�,��z�s����P�X�?�-`Դ��h	��0ޒ \:�g�n��B[�?*[�o����@�{4���j�[3��)�?��K������d�`��m0��?�6����+�vv�H��ȴ�vb��4�r��7W�UQ��ߙ�~D;u��&o&��AUCՐ��x�K�蠛�߽6�P��175��j�o2�ڇ���a��锊��y�yR_H.; 30��Z ɓ�/{Z����t|O7�#]￤'��8* c@�%6I�-���~������L�k���h�8��n\*6[&� {Z9�~��
`R ���j�̚��b ���p[]l�6!.���b-k��}�ܾ,���^p����u+6b����9u�#�w��UU�+
��t1��zz	�/;� Tד�2:�#��qgO�'�~A���W״���t��e�e]���5!��Ig��&������]����{a,��>Uz�����������w���o���D�5��gʾ�YNA��C�s���f�`a���Lg��p�������)_Ӗ���KK��$�1ݤ_�C"�ا�
tS�	X��K��s��'�QG�0�>���`��&��8.|�W;U��$Q�J����'l�ڦ��k ���PxX�?Vc�C[g��=�N�ü�`.3�v���������j�|�3ͽ=�ٺ'U����iu]Ry?<��J�����47�KJ����K��b�a������۞�R�4ёP�S7� ����|h!�;^��i?�:=�Ôl�(��Uћ�=7�	�ã��Ć@������2�\��ѵl�!�����ɢh��:K��q��:��:�{�@���*K�~~�+��ԗ_���D����غQ)#)0�0L�
Z��{'����ow��~������٪{�g��0P���9ڀ��Y#�[���~HNx-1�>\���f����7ؤ�Z�v,�a�� �Qg_/��"d�
7��<{���qA�Z�ҙ�{�n����׸Z�$���,��3{�}�0����b������{������z��=y�tA����4=�fF��L؍�(w[ߒ~s���A����x:ʊd��^�����3��O�.�kA�{�A�v_�k� 6 �K`V�S�f�\
f�<�'�,���F��iS`#Ue�A?dIh�N ��I��+����\����@f�+�
z��Ji�J/m����$��`�,���L�9p�����h|�j��a��@��$ �TDN-���}�87|Hv_�t�&(�j��M���	ںo�h>��g��צt+����_*�`^��?vm٩�g�E�ڼ��~ͷ�4e�� R?�ף��h�Ǐ�>_����U
��W��s����qzb�䛛v:��4%Փn�\�j��ﭔ*�j�JIU���^����~x���̋��HH��Q�81�&����/|��q�|��+zw�������zwE7�O�;h�t�`�$��*�q[{�z1 ��k�;0��$����3>5{��{]@<f�\�|�+�ب�d��������W�lߦ�Y�{�~��w��T���]�$��#��V@��Ie0#Fg���5��c� L��O��l���OL9��3BF�I���$�^ �Y�I\E�����lx�^���EO	�,�.x����j Rr9Mҷw����O�П��w�뷯��/�� �|Ց_�Z>{6����V��g�[�|7�k���y�m�t���@ _��)�}R�. ��ۊN�؆�Fu��+Z��!~��<�@$U��)lpb��R�v�������^��?

Z0��h�H8��~�g���3�4��H ɹ����������1^�wL��=�����{6���֏����i�M��,a��A�m�)�gJ�C�oK��u��ɪ��f�����v8S	뵽�XZ�}�DKw��%x^�jkax��mH-���~G��z��G�*
������F}?�3�
����ѫk�!��68wh�f��uW�N�2T4W��x�k�-=����r���JԜS���@_2�Cx�ςd��1>�u��n��(ۈ��3�@?�rG��gz������>{~KOn���$I�r�Y����av�Q�i�+(��Z%�|����R)�F�Ici
���x����o��lV0�Μ��rNc��'	-T�� ̥���Q�a�Ș���o�ю���L����N��P̳������؈�r9
2=- L��ޛ��K:(�`���֖� L���Uƀ��:@������=�{�Z�	X�	��:���e���]/���%邖	���ǃ�ivc��G���/������������^b���d��z��v7Oi\yv�~��l^R��E�O��ͫm[c��>��g�w�!�g�@���:#�a;I>OJ"�K��j�n\��F_4B�����`?'ZM��d)bH��k�jH� ��&�d�g�<�j�F�ӷ� X*-S�?[h�bB�;�����KgCR���_��C:G	�)��Мv�"�q�a=��	��ħ{�s̹hP��  ��IDATU���N����4�;=Y��n�}�-�����	ܶ#ҏ���Gm[|�8�m$L�v���TEa��U��F��6J�=�%u�%YF�����=\�1��Ʃ����k���Yn#�W�w=l�����i/��(��66�=��>*�,N����Ǒp`��������7+�BH�j���gSeFaNu�^F[��T_cR�8���k�a&�e5��M�ʗ���� j�Rg��`kl�b����J�aV�=Kî8��Y�V @��.@�\�������������k���_�W�����y���������$�8(P�����,Z�Z��)���tP�1���#�n�{�,c���U�uM��i�}�,9��ٜ�Tpu��xhw��DW`@���[ د�,,���@�߽ ���K�(�U<X��{r+�U*���y>��%4V9:I���v�;'�i 2����lQ��s�(�OUb�@�:Px!��j�Z�]��h�!-��� �eԝx+@���{�����O��?�����:������'�X=��F�_=oH��Xz֝:b��-�xY���VD��e��
�\��G�����(�	Y�K�T�|�(ͷ  `�^�P�4�O�q��?o�nA4����9E?�+wrI�ߟ����,�i#9�+w���Uk�km�B���\�^i{���Q�Z#�m�Z����g����1�U�}&z	,�4��3����p��Sӛ���+��/����u���姿{�F���5^�Oe$H�׌�l�~5L-�����Z�2څ���vk���l�R�[�,�_-�����QDܦ�@�jH���Ȏ`6;����5���zi��� =��z.!b4�1�p�Z� ��־ݹԞٗ
ފ���$߮B�D3�b��:_	H�`��R[��?���W����H��D�����gz��v���,�Z��(�y*��̆K�IY���f��\�b��6�ɀ�i���U}i��<���i�d�O��������fs$�i�^V��}wG�^�  l�����_�zǱ�Nt~xO��z�K��ݠg��|���0�=I���T�pm6�/H�b��Dg� `� �9yTdY�#��/�s���a� fA�����k����`��tX+��i'��r���o������ͻ:�;$��SQ?��Փ�_^������ª@DیC�-��o����
`�g��!tk��m6�
۠`�Dȼ^u`kG��@��O���Ww���
AjC�>�㒍�%;��Zn&�k���d�	Q2Y�V�W_4�<�62$e�,�k(A?ʆ�y��g�]���cݾO����g/�iϠV�L�n�V^��c�ٲ5���ԯ鏵�rF��}��hϑӁ���%3�K�o����T>z�}��~��ZiƱV_{�k|�_M���ގr�Z�c�����Yn��� �$Q~���ѝ�rT�>j4���o	����+��������� _��,)����v`)��i���QŨ~�l���$�F��>������_�Ͽ��?|�9����{JO�\��El��DJ�]�˜���|T�B�5ި��"5�'5R`�C�	x����,fC�gB���0fN1Na���'��t�� �������oN�����g�0=�q:�-��;��������y/h��p4=,?��&ޫ�j�r\sή�䂐������@T��d�@*�?@A1�
q+D�dbV�x=,�8r�w��y`ߊ䋍�i�U/���l- ld ���k5�� r'��z^�p�`��|�
���c�:��o�vxZ[=Aĉ,K�J�ɦ���+D�8=ĵ��W۴u�	 ��|���ڃ�\T���G�������+�3� ���SZM][���ݴ��o?��+��s�J����8A�Xm���z���^F���W��_��h]��y�a��������^��u	T�Ǡ���v�J�UQ�1�O-��lZ�}�C�ό:��<6�^�(�N����A�/���o��&(�=2[�FE]�hs����`̻�������	Z�� �|d{}�Syϕ���:���50R����R=rPUӴ�����+���`�1�}*i#�*�da�Ŧ�C5\�DI�8l7%pm�8al�t��@�wr����~��������[�� |������qTA΋��l#>0�9CP��^�6YR�N�,q����0��YABm2�^͹@� ;�U�����������YVV��?���Á�߳-;���p�����޿}-��l8π�ɓ�쳗���Kz���R�2X�ú�VC����aQZ�
ƕ!���DN!X.E��Jl���Ε�=��6N#'�`i�n9��ai�O��a]?��3}�����������G��[S7��=/�q؉+}�V����kR���F{X�� �f�K�3���T#m_�㚑l�ql�d��Ȅ=����M2!{�?6�-�II��1��4r5,�)���w���!���r+��x�yKD��������4�s�e�sm?h=�vC^���D�ɴ-�hS%�7"�6Y�][R.g	e���ؼ����X��)���%C�-��/򞬫G�s6�->�.�H�$l���d�C$C[�<�$e�@�G�x�x���81�(���@�6���je���!5m��Զ9����o҈�"��sz�$0���ڶ)Qƃ��&�V��BP�š����ߥ4�ذ��ec�|9&	|AL��)�<4Y2��W�P�϶t�A�������x������r�_�������=����/�, �9�|������^<#wtu���UW�QCR�ڡ	q��ҿ�r��͵���N��� �?�c&�&A���HܱݨX@$_��u��Z���P>Ntf�PR���|�_��z��W:��5�0N�7�r�Y���b'v0�A@V�lq��>|c��k�Y#��;K��TA�9^	uuhE�1��=[&��X��q�sM��{�����w��?���Ͽ���_��{�%��]��`���������� ��4�������7_c��i+>$6�.>��&}�ݑwj���E�`�P" ��m1Z�{:i������yϠ}���t݉z7:�&��_�������o��X7"��d�U���ZI�|��<��7+��~��`�6n���@�&2c_��/�����E���3���RQ~�������� OƝ��P�Ps?��e��?ƶ$_[�o][�����&H��,����o��,l��m���oH?*rY��<Εߧi�m�?��J�0� )��O*x5��ڋ�~�1�af���l�̖ɞ�CZ�Dzq�X`���Uh�k���`|B�3Xw����3���$���Vvƛ�D�糄�8��-`k�7��ӳ_����wt{}C��������%v�NT���Հ�g�PA����Z�l�ZT���>��3&�s�W��-���q2��K�8L�ҏ�w�O�f�.�r�\�v�@�1���$,?gg�*���/@�<�!<s��T�`0�G"��ڬ+`� ��^�1��g2�fൠ��2�zB�;��p��EG�%S�N*Ve�����駟�������?�Z��� F��aAͷW�CN�u'�k�b��F�_ 8�Otu֠�n/ ��;vj`���=e��S:�a���Apv92�l[^�kʱs����M�(����ʛK�#���@꒤�g% i~�a�u��G!>�_����^�:�:Q/&��t]+'�[�7w���y�1��o��u�[���+�aK�1�fu٧\��K�L������z��Z��H�n[��X����l��I�.}�۱��>^z���m�W?�c�f���[��P BP$�O�7����T>�U��N�I�0��'$�
�$�"��q~,@Y-���Q7ny�|�$���Uۥ|�B;T�N}��.��Y��[x*㉙��Y^�x'���]��:$i�NtX�=�=�O?�I
�B�w�����$�vI��b�j_�~,�BU04����t�^h�xp\?�cyƝJ�v;M�-Y{��FE��c0*���`���*����i��y�޾{;���r2Kv&'�r�(R6	���0_����-C��R�p��FX�W{	������$�f0���#�x�b��� �z��_�ի���J��~-��v��Dr</��8*�b�F�IU$��"5��Ćs,���Ic�ل(�	�՟pUJ֮U_إ�W��.���qM�e F�^H㪿�����ZՒ�|����#ĺ]�`4��\E���oO豙�>��1�t�?��#utEx�o�Ӻ+���'[�]ۿ:c����|����&_������{�c\+��J��9��G��\Z�G�����܅�G����WjM���x�����*�}�ېl87���aZeՃ����Ǯ�P���Qi|�;���h��7`m�^	�d^��s��6�/D-$���]�>��R'���o-�f��*���"��V�{JV��W�X�_����A��~paB�l��!�Vn˜ؒ�c������-@l���:.���8�8i<�򽄴�VUN���~Z@�$`N5jGr�������%�R���/}i,�Ɏ\�:�ܮq�Y��:M�� &��4�	����2�m�r� 66����]=o�
�y8}��[���A��p���S�L3���f�wK<,���Kҗ��׍��p8Ed'�=�)a�[R�z�����p'�p\ $�ǋ�m�n�_�N$l{Z����k�<����'"�b/HN5�t[l���B���o��b)M,��ۄ�T1���!5�9��G5�V�Ƒ��U� Mt:[����ʰj�y���ɲH>d�0��=3��{�Pb*'�M�ա�K'�K�Grp�h}�B1݃���yj��@Al.�ej�u�uu�Wc.��C��Pɖ�D�Q���o>Gv��^�ѳ�{0�ͯ�J'�8O��O�4�z��̀{v�tq�|����0�}�a��BJ�gۥ�% l����n��t]RC��/�-���j渧����=Ϋ�s9�Fy9��mЏ�X��1�VS��Ki��COJ�XS���dhփQ�m��̀��1�!�i uS'_x�Z+�<�hl��BԖ�
P̵x���zۃ�����DNV��\ ������,���N�?t:����$��c�J4��Z��% ���hʕ�G�N)}TmX�8g� ��<����K�Mɚa�]m�J��-8c%V�
ɣʞ�l�v}#x�����)AF�%t����kɵt�K�t�ދX�x���;+ �&��`c��+��XY����1���Xd��p�,:���H�P� SP" �j�2����]��ͭ�.�ܿq�Aa���}Wn� �z&�_�f�%_��Ug)%}�6 ?I��,|���I#6UKEp�j�U�h�za���g	!bPH� �*�
y��w� ��>�2�V�b���N�=�ߢ����X��Ɔټ��%�	[`��u��L��1�<�^�3���-�ߺ����1���g�/k����Z6����X㝤�n�[�����cQt���t?�%P�r��<���HXa��YǚA�̜:��岚{k�[0B��!�.?���c�[�q[�^{�4�µ�����L���{�5��Z� ����H��B-~ݢ�m���+�X=�MbD0(Q���فm`5��'5I�d�?G�j�حJ���d�.��6_8엒vv"o��h�$5g�v�j�����&�9:6a��*L~J>K��A "׆�\bl_f�W��8 ��g�9��$�3bF�H��,��*��$o5�*��˵d������`3�~.γ�ǳ����x":�!:G�-t<�4���M8k� xF
���X�d��4�=߰�t���2�bϵ �QC`hN���ª#�K�fú�Ǳ���9bٸ�c��|�D;�+gf��yNW����P�%��H��ɞQZFC�&kǀ�#؈�-�낔S�ƒ�հp �JI�@Wɘ�b�/�:���c@�vT؋߶N�����;$t�������@�${��7�S/�#����:c����T��h�t�A�~�銂�Q�|�#�A���I�?�"�7]�8,WR�������X��YW���R{7������^W�ѽ��8~�S�ǀ��>������z?���.����v��~<��@�%)�O��
>i}�j��� ��d�TK$�"�,����2�:�5�CNk¹���yD��a�88-�'p��؉U�-�f��1/[������p��N�{1��2��A!�spZ奅4(���[s؝ϖH[%q���Oe�ɓl=� `�� ���PGkI4>�s�$���qZ��FL�*ۯ/�" �4�8sŕ���u8-`ly�`��$~����"h~aQQi�`Xl�Η��םE�����{:V���Su ��$p̂��PN�"[��"够������#�i����?�d�i�EN�\;�զ���s�`��ƅ�\��fg(H��I���+:g>��D�E*�<`\l$JH\��6�5���5a+�s��D�K����v�� �+�Bj͟� �ю�)��D5?bG��ت�����m���=�s˪k�W��a0��	��Ճ��.(�ڊ�h�WP����}����h�V���B믞!nH6늯��\}j�O�|߷��)o�<Z��m�TG��&�j���dN���t�����^x��hP���Ȑ)���\n����d��n������ǬC�Ľ͠�C�]�5��T�uj�#;7ey�'�FZ��}Î�d��Nm�b�z?�[�����G�7�"{4��Z6q�����L S��ʠ�1��ZL=*�fq&�����(F���aO�7X���SBhp
ĥia�0{~�ޞl�u������ۛ59�$ibj� �<��ꮞ����>P��������B�{�gz��23" �����T��<�g�*dD ��v��~zھ�Iϔf<��f�å��zb�b��V��M�T�)�:�9~b@Ï�&A�|�7W��8���:�a!X�����Z<]�
�� �I�n�Ez��#i2P����$�������果d��W����x�&zOS�>t�H.q;(�C�`�jA�[�.R��j'����ʂ8/P���:2S0�q � UK6�X���|sx�U�{�����c�j��5�Z��-���{%�(���9��3+A�����-,�.9�n�p�2���>>������%k�gH�޵�-��r�e" b!�� �����D�|Q��i��O��/yѿϡ���[�ˠ��럿p�v�/{�)+���k֯�ܽW�UF~]|��A{�U�y�H��:T�{?Nw�/����q���%���B�_��-�]��G��`#������\�1Q/��Y���UL(`Q�;�Dn�ue���j`��i��brێd�~���bg��[�ɔ~��m��d�K�����iY��^��p#p̳D=&����t����g�EOO��Do�+5b���f�8P��jy��(�'d�N6�E�%��Uc����� �N�i��;���ր=l���>X�0ə���&G-�A��vǍ5��@X��i%.�S��'&\>�ݔ�c��%-`X����l�5�>�bU��~^>%}1,��L����e�VvYj���ݔ�"��A�m)`?��m�1�h���$�Y����X���9Ĳj����7�ex|�ՉuK@���ͧ�cd� L�b��2V䣶^��A���
.�P+�{�E�#�\b�
q��/xe���C�
��?��Z��in/xd?�xu��B�w�!�U6�Ww�"�92�;m�w<�R�m���,��5+��[ǎ9&g,�ח�8|�5
͘����$E���u��Q Vi3�X�����t�v��kn���m_��t]s��k�	��\����ק�,1��^A+���^ џ<7����,n���|7���u�v{�n(y3~�u��c_��^1��w/?7g<
`$l� ����U>r�[� �����j��Y�l@���p*޺�=Y �^ ʒֆ��)�JtN�'Sc���
�&���nd��qs�r�,���jȀ�*�;x�Vޔ-�ҟa��N���O�)�pU��Pl��5L��O�����
��q�5�u� l�@m�ȭIp�t���V��d�21�tF\u�z���:}xz��g*,d	�p�՚M��a��Q�4�4M��\bB��H�D�,�AI�f�G2�T�����7���L��o�� �RRbu�!A���p	*�b|� �sOg��E�#9�b�)�Z�5���b����H�Qj�-f4�Ez���_%0���y"���w�M������kA���Sh��k�/�Ύ�~�ұ�$8 ��}���ψi�����Fc ���Q7���'��g�v�%ּ$��*�4V�Qv$3}o1-Ƌ/26������{Y@�/\���2/b쉒���%)�� �gY���]���.�/Ǔ�)���u�y�x��U{m>.Z� ��	��Y?v�K�]�l�������l���͒�as;�E����ة8P؎� UbW�����K� ��>����[<L:�����{�;UH�x%�k����щ�>p��P����#�=ZX����u�]���H��Y���La���+x��Ÿء����Z�D�����e��u��p�Q��B`(��>W�~�*0,� ������߃}f�d�3��3����̱�����bPĠ���jth�S
�eA���B�������m��L��7C��`��}`"���Ǫ�Ue����(P6� ��f�@���Y��*m����}ǍȦ6x[r��(�R���� P�A����X'&P�+b��kY`O���u�z�������W�Zp�Œ��FjD�����[�w�}is��ɶ��:ZM��>u���e��E`�پڀ4 ��2W����^2�kZ.�����5%\j1�RI�|مB9!�/��̅��5-�饨����Z҄���,h/�SBt���
�ϋe���q9�-ۏL;�j,5ߛ��Zt���m�\�B?��R_.�/��&�-'����}��˼KA�s���\CIm@}�������N!ppsA8������l~���>�793;�s؄|Y��/9t��`������|<Ϡ�����vJw~��-_��e�Å���V��yi �z ��9+��q��"W�#�N':����s������۷o��A,0#[{gv-��he���֑�$W���#6�+�n���& �����RR�G�T�Ca�!�j� �|O��0��|E*(p��Q�'gT�FjZ)�y��z��^�D���j9�j�W�g��ϵLw��R{"�21�����>K�ԅ�63> s8W1�=<<4�pCǧY\��Y�3rv��ܰ��)�?*�!Z�f@6W��U_��+ˎ�8�ُV��>+83R&I�&5;h6�R}�L���2C�U#+ eb.fU��8b���^X��8w����r"��������ny�o����B4���YD%׳��J�n�x,��4t�l�S�2������k��}=�{����o�!K�We�YS�zA�0�7�Z�mv��b�['qē��V%0�%BX!�kS!> _$�!�f��=��a!�z�$k5�SͥLv�eo�)h-I"$0T�j��M b���s� Bl	�6�&�31g��B���g��~]�K�G���8��S��Z<2�%đ�|}?_�	�x����k{"w���������zj��޿}�9hc�e�)d����	�6���w�ݘ�O��M����jMjM�_`a=�+bY�v%u5��<w
��Z �4�p�f��7y���M�ۧ���UV���2n�Y��ea\�qܱ���2���>����_�����1L���k����~E#��������/{�h���cНy>�/ª��z�_�l�4W�>��)����}R��C� z��j��R�B,' F�V����V�+�D���Ha��W+ؒ�N����y�K[�Q�f�W��qAR;��q̤p6B{s�R	`�)��g+I4�&	^
;��d�Y`��.e���o�$(��ip&���^ؘ�%j�%�(zL�6+f*�p�`�pӭ��u��G]�"UІ��+�5���( 1��Y�&x�����>�h�����{z~�'z��F�|���@��n�nnha;�,��z�G��q�Lk�_������/L��G�	�W0$C�%/�;	�K�����A���/���MC5}��A���,aQ5F���3L�8%�����~��l����&ᇱ{��&��Q�#�OIV]�2�����"v�b*iZ+伏���2�|*��ZT?m��k����jgI��c���>N�s_�|���\Wl*k�]�'
��p�f����]�y��t`(��9�ղo�"����t�9J���%�bQ�s!�.o�h+X��c/W�Ӧ����j�Mǭ`UM�&�;ZN����M�_�޵�*˞֧���iX���Yy�z���f�GPq���_�xrB�2�wn7ym��n>�=T�(z�f�Vw�ظRӲ(�S�����6�����y�X��b[A~^U�\Wu��h��E��ġ�E�d�� K�֗�k����$U�W�[���`�|�\�P"�be����}�q)-U�%�0PA���1���J���)�L�c�˖�EWL�5xd�x v-& M�����J�؄j�H����<���}O?���K`l	{ܵN�����gd�d�gvs�X0�^�rt�;�^��b�H�]��_���赍�pf���w�8 ���W�~�ml�L�v���F�8,���AFZ7޽�QK|�8�w̾8�P9��P|�lǱ����E���a���!��v�^[9R���5�X�.=���6�!�?�U�rx��<�^��KϽo$J�N�z��Z�/k�ℾ�\�L;hzBm���{	<ޓ�^�/��(�?���=@o��3��Jn����k��ח(n�s_�\���s�0��{�Y�$����V�~%9_���@s��禼�Lo_����>Ot{w�3S�O��=	�x��\�X��7K�X�5��=!5�-��S ��nM�'��*%T{1M��=��o;��V7�"z�(�����qJQ��+�)��^)K�W�-����i(u���8w�P#�׆`�z�rF"�s`� �����'W-� F�T����W
��-��l�_����v~����C�|U+W��=�K�Hkkоy�vG!�%a�n\�-ڮ���Rn�.��1/-�7�)�wlݒ��F�v<����ؗ5>g��*?W��TJ@o_��~����.Aז_}��%���%��~!���	� �[-�)�@�Z������y����@�j�u3=}]��%��K��W0��[	�u]�������ߏ��~N��GY��L�DM��W����������7�h�wmʺ�p�.���_S}���d��ǵ��K&}�7�"h��6�bM?)	��p�� �r���ʌ�
�.��ݡi��t+A��|��3��u��AAs��������}�ru�����'����O��K����Q��-���U��`P��Fe�����}{sh��8h����F�@���,:����֫[~���{I�����y��^��CH�q��������?���.��c5�\m�8;c���aO#�[�&Ƙ���?1��e�Ŀ�U����"�0~�C�9�ʪ���g�J���`�J@��X,� �T|n6KD�`jjw�p��b��� O�#A_�3����Bp{��Ԯ�66�Ĭ��Q�SN��p��[��K�-2��]�X^���{�mü}�������v�-q��}�g���CC}�יP���-�J��OS��n���>ŷ^z},���+34h�ؿ:�`0,;��C�����#.�����g�.i#���QO�#���y�1� �����N�����@"��Z2�ݮbP�I��傍R��ڽ�ϫ�s[�ܤk�8�՘h�et��%�_�'C�w�?�(,϶z��R�f�k�o��\����-��Ƹ.�/��V�m?�?sk��\���f�?K����4�l�����\��˧�un��~��#���_������{ė�3�ŏNG�Vܷ��v  n�6Q|��"�4�ohjreyb�}#]gۼ(Q�%����ާ1%OԖǢ���/�b�o;�C)��y��H� ��Οeܬ�:��vY|WS3xxG�˳�����eY�mz^�X���3���]S:�d��C�އMI�N#��Q��1���!��,�OW��UQ͞�j�ԊQ��JF?A�=�����S�%�i�p%)`%0נ�|p(
]�|͐%�uz|ʟ�$P��atDD*�`�����Qݽ�N��|t� o�q�̡�[�L�OX���;�f�\�%~�ӯ
��
��Lk������_C�j�	<��ԇ��Â91ꞿ��^��yu�7�]t>�d}�x�X��t��:�� �Wh u��hwF^��x������_��9X6���1ve�Jj�� ��VHܛ��,� �(�=��%���J(�Cv�\s�m�o3��f��^&��K����` ��,��F�8�"�p_���,���F��C�\nram?�� �/y}��l㓽5�M~��*yz�w���E���~���]B�8-K,?C_���yY���<�K)�4J�|�ܠm;Q�*�q�Һ.�:%�����NJ�En���R��&W�R����|կ��-f�{>���^���� ��r�>k6eCIu�8��-�Vg�����A��Tkf�5�S(��N���ĢF�r"�x/��9��Pm�� �*�W�n ��k��I�a�pWh5>����y�#��^��KQ�VA�u#V\�\��č�.8��
����|��8��͵�w����#=��m��'��q_�TR�0f	��*1�,buV_�^З��3�j -o��OzeM�X�Y���b�h��{��t�zIU����Lـ��`���[;�����7�s����<̒6��)����U제)L�9�}g�[!Jճ�J\ܱ)wW^J+kB����2�kb��֢uq�ƺ�r��gp���c"����tm\�����������KJM�k=-���j
ە�?��&�b�\��r�Q�M��S���;��l��Bc/z>?�r�oJ��Kb/�]�����zl��V�D�s �s�!���������?=��d6�ǵ��9�{9�y�'?9�2+�������
�D�֞N��
��Z��Sw�;o�	�Y�}'��`����v�/����������K�w�R�F;�o��5(S��D�"b�:��k��9��{R?�k
�`ŁJ,��p�sU����+R�s�ʥҵe7��iC�B��m}�_QH.�U[����oy�8|z�S.������[:��p��k��tj��A?�x^�N�0/�z!Ⳓ����/DM.x](�s�ߟ����L0#�y�<����ʓ����/õ��kq��Zj�� �Xॎ�t��a0Ь�+xo*v��Z�����X�l���'�L�uT���� �>�5��k.�ܿ�o>�J�}�����&��<�����?%k\<t	�n��o����l�k�q_�#��u2������ �4��z��]��-_�-^
rj]�������X���N�
 �O�����E	����X8�X>��$�i�[�X���癤�@Z����h_��U����R��)�絽�N$Ao�Q�S��EY�y���K��U=�[�Kfp�� ����JO
�[���d�J���{zMC{�	6�
�N��nU�5�>xx%(��0Ĥm�Z%��[��Ֆ�;"�����q����~[���bȥx_��be+�3�J�]����^e�}����X͂g�2�����؊�z�����%�p3�M��x��ؿ����
(n]��l����$��ݫ7z$��y>��a���;)����,���Y3�]��\���e>�\�6�[�v������_W�?n	�eJ���e�e�]�e����6��<X8�ī|��=k�T���c��H�G��sR��$2�#��?����Fз����B	@��ك��w��4��9̅�#%����4���{^"^�-�e:���+��e\׶�3N��E�o=9A���X��-z�?�|O��dLE�U�펮z�T�wsu�6
��$�(������v)A�5���V�����+yI|_���?^_d��u�����0D�S��ĥjZ5��p�{	�g>�Y����9�����hh����0 cY"�|fY�J����D�ޑx���^k��,z����~*%�i����i �� p���,�."�5�J��Wο�*{�a���a�#���e����l+��EӔ�f�bz��yւ�l&6�>s���I��:!��씙d�2�;6E��X<�e�!��Lx����N��;���f�"ȏ-�w*8d���q�� ���^ }�ۙ�z:I�>p��gv�����vp���x&�[)>����)���ܣ�I��6g��LN��k���르��@X�C��Ŵ$�S��!5j��r�*�Gzs�������#2⼲��4�mDed�O�){Qo�~��hX����Y�E�������?��/���<�4�<��Y�g�o+��W��~�8��-:g� !��1�'�U#����"(<�r�7��y�?*_���;�iXJ����=-޲��Ε1w�e��NdI\�V�/�'�x�Tp;Rz�:��tr�'����w��Tzr�w%]GPH;�J�H4d�X\6��X� ׈���ZEb���nv`Rl}h�dU%�,���.�*os�æu}u�D�<�^�đf���0!�D�\�9��"�5�c�w���a��"�-_�R�-l@�ԿJ�\�$�e>����#�g��j�r��>�@)C�\]h���8/g�b������Y�h�K)����tHV�.�P� !C�_���u�W�� ���Q���H<��eweٹ���ל������5>3�zl�vW�ewc�8�q�.ғ�k[��7��Ͷ`��&)�iI�u��&�Ų���ne =$��K��P�K`����������^ʊ��NoM��n�gF��%�7�#J�d�d-qhe>��Y��432��j�B��6N�%�*ИE�w-u4�3��|�gf[%!^��l~�LE�
���6{Y�Q��[P6Df�mt�6]��߽.L3��W^�n�������u�0W���vS�g�^r`�6��rxi]*zq#v�nί�Ӽk|��e��%@�7(�CY@���W�b?̫���=N�h����	@x��<���������P�rt�L�*�a��O�)O��u�k�U���ԛe�������]ނ�ݬ��`Fݜ�L��]p�w�˼9�b�f�+�ST7���x�\\�]vt,1u���K�w�2�XqU���J���`Rb�<�A5
�dU9�f�긫��u�bV2��O)����uE�V�����xL�`^%_TS�W1��� ��&�aU6X\D��.rd��eB"���7����|[���K5��0.�Vɋ�qAY�ś�z�c_3�ħ���VMw^�	��7���}Rا�r�%h�5}�����ʵ�>��d�{;������������	f�꺢\���4���h�E�
ȃlj �uE�J�Ӑ����N�Yd�<o�,�|.G���$0OĚwn�����λ�ֽv�+�7����_�P�^��ڗ�(�>��S� 5�X	�R�~���� �-i,X}L��b�V�S�g�c�{)Ծ_��Ӫ���azP���>����-¿z����n� ���g��3��;�����MG>�~�u���b<۵�x��W�����#78����ҷ�'X�٪�`l�rG.+��/v�5�}1PS���k��
�8z�J%���Il����9ї��nǋ���g�85 2����C޾yC��߇��T�?x+��z�q�'P*�U0�������+�� ]���1�H�"�J��>�z��>a#W�>�;Ɂܒf�A�k���c�����u����&�I���[
�J��,�l�b�H�'�� =�� ��ی�V���n�9�Mn��K��C���E%�Ǡ�v�8��Śg=����*����ȱ6૕�W���� ,-.����6>�l���� �(�4�
����3����`}���;�`����вE�}�d,�@_c|},RH쳠�h�M(7�ͼ��C�k���V���3�aI�5���b�9�N�	�N�&`�� �x�>|�����|��8����=��#�P��4(4��"h�\�;M�F����q���u�ᘅ�� @�{�ߑ�l)���V�&�u#/�%����3�2�`[�$�'	@��O=jq�����G���Z1�����K��-����W��&E���ī\#0��k�o+<+��5VaݪJ�~�c%�����%B ���*��s0,Ʋ�$Q!'����n�>���M��X��m&E�((��?����jW7���e�Z�����>�D���j�5��ě��F�Ƞ�$S�9��]��y���e4O�wc~:as8Z�������U]'���!�l��'�k�A�q���`%��-jzXeGØ�(����I�E �1	��(�k=��>�[1��y�7#|Ϭ�+��(��J�L ���c+$�Ky1ԯ%.��ME^�db>/bp2�L�<�hdX���u��ܷ�I�e[f\��?�>��Z$ N�����Q�d��׬� W1;!{@(��B�L�]՘&�a���4yXp������z���L1���N�������Y�&��Gנ
վ	��[}��W�ml�c7k�׵��y9b�����d=u�	��!m_Iqu�ȯ��=t.Ú���ދ��q�o��V{v�;��>���n�&�őٌ��i��^w7'%wUwW�[CjZ[�7`�8��XX���?�u�>�������c�  }��n~�ԒF\�ꎃ���խ�zòVs�r?��M	��c
�L���8��}i�/?.�w�|}{�c����
g�(4H��]2Z2F~㊰���G�������]O�\`-�ZCue�0����e�\�p�]��� �sH܊Tv_h�P����ǜ�I��eWu�J	�2�Q,f��u���	���a�b=î`��uY)V���	��̭. ����X�oٽȉ�\��4��k�}<�ih��s����5l,&���$*	0��x��h�둡{WI)�~�JQ��aL�`yL��nۘ�+���ϊ��=o�����j�:0�vu�MX��_h�iޮ��c~Ք�zbJ�O��0D�jw��ށ�&�$ϧg��J�����S4����gi
�@���`�l����Gaq�
=��v��F�7�+���,�/�L�O�U$@��	��7�U�y�5ڌ�v� �!��4���t1�-��*�'��G�q�JV=���[��(�6�lۏj�Q�(�S���B��R���5��5�wK�����.�u����»Q6��RR�3Qn�^/y��m�L��8�Hy����u����K<*[���e�#�vp$."-��_��	@&�)���Ҷ���q�S����l�BI�zd�,�*��^ě�g�5h��?:��3Zc��Dx{��t�w�>�e�lc�z�d�k�`L�@L��"3��LV��J�c ��)�bd�h���;�Y{v�ǭ0Q�D��S��YN��o ,�ŰHd��]�:w-=/��~�� �D�[k4%�@�jqq�E�"�C�d�q�5\q�F�����>�ARX*��F\ӿ��m�����X�˗�`B�C�G�Q' ���h�׮�kӤo`Gj%]����R�$�OF�+�A(�1ڥq����p�Q},�_��np�j�CC���g�\��(Z[����Z�p�&�n]�e�����y��	0��wF_/��B@��py<y��)t��ޭ�m]��p���f!@2���,����o�ߩC���[%ָS�j�߃B���P���l����sn�߅@��r �ǳ�ǚ�_�̒�ݟ'"�k�
�us�VY�2�Z����{��^����]�<)�c�����&��;܍"'W5ZH��<tJP]C �Q��`��/�]���W��l����=X�V�qf��j�C
xv�f�D�\}9�$��m��/cx1��ӱv��B��#x��O��H^�b	�)���y��4�Y���ž`f�|��m�]/3��+^	P��q�������@�$s�|����g������|�$�]@�	�T�����+����BHD���!����D���&�$kT�(]L�@Z����8k�ۯ�� �?�j�k5K%�� b>Q�-Y��Z�� �`��XQ)�����0bZ|�:f^�q\�B��U�.����Ԧ|d�p}fJ6w �y=�� h/� �*�ݳA���3�(e�g��6��I����Z������B�gf�s#H�l��%�Ṳ��MtkOz8�~��胝JQ�X��	̱-l��㲸9=�du4��s3���X�w���:w�؅n�&� =P��*P��*+@ŭ�h�$��t_��dG�l��ْ�y4��2Y0Fs� A"��/[�zp��3X�������L�q�J��FQ�#�WL]Jj̉�B	���Sk�@��+i/�V�i~��������N��b֜�w�û�����c��Xn-��������|��@���Km�^kt�V_������bVS��$^$V�mDF��Ru���w {��n��ށ�vLn��>���L��������6�F���2kF��������A��k>��Ƙbv���"���D!S�M�h8�w=�Ed��d'
���rRZ7u,�Ү�QD@t�N�B2	,Pfc��8*���ta�����)�Y�AJ�K���[�A��y�18 ��05�lS�`���`��f�X�X:�#�ُ������+g��(�Q�E"|۰�
|1J�x��;����3Z|��g�t2�CXEjz�K��h��O�������(a:�R��V���W��Ҩ���d�ڶ�}m�xx���3�g��(P��c���kW.Yz���i�E�}�e�&���v8,{���5�V;Ķ&��C:���C�7��q7+>����T��x�n���2+K+�T6�;��Y���o ��ұ'c��z��{�bD��L��m��n��kjp�yͭe�����&�Q�������R'UJ�h{H*��{�C<k��x1�E�����d�����6�eqb|i禱�X������vɨ� ���/��ͫ�%��M=o!�#u<p�+�Dj��=x�O��L2ӕ�AE���{���|��$Ƞ��)u*��S��TC�S��;=)�� U�V�.�
bj��e�63ˢ�O/"�t�x҉���*�Ɨ�����<�c'1�8;[y��sd�G�z.M�d�~��:=�܎��ō�x�LM��&^��S���
�N�c;�z>�cw����q�G����B�S�	��58?�-��*�L�e���!����RO�7�h-c5H��U�5tmH�FYB�V6x���S^kȀ��x��w���sV2�ʦ�����eT�fb���b�?J�NI@0@��M!.�5��o�YW���`8�Y�:��_�2�w��2$�Y�\�:N������A�,dَ���L���hf��|>7z<�;@6�Ӌ��@�BJ�rk5�Z�,-su0�����y&�![��gh��/:+S�f��h<+gCb��E�b�IAo��O���kg��Z]<v�@��e����Z�����F�~���<ǭ�6aJ���V��H���t�'�/Z�ZBY�?X��؂0_�T��=�E2�PԔKi�%�=,0��+<�Ԣ���f��
�9;�oc�.�	�u�&�i�d4�L�f( nP)���݅���<L�����r5��	?^`�����������1�
�������6�uV�(�)�
�bj�0p!�(,]$y�J�h�����ȁ��^�n��ۢ\<1P�&�Jj�.&�d�p1^V�ż��*��(���Bg�
4�2��E�d?�F.�UӨ����:�f�V���W�=>ԜيY��i�ݸȳK�4���8�a7��ni��@��F�1`�� Evܬ���5��g:>��/���܄���2��ʚ�
�}�-/k�l]�R��q02��bi����3 �C&u�'�k���d&�D�
��,E|�j�3�nu�^�ˁ�DY��+�PK~w�d��(Ő�*�I��h^�f[RVs�ԏ���D��F�~�LB�^|}�Im� ��^.����6�İ��F��aR�k-���'��oP�T���ʾa� V���h�jNpqa��.8,��7�ҫ`bM�N��>fH.�q]b�|�Жm�����nȞ�J�Pk��R��d��P� dZ��j�,��Z�9)�B�Y�_�sE�N1��fuhA��@1�w�W<#ȴ �u2��ݚ6Ok�GV���6�{.�RX��Ǭ�Z�W��,JO��+���
�u�~|\��z�D�H1���9�C�5���˚_�t��}n�b}��A�2}��_J`�_
������߿���������Ӝ�k�X��䕃��g�O�l�x��dIJ�#�fc�pm	�i�J�d�����x~�H��?��a<� ����p� 	5�1��U�f��`����ĸ�,���MV�u���:l/3fY�:^g�����XC�9�.8Y�ײQ�iה6`�L�p��@��H��������\'F�& cD�Y��G)��)Z�ϊz���EP�r:��N�gl7��P9~qQ���dζa%�UƤ F|Ң���t>/z� N�_�9�V L�ډFŋ�O��a�*�,�X������q��w��д�����3i�\�������N�1f�%�h�k���n��[��`�/W������q���b��+���o���z��e���I.��a�2t;6�;6h��'@- `$9��o�g��n7>�����*1�kU�)���Y�lY0����s-�����a���|�qo"�j��Nw��R@���{��o}�=��ab�*�#y,؂�r:�箦��\O�2��*ծ�����b	�=�%�_�aѠ�=b�Ђ5���R3�v��
���N(�G�5�)Sk�4�Z,���T-� 5�\��K dV � �Pw]"=���0�N�y��[�_'�eA��Ќ��vQ@�kWeʇ`e�5qB�K��r���(��"!�l���d	J���-9�W��ߗ�.���_q�6�ت��� ��������d��~�P�� ��a%���K2~I��g8���~F���s)����5 <�x����@�vU.N�@JO埅�n!c����7:�kxB�N��d��}�F[�"�	� �5��+�ȭ�.����֊[��i���,^�j<��0�_�y\�<��v���-20~��.~ֲֳh��|Z���L�����fj� ���vl�6��ޜ
�������Q�[3��Ufޓ��.VPP��j�J��@�f���M W�g��H��n�,�(O1��-a�>Swb6������տw��_#���UɃ�M����d�eM�BP �1!az6�@���Wv��~��+����X��Wo�ɿD���QHz<Q���+�R�٬r��C�L2��ÛyYg������R+��_����
���i=�i
G���ѧQ��� ��4��'�(�E|+D^�V\o=��k9��;T;���
��~��%=A��f`�P�?H�r�B>��ј��{� ���I��5t�Y���N6���&m��VC�/|� /f�����N��W���2_'�;ңА����`:���b�)O\ރ����cw�0��B���@2 �A�̿�G�.���6v�y*b����_�"��A����A�3(]�H���!R����q���^�%�=��P<_�E[m6n�������w��x��p������u��ɜB~�\2tPRVK�0p��?c����5��-f\�� 3עd��zR�B�{�f��������H�U�X�Ϣp�\0-U�AC���=��V����Jq�cj l�_E9�2b����+�yh8j��~��];�0�Y��eVS���#-����Lg��.��r;44��21��b�s�x�y��f9Sj՟��eE�=�agC����b ��KE5�M"�a\G�P`���`�	�A$�bRH֬o" KT�G*����]A�-W[������4��J!B�����v�[ms��l�F�Qkn��^�L�@?����T6֤�x�d���}��� 9bՋ��f2��F	����3���ڦZN�&B�B����sc�*,��!�GZO���f�R�d|���(q�s�ѐ����Η�V��j�ܔ1(V�R; ��23W̖<�}M`�9����Z@vֲPq���s�(�ر�M�,s��
V��YM0���ek���b��	�O�'��e�A(�T1#���b�H��&��E3�xT�Ӿ̬���wE�ƠA�`N��`��l�D����e�d�oq�+H0��L�ٺi�	W*uQ�_&��LaQ-ju�z(�Y�G{_�(��-���Es$����{��01R�&13Y�d����Y^&���Jo\r���)���RE����×/X�q���K��'o�^�u���S;p-�8� �6o����������
�����*\%�`|@�Ivf�*﬋z$�B��uyVwb%ZZt�����a=�&C%C\��j{�<�[F� f��(@fy�ڦ�R���A**h}5�Г�^3M�����1al=��߱|=��uyl�x������Ӹ�n:�=����qb��Z�7S���޴FM����6A'E�ӡ��� �<+�۵gcz~!�ÌP��V��b۹����_��X��w�C��C%.����u'�(ﺓ�P�{��t��u�l�����es��l� @��� Vk��Ʊ��"�K�nDg��`�d-�ڭ������Ϲ~�����-��Đ6����@�\K�l��s<@���0��A���$.򁵮y"P�X\��Fbn�����6��j}i�K��~��n��坌��E�� Dn��)��]WX�֎���A�
�0n�:src�(aj'd��[c%�s�=b����1��2C_mq4�l!�\r��,�Gd��UV-�A��'j|��BB�cY���`��1�����X�-VKI-`�Nv �g8�� ��NQ���Ͻ;ʁ�F :��'��JU0�"�6�w�Ϛ�W �S����ɺZɳf%^�  �Z��H�p�r ˥(�p�˼/Җ��II����9��v~�t�?��8��/���,4э�ȹͥp�h6���#k�x�H�����60D�^��3S�=���)�Z7cٽ�#�[Lq[5�\�8�=�j�����`|�����"n�"a�x��Xę���!�Ԛ�dp��yb�5����=�� �0��ˠ+�"��a�����2���>�9�ȋEp�rj;��p�|�1csCg��K`��#ڻN��T�ٷ}qKbN���Z����O��$�.����K�NTgƖ�3�0yWRO�ƪX����ZR����%��J���`F<ie߳%T�g!����ҀX�:f��QTs峚�� abc
V#'���@�6��f���	�(��c_%}�N�|�F|!M&a�`��-�ZM�� ���z
�]���	��Vo���T�otK0�����`�LP�������)Pt,��%�X�Ǚ��Q3Y���e��'�L�l�il��P�*��eG7�M�9�q_#�:5Z?��Ƣ1��
��}kH���-���F3TQy�hy4�6��{��D��aR��e�b2G�)�TW�;S �EB/�c�D��A2�Tj�� ���%�5zQ�l���<�� ��E��&[�,�c���Z����*8Pqac�^lYs�cd���� U�UkK�]�  �#��v�	�����
/�X=�,�q�y^�p�b��h�RF�Fͫ3��5���x��p��%��ǳi�������-צd�VŤ�[]�խ쨽����^_`���|u|�%����Bj��d�Ö�J���$�8%{��X���,Q�_����S�(2ps&n�&E�_��q�ת�}�Z�r\���1u?���I�Y�O��G���]ex}xu*�N�|g�qT,<�7�����3&%p��y����d�S��$�ݎ�Bj�Ж��q�nV	ݚ(�Ir@�X�
�3��a��L1@�(�Pxn���<��b��1zB�
��b,%�X)�Z%t g��KhODZ��)���C�=#FD�093�p��D�P[��k�̉��0�����R������8(_�$$	��V�u��<#��Y�iC��%��p	�Ee!�ˎ����&�pپ�qa�F�/���}�}��/v�*C����3_1��oh;�, �
��e�@K�D�����167��#A�L�m�Q�V�QP/�V�ǌE��9
r`�ea�{ך�7��g+3�v�^2�s���6�ݎ���^��x�[躎[���wK�8�f���A��(���)�_R��e�m��g:>���{ZOg:���	4[���,�[f��F�� ��4gAX�$�繘�/�
�ցyW�j����%؛�%Y�(H����;�©f˼�4/jA����W���g�1����W1���D��n_XgY7��(����t�c�M�(zB��/�u��i�c�����l�j��!%(�W���U�-�<�P�X��&>I��	��Pj!V`� ;ًMiQK�3�ͯ�+9a��^�;2 U����I`�c�hhH��������AW��h<�I.;��RӮ"���;�L_%��g�e�>tPS�x؀#A���F����sSvN�Tq9�&�z\h���Mc·��)���K�>܍8$/�� �����(��ZLQ�͗��*o0���"�s�I���-bԒ |���Z|�3{>��vl�k0@%�W}]*=3]��-�'ط�����1e��j!H�X8>e.Z����l�ҭS��0�D��[�XPp �2��Z��y�&�q^&	�[�s���f�1���
�R�]�|�#!P?��[K�.i���5,�->FB*��������� ���-2��A��
H��T�k��:�Y/.���f���pm�����{���� ���V;`��
����d�P5 ���jZ��@��rr�hU\��0Ыۻ��� �g ��*�7'������(��h�Z��[������
��5z����o�Л￣�~���z�ȵ]��4јXA��4W��s�\�)yV� �b1;����<O�x�������9=���Dm���2d��3��*K���4i��p��>���_J� T�UM��KPL���%�!W��w��Դ���@77���������g�=�;V��莁�����Lϣ����y@�X_���;icr�]�o�O��'��5�ƨȑ��]��- wfY#�j�/>�geM�qG]SEa]S|͒�r�/�&K��p���ᆦ�^�.{><>j��tc��Pnod~��,����"�Oa�8aV�Kً�\���,��e�q�Vx�ܥuL���~�V�%��g��#`��J���j����+�s�e�,LrʿQ,�F[J���1a���>�b�a"�q{W˾���W���H��d�?K�,q�����LU2�-�>[N���v��CSJ_?ܴ�-�j���W������E[��<X��d�1�^'�iM�R�#���ʘ*S�*�;}&��ga���v=c��>лw藦��B{�j\]��$�25M� ���Β�x��ݹ�衟+\�n(B��}�x���^�B�p5�c���8���������'a�$U�d�3�uVM�4s)�c��$.S]e:�ݷvۻ�.��,�]
�U0׌"�*�uٌ}D�%r�-���z�'��gx�{���#���E�кn�٠���dE� �˯,���K_�5��	Kbu��G�$�L��(lG�Z�H|�?�1�(Q�n�6�~W���Fz}7�ׯ�0?���P]}b�M8�Ͷ��"p�Q}n��iw����W:~x��A��6�������;�Տ�ҏ��+z���4m��Ƃ�+�v����+u�45]���n,�����U���������ۣ�����L�ѫ6?��*���Z	n��i��؟���}1K�
�A�KYvAP]�X��3d��_TC6� ��}����w��1 ����΄�e��3�����i0����\ +')�(�c�o#GE���&�26[	��39ii��?C����H�ײ�Ei��$��kS��(��o0���I�����J.ӴĢpӡ���X�ZߧQ�6��M�z#�X�*B綁ֱH��c����0�X4)Q����Y�q�E�ZsKtV�%���G��=L�Nj����US�IkK
H�9 gZe��G��}P����S�(�
&w��zqC|�D�>$#������?�M�&�<@��]��]v7���]tÁ����eB:�&q�-R/Qd2[89�I�@�Fs��X&�����fl|w/����������^�~�7�_��+`\$X��E�"UE�E��23)�k �[Xm#�i׸8���10xc����x^�Gn��.Qq<���_~���?�"�.0<!cet���EL��Ot��Դ�3kN��Cƕ1Ю��h������ L�"�����`�^�Z�RI<�rY�sx�O����9���MK��tlL�6Fyl��H�ޑϱ\���M�56�@le�n�6�����*��$x�]�R��dA�����t���V ��U�t��]�<��pM?���!\c����Vl��@��;�ՙ�.�m����U��c���.Aݵ��b�>qg R�0�v ��ń ��R��0��U��[b�V
K�?�rFѾ�}� ��7���X�D;��7�f��xCmS���3PM��i<2 k��Lݝl4\���#:4����[�����o��wo�� ���H���)wg�5ˌ3���<kVu .�gҼ��cc.�hw:ҟ���h��Л��L;�BX�L	 0�h'Z�5[��{A�+�:�^�bѸ�aAe�hW���{����#��w�{�+>sl^�Wd<n����C[��j�I������2��d�9ù}N���75� ��`Y�!]�Z��ĳ�-ɮ���KB<�yM�L7�FOlAۻ4fK*0��+�8�V�I-� a<~�~1�yz~�?��L���?��۳��jJ�������I���U?���U�*�D%���â��y���N�*Xb5,Q�;-^��1�
\�ŧ��K�DE0l�xh�����U��쫃trX��l]L��2Q�,���-_�1�}kih��t�Ś�hQ��4 ω|�q��6���h��V�]���nO����������@�|��nnv�f���Ų�qW�-�8�˦X�8�K�|��φRC6�P������,��IE|�}�+��L��O�����'��z��̧��e7O�"�R�P��ό�Xü�߶A۴�������h��E˷v��RB =i�0���y_ܨZ� � ,�h���>3rm`Rd��������L��}{3{n����~��=����}~j@�Y��ź�ֽt� ��b�&�����oFS�H}W��u�@뽭�v?�U��sz|�C����c���O��7�YPP�T�w�	�ǹ�iW��zqm�1���>W뼸����/�&G f ���4�$�ْ�����^ҡ�ZvM�rL�|�(Ǯh�^���	���@��^�t�/th�(;��%1����%��XY�
��ܾ�y��	���X�x�Ӡbln�Yз~߷}ߞu߄����B���Z��<l&����ne^p̗1]XI��?�&���l�os�^����ٞc;kЧ�o����v*�$)Pd�g5�.��2�,QL��k]��60%��"��m�i�䳝)xQH4	l#8�g�'�����&��l�,.0m�V�
��a@��<<X����V���1i�����)"V.ag�L��ed���mt߄��-�7��r�k�
�f�=:�Q���k?p�[m�WM�}�ھ!��͢`#�+YT��ճ��j#����<�ob�;�<�� �&z>�}q6k\U7��k*P�f��V�HI5h�׳d�Js}X����;vJ�*K�O��Jr̀e�R/y���U����{�>�̀"�5��|.r����s0Zk7��i^6-����n�bk2��W��pnXcl<�-^��W�~��w���~���@��$Z%��,v1�[��_�8s��T|Js��2kQ�Z5֝��l�ƵR^�)[rۛ����^��ׯ������t`����'���g/�u���y�5��G����i�~�jY��kZd�̒,a1�i�����H'_<&i��G�)��������� ���F�_�6�y�w������7���W������D�O��p���Y�v� ���G�j2��mT�����*?,F�{�,���!��B�(�E`&I؆��C\����@q!\��,=� mĢm��mR�3�
]�����AX�??�P(��L83�cZ4����t��$�Ί���6c�6u{�Iƍ0�ev+/�^M�|ߨ ld���hLcW�R�X ��ݿ�k��(q8��`�Uvfay`��8���N�{:�~i�=� �S{��vj{�>�hy~ߔ��x4�8��iE}1��0h���	�� �{���ǬU~V�����W�΀CbOt��i{���mB1PX~)�a��4���6%/����������HM�$�����暄+!��j� �e5��[訆E��F�Ob� `��9*�Ws�yȀ	�2�Y���ǂ�"���m�^o�&��*b}�b�G�6p}ǹҮ��}6|z�����T�B1��}`d�����T[�ʊ�L��?6�}���o߾j��״�yh��u��Ю1��\=�����R:`��Ȱ����C�{��_}-.Χ�I��˸���=�����h��]b J+6m��{�sA}b660���s�[l^�gyo��F�>�5��
�q��b�u��>��-�On�R�w(�4#��{-w>ër�i%S����c͟Z����
����$`�-\�V}j����#������������o������>�]�Un�|>6�9[��fi�V,C�������������H����L��������Hi��\c���c^^�gQj����o鷿}�p�.SN�e��|V��� ���nOw��y��~�ޯ��<q1��
'jdM��"B�Z��ꓑ�)�ֲB+ң�f	�Sa�2��c m�M�15��j�N�{�k���^:L�|��5}���^���?70�����~nL��4K�ؙ����a���šb��=�5�Pi��h5pt��66J�^@ܝ���|�[V��]Qv�l �C�_f�*�q��� �5��z1p��vF\�������
�?b�ε�߉�TԞD�����{������o��o~����������u=�}�h�ih�noؼ�k{��f��yg�� ����JZ����}3����a!a��ց=�N�>6�[��?��	0��˶%;V|�d��K�E��^������u��ˈ�����9�)�b|撯Y�2�^P	)Z%�$����9!Hǀ��Ԡ�����X �P��p��Mzig���r���}O��7:X+>N����X#�"欷�&��dF���Y���-݁�F~xvq3/+(���e��D�@�}Y]��	N�IٹJX𬃶�3i��\�t�>��][����4e�ݍS����Ċ���zAMV|w�R�Z#�����=}����Ʌ}`�%��f�j��88���Y�JU'�%�@�������o����M�>>=K��qwC�������O�=2ʾPa��;RױVPh��sI[Nӻ���������P���z�omI(���������܃EXS�,m�"A��g������J\���!e��� V|_��%X,ق�n�=�^�|��)�3�7���o_��������@���;���+Q�'�����J�;���݈��PxL�vwp��/�d���`�s���U
y�[,��N�p,��ϯ���5agj�����_� ����Ml���4K��I�m�ى�j���_}Oo�~'Y<s�ܟ�8X�lY�RYKS�u����Z��W�]�F���bO�%_ǶT�kRL���G���� ����m�ҧi:HL /wb��tӘ̏���ino�w�#�����4�������Ǧa�.G�;���Mf*�UT��#gA��³C���kaFO�B8ƥ80pSqN�>�j��L
~Z�Tl0/�9�F)�,D�,�t.Dy�:8N�g�=.7y_�_���3�`"[�Xu��m�����!������3n���Y�H�����w��~�W�����~��[��ى�x|z�_~�Y2�>�'���^K������� ea����������I��`�}6A�I���H����ه��,�g�"�`i�\�n%	hߙk_�
0�5 �Z�ؐmYe?ﱶ1�	0o4<����>��[|=46��bݷ�rP;�Kn�۰��8�\��gxG;#�(���4k�m�$��%�|V+ݠ�VʑH�U�f����̆�t��,VW���T`_-���,�1g��ߍV�jF��b�!������u�V��)�r_��s��%���8*ΫӍ���&�w���S)�a���9�) �v���Z����{qW�6��ʁ,(�[��{�[�X��㞚����+z��[�{x���F�����	P�uh���d���T)?��|��bsV	�o
�}�ww���+���q1yˑ3�I���le���%�#���s2����$&X����g��� =�.�s���%�7��%��_�!�oL��y<	䈻`���Y�F�'"s�jR��KZw�HS�9��-�����K@�-�؉��$��n�:?5^���@W�o�>�����o�o������h졁�A<�RF�ĚZ�}㺈��<?s����ȑQ<I���{��'9���L?�~�,蒑ɠk���W�~�b/qd��!����F!��5(鞝W��9NZ�����J�ӱ];ѫWoiw��ߧ��C�L3ݴ����5��{����]�Y)���͛uP�*�+��|H�F�<�a� hZ�� 
2�F@+�A�����-�� �'X�f�j����0�E糘�HOgv��>���-}�6�ۇ����^5-�n7�?6�����=��~���^���Y��3�	�h��+��2�QͲ0���(�T�W�����ɰ�T��$sw'j�S��UM���z ,`�a ��1!W��D	`�K���~z�u|��a��||���:ϝ'�:N�#+$������i ��1 �,�;zh 뗛�gSw�B 0.[�V0��SjK��T�Xu�k���o�Q�������|�q]���įܐ���88>1`�6>wW$���9s؁	ڴ!����~�4ga#��k_�ΥJ���2}Q슞�9[�N�a��AI��Z�#��fƯ%D�"hu��I�	G/R��-` Q8��ƿ�0�1@��^M��d�E������ΧM���1	aO�ŉ|��9vM���ؔk��?"�^VPv�gL����.a�fi��d��)m�������8���j�Y����E�~��k��Lx��p����8&X���m>h����ʵ"9 Z\���#y)RQ��c���y��ot��S!x#���џ�5�7���VXQ	J��iT�o�:�d��L���t;n�IM:.��ߋ��ݙ���S(������>(^���/�a�e�%Vhi�2-�k��G�8p�>'h��J���-�Ý���w��I�N�)���b��a�������|C����������w9f���Y܍�Z��ŭnn�#?7,�q��K���Qb't�s�VYN��Y�
b��4 ƀ��k��UA�����>x�ҘF�RX�{���)Z���2���A��I]�|͡��+�C*���������xv�L��Uv�<�݊ 8/o��l�R��	�-�ȫ#]ݑj�<H�P� \-�C�-�l�(�}�	�,G{����t��{�,$0�Q�\Z9uu0�/5C�Xp���q!������Ĵ�������������M�O�F�4�*A�T��`�i�e,�F�4X���n+���I)>����X7[�zUq���܆��Z���gl���F�e�(�����#n@�o�̤�nS�@�x�����9�s��˯�����S�=���ꀪJx��%@S�1Z8�$�kt1�~MwM0_�K7�{ј�~Y�i����?������M�:�~�V\�T+`�1�G�)��Z�U�QqMt0A,qh�w�݉p��L�kI��밝� @�� �.c-b�`j�q�tjc��u&��mѿ�x�i�9(C��dI��0P���U���J�ԝ�y�R�L��\r��Yݱ�k��&�Y˕:R��8�f�8"��&n�6�~��ed.H@(Z�gbFn��a1�=$�"�I��V塺+O8e�p�<�ܩb.pĪ)��4v���Uսw���������z$���,|���Ӯ�X5y��� u�Ɛض��	�Ya��$;���3�u؋�?I;��V�Ac��Y�A9i�$o�S�ҟ��ykS�����Td�non�Bc�sD��;Vo�!T�V`W����\�F�((��?>﵍��8�/���?���:+]�~&�?��ٞQ��B�jlp���'t�x<d�0�D~���=Ux.�	i0�~�X�j�2 9ͬ���x�����c���2��vx?�Gz����/?�����������"�x���j�Gm�ƞ:���؀���p{�7�w?�7�~#�-��3�3<>~h �$%�xW1�a���mB�z�n�Dٝl^�"6����n랺ق���G����,XCx��{�C>
8<g9~q���#�w�}�����od�0�T��z�J֎�OmϏ��ojg!I�����@~�A��G����ڱ
D^�o17&�힞O2�q8��֯�Z��2f2l�X��@��80tZť��VN��~׀�dl�����Y������G=������S��:�mbB�"q�*Z}l�l�)�R�L5qVC�Oֺ%���s�C�
�UaA�Վđ�{�_;>�:6�%A����i�����/0�k%^�.iS��K�<��t8�]���̼�"�&�W��3YI鹰ٚk��xn��{-�������͆S�+�V�Q5=��1Bkŀ����� ��P��Jh��������%x�ok��ԭ���k��ߘ5� �iU!��)��Lf�f�"5��[�ʺ�o��̩���	3G�&?�;���Aɦ㘊[-�:��gg�U8��Ĺm�a؛-�
�.JG\g�=#�X��t�ˆ��d�O2�(��	A��[{hS��$��2PC `y�|���i�Wuָ�"b'i�y��e��n�5�[Vk�� 㪧�.i/��#)��������4Fe\\��.��h'�1����Lh�HD���6Yan{�[�V;a�,��8b�B��%� �m�[�=�%����W�R��|�}���e]��o�����uKH�XE3z�Ty���	R0.X�dEW*=�/ʀ����X;{�v|�ԕlǥ��D������]_?�7_�j�^�Ā��
�g�r�a��>�9A�i�����ƫ�衽_�yM7�gJͺ6^V�?|�@��������i<b+���ѭ���@j,V۟�m��AU�OUȴt� �E�j󪧞h`5KX�h���������4޶14�����X��D�@��y��~nH�Y��̼npa��To��!�<i iD@a ��P�P�.�jq_,�v�"�5��U9f������`��Kh��ąc@��.�'�!�⁬2�e����v�:&H	�kc���o����׆�_�q�?�������r�����zR��h������VZlM*�gG��`#��]�*B��r����K�whS��5qY�[�Dl��"RƏ>o�����UlR2��2�������bp�~�R�� ��DkL�5�@/Ԍ��4|+Y�ߨ ���Z(t��Ș����^�j`����4jB�<�E� B��f���bJ�dF����Th�Z�BcMs�,bxA���~rvK������YB�ck�W-�J�������������eP��%.]2��*4k�M��4��V���[�?pR��AU���?Ю�gA����1H\i�͒�%mBX�ۗ���%�z��"�J�~�2�b�TI�0����R�
�$�:f����
�V��1��Zq����YՉe�>j��N2���}b�>/�W�Q������㌬�I��"��P�}�q�Nd��6�X`V��*�Vٹ��ay��f�ۨ%����bEy֘a�[�V~��\�\�`ވ����)��◎�y4�C����	���+~dq8����p%�Y�{��W�����i�|�E��~HXE�#�<�D��r��,��Q��,����]�&����B�:_Sbk�H���;w�B�Y�B�O�9=5���o������_����_ݰ�J�G��b�f-��I���n��|�x�k)_�r~/?o�o���I#�i6��yn�����~�s��O�����Ӈc�K'I���[�wS�\	&׭�����	�QC��p[��(����>��o82����I0��a꯴j�r�և���|ʹ;X��U7�V|�k<�&���
2tr��m-��ã@��5|.��&�Mw���	�܋9_ۖ�h�gw��X{�&I��JP�=X���d�g�8����n������t"+� ��`�TM��Ξ2S��̪ ��23������S�t%9j�\1Y��N�`�	���~'`����}=����׷�����E�+Co�s�5�+��&J k�(Ü,�8ltbq������{��ee_w�������Y+�Dy�*I^V�5pl�0u˱�ڰ��F�xDb���Y�
�|py8jJ��d�?�iCS�ύ{߆~^M%Wϕf��B潂�F� {���h��ee5k��ENasg���Cg�W8�ǜK���*s/�K��];�f!�-a�(uVJ� )����L��P9FY["��M,S��E�W��sBz攔E�(xxx�(tB�)f`G8����i9����e��F�D��z���bX%'R&l=,k�|)��	�=����*�=p<fk�j�L�P7u+�4d	rJ0^��f[�C�	'e��.�-�,�aܚw�"��I�g���<�����m';y�JgQ:
 �v�L����<����+H���NHi��_�T�	Շy +�8�y*ޯN��u�Y4�G�$�f��m�XuB�Ѷ��*ĵY-��V���8}T�d�+�/ş�|�K))��y����*��������f3f�'����O�>��1M�f��G���ɓ�G Xrz��U����檟�u��_�qd��+q��-��5����������+v�WB��$�Lv�52&L	௻�|B�_MO�>-�x�2X��iM6�N!*�g O@��0 �m�#\hU>�-�M��YǞ�N�Mn�ퟎGRmyƬJV��1�)���H�9]>yJWO����H��P��PON�Ň-���<�T� ���R�=[=;./^��n&V%�H���oLy�U�ur'%A�+�3�HA��خy�0P�ܧϟ���W�p?��$�r^L��g��{����rywG�߽�bb!�$��g�(�)�W����?��gW����oZ���"�I,yTG�v[�Шnh����g64,������<	�ZB���V:ii3��X��������d���{���N>�L��/����G"�|a�.����o9T 9UD�ߓIY���C[JTc;���y�6��ypc`FX&y_�֯E��!Kj5��1�*���0l���Ya�A6"���3&�8a��O�5z���F.R���Z�}5�ۛ�9wen�M&$��`����sJ7��0�t�Q�ǖ�e�yf��dM���ľީT3�kSI�h����q���v� 4BS��5�dX���K����w�-�ȓ���$ٜ���9�\����(S��k�c�4�	�;�;��R�V˺HIZ�-k
V*����){�&�x����-�(�,RCؖX�P��0{��'��	�l�K�N<hJ����ȧ)�@da6?e�I�p/���(ʎ���؆ù��[��6b��c�fʜ��Ok���nJ��)�5B��7!��ZW_M�}n7�������;����C�I+�)��~��Z��DA/f�kD'`?�Z��h��y��ݮ��U��T����Oٓ{��Uw�L%��ۻ�p����r@��Q֭���������/����o~��@�r{s-ՙ�x�� &���qGf^����=Ag�����em"�0�N�`�M�N����fEO�۬�i��C[�:Y��;�$��=�zGΖ��bܣ���wZpՓg����3:+�e��-�U�#��E��K#���s���%烕��e��A�~�NO�Cڳ'�˙՚3&l���n�,y�2po!��Io��F���ɳ2I����^5�.|�5�]f!-$ʱ�k[n�{&��;N�ó�&�]Jʙ�]B$gg���o��ǟ���jK�QA��f~&}��˨L"\�����\�6�%dS�j\_u�)Mp6�vnic�XC�jɛ���(�����\�/�<&`Ah�a 1���`ǃ�7����zh=��ڗ�_r�G?i�O�)7�ʗ�V+TC�9^R�p��H.���̈́��~"t'������1o�W}�"j_�˽�"	]
�������c��*��Y� ҵ�r�\�m�Ve~���)B��͂�9�����J��V�dYZҋ����9���6�K�����(A����{�N$4!6��)i�`#���2+/���*@���u;�����n��:?�>z.������4�� Ȇm/͂�U?9 *[y|����{٧�}5��R���Ӥ�U�Ҝ�7�I>��{�����ENKhP�����5�tִ89�P�T����s���Ň��k�M0�i��HSC�F�-�٫��u�PLH-�l���}���9�=�r���\�p��<�~�x1�,Wk+�u萞,O+~F��0�O)��
���o�e$�2�F0#z�_�]V ����}vy����}���?���o�z��pPh����J�����)���5s�"��т=aTH^��:��9C�7|`�M�p$��䄶�%c�5����#� �%&(��)i��P#��5g��@�@1J�..��Y_�W4]���萮 T�(��Fq�N&�+!!��d���=��W'�5��J��o���7��|�D5$�q�t-}�\rrF�|�]A��
j<�2e�I����c\�M[-zX��ޜ�_�We���1�9����L�7}�$9U:���˹_�zF��ʸ��_?ҧ�6�	CUd����۷ʯ�9%���e�|��7_Rw;O�sl��RI7(Թ5��՝j1
�9,Ƚ&ߓ�=�o/�W`��1V�h�ζ����LY�jw ������?&��C�W�x�B>Ur!&m�Z�3��g��d�W��=�W������L4�&�\5����V�jMڦ�OD��MA\��ޱ��k�\���yU��>�ï�^P7<,F���Z��&yY�RL�D�ȇ(��s`iU�d��-N�N/+�(��p���1�J��v���Ȝ���o �\s˧	i�oE��#�-K�sn1U�2��������z��v:�^*?��,���ߡ����a�����=���@6B��
�lx_rt�hm��)��u,�6���˖?����8D#�� |��Q��^.F ]'	7��b&��Jh����^"r%��gbP�8�v�mW:�����2�3�]�L�S��0z�E�A�!t.��V��C�ÍV�xږ�N��¼C3Qm ���5�7<E�o�<_�í��@���W>��{<"���O�8	�F�z�:�D����l�8W�L�X܆׊�M�s�jr��F�e�ע�;��۔{*��=�ϧ������)<�X�[^�{���B<$���X���L`g���]J�rVGC4ի����*�hUԋE5*IR���,%��ĉE�l])�m�`	���P�������|(�8����Ph���O�6��D���&s��{w;)wj�) ��P�e�D;%���u�l�,�@s��R��J���͔��N8^���W��Lk������T��*%�D^��PM���s�[���a�̖��J��NC3]������n�����o��fU.M�Eв���3sy�y�X�>��e���a:s��,��5����Vw�h��p����u���B/]�"���sm ̾g(�(@�m����Ŝ,��l�C b�.�+���D�ߤ��8��m������_���)g�}kB>U��q:7�$���-��x� �f���V
 �1d���Cσ�L:�X�i8�z���?��G��d:X�r	�IU�M����	T��x�3���Bu��t�����`N)'ܫԷЯX�-cTE�[��Qs��KR�{)2 �Z
i��Y�f$�� b�x�ޅ$�Ir�~��{��z�>���=�
�Fג�f-(* �y/t|
��01V��U�,����ɤ�j9f��m��v��s�\-�pE*�4^Z=Wyᘒ�۳5�-�+�RTX��&��Yq���x��{Z�Vj����*��e����]2'X7�ջ�;��ͷf��1�#%,��Q/�B�n�_��Α�E4 Y_��K�@�c����j�A����ES��:'���&(Q_
�N���N��Z�C�^o%t��
C=�9�-�9���X���*�r�+pNƢ�:�s%%���������)}��W��o^�,��*�ܩ������H`G� ���K�����x��r��Kr���-T3�y���0`V�#̰��c�v'�^�S{vxH
�/./�����|%5~�����Ozs�F�l�]�B�DATAGRM�ƪ��Xg�)�x�$3a�T�q"kN޶b����$������.��ۮE�rFZn���z��0 OT�Ұ0U/�VJ�f��9{�֫;X}�+{�Yq~�7_���{���B�XP��{�!�8q/��R���H"}l�"9Eu⫎WE��
�a5Ry��ꤕ�ыYb��ٴ�$�}/$o}�l�A�7u�F �!I"�XK�aTM�(R�TaH�ׅ;�G������"�0:�[��u\�ˊ����w]�Yr�(��1�2��K��	�3�z�ؓ�mH���.���h�:��ydr�(QE�'��k^�(\�x�j=�p2D��^���ɋ�R��i֝ "PRLz�r�g�=�[�˄����*��KZn���
`	���ŋ!�y*���\���Y��r6S�T'T'k�^[���`����d�����:`z,�;f�r�M���Jiǟ[���+J���q͘����:���=�r����k�L���Gs���-���&�a�͸�2xx�6�ȥ�"�W�a�l�U��z�v�]����9-��Ɖ�k��N`�Zp�����r�������W♕��-�\��®M9�z�sb�	W�M�-U]����q��Xye��e����c�� h�?��1��#�%��<�7��>�ƐiV�'�@I�p��'�/���C�J�T"�p�x4�_�h��K/Ͻ�<�Tu��U���c���y��p�1�I�q&Ӹ���(b�"t�1	��~E�	��HG HS�:����]��<�S� \�d3��Zʣ�B�:o��`o*��IA���Xk�Qrۥ��7�(K�^�E�0��M�/�����,9"���ĕ��#�ډ��ߤ���$a�6��^,v�G��;�$��T:ɂ�*X��4�I$�={���*H1���%�}۴�ƖS�+�k�0ej�����ʄu�)�c5[���V{F~Ɣ�Wg�~zyF�)����Z]����]P��b�f�UN�F���ͅ�6ѼV�=��D��xM���T��B/�mU�p��h�_�zY� ՟�`�<�D�qb����B��}���p�����W�7���������V�dyNJ̷�$씸�f�-XZቃGX=>����EB�` �\�g_S���Z+W���2����!�i$�Ǔ��$u�m�"�l��u�9��4�Hed�JZ L�. -��+�Τb�:�̬�Q�ؙ T���A���dF(���� I�P$he��K��@k_�J����};���a4k\�N����h��52�6+9I7I�^��PRbi����@�� 0X̒Կ�<0��e`��@��oH��׶ p� vd�B�J�2X0�ʚ��Jd����P�7���k�\dHـ����8(�����<Ki����H���84<�\�������Ý>�Z�'"�M[�Aź�6�@Z=l������T�c�I���|j0���S8���`>�\��Bul�O٘GS���P���e�|���6��r�u�Gv�T����׹�i堰Z���Q�zL!��i0��n��6Cg3���-�}���`i%���#x��eE�W7����k���8a����ÑHIk[���;)��bx_�"�zɵf���ܖy#Qp
��a�3sZ�%��'�6�g�$���ƴ殃��
n�+�oH�9�N��p��9ia6y0턖�v�"`v��/_��ӗ�.|�@��)I�@xc�dz�h��i "�7��������r�)��W@�m��T��y�k�e�>~ɋe����D@�֠�p/�r�Y uAۚ�S���Z)i^J�����,�O��xvR6ɴ(��=]��� e����8�z���\N[,�F��N�a�rE��&�7y�{hl���16>!Q7�	O��ɶe���&�/������tL<믃�w��f�c+�פfxV�5�c��d��w}��i����\H��u`�ή9E[�%ҋ0z��$��+S~��{x���h�Ae��MO�����4�$)m���0�/Ϯ<l��Z��Ġ��1�yi�? ���T�	����7\�}1xnmV��W�6��8����D_WSx�y�=7PGjǔY�&�@w��S�z&Qi����ϲ#	���"��4�S�'�2��cɳ�36���KU��~ٵ%�h(n��2�Ri�H&��F�!=� �S@4�9�����4�¼�L�k���a]O*��kfB�r�?}Ԛ�D�͎��t/�K��:/���H Ѧ
��6���t�[�u� `�";9=K�}u����]�~��˺�1zlo�++=Ea�F�zH���,��|�{����C��UP� _���O�n���û�k���޽}��T�����s&iErp]CY��FM�h�\/��u�Q�#�=co0��:uR(Ŵ��r��E�o�_��7\--�Z"��x������>�5���(��Va�	R��V��$���$��
�B� ���F�ͽ�hsqȄg��tr~Q��1�U�H|���//�����gL�����2��YlU&n� �m{�V�sf�Ε��8qm!1�r��O
���q���*��'�@_E��9��;�qn˰�V[��+���"�1`Ir���Ѽ��W/���G����x9��3;R2�D5�-�d?���ٯ�>�sW��b��`Q�LY�bY~zO��D{��\P~��7�����i���P�B�m�jIƶAU����VW��ٿ?���cuU��=:|�{x�F�q�w�LÉ����L�;d&s��yR|@�Ʈ~���6l.�֋'R
2�x��4�<�{�a}1��U)³���;m�ß�.9 �l��!E0�\�(���mEXN��Dj+#-��N�<��}���,��E��T��6's��-Pt���5�	˒9��@q�|y��S��b�m�o˾(2� �+O���W� x���8��uhC�`�Z��r�D*"s�C+�I=7AG���vE�j�^N����+�wX�k�2p2��J�!�d�����F�0+�5>�$�I��㼼/�G�3/  � �(�5���ҐS��c5�yM�ٽf��V�����O�� ��0>$�#g��� �u��Su�T� (e1ٛjHx�A���*)�^k��:?.�>�F�{v��>8�ٚ	���H� ��1w& �b1��r�MO��/i��eE��~}By��������iD��'�O�y��^l�U���\R �`x�={rV��s&��\qػ�5��e\ AH�@>�p^��C�Tm
�nH�6k!��ßs.*ٲA!����̅n���*�S��-
�6	ӯ)��
�r���!Z���p�q�E�h9+��0h��n����a��ٙr�$�f��|�O��1���&(Q/��(�.	7�b�qd��?�?E�T��8ˋʂ�Q�p~��/< ��;cR�-^�������~��-ݭ�[�iD�;�\�	�u`c�ޓ�D��ʅ0F��b>���i�\佾������g�y�+m����L�͇�4CI�;�����V{�)�[X��MF�p6&*g��UH�*V��?~K�m�4zm������?q���<��>l�S�A��GKcz!�E�˪��3��������Y�ɓ./����y��D��삶Wk���
_Z�fU)���Gу����<$T��s�4�[�Z���	s�I���p��m�غ��+z�?����2�j�V&$��� G�9R&`�J)Q>�\ӾX�w�ޖ��#�?"��e��Wഗ���+c��K�������g�~�	�s����H j����B�nAu��no����#}z��67���d/�U�N2I�d屲~�\��	�<*����|��4vM�؟+�0Pܩ�n�[�0�
����N���>�BL.w$�C�'�ڒ�3V�y�%�N��˺�;�[&�����|ݗ���s(���&�ų��fjXg6._AF&%���3 �T�*� &S^�7^���{L��Y>�>�[�}6���ܣz��"���E�\'���<`}��M�����?9/k�<E睝��>�~-�`��(g��y�_��j��\��5���-]ù����JMtBx���T����1��)���BZkq����vCӹ;8�[�;��Sի����G?Z��n��ёI��4Ln|�3���Y#�Qr'����|��|/�j	� ��M��S�,C�ر����!W_�z�k����SN��q�T�j��}/������.���s���c[!n�y���^��=����&<����<��-�?���V���9���Ӳ`nˢ�½c���bQ�����䂥.�J���fEO+�v*s����暮?|��]����Ǽ�t��%=)���9�+'�'cj\L-�K��#���r�֎Y�q�<���3}_ƕ�.]?�|���!�z�o���n'W��5/72�:�j�F0��9��C�y���_IhG�V�� ]	 �r#c���m^�
��& �p?��<�0�ÿ�jL��qxRЩ�z6�K$� R峓�K:��[z������ot��KJ��"����!�I�-�3��Wk�|����V	,0�V���-�LU����� �r�n^��ӧt��7�����￧��7�mR�\@Cf�Ζ-rVl���ݚN
���K�����_���{��/��4�5<I"��~Js/^/�$
L�U����>�f�Q�¨���)p�e��y�rX���Ⱦ��i{�w֎V�x-A�Q��m1R��%���T�1j|���ȥ'ҹ$)��t��m��[_��ϑ1[������ҁ1�_�VW>�9<P
����F`чn!��j���F$78�˫<|��e���v�˕HH#���O�9��4]+ m6�{���xSxY�@�cv�V� ��I��.$��q����T.<��]}U�s���߳x�ᩙN�K�<�9S8L%�*k��؃�� �l��6��~���ɆA3��Q8^M8]�d�m3e�x�v��NQq����$_v�vX�#G�A���dL`�Ys�U�G��,\$�� |M�bBob�xD폀��ރ��Y{�p�:w�a7��^����+z^@#�$C�*���W�d)�U@�蒄lH���ˢ���H7��[6��L���6O�5Zr{�����o���m�24ޗ��7�u�ˠ��h���:��Tc����qY�+?�Y���x ��s���pRv1�&f�\4#��_h���#$�+��e��zT�p_1�� `��w��٫�51I˙�HY�	���;������Z�hK&�2lR�#�t0?�L��g��6(��/��'B�9k(T*	-eDz9C��~Z�h��_}E_�������t��	5ggeĆw�H��ʔ3P�R�@����s��g�/�~,�]��%�ȓ=�$��J�AN#@���y_��?���}�=-^���|�i. �`�C	 �i���L��?��ym�|A7�h�R:TU�I�������P�y��3�[er>�i+��;ٛ�~�=!v_�@��*�@�����~�޵�r��),gګ�1�ڿ��Fp��\����>��S�(A����M���e��C�ٳ>�q�������lk��޲c^�
;�}wmߚ!׫���2}-x�P����HG�wF�;�y�I���a�u���V=�}����;|��#h"��W*k�����<�{���M��J��̕�-I��%���C�j��2F��E�GL���5�RV� wAu�lΡl6�8M��(�y�G�x�Í*���2=c�Ү�a������se"����y���I�3�� =�>�X�� �� ��7���F��&�W ��AH	��f
n4����l�9Lv5Rz6��a�Y/�ґ �"Oy�qOT�Q,n8Wl�xH01�%;/� L�S�`���x<[��ݰ!�lv���F/�Z�pE�2O�j�p^+֍�`["�U�j-�_�JF�T��}.���x/��1D�x��36��e�.��4|1��,JS&��U��!��K^�̽�ڥFoX���<�dfR�O�L���bJ��k����<G!�I���ƚ3 �/���~��N����>M������y)�'q󲫞/d��D�8T��g/_����~�]|��'B��V��[�,�.˭~.H��Ҁ-E��;Mf�I��!�����g{R��gt��7����	<_��@��\@��/=��(!���\X�0)��&o�К����NBݞ�[kK��(�M�۱��x�k�eT d79 �ڨw ���YC�9��M�������L�������>|�� �N�P���z�Ì'�t1�E������x���C���=�x\6UQ#��z޸����D���:��(&*�{xc�}�g���Q!ٽN�����lymN�I������T��H���F�7�?�[���`Ԝ�D��AU����?�h	�ER_�OI�\˘`�����7I�ud���z��{7��a|����J�d���덒�h��LJ�38V�=�2ī:�焎>�.�X�X 9�)O"��d�p�
�|�p�X;��R�&���h��O�:�^|Xb>&o�B�6��5-(^��!	au����R��M}�Y4f����l�6V)�|#B�ŕ�����E�!�+3��q\=Cc�'��{N�5όo^y
��� tS�'S�.Si��[�c��!��+xB��䍠ҭ�p�4��zh�Y�=xk��o�#tS݇���#��J�����8-d��X��m@�;&�d�YK.�T�4е{SL��^� ��:�|�5K��
?�ȇ��F�� ���.�PZnB��^,��`�>9=���==��Ot��Î�j ��^�9vHx�1׿���M1�e�D�����?������;}��e���/^��W�}��=��kZ��Y�O�T���]��ùUm�{�{(Nh�˗���~�xB?��?�����0��p2�Bd
\#�eOy�x(S�l�-*d7G�Ou�dW�D;kc����y�^��}D�'d�v�+��>}�. �C�<w(�Bg�	8���3N7�67{��MJ?�7��هB�֎�I{5$����Zȡ���c5�;Uv�{Șs8^=�o�����#��ߵݝ���~yS�,$�h�7M='��A}sC����sF=;��m'����5j��>�s�w�����&�lXOVajs������^��-J�3�����n��k���m�l`9��>8@���Co���߽]��U�9xT�`d�iQ&��Ü�jp�����q���i��`aą]?��3�4�`��9Y*�0����d8˓�9^N8���vL�;��Q����?��l� �-�b�A�w�HK�VG�P�3�J�<*��u�����q21h��|����{�oV�BS�iC�ey�f��e�t��oT�64��
F
<S�����uR�K��f��c�����_*����6��>d��D[O�/��JW:�#�R�9|6F�/wǸА�F���T��ė�W�MZI�tP*h��^��I�XFj�����L���}�#}�mq���%߱_��B]�=�m��E��ϟ3XB(27���J՟X���Hʹ�y1��r�Nhrv�mDWW�-o\��+mP�S����%���w���O/��=��s�Î�/wJ�9�i̲{\�ڄ������ؖs]4S���$����������m��� Tea�3Y�=�d�����p�`q�뫃��}K���A��X"�42%	=G#�I������5��-9��t�;E�>�����@�Yr~ւ�J��xT$�z��s���dS5`G�ap�4~%��W� _ٿ�Ǳ��U����?�pLG�v�W��{T_��8qy��,J渟����	�� :-�9�=��☢Gv�f��AV�����ܰ����fό"2�>U�[�l����ͦ �����\�a�⒃�Ǡ#r5��hjcq� x��/rOz��A�M�B+�6��M��1���$�t9C����=9�v��Юa�=�Ur�Ѥ�b�}5�Z=2K�w/�i��p�:�C�5Ɩǰ�#*`��{��q=9�dS��%��\�ך��y���+�/��$�/F�x]�;�t
�:��|��+N�Gr���Ϟ=c��$$o3m�I�~m���QP����sT���D�岍7��G����#`,V��z<�Y~_�aMrAT����I<(��S_A�5��F��+�l��je�~�eҍ��А��1l��U���׀�U�k)	��I��,���v���v�掆sg���BքSkY>���0d�
O 1���A4떑,��03{�����٫>UK����������?�-�?�^>Fg�-�OuQ�Ӛ��\�W޼z��3|b�o��<���x����+�+ �[���0��?�* �\�_U��7���7it����懙����lظ�!����n�;��ik �8�fB�m���v����`;)�	.D��#T�ז���l|��Fu��$�P�h ���0E�?��?z+n��2����K6/:�c�=8�э�����$?v���:���`(�ŦI��L�1��-��'�35Ǳ��u{��Z0�C��u�gE�����uֶ{�s��b����7s�c�<�+\Ry���&����S�p���Ct ��֜e:mK��	q��`7H{_�z�'<b�h�_����j��=�Uf�\�np�#I�����傷� �x�O��d-I.Kk�xv�	R锎�m�rR���3,҃�G���g�^�GIj��%�MA�Y7?�`1�p'"z��#�����.b�۾$
	�x�l��⦞W��j���P��dΖ˦gU�z�6!'$���3�9��P��c���/DG�c��1�U7S=��x�9�-)"ŻO�Lp�}��k:�2���H����$�vZ��6!���!�_x�9a����i�G�
�fx���艢
v�=WZ��mơ��@�%�����I���5�$��-�|�s�'����PI��C�@��D�&��~1k�Ƭ�P�3�X\IU B;��f֤�x)�땳v, r�� �8��g@V���꒮^����w�|�s0�Zo�
����+ʠ�,s��kH������@X?ny���$��ͱ ��RE����X���꞉U�۞�@���	�<}��9�?b�3_Rb:!I���f��q�{��^�>5�(NP�9~up��D��;H���c9���4��6�8�ѩGjȮ�p��?\\�t�%ȓl�	�qъ�!�U����9Mf�o� �S��\�H_@R
���C�u$�3d%��$ �	�gx�����w@ֻ��zS��9�u�0ș����t�ۗ�.�"*��z:���ȯw�R[��+���2�9��HJ�06.����b�2�Ӛ��ޡ!b���P�D�8����̀�g:�����BW=p�P�[��1o� ����{�|���/�L�xu���g!�e�I>t�X̄?-�N��	*/��C�~/ �c�c�(��
x����������0�D�lP��������7=�1��4�� ��~~9%M��\���B���y�a��t����RJ;;R1D�N�SO��Y i @�cc�,3�9Ti��[/t��<�rd����p^���&V����)����4�ܪ��<(�Al�#�'m�۳Pe�*�N�������� ���WW�q7�=_�����ʃ�_ͣŤx�1|U{��� Q��t5��y��Ȋu�	�Y繂t1g�@5%�������)ȇ��Xlz�|8��s*(���3�A@�{%��LF|ʝ&��pl�+$� ����p�_L���3�v�{�x�nOv����0 �9M�,�^�Ѵ�0��~�� S�G�F�lNG7����`��&��Q�#��G�U���h��b��|�H6�+:���ю}�[e�c���n�3��7���V�`m���'�}����Wa9lT/-M���r]��Z�^[�p�@���g=�[�,9�c�[�>\Y=�z.���(�7=)B��׈GR8o�6��<Ǯd2��������сU��<J�MO>hW�K��W��W�x6,�s=�=0E��
�������lͳ�z��^N�Va��+�L���f}�����٨�-t�L3���,��^�~e�X�u�{bҮ	BKgE�6+ƭ �44^��2���<�H�����聲��[��1�I�dEB,��F��Y�~̐k����N�+W��`'�[��~dx�{IUM�5��A�)W\݌�rXl��RUɹ��,s��'���s�'�
�=�B`vpl�>ol'm��(�BS{���i$��|P�銲���CQCc���zU��\��~z��f&}�z����I3�cqy"_v}nU��gί-�D��"Bo�/Ķ�x�2ȓ� |L�����=h� �ݚ�Θ�Vdx��K��������=������K�<$/NO8���H;)��r`GL'�m��9���/x-�:h�k���~E��;/��_���F�!C'����}Mm�V�d�g�?Ǐ7���I]�C�ڗ ��?�Ƣ��say�l�!�Bt���-�)k��Z ��F���1��}b�&܂�x����z���Y�;�خL��\T�`�w�j��݊A>{�Q���yǍ�Ԟ�ŘR���	zΥR�e�`5{D͓����v�}�ƹ<�qL�/��3u�^D�;��йJ�K�C�O~��WE!ˀ�d���pI��4��R�^s8$����>>qǆ�����+׀Ye'E��E�rw�� ��E)���-6SNL���i���r��K6i,Y��>W5[=�ٓ�@�%Mkn=���}��{y�{et�m� �
��Z�Gv�a�ͮ7������̫M���/�_c��G�SC��+mSx[�����cc3쀓�|��ܕ�?#kS���c�Aɠ8�n�Vr�-�m����jY��KF%`�7Ϗ?���A�� �o���z�ڰ�}r��������].����g�P:Ṃ���p��۲ozmĞ"n31὇�_���T�������������q tΞ=����N�ʫ����G �<o�Sa&y5hl�8g'�Hx�xN����~����@Nӓ'W����tV@�Oq�4���ڍ�&�V��lU�4�H:y�n�c�;��R�붣��h'U@�_��
��y%* �j�<YRk;8�N/T���\
:m���vԖ����l�����;a!��ޏ��a�V�p���]mMP�+6e(��$)[����#��uޏʨ
�l~	:�|��4ܗ��~0������Ǫ���OL�S)�E�*�'h�Rd�vW+�yV8PhC���uOV*�?U���Їb�[饒�'P�N��q��( 

Ǯo ����'�SZu�lўyC�'+����ό
T���G����|��$L�DM�0������^���,�z>�Zx�7�3�U� ��嫅�n`_�����d���:r�v�07�uCj>���q�䉆�wC��m-�9���R?w/,'��W�=��A��j���T1��4jo������Qk�́�s(D]f��c��Ѫ���!��*����DK��D'�d�槙e7��l�������V籙�w!X�������2:j���GM�߱0�ퟁ��T�?*Mͳ��`2�K����|_<Q��~&�m��gL�S���<HWի6U�ǽRSU�Ҧ
&j�����U��[��/��_?̥S�8���i7¬�tv�4�:���l���(bX�D~��~�������AsQ��/_j��� mn��/-��M8QI֠�W�.�cJWk�)�x��Wz��Ol\��:����0���a�^�w�a�[�r�5'�aɞ�5\͹���i�&��(VN>v/��>�I�;�
HU�0f�����h���ߨ�}Z��%��=�Z!ӞL�<aH�Jq4;����6U�dq��`���-�В(�Y�,ǢŶ�{�(�9�^��]����ƙG�ynܟ�=��G��#	6��&���S#�^�5ﴓ{�L�9�k�w��Y
���$"��6 ���E�:k�V�%+D��2w�-�/���%������ ��b���nKF�, ����\{�a�N�ѥ7���|G���u�N�1��@

4�e�cOݾ<Լ/� ��nNP�t�L&�uxÏ_�)n�(�4���ԅ7�ƪ�Un�	&k�z^��Q��/kmϏY	�<�MB��zC��y�������=��޲�B�ާ�sK�f�P�(0�j��,�X��2��%���-խ�iI'x�I6����ٞ�ݫ�ܛu���(a���'4�hQp�9�4�q�~'��� m�Gv�����#r(�p����)Yqf��$�:����h����i?#k�A)(m<���zR�^x��dk?%��f�m�I�*�Bd�3�Ĺ���妚O��I/�p|�;&�d����7R
{��J��" ˪t�Ė���(��I�dVqǡƮ�� ��"wD������Fg������?�����{��dFl�1.��R�����-s���	r����}Jk�gBh��
V����"q�ڞV77��_�Bo޼�;��kCk̀wƤ�Jk.���8w���+	-��$��fV 1��pTv+"��ws��h��0[=s��{}m�9�P�\dT�n2��|!�+�P"+H&0oh��gz�=s9IO_�n�g��^]P5ma��2`�����i=�x�k��%~T����z����I/x �������Q<d��jP�Bq𮆎�����¸��AX?����%a�Za�`QX�f��LV���a��˹���fH@@��������:�/��[��▀�U)B���������¿��<Y/��i�X� x����Z�^;\�Sτ�[ڕ�?,���53������ؘ2�оTB�/ƍZ� �
2$MR�Ϳeih�����Ix��e�c1T�h�#0��^�M���O��ni^����}��Kg�{/�HV�T%_��=��$$'��V�΁���S ً���H|��f^�����ٴ�y�s֚8����)Vi���d���`)G<|TPf^�~��-�/t��g㭩u�� 5�J�}	�=�p}���ѳ�2�?��N��;V@ f�Jҥ ��mz�a5n���հ���	~8#O�9��_sk�v� ��3����ࡹR=�
<��#�B���q6m!T5U���I�AV�C�t��||O߽����iB�V���у�# \�E0���	ʜl�+p��RO��CC��Ak���Nl�P]���~�ᦿ ֻ����y�HۉYqU�QQ�0�E�[R�4��
f��;�LN�h���)Q�����t��\)U����d�#c1^0�|�x�µ(��b�����(�����>�P݋��;D�� f���k�B_�ڳJܻ�$h�	�?�ګ���P'��˅���?~+Dk�C-(3����_s����#�G�s�*��,�L�h��h���0V�.�'�7��ݸ���D�eTe��;���8�)��D���PCjR<8�tb����~Ka�9�7�`������É�ػ�^/i�Y�'l�e�:��s�m�S��<��$%���6lҢ�:������9�U-`�Napl�kX��j�\�6E�&���)�Vs�F*4v�ב�=�)�ǒ�3�aR4 ���2^<0��޾���޳�ϝ�ӄ�u�ɜ����{�O�O�ـC/ɐ��hƋ�Sd��9Ε󄙍��T��d7�6vp+v7�q����%JQ�D��M�>8��&O�B
���Y��,�c��&L��q)��ac�=&�k�p+w�Q�"we�<E�_�����Y�Ó����A��|IK�� ���n�ۇ����S[1�"����2���N=�6�<2�m'�d��c��Gx�'yB���nuMs�N�2���]\]�l1��fҲ���&�fx�`��� �hp��r��9�A����_���k���_ʱN�8ؓ륐�"����\��ш{q��� a��} wyA����?�z%����ap� /��a�/4^�wz��z�MQ)+8{��oL��]x5x�ސ��7�R:l�����C�q�����<�$��Ȇo�!	y����ď��b�ī�*����;y�jȳ�3���:�����#E���Ұ4!d��}��/%ʴ�0�[1��#����uD�^~����b5xꇫ �%��"��� 3C��Z���e]1��z�ߙ�����w�lȲ�)U �O9��4����f~���&�w������ ]2zR�C�_?�����^>=�b���{M5@�ے��bP���v{�6f$Ge#*�6�#wOAi���Bu�v��+�����D�� T�]SS���yJ4�#KzR�H�_>JyL��5l�� ��H�j߮9�êȄ�}3K�hR��*)<S۱{t���T��C����12�x�t`�|�6�z�k�g[Y�˂������G
�dQ���Pܬ3IR�)S�6��ƽip�:(�z��q�^Z��u�fb�9�u�̞�e�Jբ#"�ٸ�E*�s�{�*>��r>��c���X���a�L��x5i�_��z��9�����\�
*B֙�W���UhZF�5�fkk�!�tO���g	���Z�iژ���x�O���ѩ���*�}9~'�C�k�h7��>;s�WK�M�t��2�K�b@Ӫ�|R�W�~d�\�%C��;���LĚ���d&nhr��Dr�	 � ����u�6\��d�W�^S�����ⱑF��H]���a��K�
��Q�ht,?K��&7i�ԯw����k��W%,��.-��xU��*o����kxJK�j�!"���y?�{�)��A=0�M���s4�p	�~���T�8%�ȁ��|l>��;� ���3 @
8�Ȫ����<�2���}��ɶ
���c2A�FQZ勖�ܛ�]={����;No�[��uB�x�M�?����H���4[1�[��z����.O�ty6�y�.9�%+�^j!`.�g�J��n� &�hףw�@�ȿ�^`��4�"ɻGĕi�������ܚ�U���$p}�{WyJ�q�v��"c���$\ ��6a���'��g�����9�ڴ3��϶�-s�$(�� l<��+r<���:�j�"�wh%�f �+�'�:���/�}�xC;:aB�"�|q��v��}mNj��>M̙�4�~�ɑZRL���+'
��H�iJ~�ny�ʜ��m��盧�@�@�g8�� kb���DC!�y�c����e�C�U=w�}��:C�P֋f��w�s��mrx�[l�%�~/����@�v�]�獊�!x+����(2��I��7����`��<	M�-�ɸ�,�勧�(� P,Y�K�;��B��o�J����K�����ܹ����feq:�*��E���D�lE�����ީVյY����i��yh�=�!�J���_
���rd�]^�W�}G�|�-W�19dC��I�ڬ�ٕp���
����\ڍpa:�-ћ�N�u.E^��=0�d�ž+��5�;�di����Bz��^x۪J�V�﹁8<��VHS7�t����<�����"'���E;T����X9�%߶��c����[�q���g�*��1�K�D�xΐ|6�Ń�t~{qꇊy���0��1��� �tC���!��N���si���c����I�))=�4��O��sg��$�FѬO��y��3c�`�&B��L&��ڄ�5��Cc_������W[���;:�5���:�Oi��=�!��ܯ"o�޺5��@X�	���q���b�26`��P���-�s���agi.(_4?ߞ���e�8敬�+��,� �� ��.h`�TEhd���hǱ�%{�p���(]@�.!���dؒ�p�¼r#��	�����밢<�����}�4���݊���2�%r&;�Ҟ������>�����(�EQe1��x������b��"Žr<����	�^�:��	�kw9��7+k#�������V�8$8$#�������������Ňr(C��?�A���(X%�^��1+O�8̍�U;�u�����*Qj"i���I|wkM�.�H��ޮ�JQ�hu���7#kH3s�$BY�����J��cn�jD����Ԏ��r��x�@r̰����:Y� ����)�WF��jE���P��t��<I�|B�Hs�*
=�jXHIM1��^��� ��Fmu���v�1̳'�sV�����|��R��䚽v���!����1rD0v~�"`�#�z=��V�2t��� ���6���Vڀ-o��!�ui���g;�k�
(E��pV�z6�q��|P�,i[���v���m��ؘ��� 7��X�K��gO[������k�<~���`X�u8|��:8����&�#� roZ��c��Ƨ��X�GF�R��l�pɖ����{����Z�%�;Z/bC��\�0Iz����q�y�&2�����E�PAE�`<��(J�]�r��S�)r��͒޽�Do�}�i���I.�@+�Ux�u_q�-dD�d��(t/.�߯�Iv��>X�;�W<̍\���� i+�}͆b�����\dn�|w�/e�_���3kG�8�Гf��)�'Q��w,3ha�7Nf_�y_.���z�N*���%��D�g� b����a�! g���+���J�<t`P�ׁr �a���a�07�WWƹ[���iʛiYn�_~�����[�]����>c���0Y]`�~l�=/�d֓�ɽ��^���QuC�w�B�Yד	Y[�4�v��DJ��(�h���;/�;�\Ày:���b:|���1[�P��w�pH~욎)դo�GJI��V�*��l&Lލx�!g8�K��Z��R�7���X�l;IR�8Q�����:I�}�l}�]���|�.�������M�n�S������_����F�G�"��W�{��	zK5@�P��nSx�gh\@��C�@�zQ�Ai���A�1������$��Y�4rcɥ�D<�b��jF����=/ ��g���/����d
L�˼�q��"�>��f�����������d@^@?5���*��c��R��9o��I�n�vJ\�����RiX萑{���P1�&��h���@4��?���ݺܟ�?��{�I��d��|U `��l���P�*{���<��/IQ�i�yL�0/_n�bë^�� �J��tc�Lͅ��s9Pp?�B�|<�Bo��1��K��t?Ô:C���@о�����NT�y�H*�=��$���qL�8�Bβ�l��&���c溞����܂1@w�� �!ST���yG�����_�_�w߾���EY;?p)3Yr����wY��OivrN��K&*7����]���w(�vg%Q��
=L�XZq�����x_�x)�!0V��pv0�?N��K\���	=*��yrv.9�(�h�5#���9���B��-B	�W���{ID�B^�ꎶ�r�~9��*��8��PA�k2W���g�0�*��?�fe��j��ɂ@CM��9<���2���X��EI��2ځ�n���ӛ��˯	9�;&]�/9e ��)/2n`�1��R�XD�{���$�g��"nPp�ľ�)�,���l�;���h���@Pb�]Y�~oU� �}��<axC���z��[K���I2�UM(u+�6��Z7Ir��%V���0�0v�Ӝ �wڕ5��*�Ze2;+L�V^�9ƾ���2fi��s��M�W�mr2��f��0}�[6��#�_�׏���a�U�� O��a��Ҥ�1c�z�=���o6�+�g)KC�L��k�_�B��JmS!�8K��Vb�6(s������6�C���<�a1zއ�{�jR3�s��D���=[CO��-�T_�[���V?<�z�lu�� �mS	�̝���1K.,�.�9�ޯM����ԜNB�s�\/�Y��Q�|D޲����r��
 �>ZE�0��a4c�sH���kǲ4>?���ݭ�NZ#�VUX���Ϩc�4��y��e�5_G��M��b��z^��?z�}�A��Z&��W�ʮC%י�^Sy+�/3E[E8P\r|s
x�2k�΋�A!�Z{�ve���o�_��W��� �ph\�{�3���sn�ZP��?3�������2�VU�,|흤<u;���h��"c�n�Cٽ��f:%� #���������QP4���*�s�h�$�ph�Е&�U�K����m���K6�;cu/�=H�3�c�(�X�2�@�6"py��.�1.�L�������k4!�]��J�$��9O���2F�I+U�Ed$�b���𱀯[�J{ϡ����ۻ�y���}���5?+�s�.�"99�0$��^{0���uAr�g×T��@�	����r!����#�A��X� �@\ �#�Ib�~���f'���zA��=�����]�>�����Y��"k�+=�Y���f-[,��+�,���ȡ?�����W�W�;2�	W:��K������+$���+�Ly6�u:�S�%��ra3P7@�#uG���Y�� (i�H�knEfTs� �7�����/���ꂦ'�iylu����Ss*٬+��2�l'�4ENt �l4فC��)*���!e�N����3�(���½���?�#���(��S0·��9��2`BdJ��A�擳SZ���,!Q���ަ��W�։!z��Z�g�L�O5I3W����*��}��=�%�u �4Y�3^������]�����~O��7B�M��6������ u�1�벡��w�z�D징��~x�������"RO�Ko�|��7xsln�j��w;Bej��'18��GsM��*�d}���r,�����M�����(;����\I�S�A-��a4���oz$�!���c#�s.`��I�U����͋��*r�O�X� L�Qڰ�|��Z�8?�%ps"'���x�f��+��{,3o!�Q��l�U����9���c����;r

�V��RY�s,i	�5���~ٮ� A�޴$#ho��D+�tٳ�LB����3� TaI)|�����Ď��n�ܲ��0��y�䦪�4UK.�E�:c�wt�<a{�`�]q���0�����őzl� C(۽�����#�/����?�޻�[#��o����ǟ?ЇO����� j=���t�nPp�Y�X6e�|��A���9�R��D��509p��ym3g��V�0=�x��T�E���0��z�*S8��q���u��Ee��~14�=��p�n�^�\���j]�n�c�W�(�X%ZH[���L��L�_�r�H�8��y���k^��ro���"y`��5����x���y��c<��ڄ�He��z��gn+3������g\���ԯ�p2���)�:�������Tw���r�FT*O��D�����f�Ţ.2�݇w4��^~��]\PS#�b|6�ԛ�z]Z�d慔+d�t�P��|hY���k�Xr v@�`��b@sN�NV�����P�ZD-2����W��g# zY���@�)�#<��ږ<��@f�wk�hp�"�LuB
,�
��R����wB l9�D���ZɁP8��ኴ��4X���W��s`�D&��):�d�+�(J��� ��-Y`��t����ne`��UNE�3��j�O��CY�JV��

Ƿi���q�g��\&��US����"�L"6<�V#f�G�������Ǜ����:_���� �&�F��C�)���I�� �0���.ˎ�4�$giԫ�mǸ�ieϦ5B�L&�M�ɖ֐kkB]+��5�L[��RDa6���p�L�݂Ӡη�s=���lU>;q~��ת�N�'3SM� �� ��RO35����d�.�G�ə�!l��.l�`��-�U�7E؝�y��O���D��Z�+����G�Vh&���-��n�!��5p�z����[����/�/���b}O��:ἯԊ��$�E�tHfE^���h����1ڻ�)(e>��3k��)�#(KI�>��ܫ�J�����K���Ł��z��)�UF��&�n
b'�ύ�7zǀ����z��]p����$]+�����<��b�j��A�J���%[_B��qG�_6M������o��kM�L�{j��DVʘ����F���v�oxD`=G�]��$�
��<'�"	B��Jf�+{nʍ���ѓ�!T��)8G�3i��%�B�e�wB+_O^����P�@��ݻw����ʹ�g�����3z��5�������>}�X�e�o�n���:=?+��T�dQ��y>i���H�Ep[0��*�!
1�t� ��ҽ틣O�&8c�15-k�¶|rv~Du�GIr0��T��:	��l��XoQ(7�-f���ۮhyw]��	�ʺ;=���ײ�G�r��t:��0s�ĳ�T	([6�'��ɚ���)&��8g���

X��g3eQ���5+���a����4>�+%8J�X�?jA��.P5�cU�lMd��Y�e�h�>#�d�Z�F�E�Wbr5���ʿ�U����>g(��D0؈q
�Cr�=�j�d�D�"��U�{�=W.������j����N���Ô�(�Ym�M�[>c�����;+0�o��$�r>+�"��,�g�ܭ^S�x�"٢�g.��,u�d��TP�.$��P)�*k�
H����	��-k�+�ـTz��v��6����ֽ]��qS$���z%���}qn��q[�~՜Q�b�w�"w��UJ���s�I�8�y"l�y�I>�#"���ji��X!Y�dԎ��;M��[�����yC�����-B�3_�V]Ll��X�R��u��Bρ9;٦�6]��L7FT�����]�����n�<�8%�j�pn�Ƿ��{H�ǫ�0���jE�J:_�<���:���J"�ü���g+����,21¡8L��1=	H������i��B����(qe��y+�pJ S$���*�<ٸ�R|�8��g����'W�W���Vx��>K|R�&_�Y�q\�Ĳ�{�4۽ʙ���/^���+�{��v�ˀ2o���) ����_��'���.��(��ϼ�/��7�VjZW/|}��7L��s��b��>|�D�����/V��D���^���_s�j䶧m�Z\@3��Y�M����/�4#UëV�b�Њp�ip#�?#����Ǧ,�^Eb 㵝&+Kx��|/��A�Z��tN������?���@�If�b薹89�>��|"m���O}�:_��\�/���j��=�0`S���Pb���r�'޿����^�v���=��(a��y̫E>5u�*�?���E8�q�h\.vFC56��Qv�"~?����sl�}�uaI��iʭ�R+-ɸ(���Fd�n[�q[��nvy~JWgtU��|֊'K���t9o�r�s�m�j�{�c X�2�;p5v��,6B�0�E潜#KT��>7�%f@9xM#)���E�>��h��{5[���*�a��o~)�mtC){=��S�K��tb.;C���]�{���I7I��ڨ�ƚs>�y#Un��3�I��gY�q�O���Z�;ˠ�
²F�3�A��a��yi\�J���p�l:z�������
 ���}�/�o����R׀nbF��ǜQ��)�������Kz�pqg�.��	��'���a���������+m���+r�R&�u�O�V�����笗p�1��r�㌿X/O�p5K�<}�^�|���A����&xZ��Ny�mA�R��f% ~:Ge�d�p�ޑ>�jӫ'Ӏ�����n4.�Jq@677��
�s�cӐ�5�.�{.?��)����0@3��q�rr�ᖥ��^ֲ�4��'�~�+�0,��+��������"��ΰ+�	!�UYח�����|��7����S쟳��WԔא�z��]>{B�O����ў�C�������R����?`�O�����H�x������=}S@޼ ��Ty�:�;W֦���lo�nk��R��m���©&�s;12Π
L�ʐ�2U��2%�wĘ0K�9{�5�*s�Oi��F�� 1��e"��J�I��W�l �x�+����j�h�,��^�7��	� ��K��z�s�<����<��!����2��`{����ums��Ϯ��`Apo{S���! {/e����^8���v����^�YA�̥��2������z�n������J:D[��y�(D :��E�佡$���F��d��2�3{�������t}sGgz��)�.}EϞ�8�p2��)<VL��붫f��+rU:�⹴,3p��#�:%ٮUǌ\s/���9nT
j��؊wQx�dR�����b�b���o��P]���`�˨���o�t1�$8X�\b�#�0!(�a'I��7��O/ya��%�*����$w�3���Me���:1I��[���阾b�!Ѽ��Û�\<$����q�n�V&�gs
I��K�t���-��Ƿ��Q�xC�<tM��m��3���0���\�(l
B�*����+G����dsd�v���,נ.�$�}cT��Ǳ�r�Ó?0Kre0��駇��9�g� 􂨍ޭ>�G2�s|���Kg��a�d$�T�a(����p� W����y3�^^$��N�KB�5�GQ�!�^U���L��@�H#{��+Ty�D�Vpn�)5�D������N=��u- �k�Ղ�g�Z�	�ҎN���fꦔT.�� ��
�C�+u�O�/s|��m�-}��?��t�s�E�)����z������O'�_���j�T7�1n1ϯ.h�t�>kr.�=����H!��-��ȇ`c���s�u���i���׈�!�#��BV�f<�ǔ���XQn��[^Ɂ� g4�ߤ�0��Ođ0	@1q/�[CNɑ�0E��6\��$T�f�I9~^s��ɉ�{��eQ�ohy����V&7@��f�GX��м<a�N8�c*y9d2�Fkl(|yڿ��O�i3�b)�x���z��:�cn�"�k�B%�&!������\�n�c����츥*�j�ر��nW������>��!'��S��:?yp��h�]Z��ME��J��+���)C��o��F�4�x��V`��E'�n��\��v��\P|v��t~vBgtq�����(Iy��E��5�CtC��̝t� e���Ȓ�\vW�ȨM���d_L�c�R]T����b���y���Ӛ�V5���@m>���Mڔ��b!m��3�uAq���j��!�Z�i�fCf�g߃�잴ԕ$����N�_3F+�@��[��7��J6x�X`�))$���,�9� )��ٛ�{&�����~��=},7aG$�Q;�}#��(�'4Y\��FBݶ�i$�/�Bj��`D��gtQ���4Z���W:�4k���TjEF���pmSFa�Iï����`���߯�=Ǐ�fb� ���K��UZ���^�����u�x��&�H��_���/\o7�%:;Eg�i�PR��Ȕc�s<<�����z;{K��&�u̗�{�[ޏ���0v=���$���!Z��h�_ �\�~Ev��Z�x΁���	Ij��\4��Y�m9�C��\X�/_>���o�����=�%9�,A�H�TI�$��9ۻ����|Yq�9� �(�z�D���kv��#��3g��x*2��kꚜ�OH@ь2�*U0u��VE+? ��ʬ�{s=�%t �4'��ם�� .��_�;�z��<y����I�|}S�����W,weI���[�!Ɍ_�3�eT�� -L�c'�:�&�X��S�z@��c/����z�)��W59�Wb�f?������.�Iv]h�{�ap!a�P��yպzΐ(����|~�F��A��}p_�o��k�ˁ�6�:����(�S�!P�^:�ժ��zò8��:�"�#YRn�H�i��6���_	϶Y׷b�����O�8]�%	�V�I��U6��AeH+�$�J ��m�� �7���)�w.:c�c
x����\��)��1�ޥ�À�h���G�`+`��'��4� </F��Q���_��7�_�������wo�Q`c���r5R��f^J��ZW��f2�Nq��B�F|��~�hkR�����C#����v������k6�G9�<�c=���'�������jѡ� �`�3+id��������g�'"vS��B���=6&k�n������+�)�\�OD[�:�V��Jݘ�|AZMyV���q�/���������׿�Z��-C�9NWU�^ɰ��z�F��UT����Iǖ�f��M��^�^|���m?�~������[��c)�Co]��ǆ��* �Z`���_K��[��޿>~-^����-�Xb}}�A��[�{	��Nt��9r�Ꜿ���I�m�oTz���
��Vޢ�95��bH�Ʉc,�J�����sa-��֊;n#&��ޢ������N���@�/č�b� 1�,�1��=�F���[ŔCX7�������ͣ�yA�6�`�g�zU����зKP��ۛ'*�a��H�n6��z[-���䤧�U[l߽xi�U��c?u���~���*�,��ҷ�W��qP ��h�o���BJ�o���b��S_^�Cű�=�3V��4�\���<0����s�FY�7c�c�	���n'�ӓ|��T�S������[�)*��p����WϛR�bo§s�z<�����=.%����$�p�������5��@<ұ�jM���>{�w�ⵖ�ί�s����K���c$��:�cG]X����ի�\���0ͧt�o��c�����iPj��-��Vci�qf�T�Ұ��s���Q[���r�ΰ��d��u;!�.�>�Y�H68�h0z�J���eh�3���
^���X�r�y6����;^ ;�e���[����N��`�F�e�.+��2�>���H{9fkIa%�:dm@Cark3Y5��]�-Y.h'�p����)F�J=�Y�A����ಝo��2O<F����2pkB�(�Ơ����w$�Լ�������0\�[)�^��V��|]:�!��T���ҙE=��c0z7v��kz�ZWl�FΞ�G�˶m[0����������兵svW�P�W�_�Oz\?O�L/��:�JD� ���XF�K��ߧ=��O1�T�@L��鐰"�����ɬ��_�����*����1�`C]%�����lI�}u�*Nq�v�y\a��0 vԾ�g��g�^���sr]�a� �q]+�n!����r�Ӹ��y�̦͐�O�|� ˛Ou�*�� hL6^^�<!<(+�E��$�p�  T9IDAT�T����&�C����(�c��ɀ���t�yc
*��E����$WŎ���򉛎�]?�dz��vyz9dB�&�D���A����[�U�>x�+4�^|�v���ʙ6���M1���2{��ө�@�,ɪ�PPb,���7F�#���Z�o��GU�|�P���~����ܨ�M��Bt�D4�
|w���! ����CM��~���k�gؒ��b@�bm��)4h���o�u.�P�BД a�x�q��/ݼ'' ��ҹө=���,��'>��OƸ>�W�I�j ��'�f-�q����G-�2��W٫ @�9!�}+��>����g�j��ҵ	����\��'��N�����Zs�^�V�|��^�&�х�9
����p�b�ս�0̻�++���m +��-(q�ʏqζg�7ƺ :^[�[Jo��<�u��hE�z�V#�p8���W�4p��(ȻH,�Լ���}�O|���q���IQ#��,�"���0��� ������n��n �R|sL�)K
���{�����\-���y������;������cUik�ޯ
���*��*�o�~�s�Z�h� &o�-l#a֢W��X}{�Il���_��f��q܌œ /6�ö^1�pp���ںR�Ŕ s����]^G��k�� ����-�������q�����-J� _kJ��iE�[�6#�{��6j�&G��v�T=?�	�k�|W¤��]�ي�`,�l�G�(K����S
m~�
�GP�/�����{3���Wj�uX��B�U#;��E��W��x�E>���W��7��[VuR\�~���DOVG���U+�7oaQA�l�(�A����Qܣ��91_��0R��?o\�G�J�Ǆ������{������-�b]i �i����nKc����0%c �P�QZ�5=�7-pa�{`�k��<YwKZ�@�u�'����Vi�(��K�8S� 2�yc�3(B�{q'�_��W�_�-(*���6��b�a��t6ހ�^�:s�ɷm�o�^�]�+Ţ]s��O�Ǯ*X�KQ��a�\F�Cr����o�v��;{����g�a�Jk>Y�IFa�/��|\܁��9�q���1��ڀxݫ��a��t��L
@��������i�,M�]�ȝ�ߗ�ׯ?m*����핼�@!I�1�B�܀��vb%�&w�%�[(r�j(����vڰ��z��ъ����ۂ�Z��2D[1�U��H�u����6#�����_�gk*�ԇ� �{I���R5dG�z4w��C&j�i.�`9-�tڻ�3Qy����7%���V�.
H�ps�<���tDm���I~{�������G���E��t���Yg� ���cW�}E����R�6W�g�M�P���*�YS
�� ��2��T]@�n�8�����-0��P�ɗ�+���\<��mְ�CY/�5&s��g��c�{��>�/�_/4W
���z���\� �����1�(�<#��q��l�X�|oS��1�w���o޼Q�~[-x(��/��Z/�j�l�TA�a�;6K�,w�jVd�y/H��v!�}A�����HMa���v1kO��g	��+�'��\+��y�y�MZ#�!��q�}�LZu������,�u��뷲{�Z�P�M 6P0���ͤ�H.T6A	L��r�� n����������I^Up���y��?ȶ�HV-v���q]:=�IV�#�����-�K L���_������G�摝z�H5pT�UAX�{�Ʉ��i�&.=�M�|}��)�8 �o˱+��a�#��k��Q�8Wa�)dHQ�Ǎ~)[�;H�M�Ca��r����Օ�F��~/���w~�js�@
SFHŢ>�������^ܶ�;)ű�NM�4{�`e�$Ā��+'�5��26��\����Ⱬ}���Rn/�K��d�{�WVp
�͏-��Qx����|��1��uV�������qT�e��:~E��8~�0J'[
�ek��G�te�W�������ko����d�����j�G�X�
|g�+[V��d���Pn�|,�No�z�Rs�$2<�����lI����;���Z��٣�%	+�� ��SV�I��%�N�*05�� �>Ȯ*)l6$`Z�S���Ŭ���Mt�c����䌚����FZ<6
��=vJ��5������h%�5��IK��b�a��Ɉ�0� �9��C`p�?Â���:��6���S�i��Ev����n��#mk��8<c1d�g�=�^�ZRx
{@.^� �=a��N�&�9���6h�)8�I��R'O����5���^�t�[�-���W���ݥ���F�[�	�Z̥�$�Ɉ�%���G&�h��υ4�s�'%���Q%���OB��ӳ��n���(�tNB�u�t阰�����{C�XAr9�T�C��KXJ���x5���}�q��|���������ɰ�=B��<!�zu-w?�U+��޾� �nŭ1��f)�5n��
��jg�JU��˽��������r������l�oS���$�M�ݣ_B�J�K�y���C���d֧����/��/��?�$O>ȵf���=	Xs�+Lܫ�O�}�o��^*LU1�P��u�6��9ϐ~x0oa�u��K��aL�"b2��Ia��&RƺR�|?�Z+�����
���u%o^�Q�0B��T��(������SC:���ϲMC(�~��k2uH���ޖ��u��Mi�_�
��6�NUQ�X�y벽��5�jk�e���u���j�>M���~4:���2dB����)�ܭ�:9�=�������_�k/z�d\�Z���C7*�=�d�d���#jN��D������ Ǩ���pд��v�A�NY��,�
�9w����vg�%��.M6�Z͚̔��HI�7%җhm�π��Lg0P(z���f3��:�݋��Өc�X�:d�kc��p���0b��w�fNG_5�M�H~� ^<��L�q�-I��5$���J�\b!J<�N/s�f�%`��@�%�V����2gn?4�(��y�0�������f]2Xv�6��r�*�3��K�Z�Gs�0�t��ʝbw�����oP�� Tf��~��[�IS�fb846D���_�� j��o�#�����6xZKAQz��?�:W5ht+�-�L�lU���q7i�\r<�ZS4d1��i�) u����?S������3Z�7'*n(��w4�c6��5&��w��*;����[Ͳ���5�&HK��L7u������|u�W��,v���;�I�P���^g
���I��?�����W��A���Wy���{�J�lU��Ƌh��9?�|if��{�oOr��A>��|��2o�E>?ʾ�T������������KE6h�e3s�����G�7r?��^�C�?��������.�~��ac�f%�ǈ�)P��bmL�nd�kZda���́��T|��
��y�[�ɑ^i  ��8�`�hϢ�0[�R���)"�HF�0�~�����O���C��O+X��Ӱ#�>)�H��������K�n��@�z��xue���J�u�k΃�b-�B�\��H+�}Y�� kU �Ĺ��߷C�k���2��8���lq`交yW�K�/J��;R�vI|5}�0�X�d�w�Wkj����\�}�5S�.��t)X�G�K�e����^g6J	P>!�~���Hd�s�1<W��l���]��;5�����B��{�:1���A�c��Ѩ�c����:�
�z�X"�WOZ�:�9>��V�LG�'�9g��g�p�$�_4��Z	�-_ wG?A��4�B��y�^o��Z	���y�"��s(�D!e����r44�U����#,J&��(eNd���ڢ ]=a3�><�:c�q�|!w��K}3�[��Ҷ��|�r_���z�����(�|O8��=���:H>]�a%��E��s������5o�������s�P���o a�ض�x|4K��o��}q�W�����S!E�ޢ��rq�$F��w���}X�rT�<1�� y�{���K6B+��+\�_$u���VE�B�W|���͇��e��G,�������_�	�eT��]�J�AgPX�&�>�I���5���z_~�j ���~'W�^T�p/���N�ϼ�򬉥7x��2���Gy|��,������sy���G�*�*X��y�ɜ�;V0��I9��s��{�����(���/���e<�d� k`O���-y����qU? 4e����̅ŝC�70t�Eu5���Z%�u&�O03\�=��T:��[��]��U!ik�ۧ��E�}k8��M��9 �0����{p/�܅�d��]n`���-刢�lW�Yj�q�O�����J�O��XZ�=���dˁ/�H�
�������C~=+�;V|fyq���B5��4ky�0*�)�����<L��.%3��Х\g��u�x/�ձ]P�"�D<��C��T�X-��k�-
wl���G��5��$��x�s���X�k��o���R��U�ŷ��q��#r���=�b��@t(��َh���}H���� ,²tT#�	n��z�"w}:Wr�H�"��i�D3U ξ�c�e51��A,��2�|�,�I�
y;(ˤt��4��''��,��_�m�������L�@��-˙ +��A�㶩�{U�F�Y�H�[.�� � �M� G�rE߃�u�FZ�_ZWt�k�e9��|�4X���\T~`��k�Ð�@H�����`c����]pǘ��_	�X�"��x���u�W���ܥ4~�4��h㩊�K�����\X����ϟ��Ub&=i�m�7:"����Z��t�y��:��ǲ%�4�� ���h�3����(}�h�@j���ٍ��~�V�|��&y���R��o^P*ؔ:������Պ�𰏵�9Q�� :N��R4�F5��y�yn4���g���ѵ��_�]~��Or�捼������_��w�3���}�,���r��[��4��||�����<�������a>+({:ȏ��k��ۗru��t�SVl�C ��K���,�4��t�C��~��������w�d~z�s3����ZF�u���V���8��
v,f�on��̠]�����*o�^�L�J|c~������:�E��;�q����V󞙇�E�Bt�"zGF��427m�FǶ��ʹU��7�7��)�Ga8Ee����*3b ��

��Dc>�߹�oK1�ӆ��������ߠh��ϏXu��N��Y�S�hKܟ�H�/�LRn���Gh��W������e����R��Q�k��[޴�Vǁժ�c�u��^��*�^r��|���m�к'd�C��ё��{�Z. ޢ����}0]��3%t1��M��X19j��C��/�W�)�G"E
<� cKޚ�'�[� ����(��I�8�X�����D=�Fӳ�>�Y��Mt��\,��|7<i�#�i����m�P]�A9�ك��X/�|� ��0d�{����=R�����ʾ�z?�+��k���w� K��p^��bB��b��U�`�J�4�����+k}N��|DðӰc�7���^D��j�r8*�jz�F��o 0B��)��x�CGf��D��Ј?�aKv}WK�\��� qN�}��r]�S�'�������1��%-auyqK�[����Z|�Yc���6��#%����nD�2�-���o4��t��#��WU����$�e�VDI�&�報k�'tS��B�׳��d �J�7�r}}���~�zv1���Z}�����_Ba�Wh����TV�V���n&c똌�z_���S���
j'y��Q�?Iyz��?���+��&���;%P9*�!�a�=<?��w�ʇ���d۶��\r��B��Ou�����"C��)h+��$�I��2B�f���Ј�<(��׿��_�!K_��Ɲ]�jN�Y:F��t9���U�%FW1U :e�V�7K��������%�� ~�C����j8e��R�b%[Y*/�1��T&c�7�=��Y����`��_s�aq��n�ߣT�}��	�Frb^�f-̍��g���hF?6%*�_��2���m �8k��Ǳ�F���P1�G���]:%dP!4Vx��z�d������� b4>	�,*1.w�3.yh1706��{V��ķ�0b�x���1/vܠn��{)�CƧY�g{���t��X9���b���c	�പ`����8o�8-P���0�F��>Yn6<�Z�ޮ� ��ϡ:��z�*���"��m_/�ɋ�����bs��"р��`�6I���:�O�p��&��	�⳽�)������+������yO)�_��8�^�p�E:kAm�~�s �E�.�ꝅ|C�8��e�-�QRY�dC�n5䈁��T�[3��K��|�����&m5~��h�}�&�O0���F�mOz�v��	VA����U{R�/��`��˽s���}��������vLZ!�&?b����>SV_��I����N�_CKmQ���|\�nc���l�%���+�Y]��*�
��Y]��n-�B5�-[6Pԫ%�r�dh���0���.U��b�7�?p�[���`����s[�5��v9I�}y���x^���)$Y����x9O�4d@��X�-�l �]#W����;Ϗ��[9x}��gٿ������Ą~��7���w����޾�q}��Y�����/�hnV:>�5<e�<��ўd��Q~�������]ƻ
bQyw+wo^��?�A�^��-�ѻ��;dnG����w�ӿ������?�M�����W���jo����#r��9"���s���p�s��B���%��D�xh��<y��B�Q̷zA����X50�4`\_�:��*�O����#`ki����L�k��f��j(�U(��x��
��o��~�P\Z�?l4�R�޶�V'��@��(?IY�V��1�&T)+q�d���:��JV�q�
�0 �+G�Vո��SM���~��.^1���]ԦL^l-��u��w��nQ���
kR�l\�Ct{���)/P�n��ظ8�I(.�"{1��{����J}18%�jܯ��8u�Q�УV$��Ҝ� ,I,ef҅`dK�7����"g�QqDꊖ3(�_S�>lx�h^C�if��<��JY�L��SM�� ��TZ/�c��@Gs�+��`�i_LM̨]���2i�SI���)/k���p�J�lMb�LD�ޮ 	�͗Tq ֬�U�?jx6���R"���eaW���A�$f��&�G}�+z1�dT��i���cr[�5�)����>��|c��
0�@X�fZZ�=��D��0�6�|�v�.D��f���Mƣ�\*�j��V����0k��{��J�8h�A��˅`iǺ��cݟ>��N�����^x����L��,	Vk�	�>�-4ہ=�<U�rY"��͟�ثc
%BK�Z
�6{��K�G�yb�&-���r<�FOFt0������~�`ts�Ǧ�g�YWb�P.@�
ޫ�!|�ܤ0�~�Xj�6 i~z�#�T����N��o( �|� ;��(��A��^(�������Q+�������!8ĳ�+P�¹����]?����J����@���)�rDh��N���D��N������ǿ���|U�'� ^�J��H9ѫP�Cr��K�x{��@�� ^�|m�|;�޳O ����U��'nܒ�΋5h *��X�Q۪����s˫J�2��z�Ƥ���z�F�Ws����#��ׯ�j��ݳ����t	@�.���4���+�����ܓ����E��W;�����"�El?�P���v�\��FjF���~��z�7�Q�G�Y��^SH��$�
�❘�O9�ݚG�x4���6��*���(;�yf�Fʡ5���*����M�rlԘ��yr6�9/\Дnn��9g�*�`�$��z8%t}[�J��
W 7��ϒc�K	�l��9^#�d�)��| 
� &fmO,�R��ybR��}ּ<)�����9`�`��+�X� $<�{�8h�֑��q{Y�	kdٱ3S@�Xq	���!{��P�� 
�r��B���WI���@��!�hAM�D;(#�y�2��'u�i/�^�\��qb��	�ú����-�f]��n�D�t�P�fk�/�@tp7���`�cX�5Z4yR�7���M*��%�����{!���.�v�36P܀N���y���ɯZ�y���@���z�t�M�4��LXCn�>�Y�dQ����҅
.s��I���Bc�+��M 8�W	a��g����ϋ�9Y����ɠ{��˃l��e������V
�����b�~"��^��L��jBM�)f���P�Ͻ	�#*��=51�z�P!}xV���G�R��tI[~l�@M"�ӗ:v_�����iT7?==��Ãz_����z/㩎�� �ӳ��A��:y:J�2��˽��>����٫������r��˫
��j���_E>?ɦ~?l2g�L6Y���z����.��6�O?Mp��7�皭���$SqSX�3v�P�̪����(V1���SW�NZ���d[��s�t�W��{z�!u��z��#���u�N�4n���yUg���8
��]�����6x�l��~��{��=SxY+�Nr��6�{vX	����*������������C$�w�e)9��E(2��2'��b:�t{[���?ޱBݜ57�x�*��d��/���@�~�*�����vWA�v����lͯ�l�P�G7�R����I�&4Ǯ�2����i-
m���H�bœ�u�-M��5O�ț�w{GHQD܃i2�X������*m7Z[��{F��m�׼�:�ͨF'�"��2 �Ȝc�e{���4iU��1��<3i�r'��{�
�}��]+���[p��@MWfH�{jj�j��U(8�o���Dف��U���Hv�cb�P"��3�����L��p�&�Ÿ�:x��W8�条`�{�#k����W0���X�����n��������B�(�k�2C;���H��1A�g�d^��7�#"߸�>y���}�7��WT���1��V
��ϗ�\��؅�X1c�l -� R���е�gy'���uR�f��y�3�_v���'�98�����-x_�dW�i0���X�\��������>�u�L��������+rkx)�o�6tBЫi�MHɢ�q<���Z�d�:�*��$4��2�
�~��˖�g�n�YT�*0�O�>)�x���M~��Y4,L  ��D�2�ڨ���G왤�>�Gq�:�(� zx|��X����uEvo�
5W�7���y1l�I�P�cD!�}���Cެ�fA���5]ω�d��O�qv���8��l�M�w&ߑ��O�v�Eb���۷��g�DNL������}ڸ�<BbU���y1\:�v4���qq��P�B�Ԥ��꾒��f��5�� '�A���w�"�-�BoX�ļ+lV߱Z��%��"^��OHh��en�"�0�LCK+|��W14C�,���<J���G�V�Ɇge&�QC>��0��峵���I���ܤ���V��Œ]����U�����UssS��	�Zуm�.[s���2|����{r��: ���m>}��d�X��bL� Qb��)����@
�a���;�a`�]n����	�y�k��`��Х����'n
6X��P��XT�hU�Nd���n�=�BxҚr��W0�v	/�LY�� �{#$����M�rx�ޟ�|�i�-�L�8���߭��O>m,�ɪ���
���y/�Qc�`���6
�F�1r7��BI��Q��Ы>:����������8�w��
��Xr�'Ǽ�H˾k�һ��W��2gj�&�ڪ~d��`�����G�F"���2ϑH���B�1�oOE�P�z�e�Q)�uǗ��{k"T��*��U�ۚ�5�3��(������B��L��|x���|x-o��{�ػ��))<j>$��0gb_q�5D�^�m�dzh���u���\�۫�u�jaՠ�S�v�'�o����,��-��6)W漨X�)%CR�N%9�����Y|���`U³U�|B^xP�
��|��E�����aT"?M�%zo�z]����ܧ�jmox����9)0� �Ie�Mȓ�8Q�=(眳=�.h��ܕ��ɝ�"%�����>�jl��V�y!�\�Ox�ul�h�U.��Q������8Չ���B#�.
� sF�����5FN��)�<��jL��G�r;�k�ϐ�)��dF�h�Hi.�4�bd��)��a�����f]�"�DM�ƗP��d��ݸH�bo��y,�9�D�A���M`����I�)_�c��v�M�h��F��&�-^�jk�����Y>|� ��{'GP�����K��w?ȋ��e������H���f�nF@�N���Hi�*��`��&�����R@/_�.��Jak4�.���{����S|*2�u�w���)�]aG��G��7���p�U�ȭ`�!�)�k!=��&�S0G㰈uV�u�gD欈�&sA3�nA!Ia[D�դ�RE7��x+�,Nht�\C)�R�.n�Kh�V��W����0z�����͓�=|��rjt��Z�m��h�/W���A�������AFAF�I�j	��
@k��m��.���tV0��vw{��v��*�mU|Պ�tp��!�D�4->u+��v;����=M�hVP̧���u+����"�v��}"�u{)%%<^�-\,>�A����|.�їF���j5���^%�"��5F��^��MuC��y���ea�z B�K:UA�(Q&}_�h����Y��ە��/"�)%�K���:R���,��_OP[�m�](u©t?3H��u�!Q�
+�|C�  �x��|���O�C��i��h~��'����*��L��xVw������=�?���=W|.�TX��r��d���NH`��,��b1����QNt�l������*����J��W�5K��T�5���ם�V-ْ�Y� V�~�>��53�e��	V<�6�I���RM�lh�â	� �x(t��͇�z}�'�y�kJ��r�y����޼�����F���t;��"/��֯�~�e&����y%��$�ɞ�����9�~X?����`Ά��vY���H��q\Mz���#����-�f=��"�WWu��d�u�����-2踫�;��5L�r<�5ROh�+xlG�,�w�>��q1���369W�ٱ�_�@�+����A�H�6�C�Z[k�M<J������:ВET���]����<=k�c�zw�:���i�/����l��Vii��'�xeO���g��X��Y��6��j��b0���'i�ſf���H�C:��Zjh8�P1��|`��B��	��5���,��0�V�W��jVR�ڭH��=)�%(��G�|�`;~~�"����<����]���k��7o�ʮZ:ǧ'yJ�<����,o��^��Ȕ����F��Q|�};��s�Y9��{w��p�����7L`�ռ����VI�7g����[4�,���C&^^ށ:��.�����W����h��ͦb�nf��p|V��r(���J���$1]F��+��4����Ȝ�5a 	�{G�d7N����+�tOv^��y��贄*�?A��qi;�%(S7�![���9Շ�����-�\����+dl��V�����2K�J�Z3�������2��H;�p�2&����U���.�X��3�x4��A4�6P����Ґě���'�L2;r��&@���\�|X��s(]2P7��x1t�Dtۨg�X�]�-x/�YS��k.YJ���-r�h����Pm}�@�( �|��
QA0�[�6�U;CF�~�R��Nn_����%�!�c�:X��`a���\�>>������p^䥹���\X��n�N7�X��|�|�0u�+�2<�Z'��l��2Yh�D��V�v���<d)E�\H��|h9�` &��H���eҺ8_V��.��*��������Q�{�����۪3��e����j��~�F%�4��7r��VT�n�*k�6� �\�s�#,:ؖ7��x��Wm�
��������zN��F�`C���&]£S�;�{ʍp��w�ȝ�m�[�l�.=��*�Ē��0M_1a�ȕ�&2�!q�9��PY���5b���r���}5`�:��o���[ 0��=�$uh C�p��Ъ��*�U�p�}�|u/�|�[�|��0s�w��"y��W�\H� �y�Qu3KS�M��<l�Vgo�� +̓3��/>�ރ�H[��|������ Wur�=�+U�﵊kF��y//��,w�r��^�4�Gl�Eߞ�emW�&�t�n:
���v�A�c��˘gj��-�R�6�/�ǧ��������ԭ��R���<�{f
���W���1�z�jJY���Kp��R��I[U�q�N `g��9�z̊5Q.�$O�t�X��C�h�9��!¤R�֪�����v�&Oݷ_:M��y
�\|�}$�9(~N�[��w����m��[:X�d��~��]6@���̱�8�9%�''�R�B�!���s��%Gbz�%.�أ~b�p��K��v�e0�<�\��C�dpooUF��mL��si�Ä�9���/W���P;�-X�|�lU��Y±��O� � P��Z`�G��q����A�I�R�<m ��*c�dT��7W�b��e��t�?~���+����´� A!xʠG2�3礷��{��$sߧ��Vba��c��� �Q�xr	}-Rh0F�E1��y�XA�i-Tp8ǐ;O�x.Y�>����_��^l�kI/ds�&*/hH���0���]��5�Iуyn�.�e`��(נ͹ZD��� ���3����B:�|0���s�0z��[-�N\�J�kG�>bJ�����i���9(͘=����r���+�A�����,n�p^RT�4L8��I[#1?6����C�;��P���7-��(|o�7o��f'/_�a��fEq���^/(�?ِ�rf��,��cSS�=�amV��,����xD���Y:�7X3�ߴ>w���'	|�Js�A�]�'Пa=�"�L�$�f�#�0�[9a���1�����s��կ��7�j�_�e���W�7.g}��k���HI=�4:2@��"`*M���n�V`T8��@����>k+��}���ʝ�g�1��&�bEQ����|�˩�X]�(67��UkՕ��!^o����^��|N���X*�MΡ8��0<g�$��I���Ir�2a��%��V1߫䎱۞'3�@s
g�vKޱ�^0 ՄU����U�J���8�Ij�H(��z5��eTp:�@���8�$>������z����R,O/BFC��9Ow�E�@��_J�f�����xwtM�T�Z��0�ba�C�}�ôL�8Mj�IV)�{i(�(*m��F���(��)���|p�gWZ�]�K.�zhJa�ڃє���;z��"�
��:/�}^�&�sc�ߍ���(J�@ד�s�nq���'y>~�����<���]�{����a��J���p�z�Xe�X����k4�I���_rbw
����?�J�	"���CUB)(�?4�}v�e�Dm�%�*A/A/�2������L��qr@�@V�sc�͕�i_=Yb�������(q����&ۋ�s�7@r��8����Q�CU��\���F��]�r��VL�N�;j���A�����5�G*��;���^�r�BF����:�N��ᢩm8V�wn��N_�*�,�=9�f�1*3S�����um���|hw� ���k�+�vh��{O�t���$�
������{y��F^�]�� ����+[Ԋ��YA��8����s�7w.��i���j���B��2�cz�o��K�y|(7�廁/�����J�C���=8ٺ�;7�4o�+v{�B`�&Q� ��nO��O���'�5�����$��Z���k��2��2I�y<J�C21@��d�A=`�������ƪp���oc��/�ս�~v��y_��k�i� Jrq6�T�����nS�J	<�aRiL$\�^5/�:�
�|҄J?�h���-u���<�z����C=���賶!����3���n�˥sЙ�| f�S��!`�Փ����g�3;�S7��X�M��'�ا���H� 	O�2�o��ň���MU������u܈N�e(��krt6���+.�(�L�E:JЩ�ޝ��U����J�X,�>���h�v��r��͗�z��ɓ�����y�	�e�)�7l�2nP!� �
�b}{��k���u���up"��zP��_Ƅ��|bn����v5c�lZ~R쩡�'��p��ǣ<>�M��j�Q���Ԁ�U�"tm�7�Jޤ�ަB�3���d������z�y@GL��� ���VOǏ��λk��
[ACn�>3ײ�ǩ<dJw�ɋ�\[�i�<q��h���g��+)j#�վ�OV�vD.$x�0k)�Z����W�}�ޤ�(�<�N��ֹ��d9 �C�9bwW0����ZB������ՠ/C�
6�c,���Ϝ���t�Kr�"����C�>#�
��m0� 0���z_걋�<d"�4��0��ͳ�Y���#�sZU��>	���o�* �!�1����~�1��oQ��w���m}����͞��?�w��M��+Yl�Ӱ�&T?H,�xt_�k�r_r�J��0/�a!����q����L0���6e�څ��p�2aD�	$8���ƽ[���BE)�:n�������t ����H�3��u��������}�C�в��Z3x�j�2v_��ѭ���u��d�c���+����B����ꖒ�XS�.<��/�M�]1�|��Ϟ��u�rhl���CP�`���"3?(���<6k��x����������{9<��cr����%ۻ1�`��-��I\o�p<�zq�ټ1��um	�c��[j�R��]�6y-�~�x�;����`*�RbP��9%��'���4T��=�E1�.ճ��u &B�@�$y7�ʬ�LZ)i
  	�<,�Jz�F�-�}�옹"d��)�*G�l��~��Fn���
�n�a!�6����h��u:zg<$�u?Z,��.�������P{�e[���P֤�a�D�����Yڲ�p$�Z�v�,��9T���$�"�����/��{><˱� $姴���Y+*����.����κI��,��B@�Vw��<��D���Q�����Օ<�����v!_3��N)7(����W6F��5g˧��^�*6��o�	��h�p)x�Xk�q��lF+(�1X��@h�F}�~̳�S�}{�va��*w�X&(�&��UZ�=[H���;��nw���sz�#4���{��~x+7w/��GP��s��x�;J��bg�OYR	�t�,���lp�İג	#M���֋NB��8����+n~Oݑ]^K �!��?Ã�T�f��Ҝ[��F�U���=�[	}��S�k-�=oq��Q��PeV� �J��`��׍\ME�v������~�y`Ӷ���ﶉy��`A�LM�˂|�IWT����-r,:���+VOҍ侒�P(�	+!���BO������V�{��9��e��tI��Bu+D{b�����*I�k`���5�J$m����@�N��:���`��!N\Θ�:HZ�¬�U@�ht��Øi�Ƣl߹
*���¦��% ;!^_��b.UZ��gX:�+���W�S㟍�&�;�<��ō���dk�/�s�M�P���o:��V[qMq�6��#u-#����þӨ.�����d�2�?��+���A���k���w���)�Ī��lڽj�Y���Q���i!��;�O��	Pg��6cX��D��H&Vˉ��E�뷴��0�����59 w�N3��mj:�S� #�T��\MօG �,�c���[|Q�f��v���5�EO�����y=�#+�RE#f�#��d��
��B�%Z<���B1�2�}B!뢳z8�\��|I �I�X��k��^-��Ҁ�Ka�Ni@�"3̖�=�mi܋PV�@@�urc8��/�8��$0΃[��A�2���Kh��WJ�͍Ddkϒ)��-���"�/���+�|dh�<�Զ���č�Q�as��%���>��� x��n�G�7Un�"$s������e���v�������R] X@��fT;�mL�{��h˧
�����A�1�~���P�L�I�%���gs ��u��f$%<��Y��kR������c����v�	��V��*ӌ��"��oX*�J_��MU�r��y����o�wP�Pu�UD*�,*'��zc��Y��ثz� ���e&���{�s������âkPk@��7����&��}� �W��j�Pr�R��� }.{T�tяq�wup��P�R�p��=3��ı70��� ��Q k���c}u�Ѽ��jH�xq'߽}%߿}#�_��\(���u�dVщ^ c�V+%���+H?9w���}q�l�<G��&;X��g?)�k����=&a8
�ߢ4���9Q�L�8ě�-pLJ!˷� m�%�F�p95pc�������PZ܅,C�%�-D���,���l�����^6˕|����
6u�]�I��C����"�:��\���mZLI�eȲ�aX�7ch�L����D��HiJ������D�GV�(��_�D��Շ��du�x���BQ)�;)��߭@a�"���Y�|Voأ��&8�ȡ����!����Q>�(?|��]_�TςzW���8�'q��!����C9b�Y�\R�7��d��g:�k>��l�1㾦��B����)
���is��ݪ&������Q&�v������e���hx	�H��٘�G���������!v�X(TGT���@C����b��ƙIϊ�
ے��A	�=<٭h�m�N�ʥ�g@�\�h������B�`�b�V�񕗖0�]
���?��P�kki�{�e��e��|���a��7�"��� �m�ՑcY��
�������Ga��R,�뵰�A�������d{�5PX�Yxq�� ���7�����\��ݰ��L.0�ٜ}~��}���'��"ǘ><�*�oQcV��\Fm��	��E/V�k^T ��
��|n��T�H�Q�+�1�'x�m6���||x�@��|<��
a%ϟÅ&Õ��1fm����U���z<+_��&9��<c��f�Z�Œ���0�G�p��g����)��8�iS�u{�k������V�k���s}��*���T����GNf���.�X_e��9�Q�⁦Q�E:��8�@�bm�ڥ��gP`m��e�h��^�A�!t���P���B�J�iHK0��,[g螿l�: @#{�b19��������!t��}�2�^��OZ
솗�O�NC�˗/�?�A��/�"o* �W=�kO���*q����ynE�' w���*Y�X���;�W+��˾/a��m�S5*�Q� ��lD"�Y�Iz�t�Ɛm���B.�'ǂ��\��̠K�c����-N����B�.s��󮺤�&�)��F�h8V�|�C~�]����q���ڠ��E��?z/G��
ΐ�^4��HZ�>�K-��7p�0�e\�:D&Z���cY߿$.����t?�5�;W�Wzyұ{8��u��ڝ����Ұ�9\�̽�4j��h�׼�a��Ѫ|��Ӄ��흜*�E���t�yA�����U?���zx�"_��z��=6���p���JS-��gc�,$5\l�:�¢p�U0�۪  ��y��
���#
�2s�ˇ��~��g�r:�ӒfKD������#���Ҡɴ��#��?1��!l"n%����X���RȀ�&Ŕ�欜Y���a��A���B���P���%'윶m����o����7��|8Z`0�1϶'S��#���C�3��@z@3���洜t�躢�����؈C�ŹކX���[Y�َ�)J4�7Y(&H�a@,�2���0�}��O���d3mT���N�j������F��:f�;�r��յx~j��>�h)'�y_�da3��>�V!z�!=(�	ʜ���.�����O��0�vV�4~x��F��P���s���JΙ�X)Q�(��0|9��J��88���{D�q�Ɋ�dt�mO7M\�q���h�lR`�P���yr�3���!HvIP>�b@^��b��Ws�7� \D�]=��N��N��l�}�jDN��/�/�!Q�u���hu�bP"��� 3��f���~�Ǭ����Pͫ�0��l&�</�	�Ix�u��]���
$�!���'�e�_�<D�_ ���K�5��.��p�P��"�Έ�@���",����|`9t)6��C�nY����rm'�o޼�?�����/�ww����?������	^��;/��|P�C&�V������VIc��|P�r���g��)}�	Ȫ�d�
 �͙Ǔ��|\à!U+|2���;���0��E]h�Y/Rޏ�n�cH���-��b�9 d$%
Q&�r�i�|�ذ~~�<�\���s��w�W�r��*t4��
�>}� �@Aca�7�"la���zL��.-���!��	���Na�,\����qHC�Qy�=_�~���4wE����,?* e�F�d�P޽zP��v(#�${⮓xn���]<�j���b4�b!_�=:�O��ۯGy����g�ҹZ�Hu���a��>��	� !�烑��;�p�Op>Т�b���/a�Ұ��v/�Z�Ǫ��A����u�<~�M���/깰�cN��cR?�O���I��9i$�gv� ��Q��������@
�|DHv�^*������3b��C���Ӏ�f1���Ɓ��*'�"(�p˶(���CH!����Vs���An�B8��dV���~>AF�>��`d}'�7�Q�t'es?��Vfް5��M�z���C0���R��>�4�U~f�% ��M��u~�֍�^�����\5�)(J ;��L[�bU6�\���*]�[HJ�Yؤ�U�|4
x��%�H�#|<?�1��Y�Bi���2�ވ���{�4 �r����9dw��il�ɲx�|ٳ���ޣɝ�.w���P��$���Gu2�Rcg=-=��	�o_݅���7x��g�����Y:y$aP&�R�Tb�q=[��s�"=�\�ZP >�@�����=uV/��$ϖ�#�<�U�����li�)�PW��h!�\�(��������9����Y��Jm�J�h�b&��3���p~%r�1���g)�N���SG=�)Ha$��9���^#A_[p�����p{s#���|����� ����ʰ�x�bOX���%r^���'�Y��p ���%����0��ݠ�V��Ydr������L�Z��,�³���
����Y�����nI��:����`�=���=��Ą���W��O$25w�fb�C��	�e�X��+� -E���YF��g-M��Z-��E��ۗ*�Χ�~��\Ee�����Zu��ol�QB@�G��L�{�Y�&hl.�<$iU=P��W.�ՆH�P(����31+�u�d
��n�Ы�B���H��f��LP+t�Jf-�7�.�i2 0���r���uO��{P�
��̐���v$KyRpͿ��C���u>�T�U�T�/�V��s	1Y�R�SI�gX��'�«������N�D^�X���Gkm֣3q�:�hɛ���K�����H����Y�WWk�=3^'�e�:(R��g�p�*� PGki��L6�s�H�e�8�w�}�o^U(Y�ܶ�xs��Cn���!����
kk_���o<� ,Cf>bN��rH�F~@�(a�Қ�ðwL�}�+(C&`72
��� qn	���y  ��6&�l��l \��$x�z�* �{,d��@�:A�����ɼZ��ʓ%8�7��袁���Y�y�� !�0����#�_Wi��t��0'(�S��֔ZT�v����y�n9%ir%�U�#��ɪV��)�����E��zU�������y�g��$��m`�}�\��2DAi1 �N
�,݄���eqV���Mj|l���=?�@�}RJޟs�
���7,��fF�q:���.��s5�ԇ�v�h��ܓ+�S<�//� ,�N1�]Vު|�\�Vp�z�]5^���G�X���s��y�
��?Ê�klU�).��B���Jk�枨N���^�.sCuC߹.\���ƿ�����;_���?{da��t[�?���&߽}#��
�`�A���g�֑���I�Kq/U��r���\[C�2Ŧ� �Q;���#̶�c0���/��z6���{�����6���%�M��m��#ݑ���fq@=�(-\���L,i^O���g9T�d���r��0����3+JK���*u��"mL)b�|T��Gs��l��K���=Q��Ą�{L�9�nqy���x�z�Ȍn��~��|�Jq���A���Vk�w�G�UX1$!a��Һ�2t-�l3�S	��ݘwO���p����6t�� yY3Co�T|�fP̳�8Z��4�&_�61�~=���Q�>� 
q}���B�W��dZ���@=(le���@���=ͭ��zGRP}[+�¶6م�	�!��q�M�(8IL;����/A�ˊ���y3pr=��DyƐ�yDA�ӡ��I��1�UY8WWB?I��C����`�!�~�t���o����&���]F�$��;x� ������÷Xc�d�,o��f�:
�O����<��ǫw6@8T�6�6ϣ��g�g�ŉ>�0��uM����Z��uٸ����0"&��37��p��l]�U7`?!���Q�ӑ�m��'.�]�7i�6�9�t	���'b �s��r,)��R�*���fF3�����5����G�I���lF+���sj�UͨL����Y���m���C�>�?�H��#�,h��X;Bf��pϭ^o�	��Ӂi�ևj�N�g�v�����.R�S7v�o�eɴo�5�N��ҟG���h���s�;t�rF�t�^4���")%�������&]Wz49�zj�޽��x.�j��l:K+X}�U�}w�Rn�y]�۪�=���d���?�đ�5p    IEND�B`�PK   NM�X�/߻*  �     jsons/user_defined.json��mo�0��
������l�jB�M0M��8#�KJ҂�i���J;Pڭd|Kb���|�9���j���lݧ�LUݤ2˳��붡�zү�aj��|��޼��ڗs�A�hR�t�vW4)�@�'��ĳ<�K�jC�*4�(Ӆ.���� �u%��N{�l�Ԭ>n��6�-�dխ�.�y�cW/W���}[G��`=>�*��t@ǼO�ZZU�X
������c�l�P9�HY��2m0g˂94�J�[�.��eK߾y��.�1įç,��ES���u֬/�u�\��Y��Df�[!��YwC�ڟ�r齄`��uS_�75/����n.h�턶��W��C�
9����
�c���_ێVos�E�������rD��p����^�E��͇Ӄ|5���Fm��?=?��#>�Dv�h���� _��R9�yw4���v�˧��=��e�V��sgCk���[%�L�ϩk���RX�*Yt`�a�Э+RYF���Ϩ��d� ͵+=+D��� ��d�|��-_��,Ua�;C�&=x�i$�
:���&�g�p��O>ϝ�F>$�x��Y*)��H`*dw�{+k�5�� U�B���@e���wpIp'Щ���wpe7�z�T�>�=7�	�k*$J9ʩp�'rɕ����"���i�=�S��e>T���<�*��=p�@�������;�>
��T�� �6%zOl�Vz19�0��v�
Ԕc���MvƆ�"GC��ԓ�{^��J���D��k���T��Ɔ҉멏���hF=�h���]�%]�CZL�����qal�n����=񨿄��_PK   NM�X9g�s>
   s             ��    cirkitFile.jsonPK   NM�Xh��3�  ��  /           ��k
  images/3af811fb-ac37-4701-87db-865e720a6976.jpgPK   NM�X�Ɍ�� �� /           ����  images/53a6c856-3ba7-48d9-b0a2-5ca2401e7b62.pngPK   NM�X��i��  V�  /           ��>� images/c1791b9e-feee-4a68-99e7-b4273f4cd073.jpgPK   NM�X5r��W
 zX
 /           ��X� images/cccdd3b5-475e-4e4b-8694-ce23b104edc1.pngPK   NM�X�/߻*  �             ��;" jsons/user_defined.jsonPK      �  �%   