PK   vOX���l  %�     cirkitFile.json�]�o���W.�O�!�H$�wm�,z�[`��M`��b<^;��ۻ.�/I9rd��83I.veq8q~ΌF��Y��Zm�Ŷ���V�n���nX2��gM�%{z6��V�e�]��d�����w���PE����vSm�%���8�t��H�����q$+g,7R�r�f7������q����u�q�\��]�k�}���*�Z�(5YI�X��XG��d^R�R�yG�lp��#y���1��)jh�BcȕƐK�!C��\.,�^
�I�2&M#��"҆�`��Y�
�2��ɑA�a(�bc��i]9vgB��\1\�>We�M�GuY�H�"�Le��c%�T�_�1N�,�<NҔGe\ԑ�r���Q�uZp�s]1�ڐ����F����РY����Z� �]��S��5th?�QCcW�u��T ��@�"��@�C��"��@6&�/M��C�#b�0f�{
F��@
G٘������6��9fh2�@��:�@ �6fh�:�m=|������C�� �Bg!v�G\uh]'U���6P�EМb萗�ri��8Җ���Z�E͵Je�V�4��FM70�{�mCa��~��!�thea��^�>�_l���̟�)���I�.��KL�%!ᒒpQ$\��j�d��bHda^IuR��a�ր)�Æf0�U�h��A0��0��0�4l<��k;iL'��4(�4(�4(�4(�ť�c����M�q�Р�w���6��;&������0p���!�A��A��A����B�X?q��-vi}Cs��\�4�J��]2������S��3Д�y�B���g��;/4/G �E�B�e\�%MC�X�chB�|� �-h��ń�|����0saGfU��=fHvm�V�ɦڷM�FfH�\	I�%&ᒐpII�(.���!��h��h� �Y�f0�e�h�h �h0�h@�hP�iP̉,9�9�9�9�9�9�9�9����CB�bA�bA�bA�bA�bq��	��E��3$x.�ΐ�\�p�υf^.�Hp��,p��墎�<��:gH�\htt�f�3$x.-&8C��ry��fH�\���mnk�
���mv��|�e�T���:+�r��,�MY5��O��7�w{7'�B#CGE_��FY�QEl��f(e���<��
�C*��y8\w�y`�� \ச��U��(��E�a����y`�.Xe@��~�}\ޏ)��x˘�\3��S&����m�ݣ��T���Z9۔S��'+��y�wn��� �8��u�g/��P�`GGJ2IpD@K���)�J�*��˭h���l�qV�W	7�J�Q^ l��� ��%��"x	�	�(c���/ 6L�K��V^�= �h��W	��K�
�� �
^���z�/�i 
_!�|[zkh�ʬ)��M_����>�Z����V�.�5����_"����	��쯐��m�x��y�� ��ũCqʵac~�炱xgX�3,���Y�-�@-���v�T֪p�Y��cq�PO�&aa��PO�D�� ��*-��8�b�-N=�z wl�cL�$о�k��k���Q9�3(פb�O�,���e�q�
�+SO�a�Yp�*l���Va�\�
C:���
p=�	7\&�T�3� \�J(΄*Q��u�-t��^O���#v�.�=a�{M8���KcO؅�*h�,�b�Ų#U|�ώlV�K�X�;���l��onƜN�l�&9�9S笧3��8�{Xz0y�ka�s�̑3G�����]�z�[����w=���]�z�Cx�\�z�C����uw�M�]���J�bc�����=����޹k���#3��',F�46U됱��=:��/���W���84����������
~�^+���F}Y<��P��G�뎝Rԧ�%�c��5dU�8�@}�Y�;��Q߱A���]V�ǳp��c��=,d���_F}"Y4<��P�����W�+�Q�%�nL�[gy�v��	����Ϫ}�F;ia�&6n�&>n�&1n��&9nJMɸ)=4��&uhR�&}h��&sh2�&�8l<����|���`�	a�b�N��z�7UV�۬qU��v�^������ ��5k���՟��l��]U>����q�9��Awm���b�d��o�:�������>��ʎ0�G��헟6�[���:[�*۸���W�U���sM�����l,�6��^��l�����7Usn��dG1�Rfu�_���oʽ�c�/�{�v�j��3?�-��O���j.�Yt��ev����-�Y�K]2�F��鼈�''��u�J��I��^'?���l8�f��c
|泭��M�u���U�:XWm�/��L���㱊^tq ڱE����������T��`
���'��&�r�¤Zp&R�d7�܎/x��2I/�Y�����X�;���j?��r���u�b����@�Pג�e���Tt��CSgFY]�,��y�D���(�+��q^tٌ�����A��S��/����ps,��qw,Y|<�O���y���$Ohԓ��xު�x̞�<�G<ZdjI}���'*�He ���+e?�MS		��c^R=λ?�sG�������\ҟS�9�x�Ӌ?b�9>=v�O�'���SV!��Gd�-�Aܦt2E6��)�)���f�cG��=?��c*��?$q����������?������@��&�/7v~c�����M�hV�N�'�H����]N�d��D\+�TunL�:A��S��Մ��Hvǒ� ��b�ɺ�	�������H$���[��f���rȑ�
���?�Xo,e�45�S�v>٩sU	V��H���O\�6U��DT���ER���)���/�cw,IT����;&��"%�fc�a��+�+i����M��܆���S�*�����HEU��ʳ��(���\��o�ݱbl������B��)s3�~�'?-�x��=�_wL	�Xr�1�RX ��^��^�i�%Sl��䉍���I�s�B���R$Y7i�����Н��
n�!Kq2b�.a�E�����i��.@���7|�Sz��k�_Ve{oO��r��G~��G��Lra�,��[�6��������U�]�h�����U����d�+�z;�/�����>�R�v6�� ʚ��j��MϾu�U��JxVM��#�h����{خ6퇬��������\F���k���Ν�����1no��� ��=�zU����o��oL` oH����G�5��q�xWBc.��i�ګS�ϠR:��rF�j��LS����`���eW��� K�6#��D>�*�F�v ��e��J�nˮ�c�B�᥍����%�"bhd@�
��0Ѷ����}~�j*�V� �tX�ϛ)�
�^D�>�q�jZ���Hՙҭaj�~��j?˼��s�q��Ы��k������&W�"]�J�:8�0�ab3hFT!h�vBh4`����`h\!G���^K�1|@e�;p
AT]Bw4������P�E9R F��N��K)��a5����mQ�t@'ЀQ����}@��*���@���!�N[�a� ��n%�a��3��
����~�����bH�Aⷈi�d�¨�����8K�Z~�AV�N��C�
�p��1�휤�`T�@�4�����4'��K��|��{���:\�gP*gC�S,���1�e�9���E�-ء�B<$4���S�è��Ah��B�P��jRhV ��Р-H)�1Ŝ�H�Wy�ǚ�t���9\4*���|XG�;N��O8���T�<@�ѩ\��v��R�����T��UB*Su*weg�����Ǭ��U���n
v���U�c��g�ﶟ߷�������� PK   vOX��g  n  /   images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.png�xUP�u��{�;�)�AZ����C�I)�-����8��P��+�{���tw��Μ93�pfv�,B��*�  ԠJ��&��q��un���j�	 0�����z�Hj/�w^z��^�V6 ___>GOk+7>W��S) ��AMI^�/�$���Ġu����������1�6�b���w ����(:��9�A�B`hz/�抉���T�K����%U�0�2!54����+|������#�lI�)���ŶE��V�c����m+�h�@.�����9UF�*o�@��Qt&��t�t�DA:2�L��K�H�e0�j8"0��h�����A�a��/�b�V�D�o��휞�H���l	}� }L�~���>��t����|f?�Y�����0)�){��`��o5����1�䩩��-��&�{�6�P��54v�J*c�?Ν/�yޣ���;_�����WF��� �z����ܻ���1)�?�n��9[��j��U�Ҫ|[;9�K:�D"�m�R����7 쟟[�ެ�68��<Sic�"�lM��ljn6b:m�&L��}�pj�������\����ֶJ�U5�tޢL���n�l�)�ox;nx�TY �J��y�I�@��y?E�ʯ���zZ�Ҍ�w�;��T)�?'Q�63�������W��:�@��e���4�R�I`��V��ʿ׋[��^��FS��'kc��������k����$C��7HY�T���H�"n���v+k)6���2�& �gg���;�>=�y������SAJP��f,����ׯZ�:஀[�?�q���Ǚ�UGtY
~s��^�F)O�\��Ý.�`{��3��b�$�[��H�:/7(���D��Y4�zV����;�r�w�Jtw��t��iYuI��>~ɺ��%�^4%����o}�͊��!b���k����PP�N�˺���y^�i���	?	�<��횇
���<疗9ϺN�s���Y�S�nF��r4J[���松>���]!faU����3�:ːG�q_�
���?�君���g��fٮ��v*�	���P�������)��Wic1�&��
�*�QB�#}�,���Jt��Ut6�c�Y�RY����m7�dgF����w�9f`z~���������4�)�n2~��m������遡`W���g'�x���!���+�y��Dx���/ǚ솎q��0�ط��S�<�+�/@� J��,jnn6�FB�YW�1�z���0i��,[����zUiQ;�D���ϽL���HN[��|o�����\m���UU����@�Q�������g�3Y@�/���Xޏ�w;�s�n�%߷�WtMfI�0�c�IUr�{��K�����a�u:S�a�n|�IY��ARĈՈ�:� ����;4�JMP�64���g �6\]a~��u��E��5M�e)����N;�Y���@̬�{V��ɫd}<,�� rp��!wL]ה��V��`�|��L&�E��LJSKy� ��V�;/�w#����(�.��o�L*��P�,���L��f���n*��/f����k�M��C�I��V�{��f�9��e��x�Wڜ{A���S�z�}������:L��3�DR���5s���l��x9�o!�b��9�!��9�����ӖJ#v�2w48SݷwӤ�Y��VL�kR��NX�I��w�L��/�����}��ͧ���^��hx��x��|Ԗ�+�鳵�	��H|:Cu��*Z��j?|8c�{�|N�1)���.LCCSu����L���(���(]�:��@-�/!�7�?�X��M�-�p�.Jjߺ$�s/ls͂��Eg��L�8�:�?���{t	)�|��V�~ܟ�����n��Lu	�gAOB�����Դ��>
�g���xԂ屙�WȖ ��#�!��{�8ğ]�7�F�G}^���8�xڎV+/��f�}�X��}�,�<cj{h,j���~f��gi��Z�陟�`�c@�3��8���`̂܇�7�7+R)wQ6����"z���:�*��F��7�|l���nI�o;u	%�_�ۛ�?>܃�Ѩ&~�	 ��:#K��6
n�F���4epftg��(���Қe��M�o�#�a��%�:$�O(���SH\'dn��DN�O�)�Y��"<����?c�Ǫ���	Y��;���ª;�lH(�)x[t"�"G��<��㬖�r®�k0�&�`��C.�"0��<e���a��@�^�c��",N<�s�9q x���f�\WOL�F����j�&l�f� �����0����=�����	�@L�6Y�Ed��Cy]���N��5?'?_���Y�q|N!u�ʜ�s��u�N`}���$~��g��^�z�qr	J^b�e�T���ouVT6 R �zynZ�e���ۅ(�0���ȗ�<Y�/�hm�K6`ϓ'�L4a4��{�щO����������"�M��8�;>������m+2/�O������2xS_:x���S���P��A$�޳�l�ϞY�(���5��l���M�'ק*������w�}�����Zq(㪯��ϣ�,�݄1��-����E�w�>�k�O��$ܗC�@x�j�]��O��'N�TY���"\���Q��K�iJ�y��1��欎|��q��b�ӽ�#W��T�Q��ݪ�6�E�#g}v�\|)&�Π��!��S�y���k��i�$��f�*����˫"T]P2 Ȧ��$-t8�j�QG �7��XV��#�{��L�v�&g|�|�;I�Q+>T�f�b�+��s.�	�]t�ۃ�cm]N�û8��z���׈0=XX���8l����=�]��x9��^$9�m��r��/���Ɗ(Nwn��X���Ea��z/�ejǫy&�G�A�1��u^�U���e�Rv��	A���L$��t���k󴊧b`�x�`�`m�c�[m|�q����%�`���tl&i��{CwC�W���v��3zB��/�0
�}���j�FχY�e��QeUNh/�e�违:����y��',�[`�Є���l�#�w�-ܳ�ע�yRx�DE�����.B��l<զ�	�b(Ι�O���5i�K��Վ���R�'C�2��Ut��v���R-�U���H��Sh��W�\h�a3Kf"!N�PyMlOB��	��ɦ��T~��p����&��.��`�|S�����YP�H9B��7���'67���!�2RT��l�K>P�����F۞)/���� y�I���I� ݺ�
혷7������v���4��YH��V~8�(�y�E�l#� ߄ϲ�̲�'7@�eV�M �:P�����D���U9&��*(h���p��`�V������Z��ڎ@����Wu���T�xhT� � �ɣ����w|��n�X����7��`���PI�l�� ���}�wd��.�Dj�z�P�1�sB���E�!w���Q�(�����z�Y���H��-S+����D�Gb1N;h	���4A���	��73o��Z/	[)*�PV�"6ӱ1S�$RϠV�+��_��A�>��2;DU�l��
r'F����m��;d�7V�+�YW�H����4��5K�/���z:©��/ؐ�O��n�w���f�eD��<}�?�Ҽ��_)��dz����"��Y(v�+cZ%,�`�UH��(4���ٯ�P�e�+�靑A*&�4Xf�%�#��#�(�C Tq�j�YSu*r.������K�<>5W179>G��gf^~�Xݹ��������.+Ը�.��� �	Y&Ic0mu�]��;LlV���ֆ]2a.�|�K�FE[o=�a4�X85�=�%�P����V/AK�Ndb$���
���(2�R��t�b������ޜ��R�~�kbs�ۦ�]�{��&S��Rk\B\c��#��o��x��cK�\ۖ�1̥܊ou��p�rZȠ�xu	焝��9ȟާ�F��|nG|Wo�bhp�Y��`��sb+����IK�h�=�6{Ǚ:_���������ߍ����B�"@sMGK:�`P�Q��Ls��A,p|��{'�ڤW�/D?EWp�c��؊�o9M��
��M�'�c�{y�z��e�#�F�l<�B��]O��%۰O%��<r�e5C�f_��!>�ν���g��_��/gL��f�#�EgN()-#\$�\�Y���DB>'d�f��d?���@4�7h�
ǉ9���x�5�������:V19q���WxQ $���%��56��	�2��ea$�E����Ғ	�tlRh��`	d-f�Ԓu���:&�h�S�3��я.˨��v�ٜ���j$cT��	�$7~U4��Βy���&��=���Y��!1b({�o��rz3Pǌ�:֦�<G4�R<E�e�̼螪oJ�e�=��{�ތG���#��Mx}I�����G���1[g���X��p��ѥ,ߋu�e�&N��<.Y�WNH�k�|c?��M�
�t>�,�s|�2#b��-j)�������o?�ǘ�}�U�ˉ�V.f^��q�`x�9��K�!m'�������7�-�QMs�E�`λ�_Nz3
?�;�e�͊��~�]T$r�Ɗ/U��
}B^���c�k���~���7�jF�.l�g��^pr�3��+q#��)������{�{�H��C���c�L鈈�B��\�c���ġ��q���jh���@d^�Ѯii{���;p��e}w9��l�����YT�'_!ߚ;���¥HfH�+�2k�5�ASF�j�ʙ·P:{���s��	��d	��pT��!i����x~p󂭡�RS�R\o�"V�XLq/	@�U`,0�������""����*܍u�P�xC�|A7K�e#,�b�m��:��*�8�NB�������X��[���J汁w?���h��09qװ��~�g�(�5�׭�F�J���_�J���b��5Ƹr����z:P^��kϹI��\��7��������%��|�SB�/�[Q��"��ƚrK��T��(�R��T#����-K3uwUi�4_I®g����x��t�S$/�������v�"'V��c���)ʮl�R�Fp�I�xrQ'f$��[������X�%Z)	��t7^�RƄ��g��:_�ޘ�K��������.���*�|�!���K��s�?��Rl9g����fr��F���f��J�CrVZ��_�S���!�Q�̛��D'~�A����W�E�pP!.QC~:�/�y��$�c��3��4��֋��ULM��W0Q�v#�C/�B�9��q�=�݄	 S���E���}�AX��a��*� WMa��ə�qOu���EDO��k�ء��NF"|V1r�>�R�ʨ+1�T��@	'��x-x��ˏ�g�ea�{&z��6=O5���p1c���X+���cQ9bǆ�����dj���[���d-*b|Hvցޫ��i�zeG	{i�*.�P�a*`��!���]}߷NM:V�hR��~�
�v$|�RP����(����'�c{!��8�[z��!p`�����B��۟�֚�-T7!��0 ���A�Ԑ��@�$�9	��#��AV��ZO�TL�����N���V��@�2�x�M`�w����@T�'��B|�T��)��J��o��))��9)ӢD��s�a�!8t��le�%?'B��p���?�F씿��������_6_=UbkN��Mj��Y�d�_|�{1D99k6��Z8AM��ƪ�����rF�Aq�� MWZ��m'FM����;-��<|��t�mN��a��O߰�O����O�',���;_�h��u���sm��$W�S�HĊ��ԅsv�wث
�� ��2E��4���a��y��ܖ���䒺���x���X�>/�X������w;Q��kG��J�ի�q �6ǰ=��I�u��F$���س]8���3�F�j��)�/!ݲr��Ք��4��l��hgf����c�&�IK��6�!�Q0���x=��]=���,��d� ������0;����=��i�@w����sk).�sOvA�y��W��oh��6#��Mbۍ	Fm�����F�F�2��PK   vOX�j�� 7q /   images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngT|	8����R�$tN��J��%������&���-J�"KB�}(�JY��6c�!��G�I��g����*�5��y��~��}?zz[_���&&&6�׍��X?01�9||'�F_|:�����a�t����_�7-���>R��ku41�<�y�������=����%GW����������U&&!&��&���Kָ�ލ�)�N�>,ie�8z�ｰ�Q�>k���]��cr�c���e�kw1Cο�n�r�<��oL���G?[p��?t���7F��J ���}��)�u�������T���%�RtHQI�Ly��G"ovf�}��-��4(pTr�}�һYH�j$�A]�`��eE;�	��݅'�b%�ĦF�lt/�DP�����d�����sՍ�s���-�����/y �ȻX��e�g�П>�J��=H�m,T�k��kT]�t�K�H�`����k��R3�2�Y��O_�{��X��&�T���]U��+�^v�����sq0��96]�D�,潕�d ����6h�8��Z����-1�r���vsѱ��b0彄c�@��)��|�,Q����:��0�����o�t-O?�1�rͮĤ^h����#���M���@�g�p�F�(�J����pd��k=r��{ �zq��-MN[�]E�>Ò��!{��y,��3<��i8^j	G)�P���ʉ!!��[W�JՖ��N�����b���4|���N���.kK��t'w���$-���##��0ֽo��A�k��K�^/�u�w',T��}�E�	�i	��O� {���+m���.�����bmic��w��1��c+ۋay��؜=��H����:�޽[Y�^ȥ ����m�m�%{B��|F��=\��뚞vW[���.��h����?}n���ג+�KE��[l@ af� ��2_���X2�	�n����O�~����Ql���)v'A;1��7�}�Q&��&��#�d�^J�%�wxϩ�"Co���^3��ٮc�$�4b�K���#���e��ʴ�'z����f����7��f.o)��4�;�%]�'H��ĳXRˮ4�������3�q�H"��H�b�þ���BG����;���
��b(�}��De�0$��H��G��j �� ��C�*��X1��D�eE�@���]�,�m��*�$�QB�g�X�g@@���b�q����j�x�˂��ـM��BXep �r�t�ʉI���s�n6H��Xi�"I0��|,#�&��t4�/&wͲ��$�����Ǉ��T�iB�f)s����9�"��'����wB@#1�[�H�=�Ge���y���m��_7�:������ �����A�`a�O�eMS~����&��&^�N쀩ϻ�oʴ�D������$�(�Ѻ�CbC��<�t����G28�H䱹C�xK����� ��	���tw5��D�b<�ˏ����"_a�B� ��B��#�D����ŭ�~�~B�`�@|)�Y��r�L&gIϕw�57	��Z��(F��<W�g?�L���fz���؀g�]P�S��í"Fw�JLF%*R}ߤv�'��L@ri�%|\ǖ�pb�d$�i k�w1�T�Y*�,u*^��v����6C<	b0!ּ�"`K���7��C����Mlh$q��|�@�%6-"�k�OF�&�~�Mԙ]_�0Ҟ�Ԝձ�5���ќ���8vT��d��a%�8�r��3�N�Q\�Z�1:��N�䆸�B*�qx��P����t�@5?��_�0��*9�{R8�q�A����u��E�c�bJ��z�J��D�N�S.t����B�@�/�� �gh�[ [�H�����;R���So''�GqK[���51ӦT�/�����W�*4�k5���_a{H��^�(u��:!
-���Ƴ[
�,��Ä	�~X�aQu�~��p{<��S����*���詎?�A�-}ۯ4}	�S��bJq��pCLJLL�+)財E������[LA��VJ���D�Yb��������ހF{����A{d���������@������_��mQ�C�ԃ2$L��
�FZ��F���~M��q#�ā����׎�7�}�ۨ�ѕ�Q77�����mV�+�ҵqҡ����z��J�Oco�i\�ߐ��{�U�>�l��|��o��!t����������B8v "����>��jF��F]k�\�ʐf�c��1_����ٱ���K��I|���NG��1�JLn��/'�*�ˡ��5�-ڀ0r2={�,��)C����/$��v��^��������ׯ�n��x�����خ���kKۓ�N�Q͙�B��a�˟�CN>�z�Dlh\�C���nJ(Q��������6*:JNV�<g����5�Ԯ�x&�\� J�j�jltۿ��RS[�@"\k���+�Z�]i���GG��i�VG����s�V,a��F%�U˒0Bsl�!���U!;��Ш$����J����e��z�e'$�ܠP�U�Zo��jb��j�|��������9��N<#s������Yt�����B���҃Z�&�!,�(�<uj�c�8���b�ɦ���'���<:::87WXS#�@ԕ���/�?���N�����~jnǽX;f��}���	���Z�*	iދk�}��/w�r�T�����q�q%&JU/�M^��x��u�b\����QфYÄ����n���S鹈Y�Lmm-�P&+mث���x�-h�n/7%�!d(Og�q(v=��E��<AAL�ړ7�L/	v~`rw
~��ؽ
7ӵHaS-z���#�b�C�cw�%
�U�c���!����&�y EnH�GE�=�*�AA�^�sjR ��u\�0p��,E�b�v�-C���������������~�U��B���?ںfDd3��yz�*��k�QY��oPgnk�2o�	�)^k�f���:;�=�����?����	1�����];OI��5x\���������yډ��(�1ٶߔ:����,� �t�Q=|��ufu��a��]�L��/����jj9?~x�%�A��o�q�DL��=��Z�x_W�8'Q�2f	���`I��P����?��8����d#7�A�?nA �x�E���!el�%�4`/�����:�!���uZ���������ٶ�Д������D��z��g�4�l����q�Wf��?��bd�~�?؞�`��!;>В�l�1EX��`㤱��.pr>b�.�3ҵ�w�1���L^�e�h�t/�>����xezi8����KHioo��U�|09̤�T%>p�l�xk��S�#�ѣe�cɴ�6j�5+�����6k1��l!����D[�#+����=��O������C�Ш��}Lk��dMˆ�#�X���q��FN����9�Q��I���k-i�q$���1�s�q��%���2��\�6*�Z��.�%$@=�r޽����x��1_�@#�����..z�P! ��"�q,kD ��
���{��_�q_g�1�����S�@B����ܛ�Ǐ;�ʪ�Wt޸���!
ҧut(��9Kc8e7��3���Z)�f��;v��iK�{�4=�'zY����Kr��6��ntaI��c�y��?��Ib��acK�=z8��x/}^^^K+h��]S/S��7$��iIr�zE��5z����Ծ�h{���ݲZ�gDR��Ӹ1�?U33�3	����J����9���5���[��K$�Or����:�������Ȼ��H�U/�G�h'g�[ ��i�3�!,W�B�ϔ8�"�h4�=�y�c����o�)�F��fb r,��>��F�M�>�V�C�Ղ�"һ��؁��.�����8��9��h�hGק����9ɛ�2␋@�@��|\wղ�9ğH	1��l@e���Je��.~���{��)�2O;��x��n��9uXY����k��ɽ.���#��5�IW�+x!��,IP��߭׬�|�TC��~�-�а=�J/萭��7^�?^VF��F^Ώ�Y@9d@�S80�j[����̇�3H��mi*�Á�氄����/��k�t6�:¦+���k@q3����[R��:�����<=udd@�%I��ef�|DM�ۚ¹�R��TDSSȣ8���'��IR[��E�6�m����0M?����%�^�XX�#Lл<�ƔRP����O;8P��7��������m��t���w�l�^(��X�U�?)V.��@�U�c=ӊޛ��Г�I�e���m���:ꅎ�O����p�ף��*/�mi�tm�w���nsљ��OY�������x����F%��N�tw;� ��B��X8���>��K���j̵��M*Ss����+��%�.B*�3��	NM��E�C������|a������n�����m ߙ
��N���u�X�!ݒE��B���]����cZ1�=.1��jnW$�d�����[Ub��du/��(�"(Ky
�n�d8���ŏ?^���9���R-��fk:�q�Az1`3��6��L�Z��XrLa����r٫W����[� ��D��}}}n��Ds����k����R�4��vn��M>�<@}�6�4�"�~�'�z����/��OK��fwl[;G�X�H �"%5���@��K'q�*�z��K_��"�����3�+����N���*��Ռ�I����m���_��to���e;���M��
ViVV �.!110:��Hd��垆#��GC��X���X���^�/���O`2����Φ����*������D4�=��bDDc�-��ì��m����XjK�]i�}@\��=��O���S*�T-#Qu��(6��K����/ȩ_������Q�xߜ!KLbJ
bw���UW�
�����["��6[���x�!|�0gcs��@�/g���.)}��+^Xp��xbg3�9+�?��b[&&fy�r����9m�{刧�m�X�=���f�N������0����P=qw`�&�7S�GAyoO���9�FءBr#�	ai9*�PYY)86�>Y����N�q�]`���3�g)�c������x�n���R��PD��v��A���܁�>�UI	�� ̀,�Hl-{4|�(�c���lA�b���x�M�k�P������)H,,,�So���9�i�}����ـ
�C�g���a����E����vK�G���Ǿ�@�g�!��HW�R:�x7��� �R��sxb::������k�A�8�Z 
;,�ĂM		���_�/��5���i0�����UF6;�/���qAF����J�`H,TH7\�ۃ��d	�C���sU�T�Wj�R�(5�3d��g`p��c1�?Y�|}���E�@aF*j���NCخa;|r �DR���|.������"7�l]%����V3�l�]�M��\k�9��y�1��#���i)��j�%�\�Ç�pU�P��U0_׫�RW`U���#��{��M�FKWShC��f�H�x�_(Q#u�H�;��_~U�K���\" ���	eZ�\��c���0��ᶺ�3Z�����$:������8	T{�Jo��B��
��^����獋���Rrm�4M4S�h$A����
H�����/O4ѹ.:�����?�2�p��;'	+��@�~zU��5��~�r���#�.b'�A�j�>�>y�-����&^x�S*m�ɫ1�p(ۯ�2�l�3�q�o�Be�y�Q���2��ͩv���rpB�v�Y���[l'P��B�C>�{�St��.�-��!g�c�.	���!����73�OW�UlT���_��ڷ�G�ro���*�t�6V��p㳁�V�����-������_B^�MӬ��#�C#u"B�N-z�!�����w�[�0a�9t�r��l�RD��Pi����?|��g{\��WR$&7לJɣ�ベ~�D���\j��I�Ek�	�����FW����O�*⛮�nHnb��8���^��\J}��A�Cz�=q���	k�6��-x�#k[���MV~�F2��t�p��*>V�Ua4�ܮ���0-0���ߛ���ⳁf��0�p��6�mBl��q75c����M�V�o�X�v��hd@y^�U�;��)ymg��4g"m6��\���q4}u��\�V�Y:���l8q��򄲲rW$;��v1|���O"1���J(f;����ߙ�~6��E���ףX4K"��P���Ļ�d�ݫB��^؏��g�0���4a"1M�`{�`�qD5QO���:/����qqq')b]��u���H͉z�.��]�`o�-���ɲ�$�D��v��0�&O\�<K���FPc�G�C�bQY�e#u��Z�)�xq3�a�nue@<�>q$|�V�����]+-��W��a`���;*� ﶉ=��bY62b���geu���3̣�������+�ŋ�b/9WH��h��_���.�>�i�Z�brk�	{��qs%��3zz�;���˿�8} �d_�M4�����%
G� (���� L-��Ѷo���d��O5��b+�����I��֓�H��Q�B!��]�:1�ߟ����~o$�hs�͟uJ1�Yy&&Wr*Ի��Gr�f��D�Ի�:<����_�s�V��p^'�ב=rm3ǂ�cr	��{5o?�F�p�.r�R�@;YW�s[Wy#�T,}�x`��}*��%r�u����o�BWl}��+���%.y�;�ЫFE�;����N���>`7��z�B���K6���^t���y�Y��,i�s���w�r��A��I29dϖ�2'�50��P���< �$/��9F�xT&&�Y*��f�w(oa�' �oKL4z\���"�Y@C�����kmg��݉��:���bT��y�6X7�k���Vɋ�g�|~N{=�P�}f���Gc%q��@[[�+�C�U�k)�p�� �t���$��{7*1$�Q4��������x���+�|Pz\r�m*�>E>�w��X:�d�7i�3`�%�u�~�!k�^�Y7S7�RVL뒩��%�O~X2S �',Y��j1�*[`%��s�n]E}��5�pJ5��)��J��UBg�D�}q�gOA9��jp/���ID�r^<���F�H��l��'�r��+�&�RĿ�'dU�6&'��Y�\L>���NN��k�5�|�C#|��:�d�dP$1��L`~��<�Y��Q�e�NJ::�?y�U�ci>�<�N�u�tQ]c�l��§�3S��"����{��m�c>��ⓔwḑ��|��G�E�+Ĝ�l���(W��$�O��k��?�9:2��Ë�n��Q���!I���}~>'H:���URG[�\~�_�k�������!�	9.��XY= M	�!1y��x!T�L$7�����؛�>�%�k'&uc�����[%�K�~��ȑP�oT�H����1y����z�����'��eJ�4����Ѣ9��`w���7(�,��
��Y�)����k�Z����̍�-9�U����Hd���+�0 �#���`�0x�?k�4��.��I��u��e;}�d$=��u(��YZ@�_�{��kj�Y_9�� �?��o�D^�<J�V�s,v�l����I����Y�"p���u�G���_g�}��FA)�"p�Bi"�W��aX0P_>�����N}W0��kXrwT�)U��D �Ĵ�Ĥ��Gv����О�
��B:<<���kIz,��r����c錪��+��͆ʞ~��o�i4`S��~c�S�.�fj��^:�P<���<��pn[_k��|�U�K��:�(tؤ���b��	���D��p���{Z�p_��+��Q���Q���u�M�D�#��PW �Ĩ�w \V�D���� �c~\B�RA�R�J�YA
��E
�i�^y?d�⶯���A�oҏ�/�C ��.4c��JM�J_��-2�5&�S��T���퇿�ª84�=D_��ec+!�P#���;Os畁FMP�{�ʼ���hVE&���������+���FF��+�M�[�9��`�k6���cY���[�	�>n�c��G��}�ޘ�H![kW0���Oց/rNV�� )�����̐�֠}�*L_���?-���E�~������y�u5�Ǣ��$N��T���m©I�{K[�B��-0���/���{6����@��%�c�6bB�c���Q_�Y�{,���$��+u�gu<@�gǑ�Y�����c �V\c.��Z�7n���}G[�D�}Y	[�������|5�����Z[Ƌ�\E@}�IY�?@�}s��&F�#�r2�H�U��=!����z��򍓗<Eô�N�\�����.��"���Ȕ{�s��L(7�S���ؠ��?�Ϊ70=�u��#T��ЄWTp^���;��b����c�Y��-��	��̠���h�١-{$��KtS�Te���1��$
��:�"�%==l � �F)����J
}�b��_�]��z$�޷LG[��)�� ���{�Ѿ �����o�=N�b�. uۃ��O�k�Cpp'DiQV}���,����Μ	���PH^�G�e5���4N%&N�eY`�M�� ���8*�� ��'{�c�"��7p��$|ڸ&��2�C�C�l�G%��x\~'a& �ݓ c��ߛ�w�B>���x���bv�9��u�����;�^c$x�om�ɍ(?�5�5�@sUUUy�M��gD
���VZB�)���B4 .}���5�4g<�np@���α�@�7^�m������}��κʘD��2���+�u%�E2���A��bA�M���x&��2m�����A16�[P�����+;�]�Hu��u�}BK�t�9Zm5�$���<Q����@W ��_H�)N`���R�Q���	���A�!��f�/<�Ϥ��GEEɪ\�}�z���d�r�W��x]�ɬP^^8%��@��� ��_�| |�t��)�x�z,�^����,���~=�o8��H$Y�ښ�!H��ޕ���,3�~�(��#.>�r}���O�^�5ꗉ���Rfy����.V���p��k.@����γz�֝>Q��ת��jq�F�C�]1�IɅ�.�#�O��+��C�)ej��gR9���ҒS�/-u�;i>-W��[���~��m��
[��BR�ɨ)]�c���j?��N��/���<��Cl��L �����$~W�t�hеV0yc���,�`��i�� �y\4(����q^A<���᮪[WܰߞI�m��Mx�����S�z�Ma���n����<�h>Ax�٩m]�^΅�x!}��)������tB�>[��o���w�)�o+�l8�@^b����Y#��p8�8tŗ;J=S��C����e����Y9�R�>\���י^$'�S�n뀹Sz�nq%s���XW�S��x���(��|?Sc�V�i
����'�'��4����$|����giNO�-�e����f?b����� �=�q�V�����K�q �D�����!�§/��������g���:;|�^�r�p���d�#�2)|\ܪ?�k�p�0}�x�]���i+Pպa;�j�/�n��ST�q�u�iC����ދW��m<�S�8 ��b��ղ����=�I3���u��kYx'zk�#3.�u�E/S����Ew��xxy1�?�w��y9i��d���[e9�lV4����ւ�SMC���U�,�c	�`,!t�d�ᮧػa	�7�r�zU�vv��פ�������t�@��d	�Q��ge
37�d.&��:��GP�����_���������Y���E
���m�k�;�x�r'MS�kn�Qu��A��^�Ҡ��������_�׎��C�[�z43t׺�BeC�9�����yTܗf�ʱD���iy�qBxo-��{��M����+���(�W�M���FkW����Me�>��e.��1C� 3�#Z-�G�Xt2i�F�%C(!W�EX��#j������OK�ǒ?0�7t������H�Chm9bO7�^��
l���9��n&~�����Ŷ�_w=[T9_Rt��D��	�R^^�rQ2�X��c�E"S�d��_����w�r��r��9B�A��D����6�Ča@���"KE�=���F��0]F�,p�y��f���Eݛ����_1��c֏�" -�)ht���9���\X��e��w���Ӝ>������B�*S9p���
��.GL�<�@��=�ֱ�/ҏ2�DbB��n���V�Fd�������?��F�D-|�`q��x��c
���[ȃ2f�i��]ڗ6JNK�]�[|��viuB9pj��)88�21L|L���<U!C}U��Ω���~DI�
9�JZ敻�nk"?i�u�.�k��z�����^ʞ��l*�`�qm/��LK �����7�߄�?{�������������O;��b<����.?@ �^��P' k�ڹ�zF�4j��A4oЏ�t��RZW���!Сx���I�XЬ��,������K����ʆ�7zՋ�V;`{�A� �ݜl?R���H�_f����ـ�2�X�зH֓[��n��6��ϸn ��u��S0�c�WU0��)�n�'E,��]��]W�h��6�;�zh��dT�������,�C��e���lޑS7TBˈ�O�H�g(��j�r�d�?>����r���'���>&�Xi���ݱ@1���o��,*3�ѕl*���G��������p�{�Bd����5��9$	�|!s�u�VU�03�n��|�}�D�ggI�6�_��e���A=>	2���ze�g����ۤ͝����/rS�M��$���V]Y��;ԡviu�:M{^�k�Lc��a��d���1�ßΜ�A'���ڢ�{����$�hB�:�/u���@���� ��O�"}���ݤޒ��|�X��I�ORA敘k�t�^���V�Jo�t�$��Ҭl�L�bA�Jd?���5E�QH���:�����:�Ҝx ��s��øW��ᣔy!���{�U�h��\Z
�O�����OR�����h�,(p���v>S�O�����8z�pU�����hW����B��C9�"�I�w��3\W3��v[�Q���NM��yv���#:LC}�w��v�m��o8�bMB|��+\�e�̲�IS�?
�mZ�� vOf�&��Hj��-=G]���RQݣD�*v�]m�h;�]�IT�;�9�Jt}Lo~����Ӷ|n�z�Hjn��'�<���?�Z���*�wֱ�`����������s��i{�o���Q���9��>�Y$fe�v��������7�_��� *]kL���I_�mh~��k$nk�o��-���@r���o����z�����nb F*�l�S�̘�z����""��	5��5Y��㣣�A������b�]{��9Z|5��=-}&����a������@]����=��M�lt�����{o"������	�+�X�#1Wj�^��KH�P��}���>?!�7�	���f�Ny%Q>F��\@P5{�0?�����ڥ�@�4�d��Y���52�����Zn�;t�7��q�ӯt����x�+��x��kBR�bO�r��p�m��&�j���V���&6��3�,�~��p�OE���@'6�d������˶����έ3zz0�yi99��j�a�\���V�r'2@BR�\&��s?SSS'W׾�9����1����a��
h���)t҅��x{��i�P�؀faW>�^E���[��3��0���;�)�8�o�~7�O��о �|
�����x�l���,g�����P�|�i� �i�u�wR�X�A���!�D������Uν!�G[94_np�@ y�|���0�\5�����Xh���D�܃�uW
]U�߾e�͑�Fp��N���k>O(�y�~-(��ƹ��q���c��i:��#����&�sE~�Ĉz"oP�S��q�Z`m�ͱ�����������"� X.,��Դ`.����j8��Z%.���^�����m�,��\R��X�؝�B������NV���͝O�$U޳�����4��W�83��_ۊ܎�<����ӽ1�#'ǑJ2>Z��<�-����|j��<jG��ER1~C���ڔ�m�Z��>ɂ�[�pQv�1�e�D���Y'W�N��&�_�rq��]Q��u���O?�?�a��/�rlt��
�0��k��z�+Es��
���!JI�A�	���c��qrjj3���n<�@/�==8H_)��&�p�&�V�&��r�������F�
��k�v
�pB��T� �� ӊ��VYxdhp0Yr#������4�����]a�����
LqIIߋ���ѯ��uzKAΜV�j��
�I�����w��9M�
S�$S�,��_1�t.S'������T�֐�^�z������	����������+�[ih��Պ0��j6��2����D��!PM�����g��YS���EXZ�������'�5����gh�,�{�|Ҁ�xW�^��4孤����D_٬�Ԣ{�n
��^zNkZ�ƫf�/RBqY��/�/c�h��z��v�tW�������Q���WRZZ��V�0�ox�����E�֪�a��^�����\Ta�V�G>��Ê��YDݶ�7�U�f����..�箮
���7��j�s��k�z����, w5KNV��4a�l���蓶�'4�1oŻ>T����� ����Q_..Z��?R��{�SsϋSs����TيV�����'�@`��rd��D�\�����S�V�+���2s9U��x��(�����F鹽n/�A��!:FfZ6��s��q�g/*�a��������;(������H�ڔ��F*)5�х&�E{���ZYZ�#�g�_e}���Њ��R�����&{��\F%��z��J9��ck\||}:^@D%F��p��[Ѐ���Hs�����Q��n�ȣ��ô�5���q>���[)�R�#u+/e�q��Dt�>v�Xz���F�}	n���hɴi#,��Ʋy9��C���?�ySW�7�57���1����3�� �<	Xk6���hA0ƇE��DZ��3�0#O� ~Q�8=�_�bt�>�v�ADMM��+Ǟ�[K?�۵���UD� ��9H�k�W}����(���Y�ؠ�����	Y��~z�Y��\�*��"���jԡL#@�;��G�'uΣ�3�S���U������L,,^���a�J��� �����<~|��TS���VF�ݘo�G�ƚ�z���jߣ�	��M`��Z���DJ;��S���+(�U���ߚ9��My#u 1�G���))��UTT���t�X���}��_E��x> �<f�͇of��[���ײ�Fge[| vD$F�'������R��hv�De �u�x�j���j�j�:�boP�.ij��ϴv�B�E�)S�����{L��b?��x�GM+Ԃн�V"�੹{+A�����"�9�Xi�W~�������Z���9e��2@"@�9=��B��$2�}�qYÔǣ�.���yV:�ޟx(�d�.
�nM���(ef�Bh����.,�|�g�ں&��#cK���bqu�V�N��\��gqql 2�@'��[J�u�HN..��<<�I�}��Y���U\�F{�K��[��w�T�܃�s��l]I2O�W$D ������τ�Xmd���ˏX�v�M6t)%WD��]�:���� �ޗ��D�J�5�#w��ź�{�j�S���.�ړ���*�&�u,,F����"y��M|�N�`P���8�a��jPq����-(r�Z���Ļ��TaC##��{�]X�|}�0��;ø��� �<���[*�����<�0%��P���:�S��^�;_��������ȲT�Do����V�ogUz�A[RRn��!�hx4�Q�N�β�Zh]��| �X8��C�moz�{���h����k����������#�éiy'33󟫤�H�4U0��޶���P�|�}Krs�,�M��-��T|�b�U�	��B��.֞��Q�!�l���1���T���eJ�v�>��KL��W?�KH8:9�k��dikk@E��%`<�^�-o��@7T���m����έ~N�C�zQ�X��}�N�Z^����8&&�`��u���p%u��ř�}Ch��2[����o�JJ�'�^���7�#����>y�(��U]���X����1���j+xOD�+@��G!C:�����񹦔���"�NN>�W&$q�W�W'�:;���"��9;��Ղ�=��گ8<�Ijp����N��qJ���H��&$o*4�0Etq1���&A��W�ׂ�N���2�N��漇��_W��U�9Sz�ӧ�~.���ލAl_NE��s!3��R�>��|LaQ!g���HХ}�P7�A���`���1KP�\ �����,�j|־�m_�";����C&�0�����}����T´,"������^7.xF#A@m�@����G2%��
��˯�٨�h���=+�W��x �����%���(y�`UxI�E�[�����h�k�R5XYYY\P̮W��������� l��,�~5�{�_��Ƞ��_�ȠJW����x���]��ߙ�lӥ�k5�,!��Ԥw�j��1-fqU-{;����7�o��,R��ŋ��mT�,�f�Wh�M'V5S������\���MRG��95MGP��*�J�-\��ÁޖII��3�{w�Q�oջ�B)��"-99�6��%PC�b�r�2I�@
��|�@s&�G�/���1O�}!uT��(;��jPD`~��[M��g8�u)��?E�X���yg����y�Pٽ�v����A�T�:b}&���A{mmm�Y�i:�����pXk[G����H���`��� g.���[7�yy������gZ///�e=1�T����|���=�K:���mР�Q0����{�5��.+M��-&�@Rw�݉�)�ʄ���w3�d�DvRO5p���th���Uh�d��xys4��M��\>�f��?<\�]��Y�k�P���i��!�����|�}H��S�x�%��_�~y�M0���Ϯx�zp�8�M�7o�� ��L@?�x`�ϠEx N4�I`|��bȫ :%*E�M=�a��Ӷ
'-�dz����@�H?�����Ĭ�]4@�����V�A{��b|Б�jAw���;io0��x��ҷʩ}��ā��I���=-������;+ |ՙp,B����'Yގ� ���hwu�Q+´P�=�����{rRc�C�j�j+M�X�����T�k]`}>DJ�r
Qo�� 4�?O�'�խ9㶴����n�o@��^s�j{�rek�3�*���eJL�@�=ff153K�f�__��d[��1g���ރ��hW<�,��e��0(��^��_�RR��2��bb���������i��^l�XR�0�ｮv�rY�W
���	����xjb�E�����DJs���vM��S�KG`��h�/�5\Qv�j��UQ�s�W/�&s����$��׵h��ۖ1��j-#ݮ�Cn;n���xA�,?>|�I�~Q��q�$B.Rq�|��~���k({�^i|���)dė����h� ��C}�u�dŚ1��fbfZ�=3��~EC`�����P�3��D{H7Qǲ��u�Г�.��Bh��zj��h�o02�4O�3��pGgg��Ӑ�.Ӡ>�sc
`�.����h��ϾރBͯ<�)���A�*��9�'k�<�rm�:�DҀ�q�ݑ�t�pv(+-��r�$m˝<��m�=�{cN�(�f�/��@��wH`�W)�KI���+p}E�Q���r�j�R=�ԤfL]fpF��ݏ��0�_���ms �4���������1V�z��k~�qm��`�Y[g��R���r�t�E5`���K�9,D��*���n5֌ޤ�`ٝ�u�Α Y�=85�3]\]�%�e�����V谬�tE_�kKkk=�\UF��%@b�44hQ�["��Q�����ktx�#]��D��J%������ft���)'u5��+�|�WRRb��w��k���`W���I�fcph~-�����������MM���"�����&���
9���Pq�E-� vܻ@�}�zj������l�+� 3͝+��;)ꚺ���U ��*��C�
�|�d����B����~CqH�mi0�U^__:S?�+P�c#����s@� X(F��>�_O���$�}T������}/������@ې���lK+��#�5�e���)���^`	+�P��>�ޛ��
�S��\̲��Lo���T��iq��)�� ����X��6���"7�a��,��b�R��?�Z�:|ʹ�e��;)Ė;�ַ͑bc#h�|&�|}}��|��¯�b�\b�/Ў9��EL��צl(�ͣꗁҚ�a��B�7�aU���@ �$�/t�4��K:��m�pv�1���0f.5+�]����w��?�{�PTLl�qD��d��� ~.��:��,m��&?]�P�+t*���ҫ���-qҥ������r(�fߪ�x���_�~��9�Ƒ�h��>>���0>�����i���]Ɯ��ۡ{�������LR
����t��JGlV��#v��*������X@;(c�;вK�2��MǬ�5�Tr�07d����.zP����"eTY	���r$��(ϥ���={�U���>0
��C�/6�QaO?8�[�#�I7j��{U,-ο�V�_{.�lLfu�L�q��ʺ�]D�a�[q]������z�t�������au���e�t��+��jVaTM�"�N;��* �5�@���m���� ����I�WB1Z����|cj�)f�i7DN^�\f������+������冄\5�n�n=���I� ܞ���CQ��R��|�	�$G�s��0q�4��L#��qqq�++�^����ј�*���VS���F������gttל��D`�۽H\����N���H�==�C�%$$�Ӳ�l���N�.E"��|�{���.Ćª�o�;Xc���7&�6li���Ӕz@髀#�vpo(r�>�174�p�2��)j83�tt�4�T&<bH�\UY��`�x��@s�_�ퟙ����q�l� *��ފ�����MQa��Q���8�q5K �P�,��\�s�1����;>�q�/��m\��4�W ihh�'W��w���Ѷdic���������]���oK}��˺
�p�%���H�����+ `�ެr����**� ��/�QӃ��*#�1��5+ P��^c��Xh�Z��V(��߾� 겖^�g�_GT,���|}z�fhS��"�ଘƱGޛ�����t�ɋ�PYi��i]墼��|�b�x�2�<=+Km�4r��D$S��8űwZ]��-�����(�!^C��Յ��r�c�[x�j�C17�]�1䴗��m�/ի� b*���O�u�lG�5v'�9�y�����d�rs�?��t�>�Ӳ��oSX5?b���4���Ǐ�6�~���tn/�5k�;1RNkc"v��fKϝ��ȶ٪7K�,=}d�����W��`����^tIq�m[��>>^���b�X7��m5�R�!�yx�������f!;Z;��SWA*���w��/���ŃSX���͎�>~77��70	��x����B�\��7Z�&B����=��J��aT� TTwU�"��D:�T�U�"�UJ@QpE�ҥ)R#-HJ�H�  RB� B������=�9����3�<ϧ�̝��9���V����i
z� rO�X�~f~���p����w�;���acN�I�������l���ٻ��<��H��cd�����o�ÌM}�����]M��h�۷����X,/\�|c�������>�uwF�7nN/-���I��>@K�ֺ�G��`^�20X�? ���<q����o��"��{/��P֍�:�D�,>����j[X�>}�I0	{`e��|����ۡ�*$IX�ms����ݾ�h�����(erwsb��q���%�m���ħ[�:���6��Hľ�H�������$ܗ���&�]QV��ؑ��V�P*p��w��k�r0�ި�?�w��Ӹ7ο��k�-��4�R�5��:��؃��	Q�����V�N�T��U{ͬ��/���#0^c^f�O��~Ak��uy���a����7e�ȯ����XH7a.J�pG�#g\ϐ��(�����6�����O9:;�J�Wp�5iNO�(ݛ,P"�<Q�����[�%<:.��Y~~����m111	��b^~���y�zx���t�&������X��<Y�7��mT]z�a.*Woz�!����:��`�G)��2O����w9�o��t�J9[�]$v������T�ؕ
����(���`T�|��� ��,z�dR��Vu[\�����n�~���Bi�Ww۴��cR�����DcӀ d��%�O-T"���iP#=h��X�G(Ƚ�p*�4ePZDMi
�ˌi�a$��|���9������X"�%�H��I}3��(�]4>nc�u�gfF�>}  (��O�@)�W���OTA[�eWKJ���
�l��1H��_�!lRâfm�ߤ�پPߑ�6WW�Qw=ټ{~^_]C�� [3�y��֖d��o�"��ȧ��	9<|(E5#��Ln،c�$ew�K�:�,{&t�"��Ǜ6S%��4Zk�fY&�W��x�ӡR��!s��Z��hm$5�$n��A�l]���r��3)p
��|���c��7��u��G,�P5�y�8�Y.�����
�<�b��
@{��| ���+G��}���h� E�
W!k1;`�|�w ;���b���O����_�Ii�Fӗf ����h�������Z��%���[�.��嵬����gT���q^cMː��.$��.�k�v�NN�˂��y��<�j!���y�SJ﫨�
Wr�HL���/�n��M���C�E-yy��Z�4��9�/��'!I�J���r7���\!��V��ޮڊ�YX`K;��@��AN�S�r_/����?�1i�!�9ﷷ/�~T�C??U�F�W}T��VE��Ң�`��Hr���JuH^�{�7�[ec4=K%ư!y���!8{{{��R�;��O�[�c��@.)Oe���{^��fL�I�a��U�&#Eރv3@�h�!0��ɹ��|j���gf"m~[�(�u��S	�9'�h��\d�7T��-�}MH�P]٥�� HBS��d���߂��Fv��?:
�.��rf�K}_.����ގ��xy{;�;Rf�q]�,.�/LT�v@���&�2oqѩ_�{�DE�-|�4楮�jR��h���P�{[w�����I#���Q�*��J��ȍo�7�DiS|���EA�~ve565U�!�1�]V��f����~��2{�Fä,��{<����>B�g��W���v� ��mַE�- ���E�JYȺ �e7����T�.�Tٿ�76.n��#и�mN�!�W럤l��g�y�\Kk��H��|K��wS��2��<�>%.��U����t��p~���J ��յ����70Kg.��ދ4��"0"4��T*�[ӂ��5���0�P��+�R0~s�g˪���8�8��fU�V�p@�.|jM=Y��)N#E*kb"6S�C(ܳ2;w����s��@Y�Cc{����0���HaLt�k�����ꩧ�,HaA� X��_ė���\�IX#��"31��_J��Y�5L.xK�,n7�(��a�\ʮ����0K�������"Wr�Z�����{fU��l��w����D �r��Sp9�����m��V��!^��9�l����OI���4�5��˦���P�����&���d�����_�Z����<G7/TyR����Y�U�ۜ���We��4��(�a������Ll���"�fUQ�E����Ռ#�f�c���w� 1jd��~?(��I�HR��݈��Z��]|P;�kə�.@�I�:��WĀ8ڻ�/��37�N�2#�ڿ����b��$�nD.w,��6�J��;���#s������gf^����{a�
��G]�>�F��X��������}-G2�ʓ叛
~e�� ��#������e!ڴ��I�IL�QBOV뙘�|e/���	�/�jjX�;�qyV���ׯ��)���׼�~���wrh����B3��I�^BCG���19���LP�7'Bڎ��Z0T7W����>C�Z�쵢�N�L�7YG��:��\*9�^ZT�Owe_�4�3`�u������J�d2�Ex�J�T;dw��i.|`�@�����޿ln���d�.uW���t�?R�,,6Nݖ�!�$0��	��d��4f�
���{��-t�*P3V��>��/T��ۛ8�\�pe-��w�F]]�K��K�.9>|hz��u %#�U*���цz�K�
�z��c�ӄ������u,�N1�2����>H3�oG��8��e
MM0h�]�2��������(>�� CL���Ư9n�ŢS�UO��N^ɪ����^����s@��}H�ԗ��KE��{�B�Z詳bs�2���%ҋ�b��3�����\���}��B<��_׍��Ō�g~j��@���&w�hС���(�8�w��w��5L����6ȳtIj�� >>>�����P���paaa^z�v�'�� �)G[?��u"�<��T�H�e`��8�Pݮ?�H��6g��NǢ4c�����2�*Ȟ�۫o���"R�.J�~�%xwh�hHp=H�4N���ʳ����+��W�0v����{��*pL��ϗC�U�2=m�7�嬾��!�K<D�2�韮�
�{�x�H"P�ԥx����(����5�ӡ�ɀ(�@��XX���b��?#6/EC�'����L�&���E02m�����QZ��A&�s��Z�72Ҷ��2%�Kv�tt���SL{=�d%�o��Y��1�{�Ҕ�r�1W�b�k`Z��j� @%-}�H|�ߥx|�u ����������]����������L�A��W��RY�������/�G����,,�.�4�l�6��:��;�7�2���^�]
Hg�?`��m��I��z���bm!n[Ǉ6�"1v��_���#o_�Jn���/��I���՘)�BⰞ+ҩ�>y]���[�
��7>ߘ�n�e7�;b �ꔟ���a��h��I�I���F0ɳI�3�Tt��퟽ v�ֱ@�s����%�����>��v�j��N\�A�$�� G��](?e}��wg�%jcw�3�	'u{���N���@���+��6Y��^��X��ep/��X�Ԫ�E�x�O��V�M��SP14�50ԩ�<">����<{���dE]���}9����-�����`�8ϦDP�I7'���g�0��t#7~́�r��_���P�M	�V 	�ChRQ�7����?�*�I��S�d��쒰
o�U�oF� ջ<Q����uK��(�'�	��4��2Z�ڗV�)�v�Qԅ�������iC���[�f����e`e�-�c���;m�{�[���*	���������)U8DZʰ*�sH�D_9�g�跽~�k~�/�o{���4�/����y��-AYB;qnſ:!њ��q�&�]�c.�h�$�̼�rX�&#mCp�=x��?V5Gmz{/��}~~�Q��������8��X�� 5hc5�������
>7K"&y�6�����n�U��n����Rxe�1�����Ǒc��"���������|�q�x������b��(+ ͫ�a��566u�8���w%Y���7W���q��3�$��>��X{	pߕ����or���,��éd�.�����=0y���&���76�f��-&W'__#]ݨ���R=5TR��d�l���I�����jX1r~�(3%���b��9�,� ���"��Y����n�Z�_�}�N��f��tH��MOgꪶLʮ���*g�a�e�=���}�$P��B@	w�����#�� 	M���<+��/b��CջE�$%F@����CV|{p���ԭ?W� �kt��Z!�`��;x/˿&�R�x�k9������7<g~6:S�O�5h>�vFD�������y/cY�N��0γw[D���_q�:�kCZ���TwS�*�R�d��o[�ޱ(c�j=
��j�2�^<*�hJ�u����1��mm��5�p��H@��6�4[�����a����5���"��G!�Ɲ���6��2�*�
��?��*������o}���iM��%?�x��6�^�V����)�H+�{q�.�v�:�C�����~	�����^���x�UV5+���}:\�:T�9IF�����l�d��|~D��:4�r�ad;�腽`�q��~�(����P])��Ex�=�V��(v�5�~��	�,��f�*_�l�u�L�P�O��@O�� �D�E�t��	�$h?��x�Ω쾤QE�	�������R a\'S&)!g���R.ƒ��ln� b[��i��'��C.���i1�������&��k�W7NPF�
���z�
�TV�Ju9e�w�T��L�#g���ي� �Og��ȭ+�`�'ɏ̀����1�<S�|(~}C�d�~�~bN(��oM_?|�]h���dޱ����tV��x��(�=�_��0(���Ac�j�dJ�7d��]hi�!D��Oٝ'��u~����/g��ů0:�v�*�����"��
E6��;B���v���?*��QwX��)���b+^k����5�w�>�&ppk��_�J�d�*9W�%kP�w�9�?)�A�����b4r&�`�r�����h�!�t.�~[ZUQ
z�N9nv�g�����Y�$"��w�,S����s�$���@��w,��׫��)�2,I+~���(K�*��'���5%N�r	����AN,���.��_9#�j�;�v�bh�xJq�ᆠ����L �z =�c��E�T"H�k@(Xrl��}���O��Y��Ā�4{ '".
t.Mu�#�ʋnkk�1A�ÍJ�s���YC"Q(�ԝA�ӡ<���X���d2f���	Q9�#P�����D��qȳ%GM�����Kx�Q����7WO5�C���$J��mx8+�����w��!y�o�T�n0��6<-r�Z���~y7�� T8$+K�6�+����93�N��T��Z+�:b��F��mϛί�x��5����|����ו��?ip�wg?wx��c+y��ƽ�W��z�t�]��O���
3��Yf����_n��*�b[)�����"�E�U�;�"�D��5�������ɴ}3�0�7�s�����k��]�	�X��Ώq;��7(|J�6F�"��y��dd;��#k�'p�n��M��w��+Y���)ځ���;�4j����#�].���/݄�$U	U��3�,z�vic8�E��_��*��A��&e�Y7) C�x����}�z���sٞ�����bblj�~��"�[��g���o�-��YYY�R�(��`�	��/_�(݉���5
o�cƜ
�v1V{8e����3�y��������ó�����
��%����O��-/��-��$bN��t�� 
�t��s��D]B�Ѝs2h	����U�>yBN��� ��Bq��)�t����"��qBC�hu�iu�Nn�'|�S��F��=>������l���
Z��HJJ�(Q���~��+��[�q���3���V`8ۄY�\�S���&���A��}�h%Z��l���'�>}�7�$�2�n��1�h+2��%N�4*]=?�������:���w�(U#gy0����sH/Ѳ�omC����	�.m�3n�պ{*.(��n"���=��Z�~@�1�peQ㳍��F�U��t��9�,9��SA
t�8ŗ��##i�I���aFg�F��L{�������Uj1�"��ǳK�=4]fs~�֯!v��P�F��6��;W(���v�Ͻ�jЄ�0��s���,%p¨7���>ʱ<ϰȬwaA�O_:��|��F������5�vJ��5e����]5�Ϗ���5���J������v�����m�N	�0����G��GiiU��iߔ�?�/S���Z����ro{�r���me(:����;�Z9���Ռ����蝜��;;�pG�GF�$f�҂v��<h���!������E��[������(«a/ �CB%��f� ����ac���Τ@�C���(Ƨ����� M�W-���_��^P�L��X�����Ӯ4�حO��9BEo���d���������?�X����A�BCò�ڡ�Kk�����}��l0�QD;E������x�L����־}���3/3�i5����m������!�
��+��SN��5.�gy�y��q���X���-�(����G:M�[�h�/�3h�#[�:
t"��Z5?��x2�Y���ꤢ�{���Kp�yu,nWd�B�8-��C�٪x�;�M��#	�.b���5r�%z����;�lyiiԟ$`jyǷ!F�9i��&yr@�t��g�R�N���Omй�b/�Ϡ�R��"�.,z-N���U�O8	�V �a�©^�
�>�ڍ��>(�V��%;�75@5g������!0�U~�61���8��u?�lw��.ޔ��`��h��di�
�63��1X/.6��{�� u���w/}�7�<���k�����S����*iG#���A��T�=y��јV�ڍ�>b_$f�@ّ�����h����C}>��^Y"Yf�wx�B��t���\�<@NwS7<jW���S�7�J�	b�%�k��p�IpÉvНsR:��3M͎)�]J�M?�h��\k��e6G�?C����a]$�k�US����M��4�ڗ�l�M5�h���V��N�T�]kx]�Q���4��*c
�g��|<c �k�����W�J�/���/o�T�u�(��Ү,���kV�St����k��f���Z��R���#ʳ��(v�?5�\�c�X|F��z���������݇��>�on�*<�"�Ku�[����I��7t��=�[lfgf�p����p&�Z�mOƲ��T��6��1�h,8�^>��	�Ң0�i��}MG�I������̨z�$A�`�U�(P}���y�q� uH����  c�IA��M��7w�ړ�1/�v�C'g;���F�7H8 Τ�I��Ih�����VaC���-u�l_��ٝٗ�W����
�|�ƮP�j����1Lx�Һ(|Л;�I�%��k����;���}�k�j��T�ڍ8��br ��4r4}SVm����XY�3���9�P���u��^���c�tU�Ӈ�]��b9�}��V���6��ڰ��07Zҿ��T��_#�p�����>4^.n����u�w�A�"\Uov�.��h���0��>������6���@3���F��b>�(���9����-�k1�Ԫ�R�fT�eI~.�C{}����3�+5C{7g�����@����o5���0c���KM�[	ƨn�M��!�~��5Ԕ�Mh�:�<��{�M�ܐ]��k\�¯�t���ѪhoN�"z?�w�N�����T&�/^�#j�WK��j� �a��-��nf����;Q�g�9z
��n�Ãs�K݋����l2Ko.���A��z�U�)ܿ���f���*�s�Cae��L��q�^�O		���y����:��D�����|~��L+��f���@A�y�����hj�N1ڗ�X;OiX��1!g�؏T-,\�i�|�2x�S��i�6����]�:a������?5���כ�� ��!��Z~(��U���,�X�`�@�.;�w�PrR��8�k�u����o�}�
�d�P�N��X�-���f^��%�7�r���Z�¹�����C'�$C%�n��+T�Y�n� :� a3��WU�H�A4��K@Ԩ֜x�Xd�B�d��C�⟩�������m���ac,9�����m¸���-*h��^A&Ī-��fͣ����J
�,
�5��{�Q�cZ����Z�:�Oz��q����}�
�������|�WF��;TGք��m�q���FI�KS�!G[l�R����ׅ,�tn�s�ʊ�Ļ��6���)mMM���ߍ��K�ؙ�4��眓=��V��md$�ǩt�QK��?�E��2]|)�������5)��q�t�p�C­��ԡ�
��s7Z�+lH.}۩�m䏿������30(4���r���:�. %G�ם��%]�{d ���h��^�`R�TKS�5�#�9p�7�T�ϸ�IJ��!�������?'aD�h^���}*���Q(��N�*W�O�Ҷў፻�Ka�����+4��
 �ne�CG��#����� C<\5�ۏY}D
$�Xsϰ���;���T'ϑ`9,�O�TܕP��8լ:���%�E��eg��}�ϪR��Se�7�;��UIb�kk7��&��ԉ�<��U�b��z;x���N�R�3���=���L4<��K�8ǟ� MA����c��|į���ҋ3%�@ �C"��(�
F��?��6_^Y��b]i�����ƫz���^���
��>�Ԋ#TT���W���\=բD�k1�����o���g'����s�H���N)F�Ȓ���:F
(�Ui�\��]%V59���
 
I��k�+hgG,�h��M���-j�Ū^�ؠ]$|�4��{�C�tzow7H��-������	`R�:Hױ�5Uy�	��	?���B�Z�o�5��K$�_oȱ12���eQ*F���L��`�~n������й��m%c��2�nC�1s9����:@T�����s?o�bB�������{�Z��=D��@�-sFÆ���J�Hm����]�Y>D7��Q�t��d�#]��My�E)��m{�݃���s��I�V�/��Z�0�E۪l�4��?�"zv�4Ԯ�L�ܺ)�a�p �<���F�w�Sn�n����e l�wN�vPP���J��źK���&T�8�gh��C��iW�NL=���h^On��O���-��~�Q���o���j#�DX.+g���o��ɗ0���2|i{���N �!����|h:/~=�C'�`U/�U�]7�7.d��Q_`�Vگ��E��/��|�n|m�9�	�n5�FR�Q���Jm ������-+�q�Xk�J�m�#� ~j����HdHش��b"@�
'��YT=9p�\2U������yhv
��і�YXԕ��_ �z�]}ȧ�W�f8B��f�?�� ��� Mjkk������Y��}y���7�î`* bX�h�Q�$u�n���Cu�!���V�!I|(���V���{����J�$�s�x���8z@|m]]�ΰ(�fC�%t�z��z��/�޼�]�� �\�\�,]�6\��Qw�gp�?j�d��9Eg�>��YMؗ7�.��%ݱX�\��XT�%��(�/`��(wfkk�40G�9B��?�C��2�X~�\���*Ԓ/��}�]��v�a��U.�mmvG�0c�ڙ�Â-��V�<H���6aw��G�ڝǗ��.�w*�%6[{�m��"?��Gfe)��.�R8�$gx?G���|;?%e8��PT�Y[/f$%��8��޿G��Kw�F3��|������E�����PM���O�t�2H�˯]s��#1���J��P}/`PWk$(�v�G浵������j�Hf�# <�fgmo� #=���M�����\u�查���3,TF������zJ'�fV�4	d��Ɔ��?G(t*�7�n�vt*��	D��/��+<�_�{qNyr����b�1��*�Q_�[�@ɝb�c�������P#D�^�d�404O� ĴI��*~�r,��t�*v��#!G'����
�=L��mI+��g-��K�c�� ��H8Vh������Pҕ�RC�LP��fP1�%?Z�kn�~���ՅS͊� #�X�ud�(k�����[�98�,ȅ]�% u¾���� e����v��: �&��JpK$����|W<3�h%ῒ�Lp��48X`�;����	�(���a��Ԥ���hլSmN����.�h�j�Tr!06F u���<��<	͋R�_��LL�:�g@Ӣ.�Hzx�^�v)7fأc����� 7�<����|�`|i� ��̴�Ք�@��������&���;����x\�i-T,��yؙd��=p�(�^2Y��u�U7___��U^��Uk�)pZ�#�fY�ޝ|����NF}tK�a�ן�i���-���d�P U���q��������kE��

��N�pg��o�7|��N��ƕ�L�bE����D"�ɓ=w����𹅅�x��e�6F��-�>\)b|�#�#k�Q�<GhT����t�Fj�b�'�-����w��Z�?P��Bh������;��&z���+�w�Z观**^��#;��/�ɱsm�7ط�hyi�ʛ����18����
d��1�Ċ]�����)�ij�AG�>n�h��!^����s!�i�U��������M&���G6 t����g+޲q�e �R��3�kg*N3�-����9�k��������_CB7 '&^ �6����@-��T9Bٔ�lV�{<��\*����HW�]����`�t���l_��iP�ڰ=��"%U`ꢌCV,o
��՚\/u�} ���I�`"*�$T�vl�B�D����Y��#�k�}���~2����6��1��w��֏�uww������#}��q�=�ov�����m�-Kcg}����J+9e�����r�L�bT���L�����;{��uw�����n����UV~�z�Ư�=�[l��8���X�x��M�M��=��mq���ӿjg� ��@L{�/(��#B����ʽ:E�z܅hc�ĝ>@e&&���~4ٵ��	�lw��F�־B�	���tgE:����p�h۬޵e�rc3e���v�`�j�����2�<:���>���9��d���#!��Jl��&�����t�������`�3������o9��iQ�	j9��1�'�1�����"z�y�4���_Q�����{ĳ�~#�jo}Kh:�3���2677�l�� P�֐H�����qS���?���ݟ�����&��QW�~B�;�{��P7-�mycr!��71OJ�0[�u��N+����֤����`}>��O�V+K ��ȱ:>^I	�jR��t�n��r�s>�ʍoL�e�zI�^�#�䤧���3�_Ct�?}d?�@�,~N��Yh.5�1�����o�� ��wyܻ[tyI���v�0�!��-*��e�(�}���|��б��k(6�B��p�!�5���s\�gz<��h\�lܰ�j}ܗ�t<��5�#?��XcSA�a.v�:ᐲ�������:�&�ݝ+܆���������כ'h�r�B��1����hAD�	�͢��)g"¾�@:;�{x�w�̚��4o������`o���lj�[����8���Y�]y���%)h6�m6�a&��z�f7n����Y��ڞ#�%^3F�5�.��뚘�M�VJ��|�N����x�<'g�e�
�ڸ0������heuϒ�z��3c@+A����lB1��b�e�Z]s�rNs�c�������:m1cI���+��;!I}񥓢�oc�?އV_�g���1�sQfg{�����k��J1��x�X�����cSZ|�İϕ�[ǭ
��́��c��+� �[��Eu�,~������T�<��C�H��@��I�vk%���G聃���'+&�f���oj
���]�4@a����i��Ax���˖j�j������LLLjV�A�����S<���|Vw��l�b�luzp���ѣ��g)�;��K&��S�n;f�)����Ɣ��WIM�2��c�N�K!eP'$@�6v��`獵���P������#t��C��n9��>8%/�Đ��P��e}(��y��cX��뾱��}�,��Mw�ւ�U�jkE������C5��V��ho@? ��ɩfc{r�bF�c������?�RA%zhӔw��Z�M2Pu�p\`)ewWd����S�X���P-��]w g� �zM��ɃL��UT��ͤ�ٚxchtP~�66F��&3ǘ�Vm'��X��la >���8s_���q��ͅ�����Z@.Z�(ѱ�����o��ola�[k��|JLT4�~h��-�ҫ�=T�B,�9�g"ى�e�&��2f;�L`Mdl�����L+�����ݟ��+*�RN�^ˀ��d�������ag���@��@ޑ���P�
�v������$�#��tFWo�wWP�@gy��*�vTy�C��.�c4<3���ʹ�vsҁ�^�xʉT1Ћ|�ľ�؟��#"�����[D�i������=�z�����g;���H�ӷ�|�b�����+��h���1�X�ʼ�Dq�]���Ȥ?μߧ��k�	�C��&����o�Vy󹊖���!%v�����[*�U�*�P;�a S��h�Ym���w2#�����<>����w�	����$m��?�i{���E�����t$8��%y��Ob��\ll�O	N�j�.[�ݲU1%���/h�s��'r�T'�����D�]��<�>k�'?�~���꺕���Onu�&*f��$���a�?�ح[ �%�� )/))X^����Y%J}�mT���:����g��/�`p�1����)�W!*���u��CY*�c��rZ??&���8B#GLj����83t�TKKIؗ�ݫ Y-l�PIJ���!�n�UYD��8������Ą����i�}��y���0�諮�v-�Y�c����{Z�Z� T�DG1�6��O��?$�^Ze�O��k�[
�$�+$1M!v
� .A���DW�C%P 	�pHV6hqߴҴ�B�u��Y��l�8zG'73&Ʀ���ZF?E�¨UlD�rMX�r��I>��n���.��㛾c_8��=幒��fy#���])�I���T�0$������5˞�ȍ.���Š:��>p�b	D@O���H7�>�t�N0��L߳����^���u�� �cwT��G�����e��m��e}%�ɲA����09�,��o(�di��C<�ַ�s�v��=�?=\n�~�z+�~����0�G������\��\" �'m��r��@l��^
z�7�3�}�< �=d���`�,&�Ͽ�ȁ�A�qB�g>i��?�9X�{����sGGO@�k�]:։����C���CK���c&b:^7��x��B�҃�>��*�j>�%��,��ω�zh=|��`|�CB�?ڢ��w[K<W}���+.�����͌3��������ҟ�7�-�'�I��>"�=Բ{<���Pg+�1�ogGDh�S\�)9,ջ�ig{�F�
�H�h�]v�U�FA���^�<�Ψ��A�wY�����Do�@�Q������=eD����T���\�n�bB�8�����3����#q_�"@VfeA7O�}�TW���5�_l7�aqj������錇���Bem���jKLk�{6&%-`�xxx�-)Ȟ5�Af��_տ�=Z�&�{t�k|�g�=�����R�^��MF�bu��vЀ�1���ɴ�D��q���Q��Ҏ��=K����67=�Zhs �.���s'}���KG�![u�>Q��]��-���G���$H�+)x�(���f�(��)���Rn�w�)�1$���k�I�մ+\��:�>}J=�u���;n����f�� �k ��x�e� }��h�N��A"�y � ���1lw��Yj��u8���hC ��O	�i�ӵQ��&'��o7��nL�% ��rs����n#ɪYPPD��A}��� �N�:�b헀s�4���3Jw(!A�սE�\��?`��x������nx��72};���w�I���c������x5�S��޾�F���E����t���
3`zQ�����o-I(��8`lf���P�2���	��q������i����C�Y8.���Wo����s��_�2�Z���3`�<��������n�ޅz-���}]]��� �{�i���F[�@?�R��7'4Z�)���?G���g��=�ˁ'v� IA'�?a�JV"�.��c��p;������H���L�c�ss���x�Ԉ�x(������!9Lp�;�ZRR���Ϝ����s�I��f�5���{���ai�xp�i�����WJ1!��������������%�<#���AA�v�m��"�.{ػ�j�=��BE�:F�]H�����?���0�P���[d���N~���M�[������U���A?�1�$?���^�X�&A:��(Vk��0E74��'ï��.*#�����;�U�n� �j��"I��9ձ����k0ļ�&�И������)�˿tsl8�����TyR2��q1��S��y3��9�������dp��=x�\������}���#07	xE�6#����$�r�S:{��j�����;�K���P�9�1c��Ǚw.a��ۿ%u�t�(U�>���Aii���+� �UBJJ�����߱Q4:H���?��@�����IHJ�����3}���&Tp����Pu�9���7-e��h��1�}Dp/��N��"%&Vh�*y�[����ڻמcM^bLi�,��_���α��{Ȱ�#��$ov��IIe���d{;fbr�������'ؒ�xQ7�;�
{m�#���4�՛�����6���Bܵ�H�r0��/���!��vIW^�v�� g@d���e�P���" �A�r����\a�f݁2��3�	�I_@�/�߽���(��wm�����F�	@�D�:B,׀�=x���s%�у��Y��탶�l-��mHf|������j�d/x}fH��:���4�������~^��&˽BB..�~���aB\di<�L
lZݢ�-g�lы�7z��I~�g[��o�y������-�
��@��w�X0��V�^5�%�	��j0�� ��2��{���������������HD�t�޸�,��������ő��ِ��f�9fL"s&��Z[������/C��<���~l�Q�-��,�=(r�_ �媭oI��_w�t��)\D�#''g򂤤d�nw�K�1QI	��!=ՠ��{{>��c�x<�[��[�
�KU�C����/��)�;K�1�
���A\��3�+��� 6+ PMW�{zvVz)��Q���E�:�!�O�� Yq��Q7Ru�	O�&%�h6'I�[^��bKٹjSzpe����IJ�٠��鐤�r���hxxc-�/(�y�lw��B�ԩ|8�A��4�����9{DD���x
ԟ��Q_C�1C���f��15��<���ql�Qٵ'��������������0?>:��۷�P�����[����#� _�:=K'����+��6F}�+a� ��ˍ�: 髞#I4�����]!l(�:p����-�ye;L�_�¦$��f*H9��|���Sa'���δZ�_�)���de�����2eM7��x�U����5�۞��?Ѡ�.V��RKl[�ْVv���,kf��8$����y��_Y��Qʱ"�7�/N�P	�����.��1x�g���i�F=�Z�� mѯ�nzZ�fym���=z8�|&���q9"�k@q��}2����e'����=k�1��ץ͔�o]j��M4燹�1q���������:F���,Zl�wh�����R-�n���F����~v�ш	�X,X���5�z�/B{�Ą��ޣ"����\��K���� �Ꚛ��$�`�([9�]C����RGd� `�}���A�}������a�`D��F��TG�V��4�~�����Q�d	/U4z�� ����vq�u�n_�O�X�a��0&�fA����
`%�
� �A��[;Q.AC*�Kr�ah�q7�"E��=�[K"�����o��ꈲ��z�9�f�O���Z�h�"���'��;xmct�������Fi��޼��T�\22��\�k���n�����D�2Xē��e���i���:�[��-����H��"�چ�Ln�bm>���Q��y>��@�10ЀJݯ����#p��GD�P�L��O_��u�Ի�p�v��F�T
�Yx�M.�/f%k��|����\?�/���pK	�p �-�V&��j7nY\=���\"�Zs
���٪���
����B�eJC�;��0�=:�L20(;�|T���u��l�\W������a�<t�.axd.Ĵӥ�^6�������Y����ڸM�3"� �P��f�Bp�*���\����S���:���	ך�{tp=qp0	�(tƫ�Z�ʼ2<ʺ>��d l� ���%�_QQ�U9/&��vy�Ѭĸ7��{<�T)_��ۗ��S�5e��t\��s�ӌ���oY��d�����?x�Ů�y��S���%�r�Ue��>��p��`�0%O�ɍN	ڎ}ӆ�|ߤč~k�)q���?�R�9C�]�z1����'�׫z�q�l!4������l_"=��3Ր]A]��d1�n|�YVkMsn����I`��:%�mX<��$�J�t�]W��4�U�EwllL�k:�T܋H�6��9V�&۝���)����R���Fkzxx��a ����$�#q��9���@N�1c;�Ph�	�b'�Z�m�w��j�|����d)_�ܞї������pO��8� EM�$��j֚w�4���T
{����W]���~ඪ�o��\�鮚�7�:|��P|i۟v"�KP����mn�WV�7�5䏋�=='�ڵ��L#	�O����f��'��I`�t�*z�N���xn`D��P�7Ѕ#�4����H W�����K�ʪ� {"�{��
�v6}��#�|�e���ۧ㳯v��M[݋�if�ǵ6���p�����8Wk3��<D�#�޶N�k����ШZ�Y�|��3
ڙ�#�,K_m�C�����j�ҁ��̼t���{8�lvV��6�E�K��N������o/��'|��*n�\���>JY兕���dV�H�ka�;R�Ŵr�Zzc;J�J�pb��k5����`�����0��`��)�@_^����EHp"�$�x�Ʀ��v��msɌPL��/���S�8�`-���:���=d��gR
"�;��9�w�������wqP��C L�6���]<���v��I�h<m�JXƾ:?wwU���(�yOqq����2��(L�š@OV��R����n\⻎�]~��OT�q�!U�{�bT�V�(�۩\��;�Ǚ�Ha�l+��)��պ�I9<��2��O�ƞ����UJE�#$e����\���cz��m���,6���~���]t�/Pbh�[���g_ZG̙���uȌϯVYme���*��������g���^��"�B�Ԗ�x\z)�o������c�w�9{۹����ʅ.%Ͷ���ZK�*�o�W5�����M�ޛ���i��Kwy�څ���7�MB���P�%�������6Ck�����a>P¼���_���s
�]hPk�#�=�I�a�d�}�`{I��;�?����o�����h�_���Cx��<Sh��{��<�|����ⳳ���
���t
[ZW���4_��Rv��mv�)�O�e60�2%4:3AUk-�E��e���:��@��كG��[K�	��.^,L��f�n��H>?�L�Uou���O+ZJJIH���R�]��l�g�[�D!�}�"KCI�ck01J�%�c	��6���}�.W\%s��>�����rP��\�]�F1�f1��1���{�*��Q�ϛ���o6@pfB��n��:֬t���9�NGEG�WkYL���kk뤥�
��
�)?�$]���9r�Jd>��FR��-=P\3���e�~zSh�+�h��d��).!Q�������:�yI�{Y�7��`�� ��,�� +|�����u&�!"\�����5�-���_{����q�:����b8�Q[���hx���;�(���F�H�1Xz��9��s�"�����Һ�.�
Hv�������y�����`��#�D�V0h�Z ,�>��5��(K����76A��@���i���b�X�aVȢ%�N����Iw1���t�`��ݫ�,;��̻�[e�IT�� d�F����b��qɍ�K�"���]ŕUU��-KMK<���1Yw�y��y���7+���^�!�t�u�
[#7+�����G[�Ui<�6G������^�5jVἡ� K�T����1-�Õy��0$���/�l�毰C���� �b��������V��W1|mg��^���L��:^��h�/�w���,�|ͯh�N'�Q�ւN�P���=:���q��Z:Y��o���x�g�,|9���]`�������-��
y�=��ME�u�H�m��|mb��������B�K~b+26I<K��4{�ۻO1�uX�J��Ǎz�+y ���$������А@�

�u�v�. ����Vy���.�Vw�?�:+v�������ՒS��8à�\48XW�u��ߟ��$t�z�}�~ e�߿��`�𻤜xc���^��V�k�_��?ج]:ӎ1_��w/��ݲ�^��w��
>?쫝��m�c����/������=d dT2�pG�C2��s7���˗/�I�G"|b�&��G
tX��v����3Ul=�����뽏��Y���G��**��hu˭v�����|�M=R�+ ����g���/ķ�³��HW	@��E����S=�<W=9h�������p����������I�h��1�e�m���F�U*���~:�� |N��^k��0��g���]�
�w��Ƙ��=��r��Aj+s���$�	�_���y?4��6�(��%��C���4��ۚ#�ൔ�7gR�s�V����c�/�2m���󹕿o�����%�����0��36�hE�-�[��`-2,.�oWc��x#�=?r�w�Yk���΍���q��9�.7{�5����h��B��]k�Aa�����*�ߚ�u���*��|�����R6���xB��$��g�B:l�[���%���B	�S	F�z�^6��b_�G6�ȯO[���)�3R�<�����2g �hDF��?T�=v��۹x����ju�T2x4���We�{狅N�Y���q�ji!vb5+N�%�Ea	�X���ג��
;���jp������.��CϢw����^h�k�)0(�	�����x��%K���>T�s<X{��&�sސI'�d��8�/��K�z��Y=��w�}r �$zJcg�I����i��q�y!���:����5��p&��~U�ǫ�˼PMk,��x� @8�z��iJ:�J�w^9z
���Y#�����"�\��y�����h3��Μ�R����|������ʷn�je��
 ���Z�L�d6��Ae�AL4�]rnkٵ@8��`@4ud;�%pU<��Z�p�X8s���Qd�!d>�]���T�P��
r�䨟[z+����~�7k���'ૼi!1��>ۯW7��.e��d���g���y
	���Y;x;��%\Y��&� ghx���v��X��Ǫ���qY��dt!���_�<�,p!W�)  �7v~o�z����c�*��b��= Y��4�ހ*�V�A�tP��3����T/$���(꛴�膺{)a̍���[��F|SC?�'@1<��ϱp-���J�a�'V�\��Yo���y|�Y�����J���i���'�̑� �rtu���I���2���o;Mn�eGG���X�{q��牕=��J-9�e����՟������b/�L�+M���Y 0�����v��7�h��?1�W�B� �ƒ94�}|���ﰘ�!s�3Fv�#�p�E��p�� Iv巏�=\W��3K!$�p
��+{�ĉ����9+��1#2��$[)~��W�졮�Wl�E1��37S�{��l|ۖn!Z���7k�s�S�A���>��{n���ɦ�����f���L��W�ڤ�\\\&��Ft������WQ��J�fZ�9�V0V��)�]��Z3��;}?�tZ~f=jr��f:�-�+�YT\����/�g�U+YWhVS������`;����|�s�}��lVx821�f�#�",��.�/�0^,��ƣ^����;1thb'�%Z+���z�0�;��\U�p�Ω�1�F�?K�{fsss,z*"��W�y���1X��l���g\--���F��xUF�F�cU�����!�?�hQ��R��|�t�!o��諀?�ƾ��bbb�l�0�� �2��ʗ����Ɵ��������(�fWś�#�ֳ�g�;5<%�}��P׈��I�d9����7��=�bo�>Q>�����V��ipAn0�IB���+�K�-�s�vv�]m(Y$�sK�����ҹ��/�S6�ee!�:�������7N�9N��R�����NRk'��S��Y���s>�~��N�WWRr���4nsjȊ� XՏL�țl�B�s�{j�o윥����d`}����G%�x�I��Dֶ�||�����u{"ӿ���,v3ڰ���}��5$��i���������)0�C1��h�^W=�S��s�O�c��>�H���gKi�?���4Zo��kk���e�j���1���lp.�����<�)��6�o��9L�+�B�	^�S���b{�e&����Q8��Y�ɩ��]���|�1^^r����ĉIj,[n������tڜ	��<8i��-&�m���YWW#�:�ܣ��*ccc'O�Y�m�`�I��&���Q�.Kos*�jG �D�Uz�z�����!�{d}v���Xl�7n[n�b��yT��Bl��j�͢򒷗�������]�3hZ�$��o��&�C��R>�=��FaBI���H����J�)�ɘ��>�1���APr�V2���?�k{!d�{��U�ܩ %�C�÷��0��QM'B����uM��1�Y�c㤵*@��ݕN���龆�r� 0^W�?�
[ܤ[��n��RFx�c9�>��r[�
�΋6tQq���9����߾��r�ȗy���	���o���UT�N�����'t+��!�@��f�n��j�2���iii���[0e��d�|�,G� �d�8$2rǛ��~�xc;B�y�!.+�]0N�D�_Ѵ�wRCN�v;aXPW�j�4�]�u�^�}M�/?�Y��<},� �������	�X������|xP|W*炏�:��]ڰ^!ZmX����q�b���Ą�F7ʌ%������
纉�t�C�V:mSĞc�Q��Dے�ox
r����~��/{�Y
`7_�|FBJ�w��=r�]ss��A3�����n��浢�h���wJ%ee��G�N7� ��t�����Ip���wt�]���C�b�r�0h����Β�� D"q�D��Q�t@*:��ܝ��)�~����"�`Y�|΄
��֚Nn�F\޿����T�R�a3R%*�u�oy���->��1~�\���!�P�L�V��k6�'oʰA�OO����N��t
��:�nIR�<0X����kǞ$���dوf�O+�Q���(����Q�\]��DS@m�\]���K�^���%�1ƈ��jv.]	$��D��ՄL�a�R]��ع9�T[��ϒ�)�d'2�{R\q���}Лڒ�f�B�X�����_�=����&:���6iE��@�K �[!`���0J�̱��is���u�q��N�V�$u�uvuu��W���}r:��۹2	�F���.1,F���M���B��@�2� �w&�Z��8�i��������?b�Ɉ�rD�� ��ԝ�v��2�2T��������U��z�L^Ǖ��޸$��舶�>YAV=ooC�����8[c�Z��C#�������+eD�=�5����!5@�N�[�5��V����qa����e��OG'�8{�$ H80`nʞ�YdwGn�w��XB��%)ʼ��%��z�-��Fn,��Lw����"�	[A�~�h�`���O�숱�*.���ؠ���=]
����sso�u�T��!�JK������F��z�P`P�W� ��)�/r�Gi��##C�R�.aH�0�����Z���%�C�
 O�F��@���3��c�>ux��� ��p����³��p]�g���Gk3B?ѵ!�I�^ �x����3T����f%R�L	�D�Ϸ�K_�>x���� �¥$5��աX��F�j�!װ�&u]]B���<3��ܜ���)|,m���$\4ʃsJ7-1���_�82�BE�DP6���"�(�47��B]0U�q�O\��B��n.P��7�.΁�4�n��͝��K&�X��r�.�b;��&5:�FB;���94��V���eP���4?Aۊ� pI֝���pq�����������2
�����ա��dj�ND��']ܶh��y�$�ͩ#Ҏf�܄N.�G,��y�ݛ�t#��E$��Wy��嗣�=�"�(�#}����7��&%����m���b���#W9��ss�E[�{C��8��:�	=a�w�a���,���x�ދC�G"[�k��a�Ļ];t��L՞��,��tG�Q�QMw���4Ҕ:�P�fgV�5`������ǆ�ZhW�R����B����9_������vuyA��ó@>�VihT���! �u򤽝�)`�?c7*��^���#��������Y�=�,�:<��Q���r�;�����#0��	br�*�fo��˲Ȱx�5-�A��3C�}���Xc��4��j$&!?����wᠭ+�Z�:$v�ā_��220�J��F��~ȓ�V�����k ,ȗ���,B�~;4<[������ �2:��bзA��9P5�ݘb���@"��{�QTC/'ǚ�ĉ�\�M`�pE�����;���T����GNO��ӂ�WMɫ=�Wq��!�U6���}��˔�m5�V�Vx�����?�
W�ʕ���f�1%�b��sôw���j~�����;�N-��Z�ۻ�F�_�^���|U]]>�� �7�'+�1����غ���D~qII'�bT�^���{ܧ0d3C�	Z�%V���{/�o�ٳ>D�H�r�T���,elV"��>��$a����Z(\OOOKK' ��~�r)��Β�fBN��*��R��XQ��h��Ro��+�+��\:tamm!`���i�^�w�} Q�\�և�}΀��A�^��i�.��g���b�v�R�by��Y4�%�lE0�X����G�d�;����m��%?����W̑R�)�*��"�oox�������䪪���Y�U1�=�T3�X��ý��o;�A�s 갇2�2��I̍��A�
De�>,�"f��U�B�f��S���j��0�6��B�R[�1�-.t,|�?eDW:�b����U��έ�Z�z��N2��^�����{@)��}D�e͚%��W�%x� ���Xu��U)���GJ�` t�h+�K�"�zNa�W�y�@�����7Q�̯F/ '�h�,K�w�6��ro�֚m��j9�eŭW�9ݽ�ָ��Z�����T)�f�b:Pd��;���� ��P��ңV�:�'��>�y_
��H;������y���AC"��9�K��b�s}w�$�E�v���� �@�&&%�n�Ei��Z�vގ��*8�����M�������U�[��r=��<]�U��̥�얒���W�6�:���_��텂h3+���k`���rt�QLZ	�<֢�
�[{1'=��֘��?��R'&B%$�ɜ���n�O!��f���`;!�%׳zBlP!^� .�?���O���bh�s0��l�Qa<ɓ�)X{�ռ6�B�97��}�h�伛*�b���f��=j߼z%��-�Y���r}}]LD�[�=�����5gMYv����,} Q<<,o+���)�D5�MTcIi)2e8*89�����k�&�׊���Agi�ʲW���] f��W���u�-����|�;i�?�ȵ����O���%G|�76�){�VlEӒ��Eʼ:c�j'�5\�r�1�G.�&���V'7k#>�������x��[|E�d(P�o|�����A_�B�����+T����)�	Wˍ�˧��������!<� �R�i%Q���#׽!��f�w�T5O����8��l�H���}����K��:8��|]�������*y�DG��CS0arrr�ﺌ��)N��J�,U{PB|H�mf�����&E��Ez���rF�ѥ�oĵو�cf�Sb��1a:��`N���u�;��;������P�:����fBۧ���O�f%Yn�{�޿��xd�������*$�Ψ�BO�����=���T."��
�׸���LG�{�t���*3P���$�`pV]��s�]���0�˗u�B;��d�]�\(�{�6K�6s���-���5�f���kY�b�,� �ey�l��uvVK�G��:� �¿|y긹j6I�{nr��nטo�\^^^v�{W{����X��W�X�K^ޅ�
��- -�u�~N��|1�BBB����-ԧ.?��v.�+/:::�\ZZj�"D��俗|�4�#��t��X�N��)>钘��V�&�=p��:,���1E�A��7��ʉ�$4���ri	ٮ�ЮJ'�N��PHZz��NMc���P�q�v�)^9G�������R��F^B��OL�߇�"3������Q!X��j��v�눡|#!����g����4�����?C����5���/-jX��0N$=��M�{�PǀZ5�spa��|F�ِ�Ƿ���?*<�m���Y[[���~3v����*םP|�W�2נ�?c�{9=����n�X괧�)0I��������}�=ϑX;���������`Z�'�e����"�Jl�!�����<�K�X�=R�_�����Õ��|�:]\��/2��Kt&N���GG��bp��zTĸjn3l�5�����b&�¢=||
h��1$�W15W׌R�WqcR�Y#���3�>�v�L�0��`�闒�1�Mg்	��C��T�{�W*��ߟ|�d�`�Dr��Y�̸��>0�$���Ao���4M�<m �<�F�Yx`��'� %D,�R�������1�#����I�j�ֲ�+#s��f�K <�~͞#�勼N�A��04���~���j���D	ZvcZ��w�eo~>��C�K�bV&�r;Z Y�@5�ֽ ��P�盠z���z��is�Z��(ă��p�f��� g{;;5�=����&�e^ai�˸�UDH���-1H�No����*^�Q�Xx�X���ɮ�}AV�(�ޗy�\{?d�v���/�$8���z��'�ڒ�9**j&W88�Dl&��#>�2�{���VfO|̀�jhiu,ME/}�62ʇa���M�n���;ς�	@_+��@pq炓�� [Q��]R�1�U�^�NNzV��Ι��O�	3(]�N��X
h܃�n�����S�vf'���ho(����\�S}Œ����Χ�+���W\����2o���B�\�C�����܎F>�g�"G�յ��=7s0�5fB ��P�u�l(��M�XmKK�Z�F���} ��b���`�Zѳ���5�� ��_��z�%w�oq��qٕF�&;�!lQ7���ַC�V������	���K�����[�����~�ˇ����x���0R�W�3_���,����Ӆ��\�+1�#�"D�����`>���LjC$�YZ�	˧l7����$&�F{~p�MNN���r�Xzt���j6R�m��9�����T��ٓ%d��' s�n!Z���b\иw�֙39ӂ
�&�� ������e0��iii�K�Z�Kssm�Ly�]H��R��xH��y{�'��b`���na๠:����7�� �#Wc���K��B=��G!�8g�@�\F���T'=j^?�!��)��Jm�qG���5^�Qb���֣8��ք���ۜ޴�n>�`�+4"�L	+�K4�F�i<m��??��8@x�'�j���U	ߑ-�HF]���4�9x�_7I<p��Zi��\=�&==��N���};J�	��ydE��G[��i/{=`�,�o�\�{`m�E�Z�(�W����a�z����3	30�6yb�?h����]\L̬5�8�˛J� �}���� P|y`:���k�u��!>�Q�uϞ�X��G'g���$��0�C(��/��m��zw0�^���j�|L*�8�d'���2�p���?���0�U��.s\Z�=;�;�<1;77ݕF,�o6HMS�)���t˽r��C��4!�xBG.�����bE`u�(2E`)������~�G��hL��q"*�%a6VT��T��o��ך�le�$�D6±���9� 5�.���ևz;.q�Ĕ�M^��9�V ?������&/: �+��^�cvj�iMM� M��|��և�ӡ'_D����A�03�ܡ��@��H$i���3|�����@����C���~�Y:Mc�ޱ߳-����s���?�N���߷q�!QL�`��ʌB��1H	�G����!`[� �}]"���:	Eɹ���c����J`���逬Yߠ��������������q�+�G��ب�Hp��-��.W7�Be�7H�l(Ž����3��ʣ��Y�w���D�p����=#��SW{��~Te9X+�R��>+�X鬚Z$�[�++b42=+&����NWV��&�C��@�>~��~�fj�J�����7�(쟦)�?~ �F��qq ���u�=xp>g��ۯȾ���p��F��Fv���$����ɞΔ��Y)��x����щ��ݺ�R�l��g��_=+�X�:5��tV��^��а��m��(�Y- D*֚�*]�
�dW��*�*��Y=��������C�?&�D��*���-�
2
|�~��F� ]gZݷ���W��pU������;{V�6���:]/�z{��;ϲ)l���^K�fG髨��Z6f����#�����2��$i�#���1�f�܇0'�}�&�r	i�r�Ç�`���Z��D�_,�h��̙3E��Z��Yb�p�lL(�R�Уߪ7�`)��r_E
[%O��;�

[\^������ʜ��/~
؁	�P�p������[�I����]�é�1�DE���yN�� �O�
��<��H��?^v�M��uŎ(�;F졘[��fFF5��u�P?��������� ���N������?��S�G�Bq4����h�����ު�����1��JWQl�-�SQɑ�j���LKg$Οp��#$!�TH(��w�<��IX���#hi�Hr���藯ױ��cRѥ��M�������g �ݚ�_�ܽT�D����!Ӧ}���[� j�9����e8����>Xɼa��K��)d���jg�#{i�Ct���҂R��z��uz��sz���9WR�!���لh��Л�B�[�8
r;2��p���ل,qfxr,(���M ������!uZ`��h�;�i��KuEB_�D^��{�0KT���@��؞㙚����ю
qq�\�I�%&&�?�*<�W]�W?�?'"Է�*`?=]0` лp<�ւ�u%%�i
%ɖ+xl�|��''����v��7z�3%�lT	e#��*�N��l ��ӎ8~����*�;{�ZX$5<�����L��~��tu�QfJ$-	++^ ���@�J������\���`��T||���oN��8�PPKM�)� �2��	�l�WV��P���,�B8͉ͥC6����e��Vqj(�!l�/>ڂ��Zrm�+�r��ґ�����ʎ�
뽇+ݶ���!H����<G���S���0%Ƿ��ب>X�sB��t`6�e�B&tx���XOONJ-;�X��)IdJ��z�b�����*f�y��}m�O���7��ACV\��d�	�:߱5b��8 [�?_�,�ޒ�{�����2W�R�ck��V�l �D9y���I���\���L�d?M�&`Ĺ��4���JA9z��F��%�`i1�rtv6����TW��)c�ӽ����}$�%�@�k��y ș�U��� ˻���-c� 7*j�\�;V���Ԫ�
�Ð�����_6H���R��8#�"&h���9w,���>�yP`g��7��X[[��k���w;���[Y)���H�C�He�\@Nb�i�43��:��?�s�AC$����e��f�e8��È��`�Eμu����iG�і(�T��u.�����i�fck�&��fi�5��	�
�#�D�dڰ�����Z�	�����y;y�!���D�ʤP!���'����}|�������q�ҥK̓n��6]Z�I�����������=:�_H۽*%�#�����?}�]���^�5f
����uj��&F_(	�i�]r��e�צ�kK��h����#�6M��ț B��iժ2,��������-h�G��/��Z��:�A^�piX'��v��������>��Uy
kN��� Zpt�Se�F���	��u��%mٿ���m.S�2\A��������;@Ę�p��^^՜/|�*�����K�	ي��D�q}/�+{N(>��1E��-�_4(6�l:���v]�(��72*� ښ���iZ#�]��xW�dM�l��D<�fX�9ڳ�=U�/��N��3��\�ٮ���h�?�*�^�.��>rH(i��pQ�Bp���'�PS���2v|�	cK�*@V�>~DP�$�?"�&'_V�때��"ǆ�땳d8�8��>G���������8��WKHHp��= z@*z�	�b���ǎ"Lu��5��Q����,��Aw~�Zy��x]`�}�����};�㡊��$nlЉIK{�G�fU�x����|�E:��?���͛7�	I2���3H###ˢ<Ժ ���q�DɎ��˧���Q`@�~�x�1B�8������FO�s�p�^���w"�NFZ��e>VU��l4S@6�����1?�J��?��L���?�Tw�A�ς'C��
�|������{`�Y:k$R�Ģ���GV�!VwwD�������C/Oc�_���C�T	���:���{i�mN�fG�H�l]�1'ln�j��N0rM��u6�����f��1�{G^M�xIG���>!�BK(��w��o��g�N�<�����	$xp!'�F�^"o$$"r
_�Y=�������'��)�XOr�����`'�H#3~���U7&��\Q��z�'��>���ϋ�b����Y����#YԲ��i��⋠�u�u����^��������VUW=y�Ϡ8A�r����9YYV�����+�"�8���C�������yS�!���愝�לi�*f�vU�܊@�b8R��+�Y-���2A�ڟ�Xj�F����zpW�RX�����E6h��l��=�nڊT-`��|o�e��ez�/0�[�%%%�9��L���t���*���2�V������y-�IG�ť}�N�c�O�F������/��>_�|
-�_��А	�2!�22��=�	��n�=�mݍ�5(JQdU�.#����I�r�{�#�9�Σ�x~��	��,@d�ǤD��zZAN�3����������G�1ފ�2d���-���v����5r�u����MP�E~�Oډ�?
����N�#�݆������]p+%�X�,/�������TS�=M���
@p۰�q�EAU�g��&7�M^^>K����2�����_�,P��K:*T{1���Ç���)))q����5�������?=�p������	Tf?Ƚ3�_2
���hAr�QW����#�����ص����X��������Q����F`}`�<j���-������&{�XCSɚO�cT熉�y�[M�h f���Kƫ�w�� +�2����f�%�s���R�Z����(��SEqT�3A/D-��H�M1Z����r�u}�G|�"{��%u���gFbg���Gw����M�h������i�Z�n�ö��SL�?���|rz_Z�Ҳ��)hx7�Wy�`��Ƙ��##�N..�k-��Y�����/<褔+��7H�@H����=���LD���|vO�^�w�wy`f��q	��F���]Ȇ	9�w��-�rv�8�w2��,��QO��n�h��oҼd�6=Pb:D$��f��9$��$aA&L ���z��c��"����S}��.8�*-��j�-��LLV�Pl�������ޠ���<F��	�T��:uL�!Ï����g�f���V��j��,�m�7e;�i�F�333Kϙ�95�!wq9?�G��C* L� ^L�2���\���nD޹o�0r����*�@���;�{�3�:�b>�e�����ʀQ�ʨ	�޷s�w��0��d}Di� A��<E/�!�E�!p)!ezj
)Yd��>�m����q"�+����������g���9��uy�eぶ���?@VB��sz�6��L�t˚���G�]���A�L�u^�eĳT�{y�Y�^�mz���R6$�9��?N��6�|7���R6eYn�gw�NZ������M��@I�2G=�����>̌q�Z`13J����}X��S�>��mYl�6�.���ċ%�� s�����{o~��R`X���CYn��TQd��A�](6u����.{�h>*cg�=�J�{j�o��)G3W׌�o�VnRZ9���Ӽqe"�}7Mپ3�q���'���=�L�J5����;qh��o�k�|��	�������P�+�puՂ��^���6���*1�Ť�#{�����+�O�W��o��iqW�=�L%�A�y�b$��b!dupQ��v��{gԺ�.7�E��{ڝ��H6v,�Tȗ`�[����n�A��h��]�١q�j��w�pOZ?�$��g��^�[tC��a���}���69�n�������tx�DƔ����9�f�^�2|3��j��[��Q�<V��>��G(�2}��<����¢׆e�� �׍���~\��m������&w�f:w��]��{+�o߿_��{ �]��%}����S������|�V��2k�^��S���d���r�V��O�S�E�*������^iۯn����.��X}ek��=p����~j˧āCD�P��N��~ԡ�P�&��t�gO'����D[�ۯ=�hٽ�����45�O#xJ�tĊĖI�Ǐ��t��u��a��s`�5���7[�y���W������Q��Z�XWZ��Ӿx���0�!K��x�����|<=�����&��)��Yk�%r��%�q�Se�7E_}���HP=���Fߗ
��ӷEm��V�������I�b�#�y�4�Cw���o/�X�4�R*i�ׁ�;��Y��H��ȧ$Yn�9R�5Y���^J���o��3g��5�DFvh��M����15�Z�?��|�c�m�� ���soǷQMee�>[}�MBr�f�&>^o��{[G�w����t��$����ނ'11qt�ǹ�v>�۷;���)��yxZ��T�[���{v�7��J��貀�鎃fBǋ��zS�<j3�l�}W��%z4�va��/��:�7��O^y��5LȚa��^�?��|���TOXx����p��p�7�inN���$w���|ģ���4��54��1)�~���ӡ����C�^�tH1o�r~G��i��<f�r���7Y�H��gEv�E�n_lcL�ZJ�����$�n{�|n;���ܼi��%vq�#{��~78OH���q{o�/�H<�5��td�����W��_3��~���}�Q��	3&�eY�5�~�$�8�|��	��k~���J〟9��m���UEDc����W���������?�T�-a&4s)V6�#�7t�5LgЬP���&-��f���֊=)�бG-�?�<��3���Y1(��n����m������e�
�p�r��s�'��=<8�3(&33��������K�z�||�C�,�q��س�|."�R3�O��9~���QX�Ya�'<M��Oc����g�,g�;��Jw�9gn);38x�V�M�p�����~����j�)��,C3�n��1�$�3#_'6Ϭ��&��֮y)O�N���@V�՟F��b� =�~� ;�^�cn�H�:C�6(`��������� �/�B��n��((:���RC�C�Bm�Z����b&�юU&%��sñ*Ԥd�Jen�#�ee�-,�k����>�����x��sٯ��{�2������y�u^>�d�f�
�:	-���"��E�
�b���E.nn���ZCG�������u,�����lN���BB�,�?"�I���Q$�:�WI��^�ɖ��s䟉|~���w���.�
��v�w�i�w»�ˑ�1��#�N�(g��uƈ�m��	HH�x�RK�ƨܼY��}
,#���o/������g�og���A��6��v�rMH���W�Ep>�*RY~\��>��CrRz�"�a������No�J0H�hCv�Ԩ)�yY٦�an���g�޽�����fY昹�Z*˰�Z��(&���y?�y�@�:��Z |��Q�&1��|RGA�~�p����Z����'��@.����P���N���@/��b���r+=s���@��������x��]�R��x0�{,e��V���9A�Ӏ���Gz�{-1�����*��V�JZ��������?�1�6(����x��ϥy�F���/� ���;��0�fBUR'�VEaG��,�}���I��w����E4���D�_�hI�La�ȜY�"��m���u36���ϐvXŧ��4��{�b��#7�;���?�7ND�k��hjI&W���-�ѽ��[���I��	�l��K���f2x��]�y�4��K����Z_bL]��=��1��dxee�8۵0lic/�\�1�!_�^�o&ًmmO�4�l.�!�q��:,#[�����ޞ��R��(���܏�.6�c ���n�U�LJ~����œ/�ki�ڞ���Fj��Z܊k�ԗ�xrS)�jRx�36�Ѹ鷵���nxj��U�54�v�%�/��Tn�Fe��ӗ�(��\���7��ך]/Կ�`1��u�X����w�o�~|��&�����k ��ॎO��О�yp]�qK	hT�O�ߓ�\��s�2���^X𙙥\�yb�B���ƈs���G�F��E���et[c�/K�=w���1Gr}�H��>�V�����S=�p��"����	��cimt٢̽,�U���B��k�L�������a{��������"x� �*�t^$m�y�9~2*��SCj� 	ʅ�~�
G1@"��uޭ���?''�!��mL������i�������q�4�������5x���z"d�A����q��C��Y��ߍ[�T	޾����޸Al�  ��!��n�̰T�j���HLy0p���˞���u ��eއ������r��8�x�C-d��H]t�a��fc�! �/V}3g��SH�y�c>9��2��ޛ5n��}w��7�
�jHV�w\|A=���s���>W��n@����3lwo�4"�n����}��Q<��ɓ���o[;;��k&���F�[�bk������W���~=�eK��6��Na���&pvu�����F���^Ʊ�����+Jm�}m���!T�qlᮣ#G��MF����Ǻ�}?m��t^�_�A��!���Ioh�8p8Vz�ܛ^_�x�78�����h7��$�'��?A���P��>�<���-��we�%�bv�"��
�������~�i�6�z�잣�A/Gᤎ;ƾ��t��%_m��+��,��|7,w���F�ł��r�ذf������ě���1%8�SJ���]��--��#��0�)+;��y fP��tP%��oa�g����ҊG��4X�n�ڻ�����.��T��Afp���U&���W�PT�7�t*���fW�f�W��ܛgW���@8������	�,m�E�苇;ǟ?� �me̪��𫍛���I"�ˡC�����6MO\\Kmn{��������ya&%��:"{�����|��B�>	_��;0�t��Y^���L)�T&~ϣ:z���D�\��3.7,�g;~�}���mR���Ǘ��h�f74�)����o���N��P~��nΡMsҿ��b��{�,J�&c�ڄ9H�#�8��0�2#Y�?�?����y?|H��ᘻ�m-�Z�@;�IӔy����;n�ftE���4��ue���q�{�oѤ�r�\ �K��Y��@�f�P�26O޿�x��|'�	OП�]]�2\O���z\���{�贸v���H�!��u�H:��y���+@u�	_��>P�9e�O��s����/���	V�3Au���+��|D����j�<��,�O���fЭ��)���ƬE�06ߕ�t�2ɷ>Jr����v$y[J,M���.r��k��A�ϟ����ʮJ�D�k��T�P�+�Q�c����>H�U��~�@o{�FG��eT�����3/y��t�3��u>}�.�s!�����.g��۷�G��0+>ZvG�����4�����xr�Pv�p�~P �Y�o!V��q��9~e�¢C�l.5d�=���U�l��⚬j.��'�;�т٦��5 ć�K�|�y���_(1�8z��;g3�s���(�G{y����(3,V���l�&��\q�~)��6�-*�� �<ls6*M���xƳ9���z*��:��K�ΰ3Y,���_�fH��py�}����>�<��	W]�������:��F�֎0���#�i��}�^erc�f�V���m�Ko'ڮ���؂#�y�H2p��z���^9�y4�x�ax���W�%u��R�}4;{闇1]\����33�ۍ�Y�[�ۭӷn*�?�~yY�*�2zW��"Χ:�A����$Z�n�h�wc�_���y���$nA�0��ks�;�NI �C�ɦ��޽{��A� ������S I�ըy�ϻ"���d�����v����y0�$���_M|]�E	,t�n�?�afBa�t�dOT���c�c�9�t"Z:jvVW���:�2%���a��1��n���X4��9�-��i�j���;l��QTt�e��\�X�h����q1���;O�w��"4��z���!w���4��Ю3gΰ�4���b%@����h{�@�&�8�}��,9t��aө{�7����z.�eq
?�y�e���x�����h$"�5D�	���D�����cbN(�����V��!�	c/x�Tx/$�������S�XE3!BʲߦZ�":��C<�c�<�u���>���2�yi�*ZV{��F����ҡj�����)��s Mi'/Yݿ��Q�O�!�W��jI��4[!�׭�?�������W	edeoB:���HBfFd�ʖ�Yd��|#�!��:I�W���������o���ܼ���z>�������z���a�%�B >�۲����P�s� �,� !<���6�].H�/�a-���D?&���t�$'#�@��X;8���+�������������թgOk���LM��ξV��ә�t*�����ވ�~w4XY����f0�S&o�C=;WV�|�����n݂b����fnn��^�3;3��Һdh3h��8hd�U��z ��0@Ɖ��`���++Hk�]�mo�m�(��B��R�o�v�ѣ9���=�B���qh������S�z�iJ.g���}� U�J?ԣo����tV343���~L%�thH_�����f���Q����C�#uѱu�;�`0~EV���{'��~[�2ַߤi
�/�֌Y:sPZA�Ze�4���x
 8}�+�G��_Q�uw�8nke�=����/w5+���X�u�ӕ5��9V����rJ�
d��_'�re�KH���$����f� 7�bx[0�o��X�m��=_��܇Ů��o�w�z{*��X�D@u����#诤:�ܔ	z��a�NK9@R��}V�"��M"��K��'�P�_q��J��&�x)$-��U��+3W���'q�j���9��a�3�]� '����g�ɕޙq��r�{�j`c�M��Ж�`�G�NWrWj�#�i��\*!!��@s6���==�GF�o�U�&]]��L_���G�3��@%�0��Ě��b�,p���i��{�Er�l��E�R��II?�[zWS��e@�4�(6��I�8R��$�?�Er��ru(W	2������Z�}Qq�`���Q���!��7(�P�*�ŴM���ݮև�z�G�1��Ύ?	�.G��!�1�_�O,��଴>Fs�H�� �C%���ɱ��)���2��,��� ?>X���a����;��������i�N�8@��v-+s����]�����5��ۍ�Vo������~Ŝ�Jӗ/ܴ�r�q]*��˼���""�k���P����n�EtN�⡖�`��}����R���?� Ӡs�)R^�>9��C?�Һ'D"1������m�MNe^�&�A�!�����ӓH:�x����Պ�ʮG�4jQ�3M�^��+�6L\�Z��w��A�k������� ��c��}�r>>[?�ǂx�n�ä{ֺģآ���@(�l3(���1�� M�M�|������Z9+�T���1?���[l�j�Uhϡ�L�Y�h.�<��{�I��'NU(�Nr���X;���%%E0YР'����J�/Ts����Q��5���8G�I����B!���({�ʡ���%��ALq�5rC�a��T�5�&�0��A����G��"�o���ᰥ(�k�1o��GoK<�L�Fw�8�n���\�%"ϵ��ԩ����mw߁e��l�!�0�z��ήT��gB&:3D>>����oz	&�g��BCgr�\'	n�TgQUE�֧��2F5���CN�葶7��&�̖WP@���P�d%+��Dx
���z�����R�;��{��ȯ��Fړ��АL��̮G{��z/

�n����om�����C�� ��͍��d)�Q ����r���lePP T��fQ�<�v���)����n�L��p���c��&�W:	a��n�6(w���"���U�ԭ��ͼNL��Z�=����k��
�+5=;��&姅��_z�D��Fcc���,����3���47W��]��NQ���i�&���KL>��i�9��o�iOOv8ԞԠ�/x��Ƃ�`�1�c��j�i�ő�w�~`�@��Q�N[��}��z�8�v֓=Q�����
�EA�'�pm�$edex���f��H,A�Z�ܸ���s ʟ�ΐ�N��#�:�n���}�'�����JJ��[����5m}���i~���~SSww�۷��~C~�SɕX'=`�Q��ï��U{�������>�뇠�d�����re�ژ�$�&4T�2���oj:ALӥ�<����c��!i�Ew�z�%��g3��Amm׵�[�Œ�x�d�5r^ۀ_J�K	9����=���R{'�������5n�<G����+s�Lu_9��wx*�
wG^^^XT�d�;���C߀:��E��u����.��#-��3�c5x�=��}9!a����
��ָL`j�M��<%�ׯ_��tjA0�uo_nϪ��Zh���f�#�񀋋�u=�x�wM*��%z3�ޏ ,S���߬Ӭ��*�KIO/(��C�,�p�P�y⌜Q�VO��M+�vVQ��_W�}�4z=""⿁hC�@)111�B��k�!G��9���.*ڀ�	���*� U��Qg<��F�j��o���n���X�w������Q����!A�0�߿�(�[�z�=O\�p�m�!M3J�S�� P�%_F��[/gJ����r��w��hv�}xH޽�L�!����78����cܜ����K���!%
x��u@߼��Ȫ�bpp�I��c7�i[��";��J�J��p�~�qe�s���t0�]����hy�,E*��_2���'Cg�������#u�����;��Z��3�N�H���٥�9��6�$�I�2Pdsϑ�RB�QE�R�7�����b��Ĵ[���L�l׀�ba�x���u���Z����,F�\�|5w�E��ő �_0k '�%��I@nu��� H����SS�2�%��[�Y8�|J������n��q��j$~�n�/�w���j?u�1��NZ���(o�U
���ׯۜ�;j��N%''�ӑR��#<�0��f��#;f�뛍h�M��ؔnUt�lgn��,��f�?޶��j_<%�D~�>8O�[����iJ�~/Ýә�������[�3��g��3@�v���'�|�B6��hÖ)'�����������b�٠HǝN��yҟ�����,��w��x��2;ղ�{Ɩ�Tz�����/��i_����ĉ<t�UKo,�`��h0���?Y�N�0i���6p�@�M޸��BT�����뢂�<ؽ�V@,�IE���V�j9B2rrS''����+��**�>�Ds`/��'B��&b�Iy��H�
����Éd|8��$O�(�����w�.P�CQ	ķo�Z�L�K?ϯ�<�'��^��Q317gM���Qm��6��JΚC�����~h�(��H�W2�x�@�� ݫ��� '��ۤ�	�A(�$'�t��֟����9�R�x^���6H�?�00��0�!�(��?�{{�.���UU'?On�Y�Y��蘵
�ڊ1���.:��gUqG�-OQ0q��g~��C{���kQƣ�R��(v�e��*�K�Ǐ�.ɼ����)���#��e)
9v�u�I��EJL���6+�>#g��#""J��PZp�<w�*\��ל�����erP�r1ErQ�J:Y��X!饜�*��>9�UQ��M�=<�Z�̫���� ^4�D�u�e)���gdp�'�L�L�"E��f�~Sܺ|�������*�?�
'��xv�d��|ae���0�\+�Q��<�/��E{\/c,�F�WԔ�7$�E��a�I���@|k��qs0��D=������{�	"��w��l.�KSQ��Cm���K��b�v)�5\��{b��z��靝WIw���=z�?8�X~�Z�8��@��"�'/'W� g�٨H?Aֿj�o�OT6a�Pd��-�/��䱛"Lv�ަ�������]C�FC2���P�f��*R���K<r�q�7������.�m�[W ���P�O�^��>>�,Y�f�����g�I����~f��I#D�A���8\^�t��Om��`�D�Ɔ�-w~�Bssw!aa��"�o��8��%R�BB���N���G��F5�k���Y�5�=��JJ�<~e!��
p��j�a��	�Y���_�6⏸T�^DTk�0������4��/#)��cU��E����122���ʽ������Ķ���Pu�d>$�������0c�3-�P4�3A�J��䖷�׎�����^��T"۔Z�l�RR���V��yc��o���_K�K3PQ*Q�I��g�4v��u��^ryj��uF�٫=�L���F%��ؚĳ�'�#�ﮪy\\&�����Vc������o��_�������s_BZ�etTP�bָ��� Ț�M	��q��!3�)i��\y�O���d�L�\��z�ӂ@i��ݫiBr���2�&�Zװ��jkq�81 _�B��5C�㿝�#,��x�7�H�`�T���?O�ò�(�>���ϺT�4B�HE�i+Mt}�a��tI��IIo�ּ
��-=�~9��_O����`�f���z�n�߇�BC�6%���s&wL���k�NhV	s�Bx��Urr0���ZZ���6ށ1jn���&�r�8�/��{��{_?sTo�����<���#��
׳&"�Y�YyA�s���R�K���~o���h���|-	z�]T���9�>jjj�jjN4	!R�˓U_�*HBx�b�[����'��2�i��pӅ�dM8��a��;����ij	�'7�F+=�43���&����dEN�=�_���b��T R�H�g��xm�}s��=#W���P6�Mn��p�ۖɕ����Zڈ�/
C�8��y��𡰄�EA�Q�DWV��ŬF&?���͝�RX �<<|C�5��g��3(K]c2߻�+��ݎ��l��v��ݔbk�����Sl��{��鿺J(.|�o~���ޞ�-:7�1�b@K��󒷽��t<�N�j��?/,�H����i�g���q����pV0h��j��H{s��Y���uI��⫢/�ZO�C�_�D��mF<�op֞��PH�� �u�GR,@���Y_-/��,U������8!�}**�i�7���w��d�Z�����������3��753�y?�M\��c���n��}�Qׯ#�l�� ���e�G�O��/ܚ��m�iz�\K �[*x}l}q��D��5"Г�����xx`u��F�c���f�Agu9J0�f��h(��ޤD�0E����P�eQ�w�����l��oo�����0���R�mW��kN՟��%
i;)�%�쯎�#ћj��^U��#橋o ��qI������.���iC�az�����U����[���tD	9FfQ܍��j}0
{�հ�O/;�84v��adѭy�Ԑ~�,V���f��ǠN��&6}�b�@��ɤ�-|�Z��`O5x[𧪻�E`L~��FDF�����5�.O��E	b	��� A�� )�����ڜ��~��J0�ˋ�����*28<�z�3z}]��Z48V�2֒�ΝM*2"�^��i]cc�kT�G;��K���_{�Z��N��Z树^Xڷ�G>�E��R]�)k��?�U>T%�_u|$S@sae�6_���f�ձ���;��G�ѥ���BBB$zuk�CdM7 �p8M���pӀ!8Az�"at+�t�A#;;�X@'M�����5&?��Űuc��Y�<a����maL�PJ�Sa����s�r�k��'�ĎTz�'�?�<N�+VZD$��n���r����1/��dj�<sڐ��l��a��iM%w
*���a�݆�&���[�!I�8X(L-,���$����o>2�04\�ܶ���-cX��)��?��H"��o�{my�~��izU�|���k׆Xx��	e?����؋o2�.}�	TxӉ��A��0�$)�@���h�e횅�����D�"liD��hO�����3~�彈bS��߹s�$xA�2=5�MJQ�>��Ī�&C�B���W�
k�Y���ۭ�n�չ�b�}@���~1d��?����BO�}b"&���yo�,mTT��iWrZaa�И����g�f�^�l�E
;+��@:N���5��H�S�P�oݯ��#����c�t���+���,���<D���U�^nؔ|�w[1�yv����빹|@�Ǔ��� ]�p*n�:�UG-,����_{��Ɨ�.\�1G��'��g0ۓv~�74;�/��]�{�$�)�LE߫���ZC���"�#9H��7��W˻i {�d�7�5�v�w�d}�@��L�T�O��$%%��'��<h�?��-�~$��X3&�'��-����& :_k�訓�Y׸y��_�J�͕Z#w~Ʈ^BY��vui@i�X��c�t����Z�)R~R�}~p��X��P>==�@%����6L�̃��⡶�fU��S��0���h'wN/o	'C=T�}�ܔaÍi�Y�#���w�Vn[<���/���˽����V������!��6qq̏�������1�OU���Pf� <���]OIy�)�>V��k���11T(��ё\���G������m�g�n&�R'Xfh	�\[�E�Ʋa~�&m���f,a gDDD���:�@�B�1>9V�{R�������\��i��6����Z�),��9r0�&$��	͚ ��KQ��}���������,$��"�z�֙���NwD	N�qE0.*�b%��0ٚ=!�4�ޟ��qt���!���Ujj 
[�b2����7���}�#�ݜ��f�++�
�z���א-~J9��GdYY�IRmӫRR7$S���C��>����N�`����j�iT�NIi��yU8hVr;��f_�H�!���[g�R�S�QeJ�w�CP�r���v֋�n�K�
W�>�m�c]�4��iҞ�\�'�^��_����7 �f�|�=_��c2&^��-���TUUA�L��Ry����op<�j���ڜ�2E��� ru������m;;����0��#�h�	J�*�)j�i��J}�G����7�-e+��;�}��suk;�]}���� &�a��Y�-�� ������C��]5$6L�l3+�� �Δ��T/!`6�7�)pq~># D��f�]���
ٱ�##`�`T~�@[,�VLݳ"`��� ݛVy�0�ys(A(,"��%��E�Z�h��T�B�Fy�X48J�Vő�\����M1l�{1��wE�2ńU�4^��XI�9
?՟��J͹i��r��/]��&u�{����J���A��ƺ�[�0�:�i��� ���L��o⽺ T�**����L.g&����8�7�35o���
���ne��0�'G��/H��)EZ�����1�(̤��*��Bd'���%d�$@���Y���1� �[�}�E:&��hB�L~e\�8��pexE�LBa���!�0P�Q���Fk�fO��~�C��sΝ��5��?[x�}a�""�)a��@x_�����p>��)Wד�D2&��'aP�`e���r��Rr�����Prۃ+BdYr���3����ԡW��U$x�7o3�=|L k:�*��EV�0��h�У��}3��,l�į���N�?����[��"��'�:{N.�$K�0v5��@���8͇��N����^kvC����Ca^��Ҍ���%�%�7�||�ݥ=[\�����+n�������8A"p����)(Î)'S2pM/��K�7eh	�ZH���:£�2>΁`��ǝ��Ut�HG6���r����ֲ��A�"˃tt�Bt�R������V�H>×ܞ2��rRc�[^��־��7��S<�fL���a��g�O�/��v7\^ZV���R�7��J�7L,��hl1�&���,ٯ���DȡB�%7�Bj�}�Kd]���u⑾84ױ����O`�a�˻'*�f��
�y���lk������3/��Iyo1�H�QR]���$t�8�Gcd���I ���r����9�7$3��w����Xv��S�`����;*�3���w(��p��"���o"��2d@��5z!����8o��n�D��@����i�26��w�g����yWU��V�'���%��`�N�Ğ�3ɓ����E�,��ڟ��|��L){��{�%� H��f�s�-c�n��=��t�����5���k�VY�`��C9^KM�3sq�%�U�־L6٤��V�Z\��̴�u���޹g�z�n=/�?���1�긿9*�օ��:.��1	a���p)
���TW�E�b,�9xӒ��༏�ET�G1��>7X���-���0�����ݖ�8s|���Q�)�`�(���-�|�mz�EYXY�p?����A50P����\���N�#ǲ����說�������]�!'kzt�2W��9����;���ڜȈ����BQ��['N������Ρ(����&�'���$k@� :��rP��Ʀ@!���s�I�JP�i~}�H3_D�ךۯ6�P���SE��J&X�[L��z~U,�)`	Tb����&�L�̀	m3�,ņв]jņA�Q����f���<fܯ4��V�Ūh��*'L��TL�k>7[���ih�w2E���j�$��6Y�	�7v,���p�{�����_uuQZaM�k�!��SNFq
<�w�=G,z��B���7ksČ������rmꇐ����Z��?	b��% �Pd=es�G�K����������H�U6�R��,\s5�
�Mlө��/S��/��lū,��a(���TK�*�Qة�*S��]��)xWR���6O���>8���J_���fY�Nv��f�cӬ*��M�s�K��iO���щ��x��0G+K	��@�j[ �.�U����ﶴ.�����ih#q��O��"���ϻ����s{�G�w��B��1�9����O9��%������>��Bl��8�M�[�������f�?�wo�Bp��_n�>�fh�.�kH��KD+(���W�sNUM�|7h� �8Y���*�U���R��WB<�m$Y���q�������?9��ҲxC���8�@���j�ӑ��A"?�1%���9NEjo�x�2��a$�7";��mٲ.$b�XH+ҹ��3aq���H�sT�iݓ�D���h����l	p�m�,����^QY������8�T�+�2T���������� �[�8#�<�g}B��#�h�����
�����}]�����Z����+Sɩ{� F&'i�v�]R��?�U���������Г�� ΰ�:Q�|��gqq�,ll�B]���О�ɬ�����Y��{6m�KNNn���7;H���ӈsa�"�X�X�8[W��\%�QV�$�x�c�r� ͅ<��U�k��'�D�6�o����!��s������A�<�Pup�(.ʹ��L���P��͏SDP�Z��К�}�I�#�O�s��_�z�O�|��e�e�VI$�{}�.�<�2�I�p<����{ך[
K	��W��`���L�������(eS���qZW?Q�GZ��%0d�F_W|��/ ���J���/��fWa.��뾱r�kt���ĺ'�R�S�|�VW�P�c�e?��7+��IY���,�LJ.����PE��!�~`P˽�������P���n^E>��bᑑ�R>����ݍϑ�'k�!��4;+�U3�/�	,;1aJp�y$?p٩��+��gv.:���� |1;�i�y(O�I���#������|-�XH/6�H����(�y���|^y��J���ᚡ�����N��Յ/.��A$�#��W�)	�vtI�yC� W�f�jО\]'	n��{�=���[����p��ӭ#5�Tћ��ڨ78F)��f���w�&�(2��4�^sO�ܟq�w�`��i���5�Gv�H��4��TWW��(˧�໕�*�iB����>Mf	��F��o�dJ��9����;Z��/��d��Xk�6#��/,�K��!���w�1E��fQ�dA#&�#Z)�����ץ�Ɇ�NJ�~�8�4����\L�{�����4 <2�;��F	�p����җ���qy�G�|\U5J��ob��h��%
��d``xn�ğx��M��9@!�Ӟ�W񺁠8q����@MY���kj��~��{|���aw�͊�Kv�s���2�/��P~5y�:����2�'�8n<�#|E��#�����󏍇��T�a]+#օ��\��[�z��K�ꍳ�ڤ[��f�ÌoX��;���$�U�?�9��V��yu�G��}��u(r�R���{>�2�ݿS#���=��4)g�3�̦�a�=%�������[R�o_��okm�t�D@������ͦ�4�k��榦��2u1�*4���%����_��2�4�����~{$��B�;?(D#��i]��\L��������㓧c
~Q�x�U����"��nP���9;*�~�Q��N��!�����V��ˤ,�։���Ndiha�/��~�Q.��G�X_{��Rbv��"�뗘�7e�>s4&'�� 5	��%>74�"c��n��y��K<n�]^�k����\�еk��X��V��%p�H�Pu���s�L��ڻ\�W��6S��+F��MSH#����e�j.%Y���%R��dr/��_����
��Q[W]�˳��YH�6!���$,	���-Rl&?�g�wԁ:�WGQ32Z�{����w�[����ǀ_�Uv�33��d�ls�j�
_��_)�b��.)�K��]؞ק��9Ԩ�1y����f3]}}d�LD��S�֛���;9�+e��\}�"��tpp���'Z�t<��`w�#�tz����|�bz�h�v��A��%8���c0�]	)�r6�u�`hy���T�A��pJ�� �|ᙯ�Ț\����aIXq����	�↛;~�ylс�^�ecg7uw�mͣ��
<yG���5�h3Ҡ�S.��&&&�01���a�N]�����J�{��=�B�0.���U���-?����meo��%6�7'+Y�Vn��Z�Ą~B�y�Ӻ���ǯcbR*�~zzv�D�T������|����  ({~'8�W"U�{��q �BX/ �)ϭwȮD���(���7jjj%ee#;�=n@�X�渋Qu�r�HI�!��W��ʨq��X��gώ)t�
Z��F�W&��^�t����V���� �S�Xs���%�*p�n�%Oת�Ɖ�(�j&R��0o00/:h�k���;�o+�!�V]�ٌ��,��=$Ğ'���E޴��P����+�����3U�;�L����)���4��PUV�ΙB����&��G6ҽ�
���F�bH�F����W�������D��_������Y&�=�-�@D�YkU�F����c-ܡ���x0��r��b;��#��}Vw<�(�`� ٶR�J�X��������Urr�k^~��i�)v�H�<k�Dl��O{jM���U#�~�:U�������m�����d����w���,�?�"�(��+6碨
:�!���~s��b�����I�����Y\k�����Β��RR�����Ƴq�+����^2f+-��{�URۃ+W��9eՀ���#�h�V"�B�ND���IY��;=�	GB�����aqQ�f����E�~ݳ��J���R]Bc�d��\(��~`�Zf�L[��N����^`���ž�a�\�+[�ω&c����@ϟ?/��跢���p�U�V�d���2W��m�Bs=��.���2�(�z50?�<�桴1o\KK���G	t��S�1�+f���z��-�����C�%##^�d�ݒ����� d�ܮ��L�H������X!��)��:��i��{UZ940z��KetO��pŀm�\u]��6n�Qo��Y�����'V�;P��[+.h��\�eVƖ�5��$X��:9��9��o��wٲ0�T�Q���*b������ܯ����N����IG@.�����<0�̭Bdo@x�sʾ�fB�][����L�X��t���>�6I�Ut+�����5U�!���~��[�`�_|��AKE�r�� Pm�U�᭣
�G����o��ZÔ����OB+�J����M"Yt�l��%w�T�A$������LD�f���A�)��gl��)�*<������RʕLL^�?5�	��t�MRjj$���(�P������N�:��201�7M���4]�e�K�Zj�� �R��tc�->��<S��LyK���I����,H]���"�U���v��N��T�Q���4u8��N(���5���y㽟�Bn���d�x�����M���y�����6�>�~��`E�������ӌp�	�������>�:M���_���i\Z�b`O�9]ӽ��3�~�A�9R��W<}>x��Lक़�4�݀`��>2G��h�JY��i<><�`Y/>{��ԓ�I:6�=�0�����G:Y{&��9�|ؿ��A�wK�L�����{7��zV�uN����K�ld��7�9kw����#p��!�4���ء�%OO��GN�/Zq�j����a�1�B������z�� =������{_C�����4�>�2�����AI�Y\|�ך����+��W�[���O�[0^V�98R��52e��m�ኩ���`0�!�u��,�����Y%Ţ��dM[�G�k�G������F���s�t�{�&!�J�g~�FBJ
o�/kЖ|�`aUj�ˍ��������p�����^��?�֢�˹;������@a��w�o���0��K�d�t��G��D%J#_*¼Xҁ��e�Z��*wzg���sK�Z�+:KC����:}���c��C��8�h��|-j`;Wz�R���])$$'�2���LS\�ڭ��ëN�J�WY��3IC���+�{o��Vfse&ɉ2ٸ�G� s?檃��s�i%���)�>��:����/�{k�$99YHE�Q�0<����|09{�R6���9��s|#�-�t���DT�����Y�X2��mB8E� ^PL��?#x�rq�2X����c��*�O�Zy�۫1�$�����ln�9=?���2KG���%��I�G-E1�����m�� �X����t��Nw��T�kkٿ4	�����
���`̬f��|�=q"H��%
$@�-4Kُ�9g;�wt f��S���2m��[:@���7E�a�3�;����&W~�.Z��ҋ�x������ Y���_� ��>5#I_���o ��x�9
�_&�/���mtO�2�L �	*w��U5jT�%؋�J�b)��(s�8}=���}M͵���Y$:KWVN����^Q�A^��g� �0�(��7�`"/'ssW>O���e������B��Z^�>�|���,3ٛ�Ib�++`q�.E�	����v�<���9Y���E��9'@G
7Mؘ@�	�	���}�;/�@5�����>��չ��L�֔�\0<�"NB^�PMqT.�����o�[B���U22;��Vp龍v�B=�.�;N��,,T�l6]H���\�,���%w�������9}�4�;$��K_�&q�x�D9VRQfuM���[0�Ohl��+�11���
G9޸����JJ���/䢻�9]��$�y�(CK���~�.�P�?-F~u
�;5U-1ND[N�1�Ի���15�_B*�$E��A�W9Of}+�[�LML��x�IoGEG#ۊIy���ee�	֛n�]�J�#l>x�#l�2����e�����j�N5#�b�}�P 1`����D�
�<Ea)	���d)�
�$/9¸x=��n�?v��[q6��jlu����
Nzu��-������&I-~W2��[��((Ƹ3u���J30א�U��>wf�KR�9����9�0�(��ԕ+�$�M	s*�O?~�fv=�jU�(����E�$]c�[(:�'�\�F�οS��T�2���<}u
-�R��[C�=u������㩚�A��wO�޿�������R0�]�kdg�?&|kD��K |�3�z����ۨ��~��m� ��(���
˼���F�ˉ�g�����i�}�����S�
ى�"Y�ˣ��ߓ?�Df�����z;�rUG�.0�����jt�?X:�Lڭq��˝����b�*��C�Ρ��NG܄�iP���=�����>��k�֐�ly ?�|����L�+�~;T�lj5f�o��Ö|�X_b����q�����iU�}W��d`����upW��p�몴�Zj��-�~�ڊ�7��-Av�~�zE�b/$K�F�V�����ΐ��^*�'�Tdv+���p��ޘ��N@�=o..d�0 �+{d���}������DG΍���ͭ�uT
&V&o�Ӆ���^�P�&�����P{���Z݋�9����uv^ս_�W�p}a�`��������b̋c���^��ddff&�h�0�0��ں���m�J�\O
b^�\JBf�"*)),��&�I9��T�����v#4M+�� ����,��M���1�ŗUh���+Mi7y��vL�́:U�K
P�+����a����j��D�tiְq�J!d�{҉�Z����uk��BH�ޛ�p����hv�V�����.����!�^s1��#j�wpITelJ����|�L@&?8�2����C~ Vk�Ό;U����;��HzR�=�Pҭ�}�w�:j}]�'��l�0j(H�11C	�j�	Pqkj�J����{�3�'?ٻ�����˴�y���徛�k��%��{�%���_���P��m��M������n�3N�N!���C�.=�����q_�T���O˃i6�p��s?~;]�{�R�������',N�~?ZC�9ȴ��Lx������{9i�Du��K\��.HM~�a0�OF葵�[2���0�f�k_�� ��F�MKq[HX�X�B�fI���ْ�� �0R���Ȏ#��#��O;�ږ'�������_ݝ�ZF��ji7��L�,�?�������t��*��>opӳ�fKl�I�)��f�����^EX��	d��NPu��f�
�5?'@�~���'8
s�,E�ݠ�[k�E���z���S/����z��s��pRB����i׽����߃6Y��!���C/;Z_��%�X6�OQ��OQE�wģ8�"U�I�t���f�:|��g������g$�n�AY(}���@�P��m�ߢg&���Z�-:y2���aۃ�yYC��3lR�޿���V_?��^�r�c6�2�G����H{G_Z���D,q�UXb���'��[�^����hkʨr��(kk[�B�+$�Z��Ϟ2���ݒw�Hc/���]�M��l��p��$�=kGj�Uy:.��i������V5`?��ӀT3+	1+yz7>Cnf���J�uE����؃��֡�v�J����;�<_�}�-���kk���-�\��<	;��Ɓ]Oפ��x���}G��.OI82�D�{�I�#8Ů�k�Y �U�����R5�g���-�w,��0!'
==.#����	_�妺֨�GTU=	��m�8�l�?l0�b�C����g���.�����|*����J0�l�`")�}%i��ݽh�+&e��"!2��&!2��c�}�ID"*�&uz[�;c�K%��ȋ�VSI��5�P>���Eޞz�ڸ���ޱS/x���[�+���x�ض7|���X�I2uEfaĆk������raaa��9��7{�P����<0�{�sB�6�ԕZ�ʣ��
;s���i4����݀O��%`�~�Ђ�D�L�[�X����:��1�e�K��Ho�
��@!�zټ͊�σ�L�)�O|��:�o��;z{?1$��� ���QH�gĳnF��Ֆ����z�1��)������\��v�C3�Q�ìˉT
���T���z���Q�Z]��^����K��^�QB�q����v\1v��|�q0����%+#W���2�ӑ�M�'�!o<��XH�c�; @�?�"�,jbcC�l�q�=/��%o�v��R�Z[S.��:i�I<�\8�st�>�f�+6��'uk�~�"�7�d����WiR`�9
Uq�n'FK`k�uL*�-��[4=�9z�����iik ��p��w��DT�,.|Xoȳ�VVQ1�j0�LmY\;}R���Jp���	��̈t����\�]�B� �o���۔��Xe��/3�Zn�\�������~{
���gq�6]�u9�$�3������7���8� �7*���Iz������Wii%C���xh��녪PRR�:�b���<��",$Ͻ��c��࿷�֒��]�)v�M���L�M�>kv�����[k��K`�<���l.�<��q@�$������%c����yQUn�&�9���?
c����hK��?z9�@#���:���Y��[��2쳰M"��89�4���5���	@��ĘӞ�.�&K���n��.�R����݀V��F�޵B���Z+��WR�T{�n5'���H�n����ӂ�'
*]&��o:�1�4D��ol�ܓ_����\X�
؂<*yK�+sy0D�P���hf|؎΋]υ�O"������E��4
�G�M�`�"o��4~�<m�𻶥��&c<rԞ���	yx1cSΤs�^?�M� N�cҾR�%��&�bh�!��|+�W%o��Ċ�A�B���`"\��;#��g��_`0���Y��:JJWؒ_z3���J�b�9+�}몭\s��44q�<�<����9`�f��d��������h�꓁z_3����q ��A� `��-�x�NZ� ���sH�<���C�=���A��tc��M��ֱ�������Aϖ���Ť�]�jЂ�<cT\lo���勦��(�{���vv�Q��,߾��+ѵ}|y�(,��̌��g��=p����p,t �O����dv�k�r�Så��{���ϔөx��3��$��80�.�]c�
�IU���\�� �wrЦ2o \��ݳ�h�۱<�U��_�.CU{�tN�eTu�}kwwiv�>��=�6�}CB������!�w���O���_gP���$�V�9v��iy��g% �����Y��Q�MNղ�Sh�ƽ=)���;Pj�����#�n��ɴ��e�'�=�'j�����iVV��s�O9H%Sӭ�G�
zN�2E�a͍��n�n/,����BN§`�j�v�:R�P��q�^`�cBޮxH�JJz6�`�����U��k}QA~D^[%(���Ţ�QNCe-)�e��,������)3Z�4A���)�����ހ�Q9V�:W��"�}��zj�>�6G��;X3ť���W����)�ݣ�r�"��C� z����>��L�nIC"��r��du�{�H]��+>�M1v|�sL�W�4�z;]��:?���Y\F�z��ߩ��Q�o�x�{ҵ��"9�����'B>`����H� �/7D��丼��$pGHf����k��CZ'/*���s��[�>{r)>�l�u/���c	�~��h�
���<싽�| ��+�48#y��1����H�S��d������9��Vie)�;d��~C|�Io3����KQ�?{&ո���
XwS:��L�<_O6��f�%5��}���e�\ͮO����������t�������������s��iO�M;�M9AQ��m���V<ݟ�+.	~a�b˳��Թ��ͺ��ע~�T�No�p�bzv�	s��?l�9/���Ae�d���\J�����Ks�����'�i�ro 4$d�+8�Ril�6@�6ޜx{�Kct��JQ2]"vۥI��罗'ʡ�JJz����C@os|u���G2�c��� O�V�8�(��O��,�?��������i�8��&��RP�z�r�|���N�좲�Z�����I��w�[���2���������MrO����n�u�i6}��Q:7��)�Rf�$�(�������f��B����@�?n�A̩�h$�՝u��� ��D�?G{���7c�^0�t9�{Pf�$����(ɱ�ߣ`}G��}A#���NU{}��ma���;W�6����&j�O:��t��">#�^$才�Ç����� �����U���{K���-Bv�^�++�쑄�����G2��d����������x����]�z��y��|����z�^��~�n�z��|�&�n�	3t���1�5X
F��:�ʊU��Z]w㤉��ׁ7:8�A�l��Ħ)s���B|= *���(S�)5L��K�{�j.�ӏ������Y>3�s���؛JcE-����~Qo3wy���@`4�8w�V�n��ߵ�ˠ)�7�����)�-��,��7���УZ�0�P��]fH�Z��ĤOGB�㍍����Juuu@�H������^���?����1�:����������{�P l���C��21���mDZ4�R2�c�T_���r'U:w���|nre��r�*Z�O��:N�Q��.�R\�R*��"�á����l"��?ɾѴkl�{xE?>YN�̌̑,Hs�1��Y�W��uz�6���I̿C�wR�:"��h���v�.�Y�`��Ĥ�l�- S�( �x3�g~�L�#��:�����Z8c�b����'�C�����%�p� �TEm���~�O��X
��@
 �ڥ��4L�-y����g R�t��K`�9`�%ec�E��\�gh���sd�]� ��V��ɯ����.X� ��9�����]=��5D�>����t]���߱��.����|�-�睹����MMW��j'bq�s��Vō=$�H���2���=�.���s=�<H�wmep��������eD2DB��� ��,�h�/��/���|��f8L ��i?����sp(G���+d���E�����
���D�>o��������#�/�p��P�o�0?⣩���e�����ѝ�w��Kγ]3���hXb��뗙�Tʿ��XY�nk��@�NG�+)MA��fhFWhjd��"^��T���ى�i���@'H>��L-�Ő�{$,(�����Y�k��+(��������9Z>}zeii���
:	�A�������!pQ11@�y���vx]U�NI�.�w�ir̇��tO�n�hVd����҈T��֥����ۇ�[��q֓_Cer�2�8ȗ���J:��t***�?�5)���A�%�s���γ�h5�11�6����2�p��g� �ˠ����a��틍-1Ƌ�-��U]���D�n`�y�2��e���q�I�����������e͑)�H�ȆD(��َh�Y¶����Z�^�׋p�Ċr`T��_&LuV<�./���sJ��1E�����D��(��`�s�amړE�,4L�8S�8���r����#��@Ɖ,L��̸?��n� �����IZ�?;H����t��N�#*�N�>��\ %���aEjP��ѷ�m;��R~2J[��V(a��jE�6���L��3ۊN�À��],E�]�T?���?���z�M��t���Uw���j����ը����Ǉ:>���f���=V��5:Jm+�-B׊���/��)o���E��郗%�T��t
\�� $�z�#*��s����bO���u㖇��6��_3�r̦VaajC��"V|����q�	uuw��,r��31=�K�\k��H�s&7���	����EsQ����0���N	:��
�.H�r�X�께p��UņO��y��~��j� ��T�FJ�������X�k�[���Wę�ݼ/��������oO�Ggq��8�L��1��s�����Z��>C������0��[����i�������HA@�R���?�`��Բ��/ǆ���H1 �Y}_}o���(��G	JK���dJ�@�0�����C>��>0,����VP`����'7����n�<G�"x�7u�ʣ�.y`��|p/�����S� &��vw8�OGsdg��
vyXuC�K96m�ޅ{%(}4�;V���9 H���)�#�@Pҡ|���P��������{h셜TF���9���/����{�1�Dl�g>O��v��>'�}޳`�H)�{K�`@��Sr@8_�۷o�B���A譭�wX/񫫠3 ���O���X?���gO/�_��G��.c0U�!�:�=��tm��S�y�<g���3��\��@:�&*hiYH-y�"��뜡����K2�;O�	5���!|24� G�邎�,x��0e�����������]��܈9�OI�Y�_{<=b2[�z�}. 	�'Ř(�y�����@�2&Vf��F?w"��g}��#Ihxy�7Q���U���|����z��]��V���;�#-}������y
�����ҝ����/��(��Y��j�@�ͳC�&�].M��EеB
wSJ�,�ISFF^i*0?T`�ghs����t���pqO�0��!k��o�j�X�8��|�����Wn �l����C���F����'�9L�=>�À�y5��~�%Z���j��rmn��?�9u�T飒����d�>(~55QA23���f�eq�f����c�HY���[�]���o`�cx�[�������x�sV����:�Toan����^���(D��	kc��I�+�i�
:���e��S}��a�߾���Qκ�du�r$bS�w�CUaӽ�^��j ��o�;�&s�ҦL�E��\n]'������k;�&��mqqq��|�f���Κ�׮�KI9��8I�'�Y�?<�h�:����*����W ��mYY�!oj�� ?+�ٷ���)S4ظ���e@@�YR��@:r��1� qdnsI����%G-�����TW�vxz�*N�H���2!/��e�C9*��n�̨���\��o_��dk��L���)���ze+�ƭ���Έm��s������?�����(���L��O�?~�n�	{�
et �Q6���޴��9/���'���B��A��y�noo���B��LrJ;�@��!�����؆�M�����	�{6����D��G
�Ϸ����J�k'�sMinj
��/�Л+)�N\l���!�"����<���!7)fcCX����,@����S��1%7~��↳G(X�_��U���f[���²�.8b�Y���@.i�\[4܀=������2){��>&��Z��EEٮ9��s���p��s��n�a��-�dR��ӿ����gv�˟��E���Y$��r�L���|}�**�D���7&4�u��^��Qʊs�����6���_�;��.i�\�$�ɕ�_��NOO�9a��@���M	ـqS�h���V�89��H�W��=������u�J[�/��G��Xn�?Y��g�X���_�[xV)�}@􆷵�!|������!�:l�6(=�Ur�O=�x�N(+�@}
�6N�am���3Y%=K�s�熬J�f������F(C��Kե�L5`���Y�V�=!w�	�����ɻQ��_��?�Q0y�����4�W�ݸ�z�\k�Kd7�E�wnu���8�{e)�#KJn�]),����;B���:��s�HQN1*丢�b��*Љ�/��&�&m��7�"'�j����!�b��߁�����w�o�鲇ؕ�%K�bOU�ggy �1�=rx^�Z	���f+������.�-�"���m��w��BC[��=E

0k�캟����}�����,8j��-l0�G��5��Y��h�	��)-�P���bL�ܹ��w���bw������"G��1�8=�����)�Db��{��
(�ܘ��g�2��+qW��h���� ^�ҒΛޅ"Y��$��Ç�iԽ�ː���TR�%WWW��Z���Z�FG_� Q�,�!\�9��OZ�x���Z��v4.���f�y5z����{d>Ϲz�%�X�Cك�kq#)q�!gu�m	B:p�l���x���4P��-�ꅚ=%�xע���OꌡD@�#E	�Qv�O��������x��.����l���ɉ��f~��D3���P�j똚�jk�l�*9y�b��<oj��Ѓ���Ҭ�g)S���! �0�}�h&�����F|�O��z~���<��sl[KGx���5F��Up�+�5�7o��¨U��Ռ���@]X�<5/`�8)r<�7�B��|��.��'�:?Y�}�u:�%;�� ���@��O�~�6�K�!��J�i�D*7��t��uZ��˅
?�'�}�ś	TT�l\Vpێ�2L�	�7�4ܜ��n���;���ə�z��I1�4���H<h��4�XQ�xQ&�W�T�����KP�G������ӱ�F�}ij�E/l?�XU���$
�LYF~4+9"�m����ש�C���a'��0���0�e,��R�@�4�`)@ɾ�E�d���'9�|�h0��������øn��:P�����5���%;/�oM=ܽ�\��^�Z���	ʼ��pq�2�{�;?o������d-䟋B����%qiX-&�D�; �͓C��=�$��xr�}^j�5&ff�-�^?�����)��Y��r�T|P�Ql��O�K�(�ݿ��'��Н�V6�μB<�n���W"r���=VA�yC/x��W���a���9/�)+k����oғ��	j�
y�	���Ŷ��^L��(��`���o��6��rx#-Sje;�(���/4�6���\������I�tOL����HJ>il���D��AN��QEy�\\\�R����:���C@ְ3��U�1�8�3���&U#��S"�]��<ćG�Ľͺ�Q[88�B�s�ѱ���j+v�{g	2���m�uHȥ<�o��{{�Z�e��I�$ht~�wA�]��z"m>u���1�$�rݸ�����Ѕ�̡�;ZP<L̄������f㈿������_Q9�x叕��]�h	��Э #����o��gM�>��S�#-}�8���:�{su�P�К��ܸ�Ljo��8*Zu֫��g��1RN�yv�|�ghx�B�^oz�w�{2���i��%s����*=�����\���c��<(a �A�!��=��/���x�0yP���fi�(#S,R~)�	����{��A�c{9���xP�/xe%���A6���>f���%~��I�U�K+��M�J:�!�I�����z�LHXCO�/Z�9�V}%Y����������}y�.�cඉ��oK��G;w9��y�fd����\LA�k%ā|!**��4:kx�̄;EE�A�ϷI�#�Y�� �i	}_�v#VTx����g��HZ`�@���G����J��ϟa�9 �̮a��z�����W������h��M~*�S=/��	5�<y�2Ug�N�,�C��vB�5���w��(��*�U0|�pʯ������w�
>�ss����N-���hW��[{�sp|�����6@�d�tKg��E{��Ւ#^���<�m������{�A;;_QU��4�$ޜ����aw�:&��z�êo��$*�E���_��L�����HP���&�!ߑ!��Z�*��aO\�ґe��k�"��'�G��\~���^���G#yR�x�ī�3�8��S�Hz��R�a��Bj�H�O��E��~�T�K�Ջ���>h I���B����9�w(��x��'������E�؝�
���:)t���	�s���D�+?��f��IJ��cl��V�� �^\ģ��V���ua�����_T=�
��l�Ƌ���0�|.ךxv&�Ńx���r����t���P'����&t�8�������'� ��)q_���KA�'��	�̄���D��P&��1�����Y.01�$� ����X�T��@�OZ���@�ƂB^��	��B�99n�Ԏ�2��hDs��A5����,,����~w���-$�� �蠂�w��K��.x��?����=E��wx8��TTJ�xW@R���5�l[KT��ݦº�����F^��Ew"�oP����^T��L���?;���/��q�ܛ����B^&W�T�IO!�uś�%��4z~R�@��
��l���Y����<VHA�u���_�{��YJ\v��EɦS��TgζbW���:Y����*j�`�����nH�R��Ֆ߸K�ᠽ(ݧ�����Hԩ�m�{t$��m��������I�-�?wvh�%|2���Q'�ez����	��4�d�֯��p	0.P[�c�XR��Pyue,Ql�vC3Eo_JhB�j*�{���s&��G�O�~9��w�`6��UVH��a��<w���G>F����:E���Vx���FY�03��R�֖p�^���b������)7�nF���G�k���#��#�e:;7A�0��n�ʌ�+�������K�Mh������6KJ�&W��Ս��@�R}�̮ޘ�|��8[��m�QW�;��/�7P�j�R��1�-���t���'�7,ͷ��PlZ�Џ)r��~�>ˊ.����/2ά�M	7ZA�+W�\�E����=��0ZͮRSR��R։"F�JbM��.\�"q���4�s=we�z�&�����q�řĦ��y~���aG�*��8h��٩�oG#c��7u��?�(}����f�ۺ''� �$U�v��&����yNr{D�!NN?ad�?�Q��CT��������φ<w[[�n/h��@]t�7W������[^�T&���1C�t(�t��n��w�束�N�p=���d�4��iK�Á�����Ev��]@�鹽nA�gٚ�GLb�6�4[��9��&~��u}��p%^-�����N�q	�X����`e�V#������o���W`��ga�����[��geq���<4��\d��	Vnn���6��wh�`�`�y�� ��*����B��,=��,�r4���r���b����s��>��XҋI�Ƨ��G�� ��x#��9մ��+��h�N,DCHo�wB�n���4�-���������=yش��qh�;d�o$I���c�x��t�dE����j���E�:��TA��^ ��+���-O by�RI:F���a�Z�|�:�;�4����)ǯ�z�����p�q����PQE61�6y5�b0������Ǹ�:낤�ʭ�,\�8����Q'!�8�K�l�
h>��N��F��8��vu�<�quv������.G���Ø]��Գ�'
G�Eu ���DD'�o�>:�y|�ʚ�g_]S�����Vi���VWwwMuuDM͝o��5��fA�T�뤯�()��/н9��C��y2�G�����h�D�p�e�?0+�H��dH� ��q���P��0����G󾚽���wY�x/�s��Wز�ڗ���;�^���m�Y *o_>`��>����0�Ɨ���汍&���i�ts�����<�
����\t��*{>鵴�G�Y"���������z�k�>� ��8ƫ~�q��x�B�U�:��[�K��"{��MZfO��w�݋<<�
��Q��Qо��uLO���c�Ѫ@�;���s�I���+2��ױ``!��(�/4�8�R .֦�x�$�����b���̜��P���Vl����i�j[*������EZ�55
�H���r��^�ٻ��载A�T�Y��Q�zE3�m����!�3��o"���2��2@C�@R�K?��B�� r�_�;�����H;;j�ܭOn�:�_���!�G::��\_�20�ii�Q����b����`z�ID��&��g�	^��\4�ZOC�wG&�$O�5 ����� ��$B��a���m"hl�r�jn��T�����?� p��ws�AyGG6�Jd8U�x�Q�|q����XQ1�1*Yl����s�.p[�����Z�8�`x�ocZ��J�f�f�}���h:65�e(�	}���Tͺ�N��=��e�R����bȚ�~�i����Qi��ʗ��
�����+�́%��d]óm@"����H���rw���Iq	�2Y+��K��
EYRF��{5~�^�+��{�s���j�x���;��"�bG�X\%���%g�Z���h�za;�>������+����F�
]2Ck��OשB�����d�၀шB�8�!0,��B}�]����.������ʇ�C[^��[�_��(���ߖ9�*�-EC��Q++�H��<'�WQ�*%����
t��(�?�:	�*:9�`u"s�\K"�kqQ�1��9���}�]��ZKׂ��d��ß�y�������먃o�_Zg*]P V�v�gz�u�<���w���yh���2a�G��<Y}���lt��Z�x�~��*�>̇A����:�{l�AJ���61��{l�?x{��$�Fz�U@����ʧ$��۬eͫ1���4,Nva׆ �v�5h;=&��tИY[�c�t��@݊���T��ɓ,J^k_\P&��Z��׬���q?�&���%���?�#%��	͝L֣Ňn����\wuo�5�E]U"���ż9��LIDe�>���~�)M2Whk��%@X� ye���;Z!��N(�2�\�����p�{#�%�0WUt�̌Q)�B�dk�X���[�Fme�H�����A:��?��J�q��� $Oͯa3��l��ͽ~N��������Vw�t�1�r~)�����b�N|��cc�Z..�:��4x�0��蹎�<��uV�aa�noϟ��QR�����ܼ�%� }TZZϵ	$:�P� �9	 D�R���0���v����~���knS;��b��]|�������1a�d7��Cc|��R4Ԃ����G��򱧨e�y%0��d���bç�m
�-��������&z7K c�4b���3�H*8ӡ��r����Q7�+W�FTW� S���q�/n�|2����,��������q� �yFF�ی�q�y�z���.�Жu��#�����/��<��V̝��<�>��)�@��0Q%�0%�{��i��w���I��aj�g؇��̢�f���v�:�ƴ��;'�Ko-��.��/e�#'3���TC�
�\���Z>���1*��c��9�?�
�Nf/N|�2��Z�x��tR$v�'��EM�.-�9��Ң\7��CŁ��b�!A"@��KM�������?y2���j��]f!���DD����X4��a�J%W&��G@�1r!N�2;
LU�.z��v��OX��2�j�+��jddb�Ax�[ª�|}W7�TX��Q��Jx���E��x@�a��7�[l�M@�k���1	-x���Qҏ�^A��g� ���[��4u	>9U�?��oX�o�x����Q9��4u^6����	\����9��PK�,s��8��B3�]��Һ�e��Y�0ց�TnS�"�ؔ������q|-���'�/J���6]�&@��[$�sf�	JЌ@F��]��� L������akg�R*4�5���	�#�Y ^ �D��tg��)q�"P�����u�q/��u`�yp�g�����`�+���ˏ`Dި_�L�����P��慙Y�c���%P�#5Q���Dًh������h���Λs~�_GA2R����p]�OrC͞��tdk������ݦ�\Dkjj�����1�VϞ5V�<y�����L��-M�LbjjS���h����cq�� H. !T5���ڄ5@	���|=��M��� eحS/KI���e|?����t��WG>Ua�z$Q��Lͫ����&�Zf� ���F*�S�J�ms�oǈ�k3FB=����U��0 ĺ�~�Wq����>G���d(�����>%x~�>�	�L�&Y�
�� Y�#5��0tJ�/���._B"�����QR�5��}��vu6��i�g�-���'4�"��dXnecCr(Z���#��6?�U�	�b���`����^��i�S�$��NQ�M<�BS{b���t���?.����,�٫"��\�7�p��	rl�5�I��_�H� u���{��T > gi�l\_�܀<V�� �i@�h@�h~��P�Λ�� 6/f�%�%��6�w��VD_#c�
8�NM�,h�s	bN�t�-Q==7� j��;]J�ƢY$�����T���,���u]�a�� d޹��nm;U�=1!�G�����0H�gte��Md�,)9).-=���b�rH:U�ݺ��_��>{EaEA:�f��glf&��X��ơn���^�!a������y4IGŻ��+]�/>a���[=���/ŏ�b!���B�ZOL�Q|%���*��CHJ0_�J�h�w�UQ�2E�XBF��9�ZN:o���h���ޅ�߿��HV�k�OM�y���}42k&�F��ٔ귃2P�DB �Ld��˄�In�J4@�ҦU�^625���P��<(+������6� �b-�<|}���s_7��IZ����,?��c���^P����^��TvX۔�/�o�o��_���>~�B�`rn��N��h�6���� �#�w�U�Q����' h.�U�5*:Xri�� ãY=��N	Y^�(��#R� Y�Ȉq}�*� WXH��,�� l���&
�a "f��`��� ��z��`3���o߾Ex�֕M ��������_��q%�yO<y��Բ�] 2@��j�����a++��s�Y����m@y9ڊ�
tD����sZ�a9uH(H��Ľ��OzEi�y�h�b�c�Z!��u�j��}&�Ӡ�uD��Ec*1�'�E�Y�"fXo��r��R��ffe9;����_
��EsF��0c0���k�W�Z�@F]P SSS
�"p��j�7PPL,�Q��$�@>�yKH$�I�u����7�t7����￢���X�B�$���>{�_ݣ��C"����P��Y�#��J�Tu*B��i� %�1n��=Rj�'�@��5![c���|.���E�V�Qˋv��5_U��Q�\�ʚ[�5���;� �a�r��!�8"�1"��CE�DGWyz{�*p >.�����14k�I��~�%���#�;��������mݸ���&�@���1�VUu�&�]D{o�B������}vv�m�)f�^�\܍�zg4��a�e�|���b��������ݥ�*9��s�Aa��!*��z�
�J����`7o*x���yW�-� �K�hBh(�m�{es �#�{�~�P#��:K(r�3�E�
QE��B�U
�0<J;�������3�=W�{p��]�����Fr���K**H����ﴶ122
���G�A����Xb��5ו�ݮ��5wZj��[[��P�;HIE���� 8OVO*��à�����q.2E��ꌅ|p��>�jS�Y��3dv�\�3y$�%/�p���-P�~Q[)�z��ǘ�& 5��ԯw�n4���7��.��2��\�D�ݯik�{f~g�A���M�AC�$����Y>{��qٽ��f��v��-�v)G��{�������M�G8[[S��g�O�24,SZzG�u>���b��7EԜ^`!�:..�5Ů���-d�R�Qb�u�4b*+t����a���@:(Q��A�1��)b�/{?����¸N뚒�m-6�\������a�	��Ɔ��g|>~bwx]�]J����K�NDq�u�\Hb�x��\jG�� ��X_X~��X�߮c�J��`#*����n��h�WJ����d+Ɋ�N:0
�x�b "%�졻���T�7C~/�)ll4�Ѕ��s�ܙ)rd�z���"0X��|��Q4�~1
@�wAӨxZ.��< ��� ?�Wq����+$s!�@��{��l.���U䢸�$�����d�a�H�I4�l ���U_I}���%a/%�d �������xibn��t��g���=�Z������l��[�Aosr��n/�nA�p���u{�y�����-�э�h���\��5��B����/�y����4�{��&��V�9>�$-�8	p�� X�Y�{C�z�.5!@!OBd�/P0$���:�������'���b�}A�l4���4���v�`H�{��9�7[� ��T�� 1Y��rfX�D��8�9�o� ������1�R�(+;zo�7մ#��'�d����Ҡ�y7����ܺե9DHS�d���b.���&?+�$�sJ�;�g�
����jj�hCZZ*���ڀB��H\  ��\��?�=����z��z��b2 c��k�'�]E�C����dH��� �ygY3�0œ�v���hp �ᢈ���e���g�.��+�CENy����e�LJ۠�*�|��ue������!�)��Z3�і�>أ/���8)�˂7߾�W����8\X-+�,8�
�����X`��/6�T�SҎ�x⌌�#']Q�X�.ba���?���0�ǻ�&��3O����
��)U��SJ��ӝܮ<w��ڢޱԑGB�(Y�h<T�<$̪�]��oc='���䩔��~��6�",����H�{)O?��=�'��+�ͬ�Vl���u&@̓�-.^H��xp�?��B0�Z2[���ʛؕ������c�8R7�A�]�I2�J.��
'�G�T�YԎ%���'�hs�q���32"�
���;�5?Y��"��Ġ�T�d����{|; ���]�L=(��7�/���7�L�t��i�NO��7(;z�Cf�y��s Aк���L�t"f6TA�����2�E*����i7T<ծBa7�:���hq��龶��ћW��؆�nˌ8�wD��߄O�;ՇyeT(	Kx������k����_�8��Do��M��������Wb��?����;�vS�R6M�(,�C.�kp'��?�.�ך5���[+���֣#aqf�9�z�M*\!'77�,���S�-&�K�C����d���OH�6���>��b^����zǦFq����C��_��R�s��f�A2��+T�d����| ��dfib�����l��D@�dr�,���]�Z��W�9Z5����Gr?m�t���P�A��{e�Nkr���Zh����o�H<*���_�Aߘ�l�*���A  X����|�'��u����}D;�Ho��j��]��<�r[<�@MKK�M�/W�>/� �3���_��6]����g��D4(�����A�(�J=i�a���^�?e���,�a���~MS8σd��������Ө7��'("PS�ޡ'�q_A��p�,w�����<���]V 	!i����A����5��X�4ܠ��o��%�РC��ڪK�>o��	jb�;����M�ȺQ&W�&�����m�K�擗�����bT$��q++�?���^~A_�D�����}A��2�Vv��U6L�!�9g�Z�|9YX��yR��z��ˇ�::b�d�_.���iॿ��p�<�H���{�w��S@�:���.+�v;M,�~�\Nظ�0�s$��!��UN���&��u}�E�=�8HRM�U��B4�!w �uFrR2����o�G e_X��=!��6�V��Z��{�H)+��rzZ�իi��?�Ԉ����q%\�%�]$edځL� �[B�A����p�d��������r�{�Nf���e�.I��hL����G�I(��j���>���1�MBA�_̄����F�T]���bE1Ȥ�q��>gı�ˈ�7\+ڨO���@��[R�_�z�r<�w�sUmN���Ag��|^�:- ���d��B7�>O�?UI��X9��;�Ź�t������
:1y�[Vf�=�/��q�n�r,ad�+�����Z�������$�m���D{���Y�˷�_C[�|6.|� �d��޼�K�	�&n[cK����3.(�
h?`9�t.P��*Ε<�,��x�`ÿ|��,�^y��P5�GN���s�Ms�����A�7ڡ�OZի�p/e���)�a2c>��3V���j\�:q!H�:E�埰V8-�� � ��z���'��d��E]uu�}��Z�~��h:t�Y��Xbjj�Q��e�33w٩}�y��b[�˿��<}z�P�,+ͩ�]%�C�k�76����zl�V��:��� �����ꇦ��Ŧ߶�=8����j�A��Ukv��
ex�)�<���]��n,U���
i�@V�Fӆ�sv%c�{���,E�|H�x6��)�l����( ��!�#�ҟ���D��n��>�<a�v���7�Q����w���2�;h#=�[�?�-��h�*�K�������T�7���\�Z}}}�L���6����1�6�KGǫy�%G^�/ww�A�C��[�gϨ�,K���쏏�x��!Si�[�q���E��oH3����X
Fh��j�A�k��є��~{Mc,�<�<AE�|ԟT���/7�l�'��i�d6���n�]�Do5M��L���?�ȉQ�y���wx�|d�}�Hd�\�]�� �ey����*��y^Z��4��b��]�%�e��Q)����aL���{�SY?�5�B2+9���w���}�إ2u��Ʊ��V�=�����z��Ւ_��6m��.m�sq������l@楥� U�Y*�WW�/. ��W)�5p�鱥�mBV�۝���d�F����.3T�׽�IE�(������7��|��D"GE�.����xɫ�Wc�ZO�Y��%@;H��̀����R;Q������Ap�
�&&7@u>8��`e�G���쨏4��pZx��Z��e������P R-�ˏa=��RL��kC�`�Gp��b��R|������̏3��-+�(f��VV�=��11�V;�
mڥ�NA7�B���8(1`�@�-7���jRl~�F�&_�R����R`'�O��vE��	�AL�E5����� � �F\��(M��q��7A���f�`��DL?a���]���r���Ce��ޅ����؞��饋��,��g�8�_ �_�я:-�����[�>�4�ǀ�%<{aw����e���Mc�2 � �t�����_�ܹ���zw?�;�;���T�k�QiDx��+޿ק����ո�|��L쐀W���-��b�����gg2�_��
��u!U�z�7���hv�~��q�O����+�~V=Qs*+.�:R�R��t�������CP�+�/埇�;��g]c�+�l3�-��6�w,�Ot�.�$P�77J�Mp��YT`Ra���!SԾn�졁��0�t�\��g��\�Lߵ�*���g�hb�l���x��j�!������ޞoU0?7�2NS]y-َ�oc:����d��������gR,��9�-lm����_�n��w�1p���	1��Y47Z��sjj��P3�֨���VKojf���_��1��[ʠ�a#���,�J�!�Z�X�꣊!���"��Gʈ��S��e�7����*���KM�����b�kh�����i�/3%eJ���>��ۀ���{Ǖ�шh7��� ��M��8�L�Ԕu��<'j���}���L�G��D���ٶ����/��?��O>��W^]_�=U�R�]պ �v&.����W��������bm��=� H	�i)�s�0"���~�=��^�2vqu�HU�ՁFuZ���{�i>��_^�p�a������-�5�T%*��5_$�|��[��px��[gj��k�`���!*3޼�H����2��тJPE �3޾�9J�r��˂��0/(�<%�ϛC�
p~���^6���:�\�L�eM9l�n��H����>A{+7����QT��F��l\�����h�h kfN�*���^��?''E����y"
����Lk�V��~	9-�4:�3�B$�h� ��Iz3C�;q`���
@��}�l���C��b`)�'Εչ^=���2y�.��v@�7�B���*%���D"�k����EN��n���^h <y�U�X�Q�ܢ�Dux�44T�N�6�,�Kf�eB�pA ���yՆ?9���p�0F�"�pf�;�
:w��\����UX�,Z��2��x�d���|] ���?;y��{?@hC�)⿺$�%���C��ޮ��O
Q9ߓ��͔���Q~��dw�-!)a���:h )촮�X�	=>�� B�Y_��]78c�O����Ԥ�Lv�"~��͸ny�#�\�ɔ_�is��oQ��^R�%�+���/����GT��/� �ɇ��P%g}!7��A�`�V�K��N�P*^��O�i)/CL�-$�FM�ݹ5<8�Ü���n@U,AJVS[{��-��J���
�D�9�}�v�vǁ0�Q�H��5)��\_'� p�\J0��=Ϭ)q(��
�{�@�$@ہ�8)���d�	�����9P8%e�F�59��w�G!�����������v�|ȇ9C���� w�FS!R��1
������tt�*�����옟o~��Xˇ�Hˊ�n3)���)v���d���vw4	wv�Ǭe�K���z�162̿���ՙw�q�P(h���̮.�������@v��k��cuc)�^���<9�~L�o �(�P�'����؋R��X0[��5A���\�����2Kо�L٨����6O�5W�%r��Q��w�A�e<�rswV��ꋲ|����b` ���y�t��i��G2��R2����\��E��<�:���1�>�L�j�x>�x���s��sCFN� �}�q��G@6�5�����	{�u熄�S�v����VW�X�m�{2 �`mk�T2k�f�F�+��"B}ȁx{��UÃ�Cd��� dq�Z��/q��:�q�A�S���t�޸B Τ��s"�29�:!-d�
,}�u�7Ksuo��̙f�����0��S#/������'��H���
���xi��	d�z��X[�0t���<���12�����1D����M(��6p �Qm
������&S��e��a�yXN`����s��&AJ����L���Vf��W#�cВ���|i)hkt������Nn˟�o�G~N/d���9=O���Z��^�\ĘY�W��t�r ^��W�A��/:9�:���\P�}�D���m@�Y$o ␉��7s�c��� d	j�&U�O������,�Y�C>�]� �?��RSS��=qIX�犘��5᳏��g�C����ie,0/S��-�w�0�F�EC���О�o��o�UO�&�;)t�6���.�΢,.�sm�73�O�ې��'#��M��1��sUv�gb���@��;�����zpy7���ȫ��6h�1;!zPR鴂�΄dBH�����&���	-��K�V��_J[�Q�d�E�o���(��-�5A-�->�5!kO{�Z���/4���/t��d�ok�,h?��������Vܿ�p��J�^�zk�E��[[��������>D.
�fFF��!/��*Y��ch�Z���GI@���|3a��ܜS�il����>��g������&���hY��>)������34N;�U)�:�V��v[>�ܾ�HK߀�iS�7�-{X�iH����\�@�8K��ѡ��7)��Ҁ	�}7AN]���b������V�F�K���Ž{�z:-�����X[_�1���kfF�PwEK��/��U�8[��OQP >ǚEq��H�ԅ�9��I���X
}���D��d>" �1J�m�0��@���;������uR2�6���Ҕ}[�йq�g��29td�@�����9D��nSn���1�<�Y;%�(�n�	�b��;�q����̜N�g�eN���!`X�R����ѳ2����ii/��V��5�C��y�՛_)���H|�v�ʠ(��f�*�ץ]�E��w�h�0	�<$2U,h[��Y�=���,+�=zKԕ|�V|�妩��=��ɵ=��n��+*�*4�9�̄��o�Ǎ�ߑ�&���i�+��v�}�]��Ɔ睕���nϥ~�OO�����3̄�Q�\}w<����$Tv������QfF���{d&3�C:!������qp̬����~�����qz���z]�s��uߗA*Î_S�2�͝V)��s :G���	Co; ��x���ڸ�� �ǫ�w��y�H'�N�-E�с�#�-�*K�z�=�sʞ���s��N����"X��MOs��U��%YA�
����-��?�9�@׏b섳�:��!��Y�h��{��.V)U���>��T��˭����B�J�	�^���E�_�V�e|�W��=�����G; ��'-䵯�r����.!�3k�r��������Y�vt̼��R��y������/��,vq�{�sT�_CDY�a���è���HVF�����DD� e&`(Pd4$���n``�^W�����Xoq)�*���,+G��wO�D 
Ϝ�FZ+20 ��|h�CS{�G��%��?��|��P�H`��v07�����e�`��y�q�z���<* x|-j'����<��aWWW`�0�78s\*G]%�\�3]%ze~�T�ԉ�f��5��WG�W�z4�.�w7cZA�����c<�Mp��b���9��U(��N�b���������,���/2����?���"�l,�O �L��C ��(��T5&�z��$01����$��Lֹ�(��z:���>�����O��+&;^���'t�d�hbPӗ�6G
�d����H�E���N~�%�<���K����ڳF�s������݅_�A� �E�3�c٢�ed�����[ncS .�ۡH�`�F��D�yD��,X���@�����Ig��=�@�d��߆,�ѯ
4l��6�0v�G��:�ׯ%�uӳ�Z��ǿ�ml�����=��4+���4Ӡ_�r.�{ֹ.�r,��Q�Mi���D���8�VO`�������d)��JM�;��ݯ�W����h|��<3��o�Wֽ���a� �1E�ܼN9\N��0=6�(�����WE/4��]/�]	���f��Oc����p*�.Kʚ�Z��;J)f�>5�jl5|��s��p�mb�sJ@�s��yO(��/�qwR~"O��ʵ��t���I0[�����N�M��B�EDkɩp����j��;lji�
j��z��eceDZ�ԭ�Z6�$�t�{�\�Mu�Wl�^�{x���p#�cq��JI'�������A�2�<Ԣ�$��nݐ>ZIʘ���]n���k�*���ª+��S��CC�f���M���߽k������������#�1`��w�F|-9d)��k�kR��~ڻ�]Ž,w����F�S��C��q������Q�S5��� �k�'�e��hnȾ�a�"��E���'�o�k�����=�sR�a�Z�ǥ���b�g  ���mY��͡� ]��s����p=�O��+��C##�h�FJ4�N�s�K��'���:�4�u�me�DV�7�Ȕ�0�C����@	�������֒�Q5O!ͭ�?,K�n�9e:(�jE)��D�nLq�g�J���q�m��|�|�/����S���/�#a��;W1<:j9;�hE5}>s�>u��oJ��Hx�M�%	��Y
�]_�VY��ATy��8d�]���ZT���sV*���c����\��(�y��y�!x5�;��<�_�+&0HeW��y\vF[
�'^�&Y���ϫgߌ�O�'�Ϗ�U������Ĵ��F
]�W3�Ǥut�b��)_�'@�U��:�4퀽����Z�D�$9t�HʣK@����5�rNE����-7��.jj�VnF?W��2^�����Y��2�v���c�r��e���~:�\�6.��NA���|��٘;��c\�Z�z��AHh��7r���tj�Y�s�.��:�/��#�n���Z�� ���V����=&2_)P��뷉�!��C¤ �b������}'�Jy~�����*?�VTN:n�>���C��8~�%C�)����(oK,�������G
;�F�����%%J�����D���R z���R������-5E@�;H�+FHD���GG�a*-}6����a�`����P3Ƕ����UT�Dw��_�φ�$��x�p��,��x�Ĕ���vg��;/>��`۠��>��Q��\ZUh���w=;�غP��Cj)����w�����i�_��/��!��b�̒\u*�w,ohh��G��am�<3Z��̌u�<>���W(�jf���%*�!z���������+�^�O�&e����O����h���}R�k��QB���+ޒ+ޝ�������GHG�e��c�m/Q�� �^��ݽ(��%�g�ߙ��K��F��t��i����J�Zb��ƀ�^����j 9s�DJ'S���[�Ul�����;Z�ij@��rБ��7�
��������yyfQ�� d.)����s�����ܰ��u('�����9�r� ��D�=M��wW�ր�C���N���@P����`�������e	��C@&-���F���"���^TD�e�)�_g�'�F�9�ח�|����؃W��i�P������#���]^''d�̢�Z�^����]ԟ�an�OPR�� Ds�������ŏ�O
�O}�1P��j��E�;8\[���^{��iG$\C��/5a<�-˻�J��\ިQE1�{�1�����FC�� �fB��?�Rm��~��U��_�wׂ4<�,-8�Qt2KP[�ݻ���Ǜ�y-��j֮�7D��B�Ot��į��D#jk�Uy���E$'�=T����\�zqZ\����j/+Z?A��<k�n�p�9kr��8��ߝ@�Jw���R�ՌM{JL{�M��O���v����J'����is�\��������ݪ�rrbl)T�����;��=�<�ۨ�q�).k| ~����(!��E��=�����Ef�뛘���/7h��}A"��եb���j��'X�(D�:~-2��o��[v����"q�ؙ)�r��I.#��{}}���O��3^���B�~ �KV�&���V�y�0�upw�F � ��+�N�����]^����7#�`JE5�� ��W�KV��\l"^�Aj���r�ו2���b���z�� `�̤M/r���pE�4�j�U/����>a]���6[f:;��ͤ����KM��o���hxX��������2����9Y�;:����T���=;t{��S�����:��9�ǥ������G��\�] ���I~֭hJ�H)s؃ؙn�ݨD�}P�{�)c��ta������l�ݳ���;��{�AK��Nv�41͘��ഇ�<�>�C̈́�%��Tڝ��]<Ƿ9�6���SL�Mm��e<�z������f%�h���A�^�^pչ�~��$�����aj%�V� h�8�v^����խ����Р����|�.�8��d='~ [)�a
d&�7ʇ�f67M:%� ��XT�}q<m�?�	r���j�w��Ϗp����Oaj*��e��D�}�e����?����|q�~�	oڕҥ�5�_��; ҳ������,#��A{Hsf'����\#� p�L�߇�S�}^��]���{�S�9�,L����#�HX<)?$;�QJl�K���fJ�(�|��x@�,�.��_���뿥&����o�8I[�$�2�5�,��E"���48���t�����!�k�������N�X5�^=�K�b֑���V�G��_��g��yeO��Hr�:ryO�m��6���Y��j��;��|����g���+W���Fi��v�&�����E풒N�!���\k��gb��&�7�ꂃ/dkڎr�OO7.��$��╦rrp�5G %��O�*Zo�d���=�A�s�@�F{Z�}�T���㈏RR��Ώ��jν;_�R	#��t�����%�/����)�d~��fNN��n����>16��M�<; %f..DYd���=�E�����&�#��K��H+'���{C� Z|4�AA5.�S��O��+y�P���Ž{�)\�f�A�d����U���	4n��BJ��Lx���EeX�7�~PAԊ!�5�}���	(+P!�J���R��f/�fD<)$q���]5,����6'k�����л������G7ڞ���x�]	��XB/��3xI�?��V�O}�=��I�W-¶��ϟ-K�q�aI�e؟W,uu�c��g��ޑè�:�oN�Ţ��d?W�po��''u����ޙ��B���!�s���%h��4NL��%Le�w��� �X
|DP�R�6���+�K����g�o��V���$������s���8��m0)+9C���
3|�:@OX��Q�J�	�y9���ޅ�I�l_J�NB�kb�FAƦ���v�܀��~q���,Fߧg6	��b#F�u�B��BW���wg*{�#��H�(��x�9�!q�dnD��|h�݀��e�mtTDuÉ姽��.�������$���tJ���`����uꚩ�Օ�EZ� �O/��4Nt~3y:��K�e�0�	��̐3,���Y]'������S��L��D���Ү���'�
���YY���i��N�ȿ|�Ni�_�",)�8O�]\Kt[���G �:~��{�<�B�9�(�*W����@��Z�)}����Y�|�gKo H%'��Po�Vґ�J�$j�{Jdm�(è�L�˦�T�><a�9닅U��Q�EF����޽[�����m_Mc���S;�qеpܿ{��w�� F7��Q^�Zw�j�I�ϟ��&s��P�k}O{����`�rT�=y��J��'��`�X"PDiC��FEE�}^��[(ޜ�M�	�$�ɺ\��>��A�Fh3�\�����u�ե��.*����3�/UL�[F���T/�� �U씁Wj�bWW�So�.|�7�Y��x�E\Q���1DǞ�U����ɑ���D�Y�$yt�q��r�)t.Te�Rﳿ>�6)�	�y��2��\����V�.zջ�!¹��_C����G��N�u�zc<�ؚ�:B*#~1�D���u�4��ܛ޸���,y&t�v����H ��Ԋ��Fj��UK��M8/��m��z��P�r�f⇶ ���ڳ	���>V����^�z���Pm�U3[��0�����f�7�û�1�(�jNr��G\�fC�͎ �z	C�?�����dZ~������=3#o�am���vu���� A��ϟ��ǜ���l�9�3���751Qc���h�}Ë������.	f��^�WK�X*�r�Slp2Ĳ��4�җv�k��4.|�U�w0���R�	m�s��E����2M�7�<�^��e�xZ��YW��O���������	�	�Z��:7/��M��R@:���ȫ���0/��s�*� ����\�(W�= ��k3��t-�wW�FD�% v6����M#�\;~)�/MHٜ˂[7�Br ��I�G��bݩ���Γ���X44s�wה�|w�q0]��]h����\Z����:`�7�g��Q�y�<a��:�WVW7;`����5�Y]ݸw��1�?�<�\c�T�i��K[������P�RE嵐�}|�V���F�J�`*đ����XRSSe����B��q�=Gy���߻׌J���"$�^�%c��gT�k�Ɯޢ��S�YY9�db�eS��JTy]W/��
�����ꪗ3ˇ��~GQM>�+�g&������!��	�1�/Qy�B���h��'47�xRl)�NMo��5��U#�m,�� O[׏��_��M*�P�S� ���b�f��'������hs�3�Z"_�[H�H�M{z��JD��e��D����K�0����fA1!Q��4?/J�(X"y��"W�כ����8����w��t��s�WK�Ͷ��p���^ꋫv!t�� J����H̀|���g�3��&O��ʪ^�}e��8謋�(��J��w��2������ �m�[��k4������$�~�@m�Eb��:;�^~�M_��m��]���畒j1 �E/�a"���5�����c{�tLB��#9S�A�����MDX��JKd�θm;H��Ꚍ� ��o���BL��\��ۯ���ѵ
=��х��!'�UJ�n�M��%f��#pK�b	3�źF���$�4��EF����j����L7#��_�+��Y��Y��2C�^�23�zU 	��HB�t*jx|\N��������ȋh�Hmz��lQ���d� 01[e�SS[�u�O�ҩh�S��[X��ݞ�6�7Vw�9XA@�5y��������1@&�����,��S�+���1d��S_��W�#1�\�0�� _��#E:Br���Ն���W�Q[�h�P�\sy�C}������d$��2Ԥ�z%z����5%7���
 ^tRUR�����Գ���J�g�J��G��1��
���ۻ[�O�;N��������MM���KM}������V;~�Ș#�nm�2����	��qBE4��c��=��3��bFڅ����,�g��v�2Y[[�"+��W�.w��_r�S��J	3��Y�H�?0V[9QkD�>�l�ܤ�_�����kp8CF-.��YW�����ux����"�T�Wr e�W*�}z4���3�=-�z���0���-�gj�&�aT*:���*^`�;�g��E~�E�1�J�:�$���s������"��A���p��KW�r�ХP�?�,_n0ps��'�F�-�1u�G{N�-U�d��}Y��2����"�춸.4�����,d�+
/��/2�H���-z#�����������4s����4��d�/.u< ՚�9�-ѫd�>��j%�Wv��Jr?]�8D��2��+
׺g7͂N����d�m`j���܄
������@�����á�1�d�`ɉ����Kk|����ϝ�ɀ� @9����9
����f����j��2���_�T��ԍoFΨ�^�<41��%[�M����e��8E�t~�p�H�Đ'1�2c����(���	^����ش
�(��Y'm����@�,�W����$�/6���:��KY�e{!��#f6N�sX���ު��us�4������/l��T���@w�1R�;Ȏ��CI����k�8*+zc�I���Ӵ�U�/��(�a�L�K��b�nii�x�L���q�I��f����_�:�j���W�}M��,�K�u���� 7<�~Kk����Y޽{WS�4K=��S�bvM�?���eS"��π[�	�Nr;��#z]�}y�k�u{����k�Y�,���VF|Q�&5wف*P*���0�Y�#�QGu(�(p,p��ͥ:�$��Q�u�C������sl)@w�T��S���U�1A\W:K+svυ����iW3TŽ? \�q�����g��L��ל;��j��E@�[f�Е�]s��
�@ƕW�W��E��{{{�Tz��ַ�����Ls( #Y>�P�\��Y.f��;xH\ZZI!_92�,�����j����Ο1%So���8̒� ]�I9h:K% �djo  y�*���qH�����̄�?�W��L�������S�M���E��x�����a�[<Xu������,����/�lF�䙡���F�pz��*޷�ٷdԸ�HL���k���� ����#}�)R����|���tu�wP��ѕ���⧾g�8�v
z�Ƞ�%H�ߤ4��Z880���{ׇ��[nVY�o ���J��8^�2�444�^�VX��޺k@ I��6U�� �_{���0)�n��
3x�R�,N�)�}F�Hr�TI���Dھ�W(]�b�XϚ�p��S�Ì|v�נ�Y��� #0�zH�T�H�P�eXɁ^P� 4
{�OPr��T��a�zc@�Vx��P�k���Y#��seďZp��w��#1ji{�S�=�AޓrAz���]�ior������`*�$��w��|Ũ�s*ڸ�~ꏗ��f`U�P���j2����g��kD��@*�8�Rș����H�Iw:YY]y�W�d隴EeAL����AH���.�{4���Y�o��RӞ���>Ɇ��5�{��$�X+e�ue�<Jo��w�w�UDop	����_��n�L��VN�p0�0x�`"/
o�7,ႩD��6�Z��$Mm�&*���:�����7�� G��n��t����l��pBҊ!�������0N�bڪ�1J�BI�o�l�R��{�gǾ��I?>��_��l�w��]]���f]]`G�N�n�}#�Z�8E�23�<�Ia9<�Eˇ�i��U���U"��ݎ�\Z�l� ���QB���z�������X ��
��`ޓ����S<Q11v�����99L!-�R���cb����z�^1���E�s��������=�U�l�\��ϟ�����(���t���r�y��3��~(�phg͜��A�O:�Q
9��]T%��
O���mr�Q�E}��E�m��":�4��B0U�:#@��_�Y�yOB�/��i�^
��� ���u��
�#n{�������/�P$�%QWW���,x������YρϚ��ο�#:[#�W~zpB�2{�C������go/|�6&��m�w/�X�Ei����b{4_�S׹�qlL����-5����cY \0�O_ }��zqQ�TT�w*.v ���.7�vhN������89�K%B��qr%��m?�����0C��8Ӹ�X���F��g=���������) �[���	�$2�j�&(���%!
�b��}	ޏ���~? S���0����B���'c��Ն���\�9��l�Ed�M��B��4��Q��V��9��B��.�Doy~�
8=�M��\ڳ��a��$D��x�W}�������45>'�#�kU���j�I��V J�"oQ7���𦚓ఔ���Q	&��dM�w��Ltʟ��4M�̌<����Lq$^6t�ތ66��3�c���j�
��u���¢w�&�բ��]�v��,@������Xh��-�]��O�c�K�(��&OB�ë ���@�E�j��R��כ�ƺyO��h"sx҆����^�\={Y�T-��5�T�$	�_��wY;�t��o>L�-�9�+O����.gȁ��v�=/*'�<��겊?:�z�uP�&��v�6�4mv�vb�t Pϖ���i�����ʥu͂��1��|�_��I�6ϊu�kjP�L1�����m--3}��	hJ��3�%�s �w�û��kLSAp=	aׂ(�&~��S@��=�����j&�2�.�4��P`00((E�U�Ȳ@KFv l~,�]��,u�n�IP���/̵�f�z6�� �:K+A��)���,���S�C}):g���;�{ar�ߌ�����wU�q���⠒ccjܡ�sB��
�cw2����a����m�d�g����wt�b���1O������y�=~�X���.�E�z:��0A�iW�t���X�UGA��Oxq�u����s�����5��#�@$991���.��R��&Vђ� ɡh�w�#�J	������X����(c����@#j�q���[�:�k5ת�W[k *�."���i���(�2Lb`��1v9�Q{D��=�J��W7}��h[����4���)Æ��Y�$%{@W	���/ kUV�����\;�8�sz�$H�S�M���)a�� n9ӳ�?c��,���a��4�ǭ�/ƤN}��)Y޺����'�f7X��r�ۣ��mIIg���]?�^����ҿ���dT�IY�M���Ʌ��n�C�ǲ����z�&\���C'�������	�"�Ȥl�ϟ�qq�!���甾/@�R�Q�mQ�eW��b��nTc뼆[��_��y�o�`�{-ӫ�s^/��)�X�A�æ��������r�έ˓�c��o�Js���HZV��]����P�X"��� �\q�U:A�3亂��8�����u`I�c�%�T��þU/ɚ]�F���1��ͻ�2��M�{�o�OFWi�N�M���c���rp0�8�@}g��� Â��UJ��R��^�����G�<J��Jɡ�K�rN��Vt�������]��[��JF;-��B�f�KK��UI'������^�Lgw������#:�-�A���4���p���E��#�=y�qs#�V�jƦw��{�p��Q �]��t󼜸uje���|qz���%i��NM�oh9]^+X�M�91��H�J�d4�n����Fδ�J��
5�j�d��K�?�	Ϸ�I{�w����8ch4��!N�F�f���m%#�&�h���%�.t0�.�_^fL�%G��/G{gBA�	�ĉ��G#PE�V���e�/55����F.іBỻ���$�|./i	�ј�;���˳EٵU`RD͓vR�q����	ҹ��('�"���;�	%P�|�g鉰��V��+���+���.� �+5Ռ3��7�{2������?}�/q&��]s�R�!��o�*è�@��@7���p����]�`.}�!�|m�M����7#D����B�C�4W�+ot��,VT	҃��K�����vκ}.qN��KJx1`7�,k�;�ag]1W�5@:~o���o�˝!�#�ց���@'m�:������%P���]c	�+Pk�T����MMh�j�d��;wLE蓭�+,R�/{��\�{i��{�6�{�%�"V782X@Ƶ?����Y��p�H�pNp�5�*���Һ�;�P�*V�9�=���'��z�+���\�{P���FQ��4�W���J��f�8�\���*[�jÍ���RiC�Ld�Y��1��ɔ�'A�h[�q��hԜ\v�؉�J���d|���vSQ����0x����l/I�J�'�� �7���BC˚1�X�=�Ajym-���F|��E�	(k�A�����F��zpdr���R�L�?������S0�q��(��͂t�R� 	�w��v��6*�ͬߦ��c'��RȎ:��˱;mh��
�*�DF��C�̓�^����"[5�+Lp۵t�=�����beu{�j����o�r)��@\�D����T��[�,��>	(~�{�2?2�$hR왨/]H�Iy��O�����V@
cؙ��������yD�G�,N��
�A�u��)@H�n�R�M�35���kE9_RI�R^n�b{kuL�'�h^+tu�+C�0貚�565̗���-R<@߃N~D���6v��Y��A}����u�N��hZ�L�3̋�( A�54�|��;���x����r~�QVY�]5���h-[��IǴ+�� ����'Ag�0Nbt$	(+h�f������-��:���?�	1?H���:��I�Fs%�։�޽�9���y�5�B�<�0���o�l�ۜY�c�1�_������C`�;	v_�d��	�b���:L����N<~fd���h^+��K>~~���1������d��}GU������<�
�0T�А�,���ɑO���a9����5�<�-��39F
i�?�Mf��C\J�D��'���/��7h�/���"NuǄ)��M�gĔ����}��	���MӮM��;��d��II"��K�P�4���'#~"�TJ��Cz�`���]�ڎt�q�tU�,b�>/�jÞ|O��&eD� A���J��c�J��9����1Hd�f�D�vG9�9��@B�F����ꢥ�g�m�/e�bT�ΌD4��|(;?/"}�7'�K�*�>'�O�
��ݭ
ޮY���U�5�]]_�G��u��
���:�hRV.�ǡ����O�I'�IF%�� KJV�*����I��=aq�� �JCC����
�>�vzۿ{�b�$.���ϯ��/x�@n�!z9��"'ϼ��:�|���)����բ_���)�a�aT���:gAm+ek��/��>j-��}�͆L�����Z�EP4h�I*�<3�t�2�7�)�K��?|����)���,4,5r�I�lÒ��.��J'�d��k�/d����A>�ABJ&�(��u���oJ4t>��r�S��-�ۺp`�

��l��Et�\�mcly��OO�+��--��?k`xηI/2>A�*s!�?W����,pd�w ��%��ea;����`��@�_	�����R�z��v0�'�2�g��7 �9@�����}��\t�aI����=4�w�L�Z�)tۭU=%lk$�:giR�r�t����Q��^���� ��~M�?N�J@TM�=P����N���)9�`�2�J�/�E��|_��*�HU��*ް�H����ߜu�=��W���}��K�AH�D�ɓ��O��{��"n�Ѕ6N/f�G��ԍ�\�_AۯC̬2@(��S+
������!㳲
 g�~��ʀ�;A����M���w<�֠y� ����$ؽ͙vJh�ʯ����zƑ���mYIO}��E߆��ҟ>⺊f6�=�B=w��O���Ks�7K�PՆ�'����\�j���lEt�Q\����eۚg���L��K���i-t�u89��o^'gKC���'��QhR��L]>�VI��Q#��s��*����Y���p���]ÊlYod���q2�oQ�=e8�ol�i�������]"kxt�fI7��nm��lF������D�ڴ�F���mKSi�}���rZ�,+�{�� 6���]jm]]���Z�{�Ғ�н���������E1���=����������̓���&����>�8nLQV5��4⿊�ȿ����ڻ��	_������'0��fQF�(l�e�=4`j;�|�2 _�L��\u��V��7�`��?ۙ_5,#���GK��i`>����nK�!S}�
���~��3f�Uuu
�-jjjb�g@Kr�L���N���?t�o��F$��A۞��u̹�����&��X�3�QMe�75=���3ڜ�E����=7�Y4��=<���Ws�򂐑��{��)"{����^:�ׁ���.�K"r��1��O�
�\�U���\F�S�eXU���Ǵ�����sRV����X�ձO�ֈ����I7ޔ+I����D�^��5ⷱ:l4,���q�b˯��-������ӛ��v��f=%ж�}˻�%�r�6�.�2_&�-�JZ4������Y(�%v�4� �5�)ʰs����* ���v d��!���H���_�u򵡎����芵��5�k@@��uk�I����@�O�����a����B/@�0��f�q.r?v���y�L��Ռw��L0��?{�����5DTV�r�'Zb`g����&�uW���Y҆��/����Ra�Ѷ��9tx�� Y�p0��hlP�}0,}�&���}:D��+`�̼H� p��l41𡃀  (�O��8�u�(Zߨ(*J*]>���u�؝k;��Z����jP'���u7��殪ި��>���Q�1���QA�9�ތd�Oہ��[�y�i8�%��g�ԯ�*�˟��*�b�~õ�~v���O��#a���%�~7��^Myt�)���	��h��Z��
�h��rt@�&��<iUO�����K���f�\A��us6���e�r�)����0hG�R��EY�}���
��)�[=n�9�Pr��ۮL=�-�QKS�P/U����������}|Y2�z�4��5�\����jG���S.��э� o�:��ù;}�ޝ �:<$�R���3fWɭ���~�tlmQ�m����{M�]{{$	|�w%���7< �~|��"����薋n��1�7����� EL�h��}utn.�@@:��O���G]]s	V���O�� ;��=w�6��XwO�X��@���3U�=�o0?&��A�r��x@�v[�o�p3�f��bgE&U��$(�TE�"@�E�Ղ�Ńm?~�Sc�x �5_-��HlN"�Ư���tLQB�R��)J2�gv��L���y~����nD��Z�����;q���Div�9Jd)I:ksf+p����131���	Sɳ��Ŭ�9����6��R�����)O2��B#~���{�݊G�k��Y�6��!M-�=�,��/*��n�7�Q��J�t6z⵭p���c�=��ҏι8Gռ�i8T?��J	�ȰVφTpM�>��!�
�<[L�!��>)|�t>�
	��fR�پU�ioU��@��ظ�:Z�b�@�ʦ�����B�,L�K@�RC��H_� F�F`߼�腓�oK�2f�yB�Ԏj��/�w�SJɿ ����9<WD�j��"�镕�|�7fa��^(k�V�/��$%z�|K�	 �DEEo���tY
:��%#�Y߳��"%g�k�s@��=��OO_��K��Hr�"p̀���L�]6)s�d7*���D.��n��&����DD�eZ@G��3V�mK��<˖���~�Y_��C<��P�˺2sXF�i`n_�n/�E��5�~���̤���zh�D�b��������#�2ktڭK�9�Op�+4��^�
���r�B���u����o�ju���a�Bi`e����C�����,�U�=pl��]��b����8�<:��.(%��kk���3ZP��d�Ak��
�Ά����X5KY�������S���;9�C���%^�+6�F��P[�̓�X��� ���j:�׻-�$* ���'�(��e��� r�����B���Լi����Tl��Z(�viD�Mz�\���,ʉP����vtX.�'����Ϡ�����4�r��н� ��w��xJ�E�?;_��č-@{�{���=]Yo�!"�Y�yw���}�o,���1��1��� m3Y�ux��}֡F��u��7q&�����1�FcU���y�kk_�ݾM�u�1q�87����«Ԋ�L,��O���x�2�E�O��PA��EYA��6�6!�r��2��|7��K8iѕdN ε~b�/0uW��ڦ/~ʣ�n����a�I��\�����8�L��f�^��Ȳ���tx��6���1����,��6$ض���D͝.fԀ'!W�/0�xS���bY�[<
$8�a�����سT����fM1�E�2l�������
;K0���B\#���B�`��끈|����
G�{��+B�����O.;��X޼�-sTV�u]�eyt��κRh�ӕ�') �P���r�"T����DD�]�}^�*��l3.�k��Aj�fxH���5�2��J�>�d��=�G�!r�g=̗��E^��~�	�Έ0O�0�ZU��]�M����؊¿���k��\��I.��8Ĥ,�W��pa��EOB!�&�������0kP5~Q�iJ���w� �7�C�����G� ?s���Ɵno��;&L��ǎPo�w 6ؠ���(��G�
;�˩DKh����3~5�zxx�zU��N�M�]~�%���~�*W[�m�JRx܎���F�u��)�k�h��@~�u�qp<f��z�[S�8:y��
 �D/����AZ�/ȺD�
�T+��0�T����9+�V���fP�N���!(�+N�޿��wA�+�b��%Y�Zot4������uN
bC�k9Д��v��[N�q������mTuAٔ�s�����tz#<F	����V�<ޡ�!5F�0���ɹ�vA��o�E/�̂�ɳȸGԢ���˳B�� ��~h)��#%�b������F2"Y�
�1�_��_��w����Sʱ�{�����U	C/�>��^Z��F��e�B�{n=��0h��=<9��ZŃ}KU��|Hr_���P�S�Ǳ� <4w���(��i�>�.��V���1H�4Tx�t`��VX@R�je�;H�t�F��J@���ɓ�Jd}�./�P�3�eRȃD�>ϧfݓ;^�g�8I/s�e#U|	���j��}cbbRi�a�<���)jA�#�OO��^k6��al��璒�}K��SU�V�b���g���7VF�Rari[�R�Ƿ7���lI�>�Ft��J�C��/&�G��׾�<d�;���vb��;����E#�9h[@��Xb�A��3�./I���� T#�����.��'M�@ٚ����#�Ts��ۦ���s�`�K���y>�$P���F�Ӛ�7\�:ʜ�@疞6iH�_�W{�)�L�e��^��j���X憢�s�"�V�X<d[���GlTSӞR���w�� .�%���e@�_k�J��\]���M��J�,��ʱo3�,���H)�?�[|�P��&&!����s5y@f�$�#��U��T�S�X�$�3�䣨���?�}  �EL�N��\�����������9�KA�ޭʲ��
�A��|K�<�v&�t�u rY�j�� Do]Y����ir��(|�_u�I}?�ѭ�CF>pN�]avě���	'.���7���/uJr���TY�L�xf	�db����z�2l�����O:���L�4*5P�Pkg��6oEE]�����X�2+B3+�Q?؜L쬷����S�$44��p �O��	^�@#���ϼs8 Z����&�ս�||J�S[{�[m=�$W�]���5�㣩����@���H���1nZ��H��HyP:��E����jH�	��1'a�c2�K������ t�k�P�\U��U��6�:��#����z�^v�3#fSD2P��7�.�P�?��� ��S;�?C�C��KM}̓B�5:��I�/�|h�jWϝq ��S���@I�{qs�߻��j�����cwL���/��܊Z�����ɧ|4@�^m���>�v�!{���m9���w��w�USJH X�|�A Kޓ��56Q=�H�$��ԙ �0�.�<���]��@L�m䵋�� ��U�3��@mZ�UA���{���eM:��w��XK�Nb_-A�F�X[ձ�����aB�G\�#MC�_�іע����t��<b��|*�;!|�|	��!�\����|��؀VI�)"=<�JCN���P>36�������VB0T��ms�fy�ƹ���9{�Za��8S��V�\�W�zh�Oc���ny�	�ɺkqx�	9���
�sv�H[袡���c�	g�2Sd��&e;%zx��ز�^��t?@��S揫8�k��
h{�ڔ� �$t�0��S�1���.��w �@�
�RO�
�c��4BfP Z!+*26�u�P�[� �����S��¡�m�S8�Y����ָ^,�D���ja�sIŦ�u�_�|�hУ|xCgu+�a�Ȥ!(�I�6���� �kcM��q�S��.�_��r�	���+2q�����9�5n��M���|�����.t��4�oW�J���:��N�9֋wQ���=FY9����5�AAqzŗ�E���u�0��,���sYl1x���P�����I֗�v<4���owU@W��B�Y��պ��w��������Rx���.���7�t����7�:~,��p˭~���!~'[�rĺ��6u�� ���%;A���1��~e���뒜j�'[�<�z$���ɩuk~X7�k�$KGggi���{��9=R��4蘟w^���E��<)N�.�ɯ���LΆ'i w3X�Ʃ�����[xx\�:���/�C�PON�S�\R���y=d/���h 5�U����z�(���R�.�����
HHJ9��t�HI����R" "�0CJ)�w�������r�Yf��>�{?�w��
vk8TV�ʩ���t��ftx�����,�[
N�� } #��$|g�Ĭ���r�c)ly��2�أ��6=��pΔL��m�$�GS�ߋU)��i�)��T$r��[�_$c���eΐ�.��i|����[]��1��.R@g���
BɃK�j��������H�>A�;ff7F�N6�y-�7��X������4��3e���<A�l��Ѯ�� �j��f���o�G�0�_�vLW������Q�V@aK�k�T�|�ᶛ)�@.X&���N���ѡݹ� �6�v!�!�I���-�s��ܩ���k���/j����+5�k��n��Zq����;���ds3G�׽9����+���i��2��o�?
����G}گ��se��= M�o�Z��f?n�����r�o�X��;���{�����H;QX��Ύd[��}���d��pm4�3�����1�J���wʔAZ�;����n>߅<g�S��9z���W��](������8���/-����
G0�8�D�.gqH��m��U�ɰJ�P_�5j�w	�||�T����c"@h��'=!�5%ހm���7�\��b~�����X���a�V���2�QD��JǇ&د%�D�t�A��۫��fF�MY�=�j@}�e�NN��*6nF�8��1S�Ő�d�G�#��ˀ�*�T^/��F�d��<�����8 ��q��Z2���+O呕4\�����O�&������ɶ��:��� ������8:2�-�߬����<�r��9!-@J�mRq�\~B��z
S[��Ӻut�{z��V��:��ٯʘ�;٘ݘ��]{�l��d�����}R��7���B�$���R	)k C�2��8��X$��]�!�C_}��?�'6N7�*[����m�e�P���Y��՟]�����k�g�r�(�j�r��_%.��M
·�Z|��$^0ίR���Q��w�ٽc�R�ó s�����&� �͖��v�[jJ���Y��Z�����)-��T@iV�ܣ��~~Y����>r\j���s��̪�c2�e�c��2�p�n/�O�ڗ�U��M�'�Ky�*==]Q�>�	<ds���n׵��*~T	��ME�$�<j�h)-M�����2������EX��C`�S�o�$� �Fv[&<QT���"��K�<ї�	r��`��\$��f�#D��ߥ���HAV?���\�5k�5V�p�:����E���9I����v�
;���3�������p ���j�����VVV>��L(J�juO�)x-��0�^�KaqH�t$+�9n���r�=Eo�Em%F䌅"��ᴷ�UA�&��tq��#]�z�!ul��U�b1 ߿-퀘~�UBSV�)vl��Y^N�c�JI��߄e��˻�{o56������}Ƥ�[l)����rd���q�d��9q���_x��eh0������D[�1�<�]kt�ѿ��/��l����M}о0C�.���F����
ʣn��W�E���9�[#S�R����َC-i��*����&��O���%V��#JK�����ȫ�4��_���_��Ѝؾ�s����:n�~����l�J_�+Ji#��8Q�;k"&���Xx�^w|�� �o��Q��BP�Hr�c�"n~���AWW�&
��	B{8jobq�/w`}0�����dO��T·�����<<�Nl�U���5ߪ�:�;̴�M�����3��]����:��@Zh��Q9�4��d��*-��q�lj��_f��,���Ϭ����4��ci�=Gk"�u��퍾�Lo�������⌎x���3��_�>��Π� )��u������ҏ˲���� ns�ׄ��t1����-��!q��=��BQ��GGJ@d"3����C!de媡��1����~w�?�h&�&E,��G����m����M@��fM s��Ng�s�:%������ڭ�o<��ee��ml �%�� z~�6�p8"V���h@���[瞯���滈�_��r��� �pk,'�S#����\��!��k@��� xc��L��-���6P���RiiҾРl<����B��4�<匋D:�.���wp�0;��l��f��Ⱥ����EtY/��@�М��h���Ғ��������w����o�w�_A:8ˁ
�F�ffpp�����&|��ƍ�:����r�Y@'�k~�_�[�A�VIhE�];
.����us9]�~c o��q�>�)�D�
����y�)�NMz~��\d�͂o��hph*ڣZ� ���	����z�)<�eS�>=���6L\���C�@���B�I��|\j�u>ݾ�Wh��Ӛ�𒎈 Q�$�M/1� ��B2��Ǒ5���Np�|�XX=�V�k��v򆍈�������J8����щ��=qs2w�p����V1�0�]hx�[�(K�Y��ۨ�ZZx�I���P���{�k�Ѧ�R�ԥ�_o����͚��u�%5��]�h${[
3��/��J䲧&�����bh���@���S�3�:ԉT&��FfOD��C~9J�P�~��^|�D��'k�qqZ�ͫ��̓�1'7�e|hp2�&�4���(��v�m�X;���*�pKKٲZ��o�cPű�����\;��Ԋ��>(��݋�����˥�?�5E�/�+-=\-���=r7��8���I�S�d�}n�>�Wv�����1G������:�c������W���>hj�e0!�}6��8ܾWT���w8F`W(&&�4���B^'�����V�����Mfbjj��9゛��@��$��p�c���M
�QǪ�ue�D9Ą|E~ɠ�G��rn/}��g'D�u��X� �L�w����mo���|�y����.�n'J��r����*m���p.7���FȸJp�O���������C�R�um�u-?������~�#�9��{⵩�~���)"[���"B<ى癿?��zn�)Cc�X㷶 }��k��GT�����s�{����ZU���QG�����\T���W���������Yn�y�U;ق<�7[��fB�AOZf �!-���a��_+���m��X�ҫ��9���<1!�C�
¢��@ s+��su��=��'�z�^�C��Y�CW��	���o}�����ӌ���m4T��Ws*.�y�=�p62}X��<�F|�S������hDt�2�!{|m���}����4�b��|}�[n?��)��%������#�h�<��KҀ��ʨ�'O�eɱ��i�G�fEB�z�����:�"��3j�<Wu>[���)��u�G���{���z|�Jx@�}V�_���U@%�ra�k	/1���̠I��G=��8�ԅ6���w(L���`�bY�x��C��#Wl�=֊��]�A(��k�(�L�RM5��u*�_7���Aw�<��	_{��<�}~������c1��,Yv��l��4t�{���"�j��}��nB��@��2)�JE.��n|��Q�l=�4'Ue�pޘ��ࢢ[H��y�ҪkkÝ`$A����m�W�ۻ�'fm2(�͙��P��x��������OS�%��������0.�9�y��2��t�{�q.ք�q���A%[�ڎW� C�$Xp$b��,j*�{랄Ն?ܬx�I6WMF�i��LQ^�śڗ�V�g���߸���*�:�(EȌ��fE�أ�{�3������4���O=�GK�}��X�����q�8௴������^6�Y_�V�	�u �R�2.i@h5
3����7oȇ�=#o@�z7��@����:ܺ~4bk��5�T~�1��)'��|	&^�XWa^�!?u�1�;��|A ����FB&օΘb8���\t�׀E��N��nP��`�rr�$��*��� �8t�z���|���_��ڛ��_�d�=8c�A��~T(��?��wI)
��d���啕�'�k"�����k�qs��ww_IӚ��·oV?�J��_113����Ԓ>5]i1����v
���q��wu��]��w$B�p)��2`K��	�R	7�=p�cy$~�zl5��)��#^��S����j� �L�M�fb�$L��.�	4�|�;���.�XƜ%�p����Aو�L����Z���a�|��B,)�E��]�����q70������\1s�C�Û�z|ፍWpJn�;�X��������.r[=���S��W���kۼ�8g�w�`�jRX�=��/���#*w>�*p�p�`f_6��v�������.]?^B����բzI2�u��ݽK�DME5,��� / م�]�����r�;�e��L\�u�O(��@>��ө0 TV���1E~u�������dlL�Y�GX��-�\6%]`�q��$s`��L�C�B�B���k����a�����)����]�*�7��v���%� ��ϥ3[x��7e4�7���0�l�o�O�Ă9썑N0h�g�+��--x�ӧbhAҵ5����^��������g����,��ݯT
$'����%500��ev����.+�Z��s�A��N��������C�]?:�d4�p�ꜯ��QDv���Ӏ�T��}�C���#�6�(�^b�����o���vf������/��w�s�zIY(�>sG�;�e�q��q��0��׸,i�,��Xd?��'�v�*^�[I~�1l��a�[�j\ɋ����n|���Q����3�H�K�3U�[HL��5����� T�7l����F�]ֿ�{_G���#�*WR�t�` 6�`��H*"�.�<e�B�Y_�
�}
_�����Q�W���k�-E��W0L�w�@�ݱ��@�pP�k����eQ.7(�o��I�f� 1�ߙ�hVE���B�K{�zx����*yј&C�D�m9\����]�iG`��/�N�e^����S��o�oK���m� �+��4��/=��vln��O��^�z��ys��՟?[��d��=<�V�����!�!.<���|j�@>�zC����4���� ެ�N*��	IP���vc��8���cm�,|�\�R�/%2;�%�D��
E��xa�C�gYM�}Ax|�<����y�5��6�%�>3Hew‸�@���&��)	���A�;Hw�1{X��0�36q%�.�_MB�Ç��@'+~��8- �&@�>�v�UFD��I��6J�%��U5 �J�6�/_�
k &H�-����>����d�O���c�����1���. �CHx_�#��>F��11���ޤT���!145�&ڷ"�����Ąb��bw\�n�����ov0��׷���K�o�[(^��9b`jJ�8<Ħ�7��|:�w�����A��T744L:"��m��&@l6|��ر>�q�Y�H돫���f�JN���F�=��,��G4����x�m��eX�{�qY@|3��o{!_;�g��ϟ[�H��a��� K�ګ%�����rFĲE���}��\,%--_m��2'b�;�~y��'"�'�Nk��^m���22�[����\���(�3o�?�!�ӧO?�I� ��GL4��E@���j��[c�*א��L�|.k� �h��ꬻ����.��O�?�B��,�!�@�NOZ������� �Љ��dk�r8(J����Z���)�rx~{nu�W���B3ZY�!���e?������m ����(;��_��ۼ$����[��������;��8ɫ��"22o�'����G�e��'''�"'0{�<!��_�|IZ����y	S�u��f�����}���.��K]J�)���Jה��J����U1G�٣`�C|"�P�v�<!��o6��{�=�֨�O7fr��5.Q����]ܼ�LN�f��M���r7}e�����Z2&!�^oMY,��A�������6R�[i��B9զ���o��v�i.�ŞtܾlG�*B�2�f���l�?��W#�%�Qj�oi;i�`WU���Y�W�~dk����o̞K�Oe�}5�G-8�����o���̪��U#��W�"���-���"���f��ζ��}(��'(��L2x��8����@��CE�]ŷ�6~;(Ւ*Y���6A�����
���X��e'Zγ_V7L�_B��fW��o*�	�I��u%ف��ٶ��bBB�����1�~)$R$o�fV����%�Y�k���3Su�=��%��T\�rL�����M��.r�R/�'�./_b�@���ӏ�ŵ5���h":::�\9@����%���e�3�-|OĚL+�?�tR����bFōD2�k��J�Ԥ &���_iz�D� �"�<����{{��������b��{���F�&��0����VX�A�XV���8|�4�>�� �rҮON>;G~v�v��P�$Ƴ��8��d�(G_?q����~�J�Z%�n����:̡�4�/*WFӹ�����4��-K�}�?�R�w��V�`{���Tb�׶3ƌ��|",fvw�!�e��
�뻍�4���v�z�j1 �[dr2��$�7OY�q���������ڂ�&^626�y&��1�^����H��1�j��>cv^^p ,*|ိ[���Zi+i����'�[(���m��P���}u���⥦=�qq!y<GT����U9av� �DE����=����^+��2S����&6��^���k��?�����C=�Zޡ%Ξ��Ŧ�h:K�p�Q ���O�ޘoQ��41�O���N����1��
@B�8�=��U�굯���3�yP{��Fөb7T��фne��,zy	[�x_�V����,���Cž�����ag��4��
���E������\}����f����AlQ�S@��B�����=��%`@I�3GC+�Dɚ* T5��a��4�D�� H�%E�V�����%eX'�.؍~2�PiC��՝�zU������'�y������8���b�ru�`z�~N��uP��u���Ο��7U���PV���H�5 n������k��JF�4��iI�z����Du�-�������{�ӽ��kNU����g�Ƭ95��c�ۊxO�Ͻ��ُ4ܧ�%�L��˔�'#@1r~MzXc��h/����&��ft��l0�/2��ur{���66�P�I�h�q!����������w4I�LE�rrb�K+���C��/{^�l��ܳ���7x�+;/�`�~1��9G��;��L��p0������]///���F�+G0�92��n�L��C�'j�K���r��l��rx,ɠ�ig'.���V���ur+��f-����� �߱��^RAe�}��D�E�2mg�?FBt�İ?`��G�f��Ȝ�+��	ܻ�AQz3b��tb�Zة�-�)�����^a@��I����D�`�c�$f��#�.��\w�z{[�',n������ň���L�倿��'k@�F�epF��L��?|l�����J�D/A�X
,�S|(%.A^I�
Ǘ=YX���I
�E�@2��牯�]@luƚ`}�&^��q����-R@m����DDuw�"�Å�*؀�VTV>m�����5�1H�g|ʑ(Z����Tm(W1��O��@���7�t�\[#�2\*j�|�X�T�� 6�%c2�4�=�d�Iخ )��q&�@ 9Ȃ�%����/p|_�8����k;�v���4Z����j8���}��晙���j�[p�#��[���F������A]-���ל� L�ܦP��f�1��j���8ς^�o���T0f=�*�'��wTo���G�(.C6o��m���a|W4�	ɀm���"�/Q2�J��041	�"�\�΢ݱ�c��L�����v�фHe���s���J���r��T��A+�v�٥1�mG��*��P�C��nE����gS�MLL��+]x�����:coR�7�p�����BJ��r�Iti�yX��(�z�֦�4_w#�7�B��6o���'V�����/��q5i��$G)�����8X�X��"��]�o��E��R�+��苡�1gg�Y��� .��B��������W�yP��N���ǜ,1bp�����n��+$Ȅ�j��^�b_��A�Ȩ�K1�
�,W���]���_�?��ȥ���TxiCP�3	5s���jo�N4a`����tR�j������n�o��r�ջG�����WX����ZoD��� G?1�<`�:!fs`˅��}46�t�wt�	�2�����U�J0-{6���9��f�(3��k<����,O�������#���ͱ�5�N�=y�˾b{�w�9�͎�ȝ�=U�C�հ#]$�����Lv����C����1��!.�gT�*�9��t���cJ2�o:(1'ggׁS��o� "zX�e"���w;��&�JJ���Xz��EDj�W���N4Fn�s�#m��P�c�W�4P�Q�V�ܽBbbq�۴_f��W�ڄ���I#M���;C/y�]��3?��8y}}Z���{���l��8�b6�UR,��f��s�s�/7Y��a�$z�����<%%�s1n��_1�l�!��iii3��'H8�*6n���@��a��G8�_�� |�q�lj�+1�����eUlDg%�C<��Z:U���\)e�fgg�{4���|�'��Ϗ�8�8����9�
=����� ��.��c�,\���;O���9|{	�ڃ�~���� g��}Wƨ�� Ui����ss;''��^��|F���P(�+K��@I@;����m�)x俓3��}#Rk*�FՆ��f
LB9ܧ�ু�;�!nf1�}���:�_�;��G�3��uQMNZN���#���"iʭ���B2�	q�8\����+X;��\�H��[�'.�a]gQ�Iaeݸ��@��g5|��1@3���6��c�	��oqc��W���Z0�?H����^���gFL_l Z�U��	�?e�L����t��{��FB ��d?*�\�+�g&M����}����Ȩ�Q~�2I������������9���O��=I&&&�7Tc؈���P0���]y_�~q��t�c 3>-�L;��~�:\/q(DÁ�}�\���+�'Xn"����ݕҥ�/]� W���b�����{�z��*O+r�/:6)H'M��KB��h�\�u{H[M&OA���t�^�0^0��\���qo�ZEpݗ(�Q0R��緕�ݵ�3{|��XO�lDHF.ԍ-+���1��tx�;m�e�D����̽lg��<��B�C�周f���������罰�/Xۤ.���%�' ����;���8�3�Z��2̺eh:4�<���~���	� �`�Ŭ�/ވ��32RO�,"�S{{�Y<2r�>��Z�v ��Y�`���|R��h���~��KM����b�^���y���[�Iн�*��#��Ԛ�܈�+�/@����|����K+%��$tigN�/�sM�N���Ƿ�i�����l��PRr�9�=��)��˾z��eO̡t��ݽ�$Sw�ލ�Y�15�	u�� �77?pr��>�&���W��)_�C��y[U����@	%��h��+y�t͙���5#c�Ml�a�ׄ?�7tMB���E�L�+
�a�ڏs�}7qS���.//�c
N�ʔl������'n���z}�ݠx�%Wd:' ~ȶ��N��ɗ���	Ω?,����&�eБ5,lJ���ۿ��s������T����Ib�u����>��T+~�t��n�Ie��xK,�]y|�OSp��Hb-�M��,����!�͚g�9.T�Ƌ �D��*�J���-f=W�ua�'�oq�ѩ�H���"�+m����*�.�� ��{ו���N�$$%�>��)�X�|����o�ha�_�+�ƽŭ��j`Z��H$*NWK	**��;�c}gOq������/��l%�� ����V��NS3�g���v�\||2�6�a�C�E�~>��d�lAOn�z1G�,]Z������3_�xm�A����Gf�3�K�6�2�f�?D��tRWrIG'�x̉��Q�B��e��?8��0� �a���F�g<�R<[�� ������W��@��HQ�����HI!#J��7�Y���f�2�[�b����AE|��$����JET�ah�W	�ZZ��K���B�Q)�w>�w�p�z^�[c�e54Š���k�δ��*�U�Y�׻M���P�®:m�_���`�ퟲ?H
	E����FR�����Za��x?��)��nT�b�sW_zf�";u֮�������C�s\����t{��(����'AR,�h���_��\�&(\�'��6�X�pÍXF�\�ѣB�W���9:��J=)h�� A:�Y7#�<�4S<�C��q�	��~�ɴۘ���]K�țGT�����
{�� df�~k<�4��uӰz
��^�`���̳���YcG'^�*��N�OK��V��W�;�=�ܺ�=��]��F�����~�AY8v�L�eu�V�t��b�X?������T��j"�텴��$�#� V�KG��W�nk��Od�;`��m9\�n]4�>��E��)���+��Ȅ�E_>��֦���`�R+�ҥ��K���55H���Ygkhj�v�,��`���~��w(�2ɫ�E_���v���G�]�s D�&ܶ�o;���:�N�L4�������������W��$$$[G~��5P�l�鵋/5��21X��(x�E�R=.� �{y�lR<{��F��qf����K��������Y9	���_���pN��61���d}QN�%8���KI\�XU��P�_�������&y6K��z�M�)s*0�x��3Ym��7n|n,��N��;J�$����$.�V [:�����7H�}�U���m��U�"!<4��K-��Ʈ��@{���|��d�⏒R� l�r�Y|�K�r�+~t�o���@��;{@ɼ�O9�����e��Pҝ98`U|W��}Ax��
]�<��z`���Jcm$��t~Y�+-��"�P������������MQ���{,�y��G�����zO�Y�� ;��2 �X���%٘J��Q���`C'�__�uX��++W��wh��W=L{��q��&$S���<���V��I���oQ����C1�W���!��B�8&�7Z�X�dX�Ym1�gm��nք�� ?�+PR�x�:|��3YR�?v��C�]cF��`���-
/)OꉋdNz͟��jԣ(�u��;f��r �9@����ń��_iyU��J�饫k������!9@@,���X���n������vihk�͍�<����ʥ��u:�W �B���A�v�| p�±��E3����������7�U" �}a�� ѫ�����䃓�����+������a��0�%{=%ʛ7��`�/�5T����j���������8v�ŀ���"�M�"��KZ�<��g����Â�>��B�v��	}~�l�\kYѶ�B��}n����?���=޲:�a>��R0�ϟ���Um=��M+��Y�����2�eq���ەy�����ʼ=��Pah��¶��V����}�k��]C�n��8����s{�푝Q8"Q�y�ƾ�g��
['������e�����:���6���mV�苛A$r��:������%��~UD�VL����7��2�˃���|�(~�宀@��a�r�N������Ώ��j�G5����SFG�����|�C��䡀��d����R^Yi���7�y;E�ϸO�m�A��l��V��ss��cRV.�Ý�@���v�����dg�t��\O6!@�A�@M�1�0��_4�b�I���w;�Đ~?��|����)=c���5�^ˇ	�d�����de��釣0�˾R, c�å��q���|��er%�� ��[���5��@9�h���0�E,���B��D`ܾm؎��3J��/���(��ؠL�.v�<�V[~�$���l7�ᗗ7��T��¤���»��λ>��6NK�!!=K�Up2�s�=�J�C2缓@��2%E�C���K���tY��=��ϊl�gGFn	ܻ礮J�Dh�66���\��o|,�L`|Ni���M�3;�--��,����n�� e�d*��,7��Ȟ���w޿� ��4u�����\����x�5��#T !+� �U/
�#H"�����"��S����_.�D^=}%�����i�K����o1���n�,�͗��D 9�ܻ�q�l�:q�OF֧��t$Fs��G��R,�of\$��Sū����c��vKq�i*tb=�y�,
|�L��qXz�EwOD������ݖ�����14M��zv�'	��*G�/�k3�/��˓_�lV�hV��द��n|�ՃV����`��=�BB�Əy�n���Btw��9�E�l�������;����ik��?j$����iȒ�Y;�4��2M�}89qvqu��k���;�mii�GB����$�ܿ�0��[��0`���������]3�_:B̨j�܄X�c�w$UY)��e^h\Q��W�U�V#�^���1|b���B�1����z��8��A��L䘧>�a��qWy(dݚ*�6-,چ�f��/FJ'Uw��#�W�Q�0^��ѭ08l�f7+fW�r����9�g���V)�90�]���g�߈Y�&B�v�{�=�_�=���@iARN��v��d�C�/%�3��!�3�3���3��ȯu��=ր�b��9O_AYY�ڬ+ckd�UU�${���d��NW�x{��|F��CB�*V8~�mI�g���ҠJ���ߊ�c�uDȢۨ�x���?��G	�B���ܟ>}
[Y�I�'�o_Ѯ�=,��ԜxƇ�A`��*�Y�oVU��;s|L|��oJ�&�J�n���[�� %{z�r%�_��4#�����H#��>%��!����"6(��N�~�g#�R����sں'Wg|�7/�j3�	��"��Ӝ�6'�i~�k����Q5�h<��Ƶ���(_�;�R�S�=��n�7-��C�&%�"(G��z:/���`6�!bsp����vCN"K�WIIv��{���T+^P�-��z_��%�ͬ��I\�!wrr2�ћ�����������;�Vܷ�����4��,\]�gV�Rԯ<}:��CM���=�xv%�sV�~Z�����&!��R�Y�D!�g�!ߐ��'i��-^lD_t�n�% Ǘr,1֊��}�Z���29xb]����"�}�h�'���0���^�DR�g���.�$`�|�5
�/C��ҹ\jP�#-1��sƓ������	�C	.�̞��0{X=+��I�w�@V��T�Kr(�ݒV��[u%dEo��j���<*ݡVxT�r�+�\�f�yՀC�^YՌ��z����uq��lZV�� ?�8���}3�?�GnLP�Lk��$b�{ٿ\Z��"U�,�	~��T3��02>�dS[[��X[������
X^�@m �h�s��D]�+���ѥn�u3A�
3_�i*��ttwEF�{�X�=��[��������=@��҇�ݾghMO�"nʸ��C������Wk��B��	Jx���������ʗB�u�K4akDXV�k;o�-���r�@��� ��_V�p�C}���+�4
��hۧx
肍2�a����wb�������o5N�)��{P�s}[<c�խ�81i`�Y.�i��>Vb�W�.���ey.��c��l;ٯ�f�{o[�t�4ɔNm���k������Q �3W�b���+���0UY������'��rSӁ���4�Xʚ���R����FFJ%<�L�D�/�d`�g]b
&O�KF8�>A7� �4��j\��������A����i�XV����ˬ 7q8;^��U��<�]�#Q���]�@I�*��_n�K5@!96����y�	&�Wl�t�Z<-f�]׾�r;U��:.����t��J�*�m��w�uω]�(6"J��QjU%�qo${
�Ԅ�ˍ���?z�J�-X�<8Рk$-t&\��on;B��.k�(����bV6�B���}ڬ�:WW3W�>�UE�;{6Oڂ���/�Q��N���n����;z��k>�0<<�:�h%պ;����pGFCI.("��}���IIX�9���}q.M��<�Ŋ�#b��.����?����J��ޤ[�*Z1Q]�c�M)Zg,ū���J2J���i��G;��mJ"i�#?�j��t��Y���9������)��s\/�n}=�8��ס*'��u�0F�z������0t�ڶ���G�c��ԗ��4�My��Z0a��$�b�xl��ݿ�a�sz-��K3pS�q��0�y���VwOr�c@��b ޠڎ[>S��C�ʎS����nS�323?KE��{V��0�S|:�`8�Խ��OmGo"p&��;�C����16y�L����&�A�'�[�r�I_��l`����5;�+�!
C�6�^�=���--rᕌ.��Qsg� �̪nD+��YS'q�8T�q��q8�89���.���|�n�Rm('���/��\E��hM'u���7���Pj� %[��6e� iWP%��)�� ��ZE��V�5�?,7��U/r��+(�/�+V�ӽ��`a%�$�i��A�\�S��m/��^;h�.(�ԁ����`A���++N���j���΂[�:k�v4�*�������7+�����N�ґR��R�kk$�M �rr^��H?&*{Eܙ�hP�}v�@4+���pI��૥Џ�� �g�x���G�$����rk�,0�ʟ�Kp�Nj|ߣ��yݷ�')\׀�/�<AR�[�@3{o (�PK�M+o�:�P��@Tl<EL(UtA�������ط岏>;r�@��p[����O+�a�M̝��:�v���2�A���EL��b����t�$�k�&?�l�a���Ɂ����g�'�ퟞݿ�
_oS�q�I���V�K6�J�������ihb�9[�t]R���?��3m��'��ܦ��� 	�H(�ʬ�<����N4bo�L�)T�����s!j��KZ�Ǐ�����U�,�uZ'���#& �r�~������A ����zx�3����jb� 0�WK+�g��I$�E��[׊c�@Nלﻌ�c��k�����h o._�g�e7��Ł[Yp����ae����C A��MhI��C�.|"�!���y\j�e?�N�qt�e^m��0�<E�;��������v���.��!�.z9���^��UnS2��U++ī��̀~n�ߚ���؎1�vVK�K;VSu��v3��Ŋ������SF����
)��Z\]j�]S���olr�G=���~ʰsM�i/���P��%z�Κ�L��[R��sD� �ӵ���'&��3y6�߻�V���Z��ߜUmH��MM3o�֑=�6;-�<�C�Aӥ��B~B�=Q�C��Pyդ0�j��֢�#W :A7R?��i����$]Y��Qv�h��Ika{3�OF��rL��'������k2&Kk�)�C�|�޿�32R�1*W@׽c!ë&W��6��W���Û�V���.��B���N�t���c� ���ǂ�穚͛S9�f�\���w���.��|�?�=����<���qu�<姶sj�*T���2Α�T���4�v!./_b�xA�����{KIX��h��D�Y���J	�H��o��b�],Ñ444� *�wi�>pK�^q�cT�O��v�X��A��@��N�hc�}<�vY���ݘx= ��Y��{ ����.���]a��F)���1	�0N�S� D��@�➗v㤡��B�׋�q��Ƶ���x�7m�Y�E�%���&�&���4A����k\ޤ��ש�m�p��Z�u�Zq��oR?�cOp0���>����`zӆ�����/nU�B3A~r�5�i�a㮸V߾�>�Sɝ$s�g��4!}�)��fT1���~�5��; J����Y�M�@l�v���7UG��+a���c�7-���===��9��K;~~�u:��s壗�22��Q� ��_��5�+.�堦�''h~���������f�2L���r ���d�'����>�9���Y<{z�DHx�g|��ѫ7J�z��GG6վ�.�39	�_�`V..�]]][�-v���?
��W���m:>����X��e�N��{0/--E)[�
���l4��0���[���+J:*�����%��@Z�<C3j��H{��=u@�Q��U��+�ŝ��Q/,�<z��m8f-5�����6�RX���=%���o�A��R�n�{{���Đ����6���k��{��~�3I$"��כ*Ƒ�MĐ��#�g��F����A��u�razz���;t����V�Zy�� ���\M�U�|O�$�`x���}a��o22n����Z��~H(�|��&�g/_��^�M�:�h5S�e)�(V�v[6n�*����H��<T������Y&��5��31���k��;S/��Öxl�5p�_ǌ27���(n��J�9S�������%��^�ȽzuR��Ow+��4t�6�Yo�Yqg���"��C{Efzƴw�d��qCU!Ƈ�#���O����D�e�idf�cN%)�Lw�e�է@K��x��O�����<�a�����^�GtmR�>�z^{���4Q8&23憆a#�+H�� �{=������5�7k�[&�<ʳ���pw�M���Qp�v_�l�b�β��i�����Ѓ�\xY���@A�W
^h"��2z��{PTS��DY�?���vݓѳY���Q�m-XV�D�'4�_���������Gf��Hߕm�Ev˱m=N|pq����J���9 ��~������T]9*9����`!s�6]����{��+�]�ٻ�k�t*��Fp�s+(t�jd�h�A�Վ)J05�+�S�9}A]�պv쳾�)�NV�ƃ���3��GȺ7)P�[/��w���q4]�lf� ���K�D�Lc�{��O��UçOm�qqq���$(@8NN�o����}q�~ci�)"%e�����<C~:~�f� ��z[+H��L$����B2���/�N���?���3Ԍ�zzAW��q�,"?��:r¯NO�"�q�v�r�Ɯzff�""#gݛt�F����J�~���Ҍ6�L�[#��Q���.�6	==}GGG�Kr%��K+ ��[u����f�rz�Ҕj��ݔ���M�]Y�����|�yV�XI�B���n��u��u�ؔ��
�>�?���v5Rt=PHJ.��]�,L�9��_��\�+]W�&�O�{�]�����32��I��4Y��/����Ĩ윜���N�^m�/q1ۻ����ѧ�Jf���xSt���y����ۮ��{M>��3ss@��9l?x]9��͍X;O&�iv���v��h:�x*����B��!���#�Yɱ���cdfo�압d{&!�ӡc�8f��]����?y��u�������k���m�Jԧ)����"��yw�<�{�8��k����w�ֲFuR���DH�1T��������R�lT���N����C��f��X�ʾ�j5�,k���2�@�H�M�W�ډ�-d�z��Ӣ�y�g�|��]8��Iĵ;��P�Sa��sqi�Jk�a��]�W��u��JZҋt�9՜�����@VX�$�"�e��E""�&m����h�[�##���34�Ty��	4�y`}M4\H�uE����n��!D�m߾񇇇�㆗�nl0��i6؏P~Q�fl��I�+��,�ֶ�ʦ��#**�{,�=�Z'��ח���W����o������IIt��鮸ջ��θq�Dqё�M�s�����*߻)3Ʊ峩p+~:��	u�����i����ӫB�Sc^�.v�o��B�����t�N%�RYt���+�q��V%=ŠKoP�θ!��<)9S4�=�����	f��.Q�7����;Da\k��<F��9m���k[;�Sn�pYG`p��Ke��,%V�d9�R��z�<����afe�z9=�t$����:�LŮ��(�(b��Q�BaΠh~�26-��n� D3F�oA��hu��F�-���G���?UTl)>��2�@���6p9�Q#f��]�f���_����J\Gj�A������:��ƥ���
��n���xE��Ot����I��h��Z��@����ß
m����*3�'���K��p&u�yh��Y�vfvvB}���%3��8���f�̄X8�>?�^��e/�B�h	T�"�V�p�����dy�������ȗ�Vh�%�m�8��4�2�}�[ƽ��o_U��<��0�Հ�
����+(�a�O#��a�H@O�үyN�&d��u���l>�\'�@��\S5Ӵ�X�fSh�0�sM���2��ۣȾ��������O��^B��㝔i`�������@����Дd�ۢHeKK���M:��_:p����B�f�i�^�����]^P��/)2_:Z8e�7X�GEF�y�p�]$E��R���b1E˔�����宮0ꪢ����Ծ��q�v�]6�©�E�S����_嫪���nlZ�Ԗ��p%Fn~ 0s-�N�?'�ᄜ�Ǵ�!�D��jо�����.|�Lj|mo
���TM�6��k��`l�K�T�M<����̫[Zz��	�#��Xht7��e����.������h���+�&<�ƻ,��0�QvAA��w������v�a=�e��C"��W3M���H��j�{�,[[���"c��wɑ��& �!��Sh��$-7n����ù�1���?B�Fk�C���AoRp����^9�dB3�MOrt��̘��������}�|�٭�͍����Y�/|^�u�.��m�>ZT����QP(���uJ�2�K�HRSD��H�s8���q�@=[��v����!��!��v�*����!�%������V���*�luo �-��*�{�b��GoC���keP�	*	�!~l�1��������k�T��_ut�薹)f�,5L{{yED5��R����%I��dL�G䨓۪���2cC͐-���b�/�М��L=�A�o����}����`��z�TQ�nұ����m��TxhR�DP_b�ld��yH�f�)tp��>���E#ߍ��ǌ�pӥ孺D����	���}�c٪�5i������5�K.�rbi���S.�(	��)��ʏ��i���3j_dӵtg����A�+���5+/g��XR����9�Eu�v�H��`� �&�"eÜ���2ܟ"		y���C�UL�<h|��.��5�ς�p�8��%��Eb��]]���yGvk�������W65E��Z��@C��x�uXՌ絘��J��Ķ�k:H�����WJp���d���o
�N)��wG�A�:0Ӕ�q	�k�<oE�8�PS�n�Ȃ� =��^�c:a5F�o�����IRdZ{Kg�!���l�ۋ�w�*��T�<b}u��@�cx�ו������e`,�h"i�	a`�;(��J�:���jE��$����n�<�n(..�QgN�^��_�qKU_TNNď�ؑ����XJGw�D�=��s�	k��q)�������n���F��9>(Ywq�����KK�����v�=���O,w��ma���&($��Pཐ*��t�D�ľ+�8V�oZ���n�ݓ^]��y��q�8B��C���ʶ�ë1�J���@��W�w{�(��|�^�+si��C1����q����\�ӥл�Vj\
��-l�׾>���̸���5�%�G��?��h�Ԏ���5O��4o�(��:	�N2�\N{�A��G�-v��.�ywy��P *I�����L�����+M�U��my������������:Vu��K����D�#�iO��R$�g|�$Pi'��M��63<<#��Ɠ�0	�<~^��?E8Y�<w��2�~t�bP̃:�j��o��>]�@/����~��S�N��P���J�k�)xv���z�>?��.�\c��O��"�����gΠ���
�#��P�N�������&�4�ʉ�B�?���93��a�]�%�u
ݦ�-���χF��ǵ�c��qо�+�Zwň������Ԑa4��O�@lԍ���Q*����y4��_x��Э�;=���׾Z���A!*)���}*@ղ�\L������b�(ik�/����7=mű�S��T@HDTU��X:0�Dx}����9��l���^��J�>����� )�L�+Ƿ�:wr�����Ӄݵ�،��&ip�M�Y�$%��z�1)ƥ ǵ��������3�������;��շ=�Z�w��oy�=HS�V�ֻ�d!%��0���c%��\�R��7X����b�͞.i���)td�P�n_�����@���N�9�C%L��6aj�3P��
q�9��T�����
y��~���>�+��<>Й���p���ϘO�Q�XZwvb��ʝM>T+�fP�߿o�D䙧!Cڠ~��=-��n�y�r�O��.2�� C�*�ƜN7Goo��ǅ=�#�ӣ�����I����k2U�b_eJEF�t�����3SVM8u��;hX�I>�]|�=!B��A.�%-#!a|QRr����_�
"`.!��zt����Ǻf���?�1�y�(�9��^�(>����N�f�d�K�+)���-����ND��:0�
|,wo]��g�~r[���,� �}��h8�p�Jf��Q�-���+WWe�ˠ�A�vL�զ��,�J�u��� ��}�wո���*w���?>��=h����5!�By%H���{�%3��������OdZ"��D G�-BH�-�i[cFM��V��hȡ�;8 �'wF?'ٽ�,h_t�D�,IV=#���;�^H�B�����zs�b�I�3Ow� dE��3��kj)v��0�Z#8�P<Է@�X�XIPq$��R��Ή�8�sR�}�k�c*�6�����ts�"��+�'CyZ�t�t��(X��E���{��ɠ�U턜����ǵs1j��]����nn�S_	�G�g񀘥m�=#--lp��|��Y�n��(�6�=�-�,��xH�ع���T;ji+�u���� -\\��	������TH9:�	[�D &  ���N(h�?�42�{B|9�.JJ�_f3D�4;c)9W���wr�e�y�Z�Y���|򭎯���U#@Xٞ�w�a��z�)��2��V9�F�CfC�#1�����Z�G���g#mH44�����/����g��~ީ���f��������|Fژ������\��"p:�[������K��N{�`��f��@���}���|�[���I��/N&�P;|k�r���,�\��9�b��	���b�7W��;������Ā��w>�j�!? �.�gܨ��G>�b4��㡆��e�s�WRh�|�zն?�MZp�R$a�_��6U��{#kG>�ZvH$Yt�X��p���0A���/#5>��s��<��C�x����}8���p�������Ǹ�r�UH�RL�`��`�@N��3�����^Q
mJ���k*����g�[�Hķ�A@��ܑ��.z��|	��<{.�055��	���{\U�q�n?sb��Y�p��t�0>|��<�� ��dG���S�Y��
1��T�֛�6���jrh�۲��4ҧT�9w�'����;�*Dޢ������L�$��ȸ�$�kp��S!ޓ��5f��x�cr-u%~:����@�@�Ix�@M�\�u�2ի@�o�z��ғQRާ�uK�����Yg./�e+��%M˸�Cw䋮����)4��ʛ��S�l��gTԽ��١�ˀ��/��DLWpZ������ϘؠbX!а�� 4���C	�̞���`T����^Z���qq��L���ꠅ������?�Ro�Z��$z<g���I�9Z�G���4:\�b�
t)Q����"�3��=�������̖w�I��X��> �K�|��E8~���?F	������yJdh;��
_�������^�����fN��O#��{ ��������W_:����n���E��x�>���ˠ�{��MV��I+^-�J��m�6Z��<M��ށ�k�|�2��"����N��ڰ:�#l:�<Iz9x�[VI_x����u�7�o�bt,ʥ�ߠP7}���JJ�:�1HNFv2Z߄��K��������)�%%�15�y^6��^0ۗ�r�W{~��u�O�ࣖͰ�C�F@@>� U���l�gd̅M(Zk'NA8x�,���+�Ag+���RR�5R8�&�Fȓ�LFQ����i �Ϋ,rd�O'�?4wݗ��휡wʎ�����o��g<�G���I�Aֶ�AV�ʉ�@Ĉ��B�d����M��>�:����k3��I6Y��H-o�9�=Ar8��[[<)��8p�������x{�֗���&_���TR����D\A��ý�ۀ߻�x;��w�:���_Y�"Ѐ��)죦�(͢"���&���dH��
�4'Y�Fn4�'%=&���L�w�SU���zxuk��RU��A��7�_�(�1D�0%G�%V��4���
�:/�&R�`�7T�|Ñ/ܙ�l�����Z"��=�H�P�C����PS���ʅ̂�@l�u�l'�F�?����Ύ��;WMm�~����7�V䑙(�������f�,ll���A�
�M��KemoO�S�����3F���e�E��7��2���g��k�c�SH*b���k�dq�p�AS�C�DC��A���|_�6E ږ�{khh�$KJfA������嫠�=:�딀���������P�J>#4��2��v?��RzҤ�$Ǭ��%���!��R��A����a�1�q)���#����*#�B~�1�O%Y�/���}W���z>���Qndf��lBl�=�c�0aɌ~�3ʋd�+��Vp	|�d��1�E��EQ�#����ݑ̐�������g���`�"�d\������{.,�(�Ʀ���!�΄�9��'�@�����f)}�;M|!�ijn���ε�y�bi)İ�5G�wvB��YOt5*�լ,�������2�cE*�yt)��D�_���;�� [�����r܉<z����-H/4C������=�ݨ�r�ڹ��%O$��;фߘ�j�Q6��:p�|�(mB��tyX�[Ф���_�@x���X��_U��vw�`R�m�����0_�4�5i(�£�����?��`�j��ꭙޤ{��,ͧ��˹Is!j���m�|8��n3�Iw��}ĺھ<���O��śĬ�Ak�x#��ۮ�e�9p���v�+:S�\� ��f)Z=~�\3>���/����WKK�����鞒1�3�y�s);�G�uu�S��k(�b��W �ݾ��r*gPl����en[e*�x��>�T����uM��HuUCK,S���;8s��x�wq�!;p�u�%,�"�@��/�ފ������� 6^�dMB#힘&Ĳ7���}�������NJ���P�!�?�}�t3�w�y��Ś�?�fe-�~�al�j;d��v/f�	��i���2�C�P�����kFFС������p������g��0�(�|�@tpb���f�3��n����(��(P��E�D<ˮ�P�9�{G��`��w�''a�koݴ�? '��G"wTe�u$�߸
�ii���G�y<3o�%�K���HNLIq^(w�r;��I��#�d~�
��׻�LӲﴙu�N������K����7O��4�)��}T��� �Ȕy��
��-j�A���!bCF7��no�nz�ה�`�X^Ǯ�Ft��\�Q�Z�?V���Gll�ۓA�EH����X(i&%���WcV����b����;�8Bŀ��F� ���hfU�m��/6�li�C0&�QG�Ë���(()Ü�Tg�]&�`!�� ��$ ��J�(���,L��n�2IN %�O�rp�M�F��@=6�.�=ͳ�[\��x����d�\n.*��(:g�_�!�M[,Mh���$�>�?���0�D����L:S�������@�a���-b<.~=�pff����1qzA�>~��Θ����c)�	+,v���t����~ĸ�q�SS�C��/(�eQ�Aw��	��Բ�g�y|�Y�d��=��[8��u}���97��>k1WPXh]喾���M>%o�J���㒕�M�Ѱ��C*����	�+1�y��H}��kd��o+�"�"6�җ�m�&�|Gp�mk�2k?x���y��������j����:�&MM�zHr!4
�©�e�>fP<��>7���k�;��iďZ�-(|BE������O��A�.���es{���a��_�U_�FSrLnYߠb/1.5�8���6����v�?Њ���aVt'g���
�.��Uo�z��Xw�Iev�RU�����}B3B�����a�be�* k�i�§=�
��v���B�����5UvD�I��.@��u�Ɯ�_���W���w4E���US]v��+t����ܿ�}��A�mȰ�En��Puu���I|�������A����w������GC�H,����rPKqD�0f��bb�芖TϢ#�Y-�\ǔ����o�B�����k��ލ��O���_&�B9j|�+rm�#ǋ�B�M�feл�|(����6�כ��>�Xp���P���\\s��U���)�n����3@6��A	�.�Rj$��6�EI����Z�rn�|a�����A#RN`$n�N��5t�l�m���7X�TE�ƺo�zV����C��&N�h^�Frh�*����樽�G��32X��O"����o������iۉ���r�;�<��J�h!:��u,�MLxI�����wd�����[cu�^��W8��z)Y����Er��=�T.�et@Gm?tG�!�\8fd��rÓ�kHj�-_Q(�G`{�a���7��  ��}�'<��Pp�O��S���^���4�N��� ��5.�����\\o*��Z��������e:�����W�R�����Ç�;�z�w㔄-~�����i���~v;��ú����C�ml�S��F��2q�f�b����HScy���z��]���Ϊ��r��jnO�P�|�YD9�$!$�>>.�םb�C�V}�Z����"��+"%Ek+�B,q��^�^^�qj��n��G��bT����Մ#�C�����G`��s��(od�C&Q#��~��~��� T�k��jb�&H��:��#"�kv5x8���J3ā��fmӔ�J��ZJ�T��~	)G��b�w������������o֣߮�z�w7�e+�~���8�5`�|��\��
����j�h�0��B]�����}z�w�L hZ91�yLI�C����c��b��g����[�u5�[�������<Y��� ד�1�
��LDD4l�<x���}�4`c�l����-N>�����I���'�踴��-s<},��?��r�L~�X��]�]�U�T�8�v�;o�J�*�Ƭ��x����l��e���=�������.7��"�ւZ��j�i�[" .c}��-<f��[&ER�W�H4]W(�.���:�r�����3XT-4�tlE�.�M	��n��ncن�5O��޺իF� ��iZ�Ĺ������ݿ�Ƀ�(��͝�ۿ��#>$|1�^nF]*�k`�ƋXR���y��b�j̔���[�z�|��Q�Yx��;-^P����݇�'�^�Q�����]pR�?��߷n��i��W�������=�r����ǜ���A�{$��Y�6�p�-'U)�\����|��Nt�b2���[���Z[K������
�¢�}i�wJ�W�t��N�a�� ��H�d�Ι����ˋM�L��]8�T��֞��w�V���_κ`Fƻi�)�Z��+C̕��ۀ0��d��!��-.~�p�Q/�gmv�nG��V�IB���&�,��HYA:�uٻ��O���?��ʏ�md��\&H�ƜN)���6j��u���mo�0,���E">ߣ�"-��AG�1�F�fcnF��K������z� u�4-^-�AR��Cy�N��^o [11�q���b?�S=4�<`��e�����_�3t�:W*wn�'���g�R˰ B�Ѣ�/�%?	����B����7�}tG]\�>;<�_�|������:5�y�H_;�. ���"eGX!x6���ȕ*"�u%�	����@Ha\��8��]:3U@w�G��o�z�|+���9֥"�u$	�]~�ʝ�V��w�!�67#7}J�:1�A�L��"W_
��=ٔ�7�{�\�9�'`?��!4���z��t��?_Ҷ���iQqP	@�ٙ�C	�=�fzI��.��B��<�L��[��R���T`�w���(���xRcVU��f\z�z���T�����n��\?]c�S+�sH)�ܰ����Tb�)W_��g����q.A��W.��0.�]qI�E�b懲�u(F��ȗ�CM7��wPr}u����e��G V�)5�}8�����!U ��LLL R�f?q~���=s]?V"��,q��QE�$�O�ax�K�=<҈Jau�� `��p��טG�G�v��z�;Y'k�?C
HjŎl�D�IE3nŋg�6;����=��SH3h-�A�Mդ��%BSU>Ħj�?�0i(���#٫���z�%L����3^
zƿx�IU�I����1�Rv�oA+�)�CZAs�zA�n��6��Ӹk-71s��QiJ9̂z��knV��;T��c��qmU�(�KJJ
+l>G�@g�|����{ﹰDs�+��{\a�o��� �#�@;�T6�\-3��>,n1b�����i�; ��JM� �á#):��e�ML~:y�g���i��
�5f��^��)w6E ��:6/D:u��uȻмoc9)aq7a~N�XY����)�WS�9N���5�2bc#�Ԇ��5A�)?�kG���m�t�e;�θ����d�!��(���s�:���'F1��:x����zo�]6�8�3"MGW��#`3��F]������7�$/������eƤ�e Es�����edd�Û���g�G�G�����''lϦ�"�oo t���!8�"K��b�H�y��T��IPP��P�I�w�.��	��h��ѱ�/�Ņ�+��=;ğ �,x~�C�@5���䤗R����8Pz�S��[���E.�RѴ�������s����ɂ�[U^]����gV�=�!������^o�˟#>'v �{�4��))(>��(G-	⭪z�ܰ�v����n��	7�9Jw7�f���o�9V~'W-��F���*�<uy����!-�+-��c���Gm��+)$���Y�l�V�w��v}���gc]�yA������{{�u>�ƈ��<��:*ѫ�#�J[�������"��DЖ'j��e�+��v�mjw��cɉP��	.4ꥸ��pVK�b<�U'b��S
�P��?;o�k'���OACy�� �Ӫ�o���"�lR~=�~hXj��N!i��a]�q��<t5W?hߏIp�gc�}����*eoo?��؜��Ԯ3��!����wHbk;g���2��5����Ejdd�X��F�c���+�-��Ⱪ"� ,v������� �g��tt��Ș_G7�Ck��qn!��)Q~z���Zn�g�9�ɖ���"s��&�*�?47�Z���{v��9,��X�*�WJV��PR�Vq4�E94�9՜�6�{5&��n_�3��~�LO}Z��O\:���{�g�`�C����P�����6��ه|al3�?�^������I������3�;�)�(()_k^C�4�
��*_��OL<���%·r��=�"	D���#Vټ5O��ʘW�ZW�X	`fUU�P�&4K���i�%�E��S�0��s�P�0��:|�L�KK1�9�L,,��by&Tj1.ė��"�d�/�dx)�/�5`�O�/��w�/F
�C�q�_�|��]�u��]H��DT�;xQ`P��T�%��֭4-��Pg�|�0R�2�#:�%��Ӵ�!���I��@�P�,�<9� ������*�O`����b_'�E�b�v�׳��A���k��px��Wcb��d�#��lWUF�6���������>���t�aZ���@A*#�3�}7t��j@)�)��'i�XIz>S3y������1|9�F������� �Jfx��|	D�����*_�>:���h!�j�ܜ������H_�]��;	hq#?o���j��U�N��ʙ���^~�����m�}���E��^����m�
��*�q|���'�����!�&�4����Ҩ�K@��D��ԄԶ�V��.a.��А�4�&]YY��� �A�����z�/	y�K	=�w�B`\8o8*ιIS�TŠ��h9��I�b`r

���!ó@0��rCS��n�9�[ނ���[��B����wO{DV�f��q�]�5DZ�mO��������?KY�	y}��#�r�p���z�mH �����ԤW��VGˀm��8U�s43颰{�K�<���%Yu2%�6+�)�}�FKt��d4|-S����y�����o����^TZt'�$	�R�R��~����^���INj�,W��I:�k��������J��9www�t��[\�1��I�w���\޴�����
AK�5���΀G%�K��|�]j���'c�܉�׫9�4��1~�2�?�91'/n]�|��ɍ͓�c�"��~�iB�Z*|pMsꚟOFbgf���ř��Hl����ǜ@�zhF�|��O�����~I��]�g��x�|`p��]|d$�ڦ*��2��ݫ��@a&�Z��y�;��a��KF�j===�H�9��"��T���'dn[;A��G��Sw=iVx�""$.ŧ��G�6�q�{� �ԩ����JB��7�*ӳ��z@*|i���7�O���p�E-M\
�[��p����������U�5����_ye��VH��[X{�J����oət����\��\̠J��~���4��Ԥz���t\���Z�T�5Q��`E�\9�I�B�+��)��Pq���
��	�B�y��k����&8���'��_��߿�A�W07��eb��/7��e��R��1�DR^F�Z��Kr����/����i?��5�ξR?�"���P52��?�-���p�����!K�9����|��cH�6�
G��pr�'i��Q-�����s���݄uP��=���������J�*�O����55A1�0�����-Z�(�*pЂ�F�}>�b/7בmaa!^�}�s[�P�R󽳲���1�.UO��m��Gf<pB99I��x�4Q���� ���̀�u9�h'��Q�^��_�NiX"3:�����R겙)�޹R�l,w��/]^4��u��(��Y��i&>�ٱ���T��+�
�=���n���_���u��-��ݣ<"r�:������DԤ��qR��G��ח�f���ۖ��A�"��$b��������C�Q��{�0��r�aQ�����.�^�������M���%�[�hh�ɠH;��UMMןS_�"	#ׄ�.(4���75��Y�7(�צ-gfa�n�w_�}F���
��o����Jv/.���BU?�tZ�`��SDCM�p	�J��#�?��wB�w���L
�<|IuKU�re�枸��8�Gd�ڽ	xR�,�BY&4����Gh���7|��'���z����Y��C;'� �	h�+ ���J�=,���>=vL
���I�h����Es|����axw^�Ź�KEh ��&��""�X���(Ɋ��hi+,L��x>�5+��15�:�H��4���̴eZ�(�K%Իܡ���v{qw ��(���%����xH8}Rx~��b�w$[=���cڹ��8��x���u��e:-29�	�O�D�`.��Gr�F�<���C����v	�a>�ԏ8�ډ[�����m�0�\,q��)w?��Y=}J�P��:ڧ׵��q���Ʊɘ�Ɣe�aj�Dj��-���v�����^���t��%c����2˲-SSc���R�V�R�/q�{{1:#&FR���.���Ѥ�{ۦꝲ#,D��3w�Ծ��§�/��aM��^�鬟K�
�`h!��b��O�́���+�3���C˪9[��s8if��j�f�[�I�^�$��F���NN�ߪ�{`�o������ʱq q�J���{�eDR6.&�Q9J��M`[n0.[Xx\���_>�wH��M�&D�_��7�,��^GF~Ө_PzX;����S���eR"5�st$ ��\[Zbj���/�Ё�v��B+�C�KJ�e���mk�n�˻�������Qq\�_-�k⚰�?&���5i�|.Vd�5c]�=^�P����)�J��?��Kّ��?�r\�d�2��!���κqG��v������w@N����F�©�?��d�Ƭ�N��X���N�Q��a��}x��a=�b����3�G8� $�Z��{���,��o�+�d�jM41]U_���6E8B���X(h���
!�����;��jtu-2��d۷�\.(��Pc6\32r[�]3�H���b]hi�!M\�����&�����y��e8'�W���[�j���Q�6]��Vdƃ�a,�4-�����E�t����Z1�>mr9��Z`|�W��Z=���6��a�ݽ�Vʹ�v�c
^JfXS�Q��G�jk'����'���������k�	!�m�z�G����|�����K4G���@@�-�gfޤ��-�<�Icg��.u�پ:H7KqSJ����	l�ņSS? ��'��y�Ȗ1�ħ�
M���Q�,��AZ�w*Ãc�!.������1W::�	��4�[�ir���5�u�NsH�҆��e�)��߳󭕪ܚN��Q�w&r�=�)���Ż�S.��g3�RvR��7�W����UMlC��R�a	_�޹ YcN��<�:�>>��
����Y�|�I����c��{���C��/��r��l��){�n�������JJ�s@���=�i,���!����wh�WU1pr�yvK�b�l͞(�b4c�9�m,A)񇠤�Sb���=:�����L��_�aۆ���!mxl��Q�,�ٟo�ko7дC�)u��q�uSoD_�\��A�����L�Z��K�G��Ӥ�3��͞8i�{mp�3��!���.����i�FC�߭���GЛ����	SP-̾NL��`�Y[�����S�%γ�i,�P�BLX�Ga�E,�g��<a�;Q��Kz7j�n
����v&�5��>���'r�Jڏ4d�G��;+���������;��Y�0�ͅ�l��.e�� �S4�_��ABs����=�C�$G��j�R��c]��mn��"Ɖ��?ؒ�1k�s���dT�҇��AXFW�w\jU�� �=ʼ.�B�!���)v�3O�wS�R	���4u���!���~�H���F�;�/�-�fҁz:�l�$��eirg�_ɺ�0�黹��E"�1�++�"o�^6)6���q�2�Ihw��K�Z6�o
\��Ov__��Gk>�oA��TP�����q|�"�t9��֖��i^���d�d �
�9?CNFF�ɂ����yf�5�Y2���v�-����
��Qp��%��]���=%K���<$P��"��mP'�}� o[�2'כ�Q<lJ��@�k+�c#U��Q����}����S[��.�9�韭G�B����dZ���{]E{ ƭc]M���2�1����Ɯ){+��$�p��Υ�]sK�g�>M�|��b7�r�Z{6�����,��ޕj�+k0{&�HT�%nS��[dbh�����{5�ܾ]H�|� Hc�		�΀�G
G  R�@�x�3	��o<P��Ⱥ[$�,�A�km�"�8�=�����u
�F��+�f>O�f��_�Τ+Z�E���qY����Z,�mjty�**��2�Xo��o �$i��V�q��4���ͅC����i�#v��@d������M���sjc<��m�TP M�r�2���W}~s�ב>�..l�^�H���nj�$$Q�GT(��,���Q���'�޽[}.��B���r@y�MP�������֡q)�Ck��ԋ߿>�x�s�/�@^������;|����Z�e�~���%���f���tk��i.�z�#�y��g�ܿ��{N�e��*�Y2p$�Q'uom?�lè�h9��l�yDV�v��?-P�W0�o�y�=�g�k�YY��a\�Ω�{T'a��k۷�f��k��������p;�����;��;��7B0�C?ڣy�f^�"\@6P%���<s�)��h�Jp0Ć-��ؙK�l|JI1�[q�QW�x;z����>����a0R���-�~G:��gci�©]h�������� �X82uX���%tt��ϥ�o��7�6�g+nR	0�N��MV���NM�rr�f���2uH���~��w|�4���,h}_l���q��qZU����Cp��U����:~'���yOu��'�qq����y���BxJ�J�
?�XwB�?���]O*֏���ww�"|��3�V$��c��a�Jk1�A�����E������9�G]�]GǇ�jh�g�������$G_~1.�~��y�~�R&SD��m����ƀS's�6�jZ#�a��^�"7�h���a�P=�D�ӛ��??D�϶+�SL�{���d�F��<�o�ڱT��ToI��@3u
sͫ+�N䮑�f��,�Mcޝ��u��C�|��\Q���D����x���� b�f:�RO摢���3/�����ǎ���� Y5uO�Cި�g���c�����j����WUz�ȿ���|�����=z�(� �=[n��i�{�9x���߆\k��-H���r&�*S�ۏ&YL�<Q ��g�@2��`n@��:��fk[�:�xo�[�� �2�@D	�v��DY5�3 � �[b���h\4⏿"�H�Oh�
��V�S��(��σ@u.�8R�E6W�#��lE���Z�<�ԕ6^L�&��[9�zPS]���ƺ�\��)�ᑾ�7�߿ �{>���s��(!5�BjiϠ8�iVAABq��"x.9����n�a�[^î�Ы���\����N�����_"�O�C��$�F����%�myNz�70���J�a���������m<`�'KꖜL�{���r'�fwq�K��=�SIA
�~�5��u%>~4�7;ED�=#qhA�l�G���2Vf�����yP�ŉT~�ٛ��ba�"/¸|~�x�27���������i*)�6ݻpx�_Dd��ߎ;�WZS�H�LEI
 �@u_������*��2z�J��������	zu������Y&��C����L����E,�^��Ϧc���h/t6kd��ODD�r���(�f.�?~֠iĐSM��Q���hypȽ���,i%V��-���E��B�O������?z��J42.���j���i�x��@]>��h[^�r�����Z�q�1���18��0�ԮZfA&��Q���1)eX���*��G��d�UWjN��1'�yv�RW�ć`q���iI�CK�m�|+�X���
4 !vf8-�����m$j��)�f��-Ⱦ>T��}���Q)��[B8_J��4�qy��{�[6@�p8�l�{}���@�uzZZ[cVۚ'��%��֘��̿�����k����CH8ۋ��Z����73o� ]���6��Hj)����Xeq����~N���q�K�<��QFbAE�{�����M.��O>���W���혤����9�A�-x���A�O��$�#X��=�V��;zs8����h������g_�:�)��J��E�yU��<+��e���"_3ss)WJh�M�"����y�!3�%��aSo�
�.�`�{}ccg�T�*]��ڄ%�#;੟H�bG���nK���:1�|�o�3�*�Y�#�|�	���j*�55Qj��徛�A3�2v�Z�q���J�<$�,��Z��ӳĜ�$�:�K��ۇ�Kfeo��W�Pu��1��7K\���d�9��߹���ڗM����������J�:��O���N\�d|����Yk����UP�z^!�F�lsII�L�97�N���֏Q�u�.2&;��ɒ���}�N�8yc!�\��O]���%d��q8{ߏ��K0� ��Ͷ6��&�>�����W76�_�/vw+|�x�Μ��A�DW_�H�ΨN!iG�z�9
51����Qg.LZ���������˱tM�G��J�[8~j��N�*S�}�<��≵�!�؆�*F��u���x��	D�2�B#�������^2��]���h����?7ܤ�-I�8/�{D<�4�������^��F��%p��x͈{;����[|��	?M��T�����v+��������=����P�L���oxXl}*�E-·��Ts7��0(�)?y���t��rr~�c���&��3�]\�i�aw�}*/O���7N&��_�� ��X��jl��3U������d�v�a�g��������c��rܷ���%��h����bB�I}�>�0y��r��!s�/��WnG>G����|��x�G�?y�h��Z�}uHH/���������~7��{�M���kb+ѻD�ND�-D����G��-�[�&�FD�D�[��}�s�8�e<c<�^�Zs^�k��ֺM��$W�PM[���������[g4 ������kt�6�9�����cOψ�h�h�\��@'�)tR�X�if�7X2,N�+p�c��� Y^C��Wޓ��i�^)H�[Ě��	x���ѡ��(9��(�7�74pm�\���n�R�$�~������Iz�|���_�����X:
!qJ�J��,֏��2V����Pm̘k۸!f�Y���̾��!��I�L W�Ұ�S��b��I�Ќ���dM��{�:=������`�k�X�Ew,';�Qx��
��@��W�KH`��D#�d;��#L��C�Q��s;�󬽋��gZ�z�3n�8�3I�;�1;�mW>?��R�^��$�"i��pK���t��QSW����J�����q"�6+*<Z'l��`e���0���q���\��ҙ�T���G&�(ǒ[RUђ(�Ճ&ߔX��U�� -��iN�\ނ���S��b�੼`��SD�c�*"G��R�c�T�h�ݦד�ԒI&~����nlz�y���G�t���h�xң���*ݘǔb���tGg]�������#����o�v��7ˡsT�e�sM+ӌ�����ҧa��{w�'�N�bï�I6���i1��c���/�F��N~=���Kx8�?A�T �����l�������ߗ�`�+�~����;���[y�+���g��"ECz2��/��������)1�SY䐺�o~��O�}��פ�xd�z�������=̽9~����A����:��ݝ���L.o�9i�O�vk�u.�8�xB��1�R��8@���ˌ[M�J?W%:�6@7�MM��*/��:�5�7�-Gj��9({s;�'����݄;֙������M��4�i�i+�hiU���-���X�'IQ3j�HQ�i�c���:�[c/���7� Ij�c���L+0�ؐ.�0v��T3��]x������s�Qӓ����^+�Sh��s6gf�Dn�N���,�]xe�Dal<�rtûYLra�� ���K�}��`x��<�����gP��F�jλ�m�{��AKX���P�{Ѧ�
��GV0i.m���Ğm4��6��f5 s��Zl���][�O����8����ո����� 
7�;:�:��s�tv�y��of��uv�*�Sz7.�#�:C�,�u.�<oSsQE��� ����LK6GD,K�ᐓ��:�;��R6g����\����5�z�.�/�~^9mv}ƙ��ӥ�T�@����t���Cf�A�â�����6*[���mEYs󏉷oΆ����}�l6���K��5�]k�O]b�?{����oZ�q�2p�	������T��h���'�j�v^�O��2xJd���@����47�U<~2i~�C���F�lU��J��Q{�VI�u~�FSk��t�t�uG�=)�����d��X�O3H:�݄�/Da�
���� R�D5��8Gt�H�Я���\9����-��L�L����;��}!��  sQ�oJ��=up���%��2�����w� ���T�؊ê�v;��9��~��������2���=����h�`���)Ѐ��k�vt\|<Q9ɫ�;/X�xn��xkr7�G��w�I3yJ�N	K�n�
N(L��q4OM���Sl���Č��[D��� �CN�!~fi��֚4ɞ����A�AΛ�Ɗ2���c��K<�
�XJ("��v�g�t�i�f�7c4y��$U�{�/fc�S��#T�W� �g�=֋m�10pG2��_ں���NM�$���%���D�n�w4�8������QJ��ȵ�c���B��|4PȷX�|�& ԡ� #���3�9u�����?Db��_��~&� �r���I*Y�ʊ��9W#���E��n���S�Rn'��N�k�f�����P��v������$_�W�D/���0�8[�x���c5�59�Td��Ԇ��anT�v����?���ha��s�zn,z��D��x��S(ӋFP����jUlf�|�###�����>Ûvu���y�v��ؚi�-�h*?���*fi>7�V��m8����a���;�[�%bP�Ҹ��W__�R �8���p����$�}#������*�4UD�L��`Y� �B�s��M�"����[�q�KȰ��As��bX��N�EG����K�Y(p?�����۲�ɂR)�, ;"���T|D�]�?Bp�V��U�EI	7�����?�@������/��ݓ��񕑕%̶x��񫑒vY))�� m���yx�vɓ��z��쑹�t���M )�]���/fFFK��R��I�����F|��E���~s�aċP�b��~EZjꗓ��
�����=���]�)g�o�ɉ	n	F/|�r� z���o+[gm���1M�cR�׼���w�&����F�}c��!���{��+,b���e��hN�ui�B!G����F�Cz�<�C�J@��D�2��>(����h����$'�Dm@�paa�=Y�Jc�	r�O	―~����1p��C��b0KVỈw��y^��������m�[�����Q�S�o��_]�Q`5�I��r6�:�ƗL���M��3�CJ�W$������?�r��1�G�<%��lu�q榕������sˮ&!��s� ���h ��ö�N0)_�$e}5h�G��dN���X;n>.p���]����41���׵��CJ�vE���///O���q�& ��Z4�a�n0����~�@@�����G;�=]�;�>i�B� �s�������N��_NL�Ȱ��P|�*G�o���*-�x'CF^&�-������f�b����/�bwd�wvh�<2��-��rۿ�Zߊ83H0���<�9�`��0���І�~=��wvt�֗N�s�$��Ls;l1�7|������#�T{X��5�ʓ��i6�D�H���5	�M��ޅ�����`��KX�jq�u@�+���P�O6$%(i:��n	8|����ǜ+f�v�u׆�䤘����nm�n���z�#���~����
��+n����䎊�''��ι�{y�F���9�&�]X�v�W
�0 ?b�(�
���`A�W#Uo3*�ڪ:�DSK4�J{&�sx������wu���k$��ro��h��w��z���	H��:�ߗz,�� �$6��H<�>ʴ����r��!&�Ud�%���Q0�oo��آZPa���C�1�`r򉘌��-�p�q���l���ߗE~o�|�<�Ё4ޣݗRCSs�I$���o�|�3��V�XV�wK�4�j(e���u���H&��Y�n��}7퐊�.�R�#�}c�v^!:�8}����8�&�e4Ի�o�m�U��B��-T�"Uoc��(�LIM}�N�]a��[*���fff���)
p�nˑ��I*
R�s#��$LR/
K�_��,�� ����� �)�c�QC#N�"
,��"�S]s�3����Xݒ�nnx̴_�'_D-K�����ˌ��2?�6*�?k�h,$*:W���߽0`�C�mF����G�9�]�pg��A���۫������j�G�s��B��Nea��r��%��M��D>޷
t�FmH�c�ٱ�{ˌ� ���T�v���У����cct �������L[s����s�Ƅ��yU�{&�]|]
�]�����@�K8��1\�oW�`.��������lL�b�W��g�M�
��hL>c#G�r��{'�JJ��h���7u=�o�\��x�,���/XD����=�#��˳&���M7*ߥXMx�HC�"�g�T��ERcF����|���w���T���U��夘e*���R��a��C��]ϦnB�	'�y�4�_Ic���K�x�4b�/95�'w�-ڀmLΑ����&1X�j`�#>���ޜ~�ez�K}��%�B�b��ȵ��(��^�(�_�'�ݹS��������B��`T:@{	�g��Z�0R�im�C��sg
��c������` ���@����#O���m�(.(����|�nEz��*�6f�/�v�~��~���������M�Q�����KV�;+*�x20�?�&0��Iʗ=X�n�j�罯��,���Ƌ��1՘R)�ć��>��ݳR"溔��(���R�O4>��2�Kd��~c��a#�fUX͊�?'�ޡ9܁daN��r2a��4���C�� �{ﮩ}.���v�9~G���?�;"�+-�S�C�Qp��,��C����o��k(2��ܸ��}�]x������cMr�?��l�G�?VZl0��ueD]S��\��e�փ�P���W�O;/5Wd#����7..��IH��eE����>�ԕ��nN7��+x>�|�{|o����h�ܵ���w�ܡֳtY٧k��s8;{�W��H��԰"�r�{��+1�B<D"Fi�?�*�:z{���m�}�-|0բ��ՑZW�\�%�m\&�ø
D*�4��kN����G��i�=�f-�:5�$ҳS�S���y/�B�9���c) |�bꂕw��/߿���8�:
��XQ�\V��MHȓ{`�������S�����ݫ����C+)���&t���u/���M�UKo�Ͽ�����(��~l�ٮz7�n�����ѳ�f;&{�+Ū���9�(�okk�5�1���VEߋ�^���z7�Y�8[���3��140j�G4d	P��^��w��XG������S5�����EҨ�1�$_cF�d����?Ժ6���{�Ux7|å��^�5`����X����[�ty�4��݄���_Ye����J�.?���,z��h m%����%1qq2�t;��¢9�]��55���"��b�?~�4�6$�b�^�����rQ�~_~#3)A?�r�Vf��2	/t�֗���M�놡�YX�4z�X��RT�	HcTrXD�o����p>�t'zIN�wǗ����`�PlZ��@)$�3ٹw� *���O�	�nl����������\m��^����rj}dXD���Ѷ �x{pfs�$�[$i���ݱm��O�Ē��ɔ�����Q�m���'�,��Ճ�����x	ʣ�?JP�y�|wЀ��yڽ5({��q0(��r�ǀ��H�hH�PkC��1�=+���ߋ����[8[ϱ�ttH��#E)�0�G|��= �,W���y����=���}���~Q������*�r�֒$��Zq8�Q�H�\L��e�l���8�"$�5�ހ�������f"�����:�o�1',�I|������n���O�%�_+�3�Q����;G�������
!A��d�>��74"O=<���y���ku�'p%�/{JDQ�_NS��8�7_��h�=1y�@�q�w�Z�� �Y>�g�s9��%`�Y���<mYW��P�/Y����T���ҽT�5��
��~�G	A��8��߅_=�4q���]�ϧor���i0�[LU)x1�{��S33���jf��^�6��مȈ�uG���C�/+#K�z5�Տ��K��v�Q����-���������vՕ�R���GU`��ݗ����>�vc1Ak�)o�'�58�I��ͤt]�c{܇��!��4�.H%r'���G�@2����[��o�����۳��
��Y�Y�$��kbt��R��{q� $SU���m���mւ�rr�o�%%p�o���^Xu��4�����z!��[��-��-:%��2���:��=�+�{�h_���B�3��%m� "66�~�\=3���s$�Cb�O7��l�SA�~�׳[����oI�Q�JF?^�Y�����"�6M�\���L��省���y����j��j�d)! ���O}��j�沆������cuEʉ���"�5��|�[�Tnk i?���k��^��o�ς���[&�vg[q��Hh��#�k���MiR4#C�i�-2�EW���	��@w�<�J�h����\%��s�$L[����[y�BO4���u�ws���3���U���@j=�����S�Q�/�223#���&z�y���XH1/I)(�q�»B���#��������ZL+�C�|�)4`f���')�R'���XG>�ծ'p8X��֎|���_z�M�H��}� ��뇕�=�i�T�Y�8V=%�(��g��ZEt�C����ͤa�:�S�G`a\V���pK1/4/O>��8u�W�;ZW�{Pt6�F��}0~7�¦mgxuF��k����+���I�8�NNq��Oc�����eC����n�z��?{��x �\%��z�
�J��ٔ�	�]�*�����`�i�,�dƧ���ؒ��f�ݮ��b���|�#�"�B�1�0���S|D��:Q+&�p�K��J�v�}����Nʫ���/�6�.��pz�ϝL V���{��cw�fׯm�۲ӼO�W�qk�uqm�C#�휭����P����`��-鬟�������+<��8
�����JJf�-U�0���<Pd �&F�}��mr�����D	�~��f8n9������1�V'�n�W�i��UZ�!6��K<s �d(v󎌈�>��YX���u7�P��^6�@�^�>$�B��b�H \�����CCP�!u��E��,�kk��YV;�|�:(TT�	�:��íYaM���'zt�--����q�zh��SB��'�ij�U�?;�׷�+�
��Dh �xJ�-����	r�4��+I�3*�A5|��!��5aDR�H�����~r K2������9����Y���k���XŐӁF �f9|�č��Rvl�e�0/hB�����ID����a�ũ���	Z���S��Sx�V�-62���2�� '�=�4y؏��H�T��_�3�p.�B����4t�z�V���.3��O�]�����Z�I�Ν�¦�4�w��D�B�w$4��'(��j�"�5=�K7�^��$��9���ǾvW�w��ty��E�(U��JGĬx7;1�B����5K��؁����G�`�g��@.�ly"�yJCc�\�yfFoa���|�nD��/�.�F.GQ�&+~�P�:�X��|���j�Wpp���Ы.2$\{1��(9L/U��3.����W��O�+X#��B�*D��S������x&�ge-��n�<5��ǋ�>Zƴ4��Y��L��0��i3�)P���5D�^B��@Ϣ=�Gf�l,�|�.�VbB"*��^�vͅ]~S��?���2��@�f�оѿ{$�e�߇�BC?��k�|�y��[������^�4����Z�0�W�&-Q~_K�U�K���Gcﯛ��M� ��D�4��qr�7�\�^��O���@(��H��쬼D��}�+�$�srq���h)Ҝ�;S�^�,r*�8ON�Ґ���"���{�ѵ�7߬�A%��-#�������\{k����Ɋa� ��`�3ӌ��8��~ro[Ú���bZݣ�����6�>�FYޝ�>�RT{j����Wȁ��!�'� r?��v%�$r���L��F��*�m�z!Q�����7���������(�)��V#.J+oo��B���ӧ#�Q��W�%�ۺ�?�>�����ke�F\||�_���֐�ŚlAK���Hd�Z!oi,"kPX�k�O�������F�
��n�@b���=���J�SĪ�ȭ�����D8���g��(F
9��[�v0}�&�����mё����G?��*Ddk4��(e���3�Hd�f�w�9<�m�PX� U>�;a��Y��ΐL�@6z�H/A���$��K��B�Y/'��W�b�=��R��mR���M����V��Q�ּ�?����0��;��ڧ���~�7�aig�d\_�OC��W��ŗ����n	��Gc���X�����(5~�D�b~&X$65��FWN;�阱|j������QP��f��vr6�/�{�Y e�2g�}Nh���c��G1������z��m���u��4��«��e��z;7N|~������ U�mF��4���Q読��j�A���3J~��t�u� ����(���o/":��#N���
E�T	dNxP����WRP�GO_���MW���{m��X
p��U�O���tq���ɡ}�7�/X�J1A�#�������s�ef��I7�F�u�&þ�c2�sw��������:5���:���O>�(%���Cc�SdF�������Y�D���1ǺR@}#�����JJ����@���d���[M�^(�Sfo?��ini��O�͝\D@EPh;��]��[�_J�Y���\��'O҆��N��q�a���D������u�ua�K�� #�Ao��| ����l�	x�]�W䙶02����Ä�z�-i�F>%6��"�y>r�3�v���(;t��?k~|#�V�5��H��L��8u\_6pR�^9ZU��	؛�,�J��sQ��� [���>Lѩ�&,6����&ѵ�����u�ۦI��l�P}�	Ѱ�M����*eY�nxߪ4�kV�ٚ	B�	 ez���@%��$:����D7��t�nnH+�܈:u�5?j�ĸb���N� �ؓ�?h&!Ē+�7e���B�ofvU�!)� ���f�'q��v�y����PoZ����E��޷� ������ö`�Rt.�q��a����?��8�����|t��|g�g�f^���3Ms�$H�<����D	Q~�=ܼ�C���
m֍�y�e��4��@�)��=��-),�ظ���b�@�B:�cR��w��G!#+��������4O;IX�u2h�_��%�ܖr����=��OMJ��7�y�ɋ�J���Ò��v��6����4ޞ�FA�<s�*;þ/����>���k�R@��p2����'wN�lLC��])Z�`�F4�?wd�^�90� u����m��>�#{�4E#k����&��֗����ﰰ �_�pU)��77#֦�E3e���ð���ŉ	r4�_�z	Ҵ����pd�M��5o����M@��ܱ��(ƨ��H�_T䢬���~�/�/�Ș�2ܔ]k�9���J��-kW���Û�T��rE��>o��J�q��� ���L�UkAj�xziY��I�q�q��vG#��lm��%hy��s5�d�}ҭ����o l����%&Z��0�E���xfvV��*lA�#��Q��`:�	y�e�h��U>�����V mTP�$w�E��-�rj@�Z�(�O�;�Id���֯8d*�ӱ�[TK�waU�_|C��G�]�����1�0)F�J�;��&�c��]�ȑ}��Mr��J2*��d��c����h��"�,2fc\�P���'��<����#����R���&+\��桻dm��kS)�J�����O�s��@��JV�o��>�D/8�������ml���{s����^�p��eD��9�W�u?u��f�tÛ�<�?p�<��y�81����*7�k���rȠ���x���f�3���]�kH���,�r��XJt	��	����������A�e���ɴ�B���Psv!�N�	�DOg=��g�̏�����䒃T�J�f��������x��g��U]��E(��o0�D<q���GF(�F"���2||�Q�r�O� J�D�g���$%{�j9��0�l�c�\Ůէ	`Aً�O9a�YK�.�*7!�KD#�����&��e�3h�إ��r".̾[��EQaa7�w����	6
��K[�At��e�����i�=?Xɚt��᝚�W���ec��ϣ������A/��HJJ�Tļ�޸��"d��=��߁;PO?�I��P��,js-��I��AX�Է�s�.��KJ����oƿ��wz����	��%i̾�� C_��hr%(�w��/��4�EE��@A��&�:𷸟����P�k_�t�2�I6�&�۲#���9$+{6!#�;W�󕡭�<T�'X�hX����H5	�$�dL�}�8�F�����q�k�|�:��S��j�h�_hQ�gӻ���@��~${t��������\ah+�`�U�������;��5O	1�q����k�?�D~i�V�}_|K���߇e�|i���XevKmaG�܆�vב���<��GG�}}�I�R6&i���ڶ���:�y`����@�A�@g)2��lo��2W��qUm�X�o2�b�h��.ہ�R��>G���
���#�~��}R$K6�am@sc>�*Ж�OM��7��(�I&7T����X]-=2�	KQ���쥆n�GZ�q$v��$4�1ęu��R^��G�c ���sB3�{Cպ�n1	�X��N�}�%��L.�q>��b����N0�����lY��ɨ����e�^G|����c��E�n_(��aUb_�"�R=	����fc�O�f��34�FmHc[]ň���QKMyz:>.9�=���8�>|Q�P�7��U{�-}gb�{��nM[񊹻�K|{<Y���#�����oT�q�MO3�S؂�J��$`�����]19>R�c��`�L}����,�`�'�/�#+��G����^4>mfDf�5�.g���Œ"h]E�l�OE����f�5aqP$,�j �6úc����S�Y:6)������<I�o�;9:����4�!�WC8�f���?/i�ˤwG�Y��Tq�/`0�s�=_)߳����i煱2��oi�s�@���G<e�	|Y����}�r��`��MWW���z	�ck^n*+SSR�|�
T���Ǎ'/4x��^����O�t~�|V�q���ɞ�q+9�*�a����Gl�������!��=�fW����@�c)y9n�N�u/�0@� �G7�|��m������QǺ�k�Ƽ���B)� ���Lѫ��Xc_�g�0��fY��|)�&��w���3;v�p�*�p�^m!�,��J�]o:�����Xw�l/�Ј��� �y�>�N�ƕuk�%�S8MAs��{�Yf�WNBП��������KSb��^���M��MO�Ɂ��ŝ}�?�����H5G���$+:ÿ��P6���Dr�2z��ѐBw0���A(a�\ ��V��c]*���/��:	�b:%��t$�s�x둝����\�;�U��G���߁��y�������!�'7�\��fh#Q[��ve��j�!ܦc�h�ʲG��D��	�����)]I»\��������`��ә��nړY߾ 0�96i����I�R���tE ҥ�� 4T�a[�+XR� �(IѲ��㣵����8����"�e��C-��5���e3l�k�Muj4�����cy97tcek�I4O.3ytOէO�w(	�$$>]y��91IIa������P��tшA�c##jNb�+c	�ˀV]���|��^�S"�� y�`=S�z�w�_�٩��</u�B�)�K�2K=��'n0���:�:��.8��"�΃���f:�j@n���?P�L��H�����C[[�w�<24��'�D��2��xY׮&�xD"ɝ�%�;67~A�̠%�=��y�8���I��Iu764tLֻ�B}��Ы�A3���@�,��pȊ��Y��DƣǏ�
Y��m��댾_��Yɦ��r�^g!��T����265�Ao[���4�iD.�t�O�(P������C�RN��#�~�Z����4�$�P�o�V"���m�"`rg÷bw��1��!�-u:Z͵��#�/#1��{f������I/0���5�qm|u�K&��_�� ���?�E�����A�.�Zk��ң�#�`�)�YC�6����5�>4����x����,66��"�B*�Ĥ��+"��Oq����t����t�%���7� "	a�MEZ���!���T�5)$���=��10��z���Nߥ�����tm�֪����p�Yォ(_����^v�ڄh��ީ�:�EІw���pQ�������*>�|�߶ߍ��FT���5X<���H�`���J�k����?:~ed<��Y�%��?0�3ߤ��rlL�0�yt���������] �?j�|[�w&6I�,Щ�g�O�dH���0�)O�)>��0�����g��8p5DRC������3�:x�h�/p����aqnBC?� �ߊ�/z��~ YJ��J�����:��u�#"���<�.K�(��cZMI�Lc�ZN\[AT嵭����
,C��<=��c�{��xn&9o.7u�2BY���\4�����?_`#�ɑH�cBa�^QwZ��3[r?:_��*�1�<��f�7g�}�k`YRn�����{lB�1�m�.�w�L��l�h��9�V�@���
[�a����lƸ�����G؛��楒�]\2���4�4H���-%��_�񃢑���"riO�bJ}޻9��S`�<�ώӞyy�$����A	�i��=%v�v(�S����]f�ꊡ�2�޳gϢX%���t����*�\\����p5-X���s���^`P�,}T��fZ�)�x��������qz�x�5pS��|��1��������� %C�	: ^�v9������=��l2��--�2����칛�y����C��Q~\}���ǚ�9<����t���������q����h�>������1|��
���^� *x�T���D+�M��^ sO����������(���j��k��{JM��@] �d������ma���XX�;�;������A�]��r ,�oơ�(��T�?��`7�+6������1A'Z	�M�G&��2!��{û�K�^M��u�v7%�+�gk�����]�ul�z=��Mz�R�v�<Ffzu5�w���>̴�N[��D*�c}=����%yk *gs
��\_w�^#�����Au�io7fNN��K2Y$��"���PM��k� נK���N�+�	�-��M>dުC�tDP&��餫�¨=B��ˣD�Ք��'���>��ݓP��P�]�]��Cm��kfC$Wm��c���(�q�z�o"�ڍ�<������l��Au� �aSkJ�Xaaủ�cyc+#ǁ�;[�e��h0Y:���Ι��d�7����"ꊇ��)�[�R<��3��ܙ��\�:����o�r6�A���n�����}�t<��'���
�hܮ��������g+P��x�5/ҚL����,�s��cwH7/�Ytd��0T`oH�b�|^�4O�\�N%�J��<���G{�\Z�6sMU��6n+����N"VPK�l{v���ɶN*�_1^.��(+J&)�kɪ����;�������n�qA9�p��]E�Ũ����⏬��}4�R����wa!!����5��@�h��E��z�A�E�3wnj4���L�Q�b�?��ገP#��D�g���w?v���y+BR������uT���Ń�X%_,��������3�v��?����h�N���Ŷ��1���p7/���NP�B���5�#�WQN��D��ߜ���2�B��y-�����'zT&h{ěۤ�r�N�-k4����y�[� � 1~�/�7ʾPc㪴}��"H��R��A^Us��.G"�^ ��=�:#�	��uV�Þ�2�T~�t��簳,�0�d��uLE�F�F�[���wI�(�(�����r��� �F�u��he:k��8�O25/!KN3�{�n���>2K�g���|ӿS-������1�^��6wת^�M��>�O�^k��,=��i��Ͼ��}?�H�@�~����GxW�����2�hr#{�1�)���^I�<Ylm���fXN!&��"�����Τx�=u�%.�9�k�Q����Qd���C���F�r�����Ų��>Ǌ�[�e2�����D��]s�,I��W~��Hw��7�����)$@�0�)�TF�����[
!�}���F�N	���R����tO���waŶ��"I�:Pu6�w���p���>��l8+��M�*�+=+9�i~-����;��Bf^2�a�%������V���iNS�9�i��ޞ����Z�x�"�IKQ�e��M�͆���1�ԮEnb�yЩU3x����HZ�ظ�,�n�d�FE��E�v�V��IC��T ����l���O}��7���Z�N�x��W��8�k{v!�<_8����wP)�C;��BT�P�Z-���ocǵ�ܓ3NJ�=��7�p��D��V~�,	���w,Z�����{0/�O낱|��������<{6G��	&��(f�������6�C�ze��H�%�FR"< ������A[��b���U��7���j�y�����ꌨ���n�z�!E;~�/)�e�������|��y���,��ȭ��$~k��w���h������zM�H�^�H\yH�gU�UX8J�i�:�lH�do�r����/�F�.��s�_�wͿ��7��:�v�c��i�4�O�#��~�?���](%~:���#t�w��;��]܄�K���#/�4.ѿ��Fq#U�[W8�����5Qq�}��M/'�1t�l����g�wN�#����vv�3�"Vӓ���/+F7㙤�I��x�����K�[9�����,>B������3�3m��f��;����W��:{� OV��k�z�O��Z�j���� 0QK�I�#�+&��όX2����70x��YnҸ�J0Yz���қ�a4�C[�.�;*��'�A"de8(2 �($�nOk h�'���t�P:�����₠/FO�M��s���)��6����eNsN���H�+����t �Un�{���4��[�u�o � <�����Կr�/ٰ"%#��ޏk�`Mo��ӀO�Bwq�,�����"�s�-ػ��赜�MA�J&�d	I`8�X��ӗ�1��5�p6}�0t�`�ÎO�7R�#}�(����K�(Ⱦ��
ߴut$���'�,�FWXD���e{��}�v ��ᆔ�L�@�����B\l\�����֡����q}}}u��hccc�'����˽}}Y<I�s;��p*���8��,�%R�D-�;� ��i>�5��@��Nwx:��J��772�����B�xS[�����$�3��_H�t�&p�y?��Rґ��qo��~m4�y��#}̨@�S��PB�]dn�q6���)��� ���x�iF���<#�C���2�_��W�'���2�����W�t�ᓌ��LNN��>���b��[��YjF��-�V���զ��t��k��i�s�*�6�r���Śbz@oN��
8�T@k&��d�j��XN8GwB.�>-���umb
;
�,�:bSJ}�֡=�;�+��0�Ww�T%�*ec���}�!���Df���[���/�3R��9���W�vu�:����ۋ@�N#Z�fڂ�4<�q֔����|��*�QP`5	���Ҿl&H�ΐѕ�J��Z��'x��]'��(0��Ug)�A�=�n%����D_!+������0-U���N�E��,̥��L{s�?�9����tm89e�Z��5!%�,!�<�dl��b�X������u��^ǳV��w����X��c�'j5X쫙�����?^;C��䣷�W�x�o-����(_JA�f�����a�`Rؘ����ޖa�־�!�X��:�`���R�*�jEB��5�I�6"��n�x���7g�,CB��&��*��X��##���+82��MI����`F�'���nQK�,G�z8q���D��7t�-�v����űc���}�(�7n��R�#���o`�>imj?�����y�d��T�̵�~��y�J��g%z��^��J S�C^�9Z�~$��"��2�1w`te,��Q�Va�3�a�x�3X%��}r2iU#{��&��>$�C�cza�����ǁ��7��
jV��S�X)	�lY���;�K��
ᔕ����s���p~I��X��mk�vP��20@�������P3u�?���.nQ ��I��Hcy&��	:;"2���փX��ӧ�u���r,-��r�\��cS Y9�"����1��J��7�'7��������Ve]۶q*jB�@�|��*ҋ�r#����%h���\2���� 2Z�ɵDi׿@'��Q��¹�lYkW]3�c�����'w�Ѩ5/�Ҿ���G>U��;�J<�^��RcKӗM&��Д�Ԃv��>�/kJ��eΤD{M9�&�~,/!�T����/��`4q�p]��R��o��J���gn:�:D�(�=����C���&Ly�Id�����^��O��$�f�hL��}k��=W�,)\�	lT �db�%Qw�{\�|�=�s"�4����Q=?z3��Dz ��GC�6���K9k�6d���wH�c>��$ߒ>s@�OMA	�^�h䫮&#Ŗ�����~/i5
������W8G���pI5�����<E�i-"ݶ6Ҡ��E�wˮDV�Û�ßX�p?��K�4���]�5��-F~�mF��G#5<�ڂ��b�#)���-s� ��Y���o:���5�J��iSG�b	��D�u�Hd�`�#c�bz��޴*����Y掩)�E�:��A�pF	O����L���==�P�!�����$@R�L���TdUӟ��L�f�H�ݞ�ꩍt�^��(C�p�;�W�`
�Q ��3�C�U@���[��tK��'�n���&j��sGDH�ކ]�v����p��N�$�;�Ǚ�\_7��N��&40�S�R�Ew��-�`�^8�|�~�Att�H�����r���ǖ�-��-5����iz�e7����JY�r0=?{�#	�EU|�=����H��wz�MC�m�a����!��v��3ц'�v�M$�R#�<I��M�	߬>^v+wqt���������/�|��XX�.JS�e���@ݱ ����hAV̻T�P�l��.q:,|TY�����ܕE�N����)R���{�=��5�W%�n?�)QZ�����}��m�'�NQVv����ݦ�蕍XE��\	���<��k;m��4� ��]YbɄ�盽B��l1a���J�R�E����dx�[�i���%B��V�)��G���ל�.�g~�e9�xIH_��}��d�__�"v�Fu�#�X8��q��w\LU�����G��1Ҙd�\��F_@p%Y��x���k(��Qy�8kr��	�)��7S[݉7�]aʟ$2���P�5���Pu��T���?""�ұ�U�8٣8�3#9��(�H������22BV6�J��3�w����?~�[�ԍӹ���|<��u]�Wγ�ַ�<ob'�vF+� �m�<�k���R��@ʝ�:����"\Cګs�7r�X���*C.6�fN�� y��l}�:�IO�S�2o����R��F!��ռ��Q@F⊐�u9#��F���hV�h.�K
0Y����V�)�V5�_����%��O��3t͏t��q<ڪY=��c�#��-��gX1���V��w��P��2�����+Ȼ�z�	�>벢��z�����[��I�3��{@{څF��\�(�I���y����VYuh�����8��l����J�Zg+^��_X�1��_= �
2~�D��b�A|�̢�[�յv�$)�ӬXOㆉx<w��e��)�4+��e������W���uiV���[&u���Ra�=,{(���'jl�Qe���kn� �������%ý�%�t�ЙtޘC�ﰹ�z�,#ic�73�u*��e�-Йtv�!ǝ�q]8I��L�F��v�ߑ��y��C�E�����6�P����4�Y��W����)",��L��t�Y?��[!�$����y�s�8��Wj�]���6�њ���RKU6zѫ.e�)}�M���ڕs��X��/�;}� V������m�߿�KN�=緍Cb/�fЍ�D�_I}x��K��J�i�y���tŘ�dt����)�S�*f�G�-܄���P�^+�u�o ��;��X�$������#W�-�$�����͹�\���;.���ƺV��٬����z�/����"��4*����$լ[n�X��h����Ak��F�?KV�!�q'1���P�+��*C�"��r�6�����2Z�� {�cc��s!V�OB?h�1��I/�#��}d3�/g�`3��N�-��;ԏ�N.��E��a �$k�t���R>���Y��1�2}X�W��z�&A���ѯ������tҴsmOr�fi+V�^�B"r���ik�ZHɩ]*���;#�~�GS`�swY-;mHd���L��d���n5�Z��=[[(벛y�>,,�X%]��q����[y����irE���ٽc���9��hJ¿ou��b�Ƴ�m�c�
��z.V$��~�D���Q�(�F+��y\
H�X3����{0��p�Ha�snW���h7���	G��Ɍ�0hJ!
j{��_}D���f�<��f
�V�s�E�<��u/^�3��o����:u�}�����U��ޑߏ��t-�+�=�'�ҿ������d;-����n�9:�yR�뗗��Dk�+�ѧ�+$#���D$�j�Я)7���dYu��nq����W�A�VF�-+���cP/���9;\�S%j���|���&�Y�?�X�O3a���'ߗ�I�057o����6e����}�n�JnM�� ZG�	T�/�Ɍx�F�3�4�fOڀq�(n���#�5<��$�F�k��~��+iLV�W�����V\;�)K{:;-����z� ���`��QF��u��3 ������ɝ�o�$����t���d�'hTX��nI���δ��� ���]�����GT���O7���M���5�|3����; ��<)�S��{���u�2��nթ�l	�����s��|��&��T��;����j���L����ҫ/�2���	�ͭ&R �����+#��x�e����ڢK0͊�b����T��h�K+PI��S�4�׀|�)���"�m/1�H�`��%�>�_�㭮hg�I��klW��I�ۅ`��@�S�ݢC8��N�o���m���L�?�������{!�Ҁ�z����\\:	�q��f%��ȶr���]CP�.���!�0	��&$\6�k� �7up$J�׉��Y�����'�`.�����gS��%�'��2��?�D��N�Y?���H���?;?������m/��G�)��X�ʱϏn��]�b�|)�}��~��E��v٤����c���+��F%#����i����ۮ�!�I<�h���5N\vְ�>D�P�z_���B8%�eM�;�����r2Q=6�0��}	+8x��QGl�`u���NB�͗�	>&˘��A~ͱ��Ԟ���y�X��e�]i�jo�G�[*��-π�a�������4tZ̪��R�-^�����̩y��G���M�B���ʂ�Z}aa�l�w����e�n����'��J�C���H$�TAg^�]�~��5@w���H������w�sN�/�L��"ږ��iپ��z�7����3��^i���H�2�.��aD�t��#�ҟ"��k�4}�E㕡��7PI�
5f�H�G���!�W�/��Hר`g,�������hX�=*������V�hc)�F��_�grgU-����&k�1�{�	$iؽ��3�0i/W/`���r�C�4���A���&� �0���V��3ir۬|�@����Is\o��T���3�6�$�'��rzl�X��8u|��߰��NE}�
�n���2wK�Jt@�+�3\���쯨��IL��w���N�c�O�G����G��Ľ!W����cͭ����+JFn���X�~�W\0����EQZN�20��j`#E�?h��o-�-��DSL�|�J����F,�	����;V�m!���b��}\��fp���ͺ�)�pd�ud�+�c�g/M�e�
�I�Ubo����M��}ۄ��\X(�(���X��g]��]~	����ͳ��KM�iΣ�o��Etު?g�x6��p���E��W�g+7:�;��><3���S!�t�~�p6#bFjj�M����
�Uе[�m��j�>~�حH��߱w�@�6S9}V�c��҇~P��8��e?�2_P��4�[2�y��aB��ƭ���m�D�7H�lJڹ�>}���6H�kƍ�\�X�t��оTފ��ă��6Nt��J���X��M��7I��$���E�T�+����k�%7������~Z�\\���>`�V�P� g�j}��X� ��Q9˒ ujW�y�;�W��B�*�@���`���_Ǯy��2}�h{bD '̵G{l�:Lsp�2EHo���{6Gk�]�d⓻�29�ႋ�{骏>tdg�F,d����:�wչI�z�ϋ��u
��u���uNQ#�SyB1V��!��c���8�j	Ų͍�[�2˒vrw0A�mq����{�^�ƃ��]��.7P:�`{Ȁ��/�my�|
d��߫Y�,l�-���2����!�V���'�.�L�2~���
==υ������ �L<놖�7�ێ�6�$tx����c*A8���!dݒy�)P��#��pI�RAc$�Ї	�Y������&��e�]����LT���<�C܉�R�9�ߘy���^F�'�G �#�ق\|Bm�9�:�ӟ�S7��Ҿ_`�TX�ǡ�~�gc�pE�s�
\Fi�P#�uA�$@y��W��JF`O|�~,�>�Z�����9����2c\��X�r�t�������; �UV	}���H�+�g����z-�����B��I���^1v��ؽ(�=���j&+v��9+�ܫ�[:���$��<�s>f�����?I�߁��vx��7Dk�.��7��}�uI�rל����`�nʛJŒ*_:� y��͂����`��ۼǇ�{z3���Iz�$�yX�ڀV2�sv�	:��=΄���(�M�Mm��B�R�kAb?q�ċ�����3<4#��5�!M�KI��N���.N�����H�	9A���0H�T1�=aX�����v�魼A�?�5�qwQ噤�II�W�x�P���e2�>����XA!2�yW6�/����s�d޽�BZD��*�i�H�S1�1/p�/�
��+����m��;!�V-���b�p�N��*׳���N������P��C�^���O�5��,�->�A���N�x�F�����] �|�τu��K�i��^X�:�e�Tl��,�z����"o/�y3�r�L���.%<r����r����&KM� ��n��S�M̶�ir.v��qmT[h�>�<	���QLi����i���EFYי�0m��ؒ�nJ�(�Z�*_��1 8�*	�&L�X�i[�W��бe�`�>{r���Mi��R�� �K
�*V3崜�1g1�B�{�5��1Z������Ug//��G? r�M�����yjʚܹ�0U�QT�&S�E|y�='���D���?�c��MZ�)��x���q���c�ǼL�;*�n��mn��${԰7�24�XYJ�?%�r�T��2	3�":,�����땒�E�@?��Γ��Qg'^�;V1��z���ݟx��q�T�ʐj�����|Z/��2� ����������P�"yHl2iJ�و�h�:����|�D�@����E���I0��cP�`��ڀ���]��`�q��ɒ�ڞFC�`΁�U��W����m.�ۡ���/iVv�~=i���S�F�03P�83�*�֩���,(�B񬻒�)��Kߍf
&����+z�Rf��fQ��޸���+��Z8����KV?��g˭�f��^ '��ʍ��u�jMѢUb��X�K"������l��:2Q-�StYBNꚺ���A���
J������bx(�����嵲B���9��馐�]�=�^���W���� ��X�%ɒ�U1���.�/�x��!��N��`���Y��E��|�_�Ы�Y���G ���+'A��ȳ+,�*Q{����a{J�ǚ�ux����a��vv+#
���?*q0x>F�i8Z�N=�\���r��`���E�k�+2����%Lt��W�̈́g]��L����.�?Ҋ�4��s�[����hl����[T �O�����1���w�����a�`�����Z��	��\� y���T�g��G~S��ض������/����6(V��w���.�E}�g#��n2�4� Ӆ\�5T�j���;�J�Uk��;9=�J��O%[����_�#d�6��[<'G�j�L����4��+P���z.�`y��"r�9�ED�j�Ɂ�f��Zӷ���=�����0���_\���M��|]�r��2� n�B-]z�U����������#�%�xr�ܘ��whd�OJW]Fy�}&�j�g���R����0{���Ot���9��2���6j�v�_�y��Eͫ��\0�s,�暦�8㳄<؞�]��^`M�2�{����6y��e�nH�]�������ݵ�w�yi�6w�F�@찕]���/w�����,b]��GG��'
�
�yՌFkv�~@� _��>�*���O�ʝьqެ�����^=��`��Wߚ*�v��w;L�l��.�2OA	�9��͈xl�#cc�I�۱�x��>"�<����9G��Vo��O���a5���ӃĴz"��u�ܕ��mDG�k��Q����30YJ����/�}q�5O�x�U�S�R�u�����.H��ѿP�Ԍ��hu�4쯞e��0�Pף�����L���q��h�M�޾4읏lȝ;u�ե��Ti���K�����۔�+?]��!}v�S�rNIXe}�eS{�_�������nwF���<��͋�������e���P�{i�D�{�e_�P�����c=q��;A��9p����z/A2�\����rz�Pc��mRc�|r�ax�Y�"l��w}��Ŧ�m����s��8���v.%�O�F�.��'���E�d���2�v�������K�rZ .�Z&}h9Mw&�������!颹 R
Z�¤�М��Z��(^ �C�/
�g�N���-���f�]Ÿ�uv�=��ec�������˿����Ț%kP��W/���юsT��n�ۀ���fP�����n��J�H�q�u��G~h$��:r� s�����~����3$�Łb-����A�����̿	���׈*w���M��װs;mZo�%j�Y�ԑ�:V�	��J
D�dO?-Y�����jiC"�3cw�|�6��O�/,CY�-X����?����h�������"Ra�����
��"m�%�^��߼q3Yږ�g_	���-�ue�^�TW��dӔ��������8&Id�bA��_�U·����h̃7��H�����=�2�����ꠡ#�uoh2�O��e��0�q	5N��՛آbڬ���9@�h*��}�(*�����O�g=��I)��&M��p��FZ㕉!,c� �X�q�(<��D�~�������nE�t!��fǭ�y�1��q/�,����]?~��bۘ'̿N�]�.����ej�r˰��|	EG�x�؅,=�M�,���\��){&�K��[�;I|.�4�W�H���I	��MM�q"
�8cv92��A�ߒ�v���|5{�'�o�ԩ��x�$��%%v�����!��g`66>�~ν��´�e�b��6�-)��X�1�)![�o���y�=$Ĩ��?���J�d���u^0�����7��)��9ɺ� 8��:/�
WW��r��p�{�MQ�����h�dL�t>�'�����
<P�}��$�ߤ[$�xՂ�E�M��� ��Y���I�.�-3K���Ei�`�-Dy<��RBvnmw�M��E�&���m�(c�z<�w]Uno������>�.뛢M�J�H�v��,��.K8��h컸8P��P1jRV��+��^Mc�˲'A�f2v'�sN��$Ф�?D!>�&�o)ǯ�脗�s\�a�������ܛ���(�|�~&�~�sl-f�=}~J��'������4�4��"��o�=���*�ƨ3��>)�*�f3�汌g��G"���`_i�t�[)��Ő2`�O	���e�A�������A�������Cƅ��s,*IW�x�,��YX���Z�e�새�s�2����@��VAW�e�b[U�A�%gkiI�>��7��:}���^Ún$�*�Ә��7~Pajj�<wh9�o��ɹ�����Qby<Ww}`��0/ҷC�z�;M����(9)�����W4+nXB�쫦ᳫ���#�+��.���➝&�y�A��'�k*������zپ�v{?�����U����jS��ݽ�/�W��7.�Lr�1�����w�G��e����_-
X$fda/�d6g�ͮ`������oy*��hp�u�v�;��n�L�%ʾL��zy��q	>�:�~O�����9�
g��/���a-o�������nb�2����su��"�`!uַ�'Iy2>6�-{"��P����^�N9<wLjh4�M��s�U�"�_��V:G*au�� �*�D\P<O�0cՌ�x_�dо⧭(U�b�w~[�s
���X%�z �齱��H���H�_ׅñ��M!t�yt�ꎽ4�3Bgw�eJ�I+E��,8�p!{�l{�{:���d����@�Nq�s��GG�����u��~�C�=�m�˲�!���L�ǐ>�;��B�NK��ٗ4]c�-$]��א5��,&���ˈ�O�����ޖ�}A[_����%�WW��1c�|��`��W��&T��[ҽ߻=�����}�J')s�<E������K�-�Ejj嚼�Jc�lw�J�߿�����u����&^����5���g�0w�GS�U�;�x��<\�2��
:�����Cc�����f�����Ph^�?c���=/Ӈ�E�A5dZ	<3we��]��t)�!5��r|�[�� 
�_t���.^Ä�V2����j�^+u����O���~Q��I�V�j�g�7|)�;<,���?jNr�b5�^���$����9���d��BU�o��ҋ��dC*<�z)�{�g��H�i ���֍[��
�H�1��U�]܈���l ��CP�6O�-M�[���]�����!�,�c�����A&]CX�vh��_mD�'�f3?�A!��"��T�nN?��V���N�K���He]ψR	������2����Pͨ�$�i	ı�Boy�Q��~`�pA��s�p&|Ȉ"�gHm�O����B٭
�����`ĘZ0 ��VGR��\��>��"�߳�H���g���{��=Lf��'�J���-�����<�@�����2�Ր��뙇}�n�Ή�=��̓�8՜C"�����
�	[	[�{>���"�w�-2���5l��J��|�Ps�g��@���*�֩ss����Ϙ���U��+8N}�{^U%Q�yq>H���xM�r��&��rB ��l���=��5���(N��72�o�3��ٙ�#R~�)w��
���������ζaQ���k�s�E�"��D��`�_��"��(�M����U.,���'� ̀b�������{y�6��i�'���aMz��d$}�FRWv��(U�s��2�	�2=�� O;k~N��.v/HG�Ũ�hN��5S�
�Y@t�AV7� ���lU�;�!�k������<-��E)�� �iƘ���y6�͟o�H���	�nQx�&�wҒ���Rɿ�ɇ]~Z�a%�Fd�k�
sO��<�������=.�kl�;yK=۠��L��}9'��X*�8�T[�:���Ǩv�'^5ə�:�P��D�ǈ�o˖����ʸ����zJz���kͩ�˴�}ח�n����`�>_KIpZ[��9#"��J�F��ee�txϬ���*}#B/�[��L�SjI������L��������-��;���f&$
<�L<����������@X��BR�Ա{��64+��w~B�c���ԓnla�]���1�-�`g�Q�D�)tsJ6R�x3�%f9<�&��6�'�V4���� P�J��>��'r_��)�K�^�w�V����Cܠ��*#�ޔ������A�٧���Ʋ�1�y.����<�3>��Ԉ@U�Ǫ^e�wcZt!�^)���̆s3�����(�|WT�L�~0��$�'�P��13',kTy3��͡UKqe��՜��X����}ʱMp�qsCe�R���s���7���.}6�$s����y�t���(�Ɛ��P*��N�����gF+��Mޛ��ۑ�d#�%����h���2%�4����I�2�>d	����7"�	trk$���ኧy�"�����*9�3��u��H`�6R�MG�c^���܁pE��+W��P1VV[�E�a���}�
��Am�&_Y$�5�2��iE[Nj� *D�/}Cބ�7Jc,N���<�����M2����>�R�Vm�C���]��~�0{\C��x�����s��bR��L�}�G]~�
Oe���jjH{y��x�^� U������N�}�<
n���p�����
e��{qG��\ǩ��3f��#D��"����72C@m��Q]� =^:>�)�L�d��"z9��@|I�b��Ǡ�rH�e�"w��!�l;ZT��[c�ڷ�<Gv�4m�@����DY���i�ЬtG��]���΀��џ#k�,��Bl�r�J@�eWg��G���I�Xq�-^����w��&�����w�P��e� �w�	/+�z߇}Z��J驫�-p���g��U<}�Ue�_s�='(4%F���=�4�����ӄ�3��s�,�3��n����7�B`�D$�n�%�\���L�(�1wV
�_@�~]�#2P7?���O�-�6|��ֿ������p�[�uUU�?]]9	@Y?[9a45guv�"X�/C-'<wT�B�Aa={j�IOs����Pןb EF��j.X����}�I�X�5.���\�GQ����R��v�x��8���Z`4-cQc�ճll��ڨu��x �
9W41'[<����f���U@I�`S�IQ&���Ԓ��&��=���]��|d"�T�Xm��W��Q^�p~�����E/�^�=����9;�����y���2�Z��;���)p0��Q�nK�g���yga�7�6~�ԫN�}-999pj��#r�����q�d��G����#�۷�}�� ��p���O��jLN-3�,b����9j��jz+�v��1oe&M�`�o�e�'��*�N�]O���[��p��%ٙ��3��^���	�R�zn����BH='��~�@���~��ĩ��'�����t��e���^��D�K=d�S��>���,�5�aH�M����NE��`_4�e��L�P�4�Ȗ��k��&G_��Nņ�oH��\�=�&�I���Eڄ}�ѷፃ����8d"�C����{��e�V�Rt��ON�xi{�D*��P7�
1���9�� 3���K�P��ܝ穰 �
Y-?���3x�Ѻ�����7�IT@=�O��;�;�A*�KxÙ�}\�js���9�r�[���L�3���G����2}��E��������?Ɣ���k|��%�-�O�ZU�bp�8���k�I�yq�� =�-�����k����t�rX���-�yJ�2��l�C!H� ʕ���6�Tt
[���=�S9�S��i��>���T����o�e,߇�ډfkqe�BD���3��@)K8T(=\�a�>���a���c=��u�̞�{�_��`���H�2��o�ϵ��dr!_h(�7\%����_��r6�EMW��F�'��9�';�Y_Њ��ٶ:f4�t�֠T_#���t+�f�{�������/5&����,B������j�Ơ2of��d�Bj�,�fn�7�n��1�\��{k�~B�NNŮ�([R�4�s�Kgo5,ԯ�}��-Ɓ��#4�/�7��E)�fvvz���
�T�A��;Uа�]�_���W��\��^Byyy�ؑ��Y��S$��q�������zF�����+ԕ��rP�X�j�k���`~��<�I��_��\��iK,e�����0LXa�]�[$�D��\��h����}ؾ�Ƹ0�)!w?��6�%u~���F��?����W,�����j1�\^�q<�vp�aJ�iAaN��ѪYUR����`�ʻ���5]��!�s4	6o��g�"P��AB�tN h��h�4�FQ���0�|0�3�p��ƣ�0{�~_������U�i��R}(�ޏ1�n9��&q�ı�����K]X�sR�C^��!1�WLb���A	����F��S�Y{0Qi{��Jg	:Z�U��oy��ԉ�ޑ(b�"�%��������>��k�4���l��#c�d��r�V���.���y+����]}�_h�n�KE'�A=H}���<l���%�S�y�ա�&�K�"�J7�kn��y�ȥPŌ�t���o��_6��h���Y S�3��@��`�0�U���Q,�E ���O���x��g�Sl��l""%ޯZ���4������CP��L_w���BZ�.�Z����<ꡟ��[#!�W3�Ս�u X�dx�����a�{��H3��N�PIm��,:�N�X� /�o�_�ξ��hw�Q_"X�-odz�ש���0 �ga�a��<�t�,�\J��Zo��񵪈��-�eNk�$����ZbB��f��K�����d��1�w��C�u��_@Ҩ�	���)T�lEc�d$g��%c���<�m	Wx��.�����O5���U7�|xb'��<��y���0ʤ��#E�z	��װ4���rS'��s�4�Wݧ"�\��D&z��#�V���E�$߇�%��ME}�A���x�� �Ș�vXa��7��p�?*�� �z��X7���e��r�8�[��Ed�Pqb	����I'y��+*�K�N}N�5HOn2�<��|��}��0����C�$&Y����,l(Q��y*f�Ն�P��̟v���WҖO�� R�}���.:�l�%�ܶP��������]4z�|UIEu��?����ΝHYh�C��P��O\&�;V')xv��%�f{��m���M�t�H���,Ȭ�J�%�o'X���#��ny<�%\f�ƌ��q` �[;ڐ^��b�7
������YV`�]�@1pl���޸��m�Zj�e�P���>u��ct��JR�ƣ30��>H��-�2w����h�k7Ϩ�r_,�}��@9��[Af4
�7�D��������7������E�t%EO�T��Ͻ[�a�8��dOGݥB��<��?�f�/�&$͒ݷB!f�����+~Z���*S���?yE�3����W-
ص(�1��Pz�����_ !x�����{[��p�]T������iV�-m#��]j�Ӌg7��T�y.�g���'��!y��E|��N���� ��jE���k��ę`Q����q�,��M��v3���w�_�]��C����}z�{��]�d(w�܃�݃����V�~�ﰈ��u^й�u��0$r�}���o���[:%�`u�~�������Y4�S�
b�m�����8kp����x�����^l�6��^{
\��=j�¯��L��/���rw�>fP��㒺����"xb����գS�آT�KV���=U�ˮ��U�5�3��T����(Ӓ^�t�ъ�(�ɲ���%�4�_?�mZ0�$������$�O5���U�]E�����eM�6����Y*x=T�b�ra\u�v���.K�������*`%M3URP�~��b��������&rW�V�����e8a��T�斷D+�I�/�2x��un���$��v�ZF�^��r]����2WTǲ�@����7��zq}���H�01�,�~EIII�r�j��&���ƲI���yF�Pi�~Ը�,�cy��GK.�fQ�[�n9���B��+�J��C�/�|P�خ�O �+3�ތ'��8��)C�,�� %���϶�54:��1!`��m7%�fZ��i^	}������oV�]A�9J�l�EbF���jp��$I�����G] 39���suc̿`�B_ƻ|�rKO�������0 �N��C�4b�k��3;;;;��q����՘��+�^y䵐>ʩ��XU)ݮ��_�� '�7���D�\���1 ��#�V~`)��iLJ0���m4�X3!�8K
��G�xF139���"�h� a�V��:�ڕ�m�*s�֚?�V��ݾ�?>2�@���I|�:*5|m�mT�����.Z<��k羄�<>���I��\�N&��au��(#ߊ�S��d��n�ܕ-������
��7��u�w���`<���F[i�|e�U�{��H���;|����N�x�=�&{��2�
�L����DUs�~�Pz(���=�K�_u�����o�t��I����CUF����J3�I�N@c���\]�y*ɦ*\��}d_�^��{ �-k��SkwG��C�^ޒVt�Ut�ؤ�6�*�sm���]hèW�Y�ӏZ�����`h�)�����׆g���Ӕ�4N�au�ȕ������p��ka�"ǔ��q��㖐mb��<i�78��:�E_F�Ph�Db~[?�;�N�U����ӧ#P�	�߿�џtL"*]�	�V٩�o"
�[;�m@�������"�� 5鼓���h��<l�Rt��<�}��UWP)@�7�m%x��ѕ���R0V������7¦�j!3�J��M�����G��=��@o�#�@�](�M'ݐ��tB|�Rp�Pts��q�{���r�r�xi�����@M���n�q;�۱z�}j6�����N�����o^������Z�3�M��˓[�Pް�X���*�2�q�y���511�L':�z���N�z�)�ژ��A�Lh̯�X����!חMK�!h�f2��'o�Ki���U78�wZ��!�9���x�
���I�R�O��S&#��a���5�Վ��n��^�Z���&��"�i���*��8�E�_qqqPs���`=��7V����/�� ���B��Ï���{�bf����6V!!eP��Y����jz#��Hy��p��V4���1�Sb���8Qʅon{D�ϯ�a�K��G�Uz���g���Ѐ_�i��J/w-��f2�6OT�:��Mh$����^/�5աzOQ��/t��9������Vw�q���S�D��2�7�P�����O���S*X�	�K��$罬U�h�F��u���L�a(E0o�ʦ�h��ŏ�ϼ_,���U6������Q�� ��Dn\�K�nha��]�H|M���2�tY{����!h����kY:�ae�q�'�B�����:]3�^�.���i�W@}5>��#��������[�E���㽾Y�v��9�~TQu��ZP@�|��Ʃ>�U��
o%����500�8�ĉ���[��V^-�)�*j9�X�)b99J{r�W 4��M����A���
���,G��xF#K�\?�l�^�'��EX����ʄwB}A�@�y1-=���D�,�Ím���w�Ըuf��^ ��0��ݟ���!l�6��Ч��H�x��n���,�L���_O�s-S�[(��At	�ƫ���X�&{j5l��J��t�TI���>=��j7�v`*���l�[0f�G.�%9�l-J��K�����>M�&��AM������?%EQ�`R��� f��4@��c��N��+�'퓯V�akEkK�J�����F��"v~�)� 
���n��㾻!��n-���5r/7��z ���6o�a���8��q�|�ҏ��`��P|o�y�7N��mJ�?{UÖ��^��e��|��#P����
k��#X���˕k��M� v5��S��(0�I�M�z��%i���S��D2�W������-�����Y���N��ʂ�(ɚhM���S���U��N�:rE��r�O�����ȾIy-Ol�LJ����s�Oc�\7�^s�_P��A�W5&OM��r�ܠ�T�z9���g�w��hV~�Ȧ
�9���r��)"�oX\�r
O$s�Ûۘ�NfF�%*QWG)JQm&�t�CoI���!Z)�f���6K}��Է�G&ZL�w}�8㓒 JI�ɓ@��n���/(�O�r1R�s5�76�|��n��x��]d�����G��A�k�P�S�������
c�� N��H�A�{�34��_Zoj%����N[�Ua4+5CD7O�d+��9
�� BO�r�����l����g��?�P��s��o�	g��y���j�M=}m�^)fLk�F��r�!�r4]2��u�[��և�y���j�L�}�����v�EL���l7� �
��ff�>��59�c]�P�Ivc�
b�l��/�Uf�x_J�T���l��J_���9��v�>v�gJ�v�L������$Ұ����"=��r�v�$l�����g"}X�؝��g����1�������K@�Խ�$��eM�gM���Z �&���I���B+��L\m3TC���y�z;8�P#��_�-��Th�Kզ��^
�GQ3A~,����:��9�jA��ż����}[��,a��e������O��M	�9!p���|7V�r����J.����r�����U��S�r��Y����x:�t�sfQ�b��#��h2�������H��54��o��*��4d�= }�u��
[��{NZ�_��(ȘZ����m�<[���׶џ�
�-.ag��;�Q�1��G�d-�1F��(�_�l��X�Qv�%���;h�����Fd��4+*0��B^*��mՏ�T���3T�ZP��R<uN�K ��,)}�iR�0�i����J��[�y���5�����;�/���	��_����ݝ��(<<}�}���F�+G�;�c����� u���|������y+��X���r9��Nh�j�g`8�MnCrpxd�D8��j ��=�XI���3�����^ܗ�ĕT�g�tm �pj\w�YL��!hȦ��[�{Iy����*��(g�|	.!?�z8��;��؉c��$��?�������A�//�I�v���rs����.O�$�l����4cw��2��8qjL?�2��L�ݹ�ǍLl����|�'��$���e"<[�Q��Z|-/+-�%�1�(��m�$�kY�k����OEh�ym��0�B���R����N=�뉶�.��uƅi���p�9'�?��}oM��>q�fR������~|�EG8�r�ߦ�cY��t����Ih�}&��jP]��2��^_.��j>��K��6�+8~���q�(��uEf�a`)5r�<��QW�Cڒ �cTqq�� �FS��/vޓ�m��p�z� ����P#Ҫ[7"��w?�Xx��u�JA���h�t�)#6�
H���3�K��u�R����a�m�����D�U��ՙ�p �7>8��\��tK{J/a��4���_E�dP��=4rZ�Zt�1}����q��>� �!��!O�?#�o��O�V���0�G��e��l�yÂ��f�^�m���RFފ��ips)usD:h�+��T?�L��T\ou��ON���l��h�� }x�P݊��a|[���Fܬ�ɼ���J��y�����y&Dʖ}�2aS(釀-��M)�����xJ���ֹM�H���?Gh�7�c��O��"-�G��e�����=<�t!�p|LT|]A��۽�C�j�o��,�A��D��ā�-���@��>�э�'�V�(��=��#���R��W��m�K�x�j���~��l_�
�N깺s�睠]�`��l��>͢KG�+�_��m����.Ĩ�����{����)=mj�a��OB&����`&�;f֝��� o�NQ3B�c�|���[ ���	�����pO8�x���=;�$u������N� k����4�m�n/G�,��e��Up��Y�T��S�[_L�~���Sj���6�$�z�P����Dl0ەw����V�� ���h��Q"A��LPj?�4��?�4�F���3��c<�#�ſȀf� Vە%�"(~���2���nd[^f�P_�&�u)�jxA�],)W%�đ�d~���nM���NN��WM�=}���0�Dr
#oiݻ��C�Wj�\)��?�������6I�&�k��d��D���Ԅ����j6c��}�����o���!j��/�.1:�{�'X��1�<��3jC���ݔ��uErN=��r�[�ˡ�����Ę�5*Q�k@������O���*GBd3y��˲�>�΄��q��cPe*�]���0�-Ķ�P��[^���t��{f����^���m߭�KJ�d�.�+e���h]p0�5�({꣈V�ʓx�r�X�"Ů���K����hn�ո�vi+�vL�X�.K����'�d)��:�ޫ0�������?9dS��ɮ�tdD�讄�d���SVG����EQ�l99Ƒ��BV��d�C���]o���{<�'�^�k<���N��2�g~ӯh�qiNx��R�g$��>��$��37�#XMuIa�M}�Y�^mB���Yy�~K�ːӔ��?� x��,Z���{�XjA3u��ro���{���F�T��(�<�m��}���i+?���:����n���k�v���B�����0���o�,��B��`�=-�;v��ș�e��m^���-�Њ߶�z���jAȟ1���c�OoN��� �i�q3_e�0q��L���ֲ:��%���������},@�z���%|�gpp�kx8k�+A�4Aڠ1Y'Nݼ�����=%<'*T(44t�m��Z�s�q&��	v�ƺ��p7JN��9 k�Ue%{(��� �t�Q=R�6������q�F���� ەo�ׯ��jjj�_}&�8��օ͗A���33-w9��'vT�~5U�q+mK�':��G;h��J��=��m��)^++ny^��M�����KZO0��s-n�ЃNyq�"K���_g��F
VPWW��q� ��03Lޓ��u�EԚ�u.W�Z
j��OS�Z�0�jLLX=nk}=8��u����2��������wɑ'^�|��e����=�%txE'�<�%�5���S5�����Ur���nCӱ�A~▽VXQ5q�0��sm'"x��˃�z�+����H��X�nl<���}a�޳ۥ��y��l|Rj��Kv���k�ќ�S��a~N��-}��:\37�X�#�)?=n�ٮ��p�F��+}�J��7&�i�􅋕Y�Ž�ѐzd�z%� 6��U��Ǧ��iȧ?�7���I���Sտ�C�9jUA˼{��j�%�Ec`_?u����@�7��"�h�!����'� ��$rL����#ZI�^����JW�N�a��4>8��W��A��'i���NL0ϖ����b�j97�e�b�L�����|о���(]"��S���p~��ku�]%%Ogg��С��̱�Dm��Pm7���{��W<�OM1��Jc^��$���ʲ�'��g����s�R�!����!�&�G��j^I��O���b*��ia��ӳ�f�%v_Yʟ��Y�Y�q��u��ͼ�b��]O�ۭ.s�6�555��v�h��\/��EEY
�m�`}G��'Y����72��yE��8m����=&��x� o.pM����P��ɦ��Bp:o���(]����w?@II��zr�I��tD���/)��+�}���}*�49Z���]���(��w������lV�`�A#%ޯx�����UE��N����Ӑv�=c��J���H��+�����D�Qć�⯛����C�I���J�x�z���>�V=X�#cxK��XS�
��3��RN��`���NE�U>�F�9�l�)֎%���Byu��*PVl��ȕϚ�z�h�c������'%����	�F�`?3���e�p�c���5�ϲ�z�x��2Tߨ(�>��������+?���k��S�E?Qǈ�V81���!9��z��v����z����ыd�2)j넄��L�g��h��
5��i"�o*d]b�N�!G�Dd_��x�	Ý�;����$m׭�	{�VZ^~�2F�� �|`&�yM�N�Q.4�^%_�F�7x�x\��/}��_Y��W��b.�[n��R���]��(��瘖�h�~/�w��g�=Ŏ����?��������,��OM��H���f�)���m�Ճ�|���Cᒔ�]�����6=+.Zb�G:�F��_#��. �C����x�f��9i��9]H1	��?�������1��=�> �PȞ�*IЗ	\H��{�cm+I���	)��'骺��UUn>�~qXwyk������������Fp�]�	i�r�Y��-�Я��x͟�������t�dW��qT�� �ɷ[�J+** ��~TĒ��K��7��D��Ԡ`kk�ãzb���`SsklD�[�34n��l���O���O=��l>��q����g+mi�d�jƏ
�>��u#�~���'�˴���@�ͪRc�=Z���������_�ml��,wz�E�`'C�&o�A��p3�f!�h����?`4^����'���iR�Q$ԭ����&v�+^ԫI�颉�Q�0r����>炶�	y����a��΃lD�)� �2�&�o1��2Ÿc�ֿښ}��(Q ,3��ۛi-�# G���)����Q�V���M��Y��Rl��v�==�Ū�K�A{=���0�*-t:���,U\.�H���a߉�J���"&/�Y�u8ꘙ`2%�?;��F۵�X(�,��t���QV\L�� ��W3h;��í��W��`�w�$�u����@Z^~S��9Y6��Ca������+L���f_�L�W�c{V���ܳ��&��

�֏����&�ߓ�X�������'�/����T�ѻ�G��f[��.'�/6 a����M���i��Vud�}a�;��&ݣ��зdt��|3��	�am,�%�P�=4����vS�o���ʰ��j���85a�@_��֦�&��m�ǩ����X��[iVb^�Q��
���hN@r\i��d�5�_�S������C3�����i}]+56�B��z/�k�]фl����OV�:��\5a���ړ��l��0��0�B�0�_JyM�@�qz%=�JF����vpx1��E��s�F�qvmD&P(7$��R�	h==K��~S�Ԫ�m�f� ���J�9,�����_���S���vW�R��׫5�$e�t���񲲱au2���?X���$�<_����h7^O96�42RN�iS� �D��3D�K#n�f��0�[����ֱ����wA����y��>�'����#0��$�������r<q*�>�2�GX�M�/n�>0O=-gQ�}�ڵk���Wն	@�$��Ss��2^��f�[bp�*5�F6vr.���e��<�u�H֒	���f����e��Q����TK�09�<7�^x���ԯ�ȫ���	�_����6~�Hz+���A`;6":�7��8��e�����YZ���[֨y�r�~��o/a��U(�O�y��7�ۏr#oHE��Q��6喅97A���k�N�@<��i���8b�_�����F���>" S�K�G����/��<�8s�!$�Ԉ��#2�~���;��ȾT(��i���+�#�0�T�2;q+`�����ܜh��r|��4�?؀%b��$tv�$&�͘���uԛ���ܸ}�v��[b��|&,
���Q�|��sk�7����2�?�йq����ʕ��6"a8fO���E��.���F(6���j(;�f�$n���aᎵ]yU�b�L}�-��,�Аkn����"��+�.��*��u���3�U��?�ؚ�32p�[��r���b>��R&�<Y�P��G��[�O#r��J7�^�3�pJ�/Mоw��%EE�����͟{~�2͟���6X�+��)��nl�Xm��E����j��K�h�dLFj%j�4��������13ށ�`��`����"%����҇;&�Px�_��V�?x-����W�� =rn����NQ�A�}	���aGBr97ʁئ�A_Y��iKȐTza����Ċ{�l k�*nO)�����a8nLHz��-�]^�vw�F�tPj�r��۰I> Zzꑍ����!lp�V9��*�؍� ) ��z頋�N=>�U�8]t�od�sq`�ݲ��7u�����;_k^	l�,��˃�tuoFV; q@��p7Z�����l>��>���0^�U1 }v�W[�s"Ƿo����w�`�����f���l��ӣ��1��	nA;V�nx�R5x7�������ܬ2ʽ �5�Ǽj��dۻ�a+�U/�C���Wf�Kʦ��I��N�e�=Ы�֏�.��>'}�Nl�A q����θ��&�B�w_�	W�"ޡ,&���|� �bs���gI�߸0P��R���&V&�c__@Ӡ�+9p���0��+�?N��S�������2C�ih�ӑ#l�7�n����c@������� 2��v1��Er�S"��%�
h"3��5��y纴��L(�O�ssHC�w���2�?�;dWZ��ðy�d`���%4D/��#�3(�)�%��M(]@U��]/����X�xAB[�kVV?�5�Q���b����
�
ac���4��I��Nzaha暎A��IX˱��}b�6�z��qn�0��<7��4.��H��0�}D=��R��7�
�^ �U,�=�m�m���������K���OT�Q[�k{�5�qP^Y���-u�[.�F������[in��Y6q�zdfhtD�����SH�_g�7�,�gJI�/^�|5&�`�����Lk{���_�0�2i��eI�vl���tU�GIc~�`O�Y�����p6@E�C�����C�S�]p����(`v�H���jLM���N�iY":��s���3a��i��_=�*�7\\��Ҷ���,��#������I�9Ɩw��l�VSgN���?�z�87D9�#]#�g3�e�+��B5���^l����n�_��X��f&���ي�o"N�e��0�����8$��}��y�Y�d��=,��e���vb̍�0�S^K`eR�\�~o���F��9�g�B�#�pz��<񔀂"P���~j19-�P74�n$�^�\�s�����--iZV�AbY-�4~3b7.z(s���ׁ:���+�R3`'X�ĚFG_������/;��4��ɖV��Y�6��ne�V%8��C���[W��ސ�X��T�&gg�� M��TVT|ו#P�"�N�ƕs>�%��Y L+)YH-���T�i��X�\��ȥqeA.b��n��E&nE�1�K�[�Xoؤy�X��jKQx1��NSS+(��ƹ��v��S}��n����RPRB/��J���t^��x�����Ye��Ҕ=}�^��ުl�(��NVfwK���@�z$.T(Џ�a���>(���uh1'�2_tm��P?������/<3��}�Fh@}ϕ�������Ձ=��:;��OҊ���I�
3g�1UW����8K�89����]���L\����|Lo}8(&�}c Ia��*.����n��u�R����vjMxhh:�QA�u�����{�P!&��5�vևրQ=|������xs �� 5��k�}O����Tu����S����ӫ��t	� w�t�t�[5��{3�ޚjSc�P��E�2��΍)��f�Wi�!�ӏS�l�cx����_�ul��O����?[ݍڞ�db���T�G�G���Ɪ��w��vWߍ��H�s{e�s�$drf�z`��u^I���j�;��bb���������7��45e�Z;#(���K�f�����{�c��#�/��ޮ�P���%��ƲR���V�(�����y3֜��s��H�Ϯ�n�d�92�_�~��s�'Q��G�[g��ԋio��{j����˳��:1�̙�-��d�v)���f�-�WJ
����:iђ`����tǽ�ິ�Sd��U�����2H��M���1P��Ir�SiZ���r��r���ai��#�j{%���Q�t���Co�H<}Z��6<��vW���,*�>x��2!�������C�+���;�m�˹���6�B�߮q�m�j^+'�g[����/�z��@N,M3�QO�Ac��>/"4�p\��p���"���~0�c�W��cg~�LVĆn��\�^��Z��9���ڍ�g�Oas|
����Yp<�A�9>Å�&�{�c�gN��h�~p3�����+=�a���̓;����a4����z�7Htwt!{����{�]n��F������kc��Z��c^ ��\ �1lm��C��\�	��k�=��`i��~*�T��5�Lpx�F��V��5J�p��\��\8��=8�}DP��(XN"}�:��6������Lq�e���r)Z�z�}�=u!΁���J�|~��ծ�����F_d���w�P�2kl@�v�YE�N�E�Lp:�ʸ��6�x�?5׻]���U�+�~[��&�X|�i��JoyL�p����{�O\�(��XD����1���?��uߘ���.���%���KHye��}]��xYi�(����NǶ�R/�nd�|@3� 3�z�M����J�Z��9���H�0- )��S��4���O+9P<Ի��À:gA�O>v�����������L6+~j������'w!�c��W��C�7������\�N��0ڍl"�#O�f�CY����a���d����~T�q�vy^]�m*����Nݵ�"�jS�T�LM�lO�SeUϬ�/>M��ٺ�.��׵�m�������u�YW`���!��f�BBDGL��0�^���)'���k
��<!ٞ����D|E���u�&�|�%f)h#���[=��,���!%�e�`�{�Km��0��u�3g1�25f�1>���h�ދɛ��y�Wd���%ج;6�q/�:y�	�N������֝�(�c��{Fx]��x��N�lI�<���,�YZX!��n޻����U���cS��M������{*P����N	����v���(�a�W?t��9�Q��,���W�������9�GZ�m�KD�M���!�t�lRg�݆��<%Eˊ禧
��wK��/T�v��i���z�*�n/u�,�����;�Ζ���>�hi2B�_
�J�[���Қ���?\)�s�,�u��![>t�ݘ�.�1P�E7��Q���A4�לk��7B���<H�%w���A�-Iy��H L.��:�\�M,�l��)b�;nm�jH�wePÎb �Z�Y��@����ҳkՍ��������:o�]�M��e.��Y��	�B��5
7���'�m$9?��~]^&<?ϢQQ�J����Klu��8ۭ�xD�.A?�c�{�@��WF$7���m��Ŀ=��g�������rU0fĔ׵��*����8r����yv�gU���u�'����V	�a��\.�do�����<�V�|!$&�U&\��qA�W�^���忱x���!�����΋��a_U������v�'�\<1sJ}8|-'��Q��ߐ�2�))lA����v�_'E#kj�SQ�/�Gb?�x�4s�w�
R�eqrph�%��s�j��g�_Oˡ��+����7�x���Q����#���URY����C����{��ث1�X�-! :�n���SU�V����u^�Q�,LCj��M6�G[B�j������ݏ��h�x4������n��R.]�q4f��׍��3�,���fM7%rX�J��s%&�;��]��H��+)a�]�a�Ar��ʏd�zZ�f0;LEM���=�c����� +�Ia[��d�O�����<�4�&r�ˆ��x��Z{���$W��
��Vv��B��ͻ/9c�ٻ�����#�'i�8ɫ~�����JOǙj��E�'�����řN��N�`�>��ؑJ�b:�[��;0�Uֆ�84S!T��u�XVTR����k},*p+��S��s����n��Q[q��\+'Rj��@���>����g,�J�%�
�Ŝ35�t=M���,�e"M@Z��;�+hik$�l����l|։{|�}��`�o�joK�Ӯ>�wX9K����QN�$B���ѓ�a������[A?��b���2)���:�C^�%��	ti��W)�m4�J111^��GX￧J�Ȳv��>�T��AWW� 6J655a���|������z�nd�M?�R\�	�����?t�N��Y,..�y�pa�
�����5'�����3��� >o�)uzĞ����E��~���;�βݗ��Č܋�q��LfG*�>�	�����w������&-��%�,��P�?p����ń�W��K몧"Y��g{y��Ps8쐙KLa�7CCM�@ch�+�o��-lSB�u��F��m���w��YEf��K����I��?��\��k��_���۞&���/��������;n]��D��Ǽ��3��ǂ%�<��&@W@�U۱v�kR� 뎮�������#�H�� ��aq�Px��X,��' ��͏fCa���G��B�3��~�e��&�����.�w�p�W�a�XE��}'B��'�p΅��F�W<�ǣ��u�	��Ӵ,E�T�IK�|隋��չo6����GHK�r4�P_Nq��RMC��~`���}�����sU���fl�:��7���ފ#�+��N�
tH���C��|�B�GOlWW�ng�
> ����Ü���>�j��#�HDw)��k�FK���1�|å_1����iPc$%r��Ng��+�r�<��F">Kv&�E�$BS���jv<���N�	`A��-�kE�Va��b�[2�u��Qx��/�ѩmv����I?]���ƤB�,b/�\�bJ<r^Q�(������.��Gi����4������t�0�2]ӵ[�����6��n��������s��?3��!-�i�G�Q�3�D�۬|�7����0���Mi�[�Iy<�,�S$�O�F���	�9���LWV�d�-��[ ��GOZ`��w�4)�y�\7EHk%m�2;�=�ug}RZs䯳}+�程�
��C�7H�jl�J����X�'�Ѻ4'�LN�(�ܯC��/,77~��E#5D�~2����.�b��!�t�f��F	TUlJ�*��Sb�ώ���f�m�i�A�КNX�U�9���'�Ze�}�/e�BM�u�[�d�dj.wG�MԾ2��>/V�J8�K�������CZ�^[��*\$�#���3�ϩ\j��_)N���ש������WYe�8����k��Z�����NZ��V�������	I��6��v�L�]�C�v���S#��7���8�`x{[�;n� ��>�� 73c⦟�g'��Θ����X���S uY:\�&���iݫ����J���!��[���S����џ�_�u�����Ɗ��`Z���D8��	���1�[���ڽ�ne��0ioY(����.+�t��Sct��[���}ԅ�V��qa�X��{Vw��oUX�8�bX|�r�e.����y���n?M8|������V[��=�d,�ޯ+@��?1�,�s4M�A/��9s�4#���WEA!ܾU�A�r|����:����/�	{dʽ	�8���:��)�*�*��g�SS$�{@�c2=h���h�|���VR�B�0?���ز���wa����7>��<�.�6';"����a�\�m�n���OL:b6�0���lJ���5�����ޞqįD��6K�/l&D��)����:��0��~G�4���|t��m�w�g�.�B�;h�  96M�S4���cy�1��L���a��GG��CI8t�����FM�r:@9����wV�p����'�لL3�B��lӂ�5��I�Y^|���� �Č)�f�u�ߟ�̬�;���%+���)����9}�wy����0�`�9�9��F:�K5��zIfKb<Xq��H�٘���Y���q$�m�+�e�?9�Z̟�9�PB;k&��r<�CĆ��Ѝ��[�&�2��.�Z���;��`;�sO���7]~ͬ=�[X9Zמ9޺�(���)(`b�ګ�~�KryUPקE��!���1��I	��I����d�#�v�H�ॴ���"\��q�� *~=xS�:tb>�ku7�M���D�u��?c��[������>��A�1mZ�X~�-��5�Wt��8Q0�����ҷ��'�����?�H$)5_k�on(3��:�Ǩ�!��b�jo�-�3��u|~vl���mf��X�6���o�f��d��S�Ҟ9������l�Gi��oi� ����an�+j@Q���iH��zV]~�EN��B�Oݺ����cz�H�@��I�O,,K+x�{��"��ne	�����6�*8�+^ـ�S+9��$�ZgA�3�����J�.VR�v��9�.�R_R���R�A�uj��D��>F�TW7?���q%��o8e�1��}�G}e%:� <B���y�L`n������~�Q$�Uۇ�w�P@�Ը:ܩ�����(����J����aFc�!9Po[S�p���Bܖ�4ŕ{�1!/�+L�����Ջ�:q���V�T��&��&��g��U���ׄ����������g�u#S��*�@7)[�݀�~f�ObE��(��h��y;}4П��+��o�3s)6GA��������̄)�6�o�5ٞMVJ�\���(��)C-�:�U0T�����C��ּ{I⽫�_��4�jeE4�]��լT����?Q��	�����,�A,��K��v��1�$w�mEb��I,N'������ �K�"�{n�(7)�6�˃�z�LW�� ���&�_�đI)�o�M^?���O�%y���G���7���H׻)y�EIl�^���DM$Em�"��F��-2�n.��C{��&
>�~�b+od�*n-����;"H}���ov����g�Y�o&�y6�����q^��]F�U���w����V�1-A]�����S�+��y�xQ$�o@P jȼ����Q%���u�s�?]K?�t���Wc���w��[en7+��I�_�����R�V^!�쥙~/��4��&�t�:��j����IT��FEEř�t�}��QԷ�R���"{A�j=���-.IJ������1�Xh���Ť�E�1��ts8��5B`Y��g��k�x��6����y�����a��ȿPUP~G���n, ����y�� �"���8����qY��4]��P�����1�P6+��;��wZ+�O0�����"�z������;�F	���Z~E��!4�2�� ���*���T���FB%{a���ȣ���=DE�V��K�W_�k��_�mhOt�n���Uٴ���:��%��q%����@A�UnУ�
J�LX��K(�p# ���S�b�����Yϓ,���f�R��֊�W�n��:�/ũ�dBW~����	��Xz����.C���g��=p�(1Ff�f^�ҷо�/3k�AB�md ��2�E�Qи:�1��)��f����P�����\B=<�t��D�y�m��D�ʐMh���~�]�"�#���X�_�ޙ�E��N�ܮ��8��K�,.�`�%y)�25��|��e2GM�H�mB�c�=���Ր��(�f?M�<�s=���\���aQ�[����4�����Tf2&��<f)�7U���bl��4Ѝ�����f%�s㦦AȺ�P��_�M��d�߻����fe�C �y�y�%3�阇E�ܹ��;^ vOW�n�ΝD�MŠ�y��ʈ���� ���;fD=ۺ��W�OL����6x��X����ĝ�]�=���s��R�9K�/t���B�����:5|��:,_'=���Wt�ǭo;m�CN*~�	��3��F��T<�$�gӦ�Zs�ܫƙ�r٭4������t�F�jc�#Il?�t��@�2	�O��������\8ﴮ��焯��Z |��B�$-���1*�hE�A��W#8t3��3*�BV��9�ʰ���R?W���u�I����.~�3E/t�z��m�sj����!��Ԩyq�;h�'z�� *���a�����!��~Խ�67p؋�K��������.g�{�i���;�_ɱl�
^�e�ZS�4}%���dO=2� ��~LV���V~����5
�*V��4����=�&Dl�Ww8� <Q��$NͯP]���n�>��+`�>Jz�0/;�c�Fi�=ˉ�|�:hS�k8�R퓝jU0��l�J7��j���{�x�z��� 4ݜ�z���J9�s���*�����~�.V��������!)��A�1�O)t����Y���E���L�g4c��`�g�!��Ѣ��gZ�+-��6�d2�ئP&�W���ș�R̬R�@�r7؆9eĺ�	�M&����8 t�nj�
�0K	~ڦS�ș�ӧV�� �֟�ӾMIk��}���Y(�^��G�����Kn�X6~U �o�`�V�0�R�P;�k�A�<"h-��ͫm"ٴnJ���J\/����"T"�^�&���SV���M�z��Ȳ�&љJ&�Ն� g��B80���׶Wt1�G�g�^іm�AH����ٖ�u,T`�:7J�̖8&P�K�6~��*�;{c��NP`YSǯ*}�es�	Š��Y�cA�$����9��=*��J�����O`����~Z?=�j	�-έ���F���� +�J����mm�Y��
z�gP�8��KD�p����K�di :��)�_@�3��t���g��G��_K�S��R�]S��{<��&K9��ݐE��N����4p;��xb�21��Rڐ�6�W�U���ՠ��#�3R��0\���G��-q�B�1�[&�����*İ8 ��6(�|�a������1� �N,Z��ǹ�Z�-�S��=! _�w��q���V%��O�9�
��}�p�u������&��yqhP'�N�|c'f�4�D��������#G'�_k��D��cP���; ��ԑ��0�ʕ����rm/�Y(��oefV@=�zC�.p:To�Sf'�$��{�T�P橺���V�6�D�����xF�����H �Ǚ�4j@���ȫ�l0�����PasLI\
�`eflv����<k����_
r�0�艀44�˄k�>.Ëߟ�?��dҝ� %�j�i	���NZ����w��u��/w*��a�����g�݃��>��������/�0K�~�Y�Qk�^:�n�_\3G���XS ?�$Ǘ�2�Җ����ʹ��DGr�������?r�ey-:w��Ma���q�[�_[���ɑ�^~W�,�ѻH�1;�}`@s�m���p�� �-m�t(��\?��;�에�7���Q���f>�	\w.��t}��J�=-�E�L�����a _�:��������c ��u�����$'�N[t���<���E���Ō���=��ro7F�,0Q}�|���A�������~��v�w�a'bC�g�G���cxi	�y��s� �8�w�� b�	�?6}Jz�*H������T���lD��=@�PF6�ȩ	lQ��C�K�j��-����p;�u���H�b�gL�&(=��G�����0��D�: ��q�@�����=��#��GI�8�_q�Ys.�7���RE��h���:���_¡�q�SS�3�;п��}�Z:7`3�����(cr�[�@�f��/�����v��G�s}�����h����r`�(&Q��ɱ�a��0�@ >~����Y[k�]��%��.��%���',�-��/������A\�'�_����A�bͯ��J	J��<}_x�ȸ؉11T�i	6��dӼ
+����
|/*��{���/�aϷ�tT�s��%uQ��CKe`��W�G��|~�}��L���=�ؕ�N����׻o�|@�@���J�i޷�v9�7�ԅ@O�tr;
T�>|N�LE|�x���_��C�,�v��M�gdPHR�&�r	��.�{��ز����y�N�+=�N��8���_�S�ܰIwݿ o]�N�+cb�_�3v�Kڧ~�/�1{�`��Y�Nr���.ՇE�eڱЍ"��a}7���B����LX����.RP+_H�f�������N��2 �.�3��a�Q^ϛ�ĩ;���㥷���O�lTr
���rf�y�:I�ΘcȄK�
�S~�����> ;@m�	(��bJQo����w:�S��U�f"7����M���=��nS�X{�Ӆ��>�"��/��<��Z�;�q�����(�wcP�,���Q�An���I�*�l �P	����J0��=|�$��d�h���ǾZs��UA$}�ц��-y�p��(U�;/z�!��@��G�ʵ��2���r!��p����;����;�*&�Lu��2���U_�z�7��A�v-��L؛�6׀~}�*�3��AJ��,Ԋ�s*��c�AuN�f�����۸P՚
jc�j�3/�ʄ���I)�`�u�t�����"f/���2�D���8 N�������j`�r���Z�t���F��g�Kb�m fRϵiJ�!̎���~�p�7|-�M��b��L.�Fj���^�6uI��Zf�[�ָX���@�^Z���<}�U�Z�˪M�@#)8݆�8k���,��Y�|GNO1V`�]M�2�Db�ૺ`}�>hx��>k�Ʊt�-IC�Gq�N�$Г�Tgi'��a���� c�I/T���/���x��6��� �٩����m�BR�>�(3	��5���$�^6���w��D�ۑ'�0�����
�pERPyL�(�D�65���/C�$�j�
0���J)����߂�E־}y�R�,�KJiٿN�d�g���y��s�-!�����^}���r��`�[�1�e/���-��7VX��0v�{u9o��?z�?���8ٵYa�ͨf���p����ӆ�l~�(gmI�<��>��;
��+P�i���a44�,���U����Z�62Pu<1�|�i��-�;�/��R�@w���4�w��9^9�M���B�2�s��
�e 7Q��Q�U)w��� pF�`�����]�Z����� &4�ŗi�l��+K�F~�{y��C�-v��y̅iMx_�k+��BF�u�<�q�w.��o�=�@�U��갾Q�W�Q�8�2��7�g}���$�.R����U�����@$O��Z=mt^u�V��/o���+x�l"լ�wI3_�[�Wԣ�/���+_5}�D��C�$����▿��Of�(�u`#n�O��9��W���g4�)��2N���{*������X�J:�����(�d;�J����'^;z�K�1�~�� �Č��	��r2�' 4�c�$q(����#�^n���%�Bhjن�>�ϸW#��"i��c��������5J�kJ�5�(y�6-�f݃�W�cb���&��G��J�m�Gu�)����V߻:�=���v�%��#��6�KhK	� �C�u��85��u���{	_���ɨ���H�^�&]W�/�-=ŧҤ[l�f�:�i�N-f��GA~q�u����7�]i��I�*�K��M~q�^#5�t�������	�y5z �@� ���t)(�c�ێ���j�J�P�����oB[d#8LׯH�⻼�8{�I���yl��2˒��%E&�o�oK��t��ޮ~X�_z�8�|�d�6�Í��PW��1\��h�۵�漦���\�)����w�_�c�"���B�va:�� �2�W���';	�~͟����
5RE�dJ�����ZK+��`41EC�%ߺ��k_���^��1�D����!�G5�͑'`hs炠3�y�+l8۱��������[�/[v<�!k��Y���T9K�k���'Ǆ�x��J�d�8I$�NU�QA؇Jd��6�:6�����(�l���}��n�W�l�JVOݫS�n�Q8L�K�&ĔA{����|A��
�>k6�VLNq���*����x�#���b@9���*����i2������<}�mF�ة����U�'I��#+{�L�P4}�+�������268�)3��:(�-!U��^]RcC1�F��lƒu�$��N��A]�������D���W������S���BMw�/1��I�I�'h$�|:鏁�����G�[������@�O��~δ �Ҫ!g� �4�Q���~F��/��E�\�'�W�),���J�2�u|�Q�j<�����͜9:L7�)U��	����5��/��}�ⰾN���UL,u#�'n�g��g�[x�o�ˇg�m:�OPq��Ԗj�DY�����ӡ���� :�����q��
�r���0���[NP`�������"~J.w���)>�~�XpHeZI%Q>�F�%����~N��f�hx��S	��a��[��|0ܦ��0�|���c�1*B�?�XJS��,�/FJ��Q.bp��$�8=���h��i�oD�σ�$U�.  �W���b�� ��FZ��O�9�=
�sʸt{A�'	fy����O�����a;�&bX�{�-��~�#({e8̃J�!�r�P6;�@���aiQƜ�FxT�����v �dw N�}a�3�6���^����
���%���tM�8�6��b$  �I�V�9 �F%X@��E3�%������]�DY��J+T������S��_Q��1l]L�e���;�
Eנ���kDFj��d�/Ϡ��@��Ρ!!�n>_���	�r��5]�H��\�b�|�̢(�0X�S�s���F$�`2����{Jk�ʁ[6��V�zH�y�=��QP�!
� ɻ*��gb�-����-}�?�DGX�oc��
��F��P�W�o�h7�m	�e,�b�k��Ą�h<%�������ʶ�<Q`���Z"/�Տg�0^�{���a�s%���l�������Q�P�"�ߛ�R�
�լm��"y9A=�@xb��
�;ٶ��#�y��,?�r���lBS��f��9J;��.�k�埰_�yf��\��4�g=s%���
,�D�ԻJ���d��m�1N��k����k������;��~"��6��l��iD�}!�qE�����S��5�����V���ب�A��%���e񺯊�YK>��N����D�����B��(�14X���Y�i6����F��s%{.3ᚏ��������0�f�+0�~���:�9����D��\�#�R�?w,�j��l�P�/l����|� cA'ЦG�{U��X�Z!&=�^���\�,�WH�Ls;9��w�Dn��sC\��LH���Bw��T��5��H�4�J���r�+x*ܬ#dl�,�S�k!���_a��O��5�S�"}���vL�	r��ï�R�������P�ǳ���"�E�{��i0�A��=��`����U�59KT+�H� ��0Uf.��#3	�����]��F���P8���/��{����%���fC�ei�}ɾ�]c�¨�-%*#�d#!	E�6#K��}_~����^��ԕ�>���k��y�i,l�E��p�h�:�Qe5��4�Ԋ?ߞ�mw*�t����mM���DYfg_���d����O�u.�J���'r������bA�A�js���� �Ӏh5�SC+���ʟ���8���Φƫi>H�@1ʽ"Q|����k,,�`�$�� *�ߒ]i�ʿ�~J���S�м3 �YF�+'�����`RE����>���H�f��B� p�;��Bo�vwQ��K-x���92w6�Q �,P��u���K��A����i�)!��C�3!�:��+��nԠ���n��ݷ�?9�-!��;43m�s�V�.V�AJ�;�"����]������'��� ���n�*��#�S�M�@��Op�Kp@�ټg���nnZ�w���/���3xV,x�fyl�-��R�����L�$P.�*s;�{s�(�s_@o�b�����&\����}ޠj	{Z׿�ê�.`��w7��{l.��ć�,C��O��c"}80�aնH�@_���xm�A���|o;$Q���r�R����'�
��N���sq8I~p�P6I��,@D����7;)�^���r��u��y��Yz����Yi�awO=D�P0}\/G稙AV��VS[����n��J���]�*KMBI��9��LJ8]���<��31��CN��N<
�+@���Dۄ�|��+��m��7+���W$s��W�5WQ^�ʹ���A��7\���Hh���f�d��^V�qm��^~ {}����T�+jmQ�<��'����� W;^�	Oɾ�u���jw�m���1�p�!�+��#���Ns��'��;z�s���������%���K'��{zz S��P�K���"�7�i��q�ҽn�8%�7A:��M�j��!�:�;��*��e!SU�	\��o�9f���)���u�c��R�#3�oF� �8������@G���-�ꑀ(M.f����3$UB%!Y�C��|Dn�	f��j˭���왯�6��a��7L�DlAy^ڿr%�\.����|?���Jc��M<%^�m�^�ؼ
 �4)�a݂�FN}N����a��f�9h+=�ҕ�(��R��|>�*S����ࣰ�\�O�{W� j!� D��������]���SBJ���,?G�܄���'�ɒ�ơ+��ӫ�n2��������"獀�����ujN��>�ۍ�X�4�.To�м��r&�M��їV��*tQ���@�e$k�2��Ea�j
P�q��y_����X�{-f0��c�����x	��ᖼ�eEM�BJg��!���֗i�� �~�$�R;���=����'?���
�>�����|�j�Z��.Q�D��R}Z�͖'?��>�,e��&
�+˛v���)n]�]-�����D$'z���y?<_x��C�X��]HyEj�2�,�`6�7��mM�����d��
�e�4���ܦG�o
�=x��r�	��TN������#��@=�r]L�>/���X��隇���,�QdzUϸ��e��@ ���������u!��h]�0���"��	J�zru�^:)J����|�f4�g���ɺ��W��,`�⽻Pc��NA=1��ح�����'g�O�@r�T��?���F�?�~�@�b�=�T�6DKL~�Y������5��� �F�ų'�e���ϟ!F�=�T���P�:���{"��|̃i>j�Rb��m�}Qjʗͫ�P �
�J ��v0��2r���;��r[bZ�@�e��ua�.�ToQ���D�l�Őc0t����jPҋ���&�d���!�H9he/��`f�s��>�8�/�,��?m�FhO��D	��v�����dʔyv�/�X��La��k���_K$�RV��x�IYEW_u���.[Z���Q�3^R�$��]=�=�҃`?���̾��3G���P�;/��f�(fiN�?SW�%N �j�����^�d_�5F�1�Rs G���S����9>����,���y<S�QKՋ��yM�FMsy�;'��#]3�7;{�u]�:��3_H��'%�k�\�t9�����RF {Ӹ#P. �xx�n��Y�e�
�~�,F:"LQJtCG���������ј��D!i�ٞ���:�&�܉.}!�w�>�>���.cn���ׁK����_O�l��o7���X*���8��%���mW��,� s�.��<�n\r%Jϯ�"�hJBQY�l�B
���t���)8V���f���ḻ���{���C{UlMG�M�i���}G�y�)��0�a1U�Y+�ޠ1�б�RA�fd��i8�G��1䘃��7w��i9j�dQ6��aє۟��N;v��?���Fy7�	���Ʒ���E�;v�z�����;n������x�K����--d��	,~��,�g���/�%TO�&9��oe��G�I�i7n.�p�wd��AJq!3���S�6tU�M���hzb����azQ� �7'$���r��qE��џ�����},�e���[�t?# ���W^QS�s:yV)������l��S�Y&��^�Z�7�hXIY�X��u�"��J�P_
n����#�x���'��sTr+������8HE�9�|�5b��$@8/er1c��(��|�qIk���ZW���J�$O�h懓�8iYI��+,m���o�/N�@$u{)��X(�p�b]Z�CG�cs�m��J.[Bx�?��"ק@1����KԈv(���XQ�P�^�W��ϻ��5(��B�Y����i$���E0�����g�*<�EVY�Wϳ�sS�_��3::zT�^#�ǦɅb�;�QjX��%���Qa�D���G���cJ�TF�^���d:�I��P�>�u��̈��U�@��p�෼G�ۅ�P����x��z?�9�2-���T����G�
���b��ʖ��B�k���v����}�@|<Aj|��	��N�s�r+�1z'a���"���m�m���"Z}�&;R ^�� ���B��Š"�s<[�tb��^�B� �>^)=�C䝛� s��p�2Rͫ�i�BT]���xux<HP50�ve�q�%mM[�W�^�Sٽ���h��E	Q�Ά_�ۛ�쫺��L�$�Oz�a��]�y�OInM���L��:{�*7��Ř�㣡0@�����R� a�8�:����])����"YV�f�Q:)0�!����OC;�dG�\J:+U�q�����(�[e���ӣv�!RS[�~��l�K��/$�u�����$$^��(�$�vx����♸�>L��:;��5��p���>����Dw{�I�  aW�e\q��xa+�O�?DKЖ[��l�������-����3�u4��)%��ב-[>�Ŀ��լ���x@6YmM^�fg����ϥ�����_K��d�ypZ�Dqril����j�Q�B��ӊ_��/�typ �2���Ж:�a�:�'0�N}��D�$����c�=�����b����D�6m�Mhj���Y(Q���p�)P }±�7�u�ӗ�5�5�*���X��a�x��h�ۯ�_���%C�Pt����`�"�:E�Ly�跂��"S^�s����͗�	�X�#9H�w(E���ZJ"r�"�F��:�pV=���n
"ݬjN��w���T#��6�8��ٰ��G�K!j��17]�9:�Z�
4��׮��Te�9��������wfbS���J��Xi��'�&n������֗�B�?�ٵ��J�N�'��� pv�j>��̸"��Y
gu��<�R�Ͳ6L('��a��%Y���T9���p�ҦH�O�e=�R�aQq�v�"Za�
���3�m嶘�A��k\��0eO�]b�NÔ���:vh?�e+Υ��i���|M>Ӈ��c��Ē��t�����>�,��q��ocϡ0��[������_��R������,�uf�pַ��|:A0��CA>����Vx�maz�	��x�MD�*H�p>�/����}V�٦X��\�VU����(FcVr�l2nK��@`?n�з6�r�4.d���%�j:�%tR�*ƥ~V�S��D+9�}���g0����{Z�6`�
u��BI<������EÛ��hnR2n�����8�&/C�b�H�(�Q�-����oiM�%T�ky=ۮq��(v@.^Ӥ�:}y �V��.?1���� 9���y�<'X������>���Ÿ��W%��h+�oj��2���ZC�N1[��2���¬� Lልo�U~�c7�h&�o�����B���L,��ن��ٺ���EZ�r�&�;$_��o�2�x�"����y�#�'�mRu�֎懎�@1�𙔺i�On�\�0{���LE/MݯHЍWc�K��
BZ�p���ᏼL���gwt�7��`
��;i��fώ�k��O�jbY
����-Yv�1$Yܐb2�
$H�4~��!O\^7������<ֽ�F�3am�K� D����>�;�ZPm���3�kotE�})>mQ�4nycn$�Q�vU(wh����VAg���?�1OJc
�A�=H;@�u��X�������=��SE�q�Iiۓ;���!�r�*��Ƴ�GM�����ulp�	 	_�4�(R6��(��ǎd@�����mb�U.|5�
mO��󖦚��J"ذ8F 2��z 1�b/b�ŧ���O?z�$$�Us�&{��}�B���ޭ�i\-�5a��s���)D�a���8��!��z��-K�<��-�W��#/�G\#oTbY�����F@��ý�w�8](��7�J0K�ݪ�w��3'{�)ϻ�`�K~��z�Qw��/�� �R4a�駜K{��5r��vM! Z+�p�������ӈM��*=�4�����&�O���:����?��{�������3��<V�Y	�����]Pi�����4�U�Ƈ�LZVtitF�XQ�d�x�`�
��)��<��z�	M�]E��� ��K�"�yA͠s�z����:�b̰���I�i��w�,�dU��j��F�Ϊ��`n7o��^��5�qO� I{��j�i<�F|��@�j{���o�Z_��d�H�Ķ�Y��������k\x�w����K��d�>+���.��vHz]�:�vO�B�H�2����S=*	�T0��3-u�v'����7n�qwY����$ z�ޫg�һ�ݨ)P�;���W�n ir��<u��kT�+��d!�b?<o�`ꗱ�T�p��{���|������E���oL��k��9�-o�hStyeA���LtƦ�P�j}��!/ͺ$-q_��c�IH�C`��i������	�)���iY�f%�����zfQ�F|Y��\FE`�[*��"�E�.�èB�g�2��b���'���cG���`��QBp��mH��>U��2Xp��ǯN�P��n#k��y �d[�3-�iJ:��"Y�4���˂a������g��=����*R����yr]���*Yy`�<`�`7{�� /Hy\�a�Ɵj�Ú�}ָ:Pt)��,�=��L�
?����z,y��gf�~�D5��oofy+1�3�yMӡ���%�Xn�z��ʚ��ˮbh���b�O3h��%^�Sq��	a ��=7(�x&6A�lT5���ٽI��ZBV���H�jͣ�Y�>��AQ \y�P�]���3S�������]��w�R�e�J��A����V?�:�5�rZ����|e�[lk[���q��iGܘ��'��;���2"���P��1����3ĳ@�>��k�,�\��pEk��ф�x q�4NKL��q�/�0)Ց��"�)������/�$�Y�ƴ^=A��z��U���z�}~�q]̡U��d�Y?�)��Hߺ���y({�8��n揤:�tB�_�(�L4$��<�O}�E��{mﯰ��`�y�vv��_Sϖ�`��1>[Z X����\�H�|,��k�'��y���!�6Jv�;�j�l�s-�7KI�XFv�
�u����h9���X�>�+Ϳ'@u�ɢ�UQ���Լ�[�H����#���J_
G�=�DH�]���i#,��k��q�h����gP��I�:��A�62<��&7���BI�Y���A�Vt�P#����bo6�	n�� 4��Q��B&��&������EK="2�W,�~N{����m�A�)R�����0��?�bM�@�|�2h0�o��\�ȑ�A6@oO�`����^��}�����u���w3�x4-b07��Ӝ���e#'�T��gu �*����Zg�_���O~ڐg�j��<�x�q�Ao�����y�j?0���Y�z+�{)8��,��x>(L ��@f>� �:qI./��q�a{�l�>D�:��O#T�P�df�nC�r�]��gI@�&NMv�@�F"q�F ��7~z�i�ɟ`P� �v�n�w;T���)�N�y����#-G��E`�o�+�` ̟�>{4����>�H9l]�A�C�l�&0���Wn�a��'�+�^��iG����F_�g'3����p0�v���j{�f���Q��I�P�i��*HxՒ��hc*����~b+��Q��P~�T���W�&��H`v�4VR7kuҨ`
��{����_gP����&�s��E�}>O=yȲH�4,=�@Q��O�f���������oщ��*#3a�{n�=�sh!;�x��_�C�"*�Ť,�w(Z�T�;�	�2�����oB��#,J��h57��֋�$?:=�F���y0��/T����l�D���"J���67�Hu�[�@�7Q���7��+i(��;r������W�;\4Ү?����CJ��)����jL^+#�v[C�Pfl2��5Pi>,/>�_���B ���R~۾B�p壻��iӸ��5����PR+kQS�n��/Fn�B����1}:��ӈ u/9�K}��?�L*�IB���Uw��Go$��^���̽#�0�ϒ���_l%�#A�g����E�:XaЀ�}��������k�g�r�Kg�VG��5|m�2x!��5��OR�=md:��{���%~�dkH��	�#��[���r�_�ڄD?����l�( 5p.$?�*9ѻ��Ч��Z�����>��veϋb�\v]0[����V��Í�5���=�20�bI13����=B��v�$ߡz������X��ca>���
�Pd?�N�3�u]�s���H�xZSo!��=g�vstz��E�����`�Am��@z3{GE���%h�FM���w�3��+�$<���{�:B���_���@ӡ����U#鏲�3�V�Ԕ�����2�&�r�&7����ѐ���3D}�}!*K[���Kʧ��#�m{6���7��3O�Z��kr��gO{���Q��, 
��y:�7P��Pc�+����45~p����mp�dme�5%[Ce�E�d �gbRa\U}D��bTN�j����R������8|������w�8�j�<[-ǹc7BYO��\�����A>��Z������k�f�\� �I2X���y��.w|�)<��S�������
��!0�E�������R�_��|�W'��� H�2��po�(��x]#/UFʩ��V�̹�"���^�+ Qn���>��{����R�)%�7�֯+X�#��Z0T�U��Y�}�S�"D��a��^$�k�E4�v��~g�у�bS��1���RL�Y��g�ٻ삉wv�0���<m����4�/K�9���J��R�8��94)����Ũ�cu{��~�ә��3���;s��\�%�^L�� ��bWP5��u�Fz
�ǒ�j`�d5U{�F�����O�zg����&�`�9�p�e���j�d�Z���1�cfӟ��p�o�2�>���)i�_�x���X� � ���$uzc\�)!9/F;�jEgqa��@3|�&x9Tvn��f�w�i���	�l����Ҟ�0�Oj���y�M��q���@����I�m~w���Ց'X=Ýf����Z����7�=,��tMѤ�C 9��5%�c���un�)�Fw��}>�����܆��w>���	�8Rd����d��Chq�<~Á@%�<<t��DX<�HI�#���5�>��$.��<ñx�[��龍l�Co:%���*���$ HF���?��Yޕ��K�����x��:L.����ЄL&��7�:�Of%�fM��2rT��@n��)���0
�Tm�����sj�����[#���26�����e�l��q�.G�e�Bȳb$��'
��Nу��n1i���ֺj.���X��$�� ��nsk6L�2��_� 8_h� ���:Y)v@��s��x�JX+ʳo111�v�^�@%�*5���3���p�c��_c���\W��5 qu��s~���'5�e�"��8Π�[�$9��/v�ߠ�ђpw$��H,Ҩ?�Q����ɺ+�>s} ƍ*��E���0ﱈVo�P5Hg���s�:��A�]�:���+f�gg�E�6/G���_��m9!EE�#��/"is^�{�sѶU��e��E��*G7��)`�@EձI�I&M9�(7OF2F�]̣������X�>���c�˾.<Q�[�L),�?d2{�isc��!������*�16�]k�P���̠�cpaq�hƟ6�jb�T���T �fy����f�Pԥ'?�~`nu����%�4��#&>������ЋP�u��X�M*qN�!q>���`��)�ښM��gE���Jg�m�ͫ%i'��p}����:knV��bO��Em%[��4n�+a����>=���H�nKG7�ڪL�h�C�5��o1���b�n�ׂ��TU�=��������(��
��%+�i+&��7��h�a�H�0k潻J{=='�[E7ި
�[X\W���.ǯ|�Ak
�Ǚ��4��������*@ӷ�$%G�$�b�ڜR�t��{�ڄ'
���!�W-@�O��S{���~Ku)D}�-;k�*�m�����Ru3BU�t�c��i���>��U�RCk���h6�w�;|[<�L˾a~sYJ$��P���6��բ�`}x�fS�V�y�Fk�`7+N�g������BN)r�p*� a�{D�����o@�]�172��#�5����z��#yy0U�C��vZ�c�,��*�є�l�ە���n�&�F^�_Zpc�G5�����^	���Y���ɫ�r����FX�)уg��b�ŅL�&r� ������D��H��
�O�H|�e5����WY��T�N�4�ą[a;����?������yE�1��H�Fצ�r���M KA��i˄Ռ\ڕ�Q6j���YR�Y�19��K���hf�b�NYm�Q��/-�����<�C:�iJ\�[H��FB��/�˓��4�����Z����bIQ����eY�Y嬀��<�Kk2 <`*���W�4����l��}~L�K�_Ɠ
]�v���of�#����C�P;5ۂ������u6�!>�?�(ٔ��>w����M��+b����V.�HJۮ��@5q����]�	��qǸ!P��P���[w��� 
��Y�F/�ا�����Z�>��_w���oi#��<{G��&��1)���u��]B�m��	ּ7#A*�-X�U7���V�9u5��y(4v�ă�C��v�\�,Ԕ� �c�W%c���
�-���Љ�3O����Z�|���v��fo.�����>�M�x���&�[y��f��S�M��.�����ZQқ���#5ɹ�Q.����-[��� a��Q��5��#�#@_��O��,=d�j=��'��oƺ��Q/\j�O� �{"�D�2����/��׃-�����Vb�7�pV�fv"
�-�ܑ�[���ZS��jҷ</7wGñ��2�Z_ RbN����cK-��t,-*�) �ӻg��jMv}R���J^=�]�ɔ8Z�d�
����\��R*�Z"7U+B���If�U�f�{c�C�{����Q���@��;��
T2�l���*T��]��a���ތ������JᑬPB@v�z2f�¼̆�R�м��V�}L��q�5��ٺ�F����<,[���E�=��	n�"ˡ"�������( �K��G��C�幥��m����"�����9!��|1ȑYf#��Li���*��<6�V��H}�Hӻ6mj-�§��jBl9�Yԉ��k8ܡ��ы4Us<_v�%đI���R�����AG��-LAY��V��zŭ�3\����þ�m$��{�����z�e:#�+4v�~��[�m��!��;'9� zp�΃����#;�e��U���c��uP��g	�LC5Q�-��]��jp�Wvg�I�U�9u��ï��z+5k�ut����1uu�půs2��^����DX��aUڼ�ld�鬧WҨaE �G��x��������TQ��1F��{H"���4���+�o�P�������/!�'�o-�Q�
M�FT~�}�y��sU���8��(f��`�."a[�t[j��������T5w8+i�U��]{4��Y��ƾ_vi���? z�u���׶��_���M�ҋE0��x�oN�/��>�� 7:����� ���׈p=l�����΀*g[+��(μ�.���7�:�N�s��}�����V�A\�֓��jd�pgVV�����a����=JCs��Q�sf0��Q��#Ì�?~%���+���3;���}<�����tM�cy����A<$	_��xgu�z�^�*TPϲ�Ok��&�l���>ͷQH���Y?�d��v�}r3܍Bh�>
��+i�/&��	��Z�<��\�?w�X]t([�8��`����Qlf�)�f�3�B��#ic������n�on�(7g�*�G;?<�whqGJ$Ǫ�qY
���<����N��)G��{׼{~D'+W�΀��
��󀟆ktu5im%��Wb�]-�۬�֟?��/%֓����Ê	� ���7���i���2�u�[P����j%Q5&;�J5�HJ�-<�a�|����'5��cr-]Gz�B�X����hX��!�A�7�%��H�J֥���c'p
����Tpb���M_�[!h`5�O�f�MF�]t����|���]���ӳ��c�K���z�^�~w�I'��K���c����J��):������Xz�	�����6!�?�M��6t�w��-3��I!v~�v2�s!x�/�+2�����3�g��i���%��;���W��"/ !Ժ����3Z\W�E g�w;6��bJƖ���O0q��T�jo/�!������Hn�j�+���/�V��k$���f��y ����<Kq�Y��.�j"����t��L2���4+S��|=jo������D���?t��N]?�V tZ���n���Y�&<\�|��'j�����4YYh�(|�3� x$��P�����
1J�x����qJ�FN�fH���rt�@�\>di+�A=�G�Z�_�x�_�UM���/��QI�� �;,�UVn�Jc?�l0/{�r��Y8kx�mt�Z�6�)�>�z��+H��M��S���}=sŲ�,]>�m�kkk��`��VW��y�Q��1��6��H"���	W/��hn6��ΐͥ�
|�.��,|�\K��z?���b���8W�ҶPp��U�������RH��\2�b'�����Wj���*�Ԉ`��Sx��������f��(.k��yb.d��尮��6�q*�,�yK�_HM;��K�qo�sߵ#��@��R�M#��Q�?�uҨ�����ed�Z��C���p�aYA{�m9��B�F�Q}����o�hը����'�����>�	��1�٥�JC�cXQۚ0��ѻ���x��T\�H�� oX��N����S��?%��UT*�㭕#�q�����jꜬ>n5��mO����Y5L�v�@êjj?&V�|ˬ�[�������1U.��q0�O~�Sᡭ��z<n�����`"�����t���gЈ����Ua!|�x^��7i����8>�,����y�vA9P@�z�׬$�j*�
��D�H�����&�~�l�|V��@�~㿄�[�`��O<�(�d�߲�Dv]F��P
��B��7�zX�,������a1K`
_�����4�u���N���ԝc���K}�,r���~u���p��,�}�e ��o]85;�Ĕ�"�@�K��bK�ɡ�죸�e���N�|�J�3n��r�`R�صnmc�iW688t�kCOO=[�u�2��p�x�K�؇��|\62Yl�O���0����]�fjʯ��󦿘`hX�~��G�p5�i4�]=�:��
������:F�^?�fNn�t�pIG"ǹ�>,vo����a��?>�[����5�PJ��Ћ\}S�����	FE��cZ�s�[(b:-lG��]�艠#��/񷜁9tX`,��?���>�4�i%Y� h> 1ZY��B1Mݥ��R��v:�8SR��F��Y�~0���mۨ`@>Z�ٙ�s�<񭭩�?�J��m� ���gve{]���i��ͼ߻������q)V�5�A���#l�}s��"�W�`��s��,l�;�c ����]�kdK�k�ǎ�.!�;���\�hX�8�/��6^^
�eg瞮�2���S���c�E�s��JM�KAHX��߰αc�ﾵ�{۴�&�jc��b]�Kɤ��9k�R>�$�k#���+����#M LJ�����ƞ����V8tc���A͖�>t�h����#Y����k�xl����v�w�����Y����ް��s����;��R��'[��䥜�k��X���/��r�]�ģ������^���`)�	�VA��Yֲ��׳
�߭z}��}/�bh��W�,y����VS��k�eD�����o�7[/,	A��n3�NO�9��ïBWy����G����Ѧ0<s��(P��Hp3��X�\��`�L���A��J����`%%H��-����|���]��[�粨ۃ��vL�<�1Ʒ�L�6��?̵W,��I)H�\7���<_���0\üԥ��ɝ�k�S�E�.p_۹V�t�C�΍}��#WC;��']W/pN�5 ��#�Շ&��cgd���`�7n��4�����4���>�
��i����v�y�<�]E�y�^�x���B��~���GT>k�cV�06�~j�s���ŴlP>�Ý;[Ŋ,��"�C�g�.{�~\ы�(�%01ݥ�T7���������ū+s�g��p,b�rҠ�����_	QF�{�1���&n��6�I1¸b��������, �f0��S�_S�&�:�1�;VwP��^�@�ha��C�q	9���t�������F�&���},��u�C�n²�R�t��OPY�U�U���K��;v�?TM2����y�Pw}������-������,¹	v�rɫ��)�@����K���^��i3Z��A��v3ͭ��}�C�o���k���k���4X���뫮#'���1W�5�x6�� ��ܼ�����˓m�e�PF�����z��ʍ$��7��KJ>-#��=��i�K�5���ԡ� `n��K���k��B7�K�KK0���b}��T}\��7�6��-c���pw���e�� �?Z<����5Pn#~|����vM~݌��gS�`�Y�8��\Mn�=gZ�aչ�RZV�T�D�#������7�x�0�F��wv���N}N|\�t�י)�o�w�9��cc�I�_���c���_���x��8u��6������^�S�98�"D�nQm�E:\���{i��|��O�^g�~)J�S��r�K!�=���S��m�K�8?[�G�/��:�E��`>����>0�� ~��A���L˟��T�>:#lI��D��l��ͺ�1��諔#e7F~<>Gx�-#~�Rד'4�R�:4F���̓�Ca�;C�^�~E<�2m1�����h'�Ӯ�T�o<�Ɠ�[�D?0`SU��Y�n�Qz~?���4c+*ԡ���A�ǃ�h�Ɠ������}�q�hR0t/%�!�������i@ּ�>;��}��V7+	��ƚ������w<,�����Kg64�a�`R��Y{S�������wR�'+�[�'�`��et��*-̍�咱�����?��D^�(V���v��3H�z��2�T8Rs|��"�:���ˁ�kg?�D����?����{���O�X�#89�M��Ժ��WU�G���T8��� <�+�,X�'��ݮ�[�+r�K�A|�N�>y �U{χ�Z��_�2�h���k0��O���/<aDS�U���������Z�lJ��ol͏�m�U���V��Vmɳ;�����pA��m��P�/j@:_�'so��g���54��H�ռ�F���nJ��<wO_�/Vgˠ�a��.��J�[2�ZY�l-�h ��
���V�
�32���T��$��M�w�G�`�z   �ݭ���f�7��&�qz���r��/6���я:򃞃�hk��g����NNm;J時�Nt��Rn����Ϳ�*�"7���"�"N�0��s�,�LG��V���/-ۨ&�'~>�;����R�Q��H{bIN���� �mG�f���*[�R�5�Z���K��i��!z��b+e��;o��x������$$��0�)t^���4��_��+-[z�5��VS�wW��ʑ���x]�;��2�@L�D�?R�����*e|yrg\E)�x��)��DV����������bP�p1�����U0�N�����q�̕���ʷ���0��G���F"Q��^7�a0�^@t���%��[�ԽN�<s��	kߨ�j�J���dM�S�����d"9�����Y*n m������l���Gg/��mZ�f�6|����N�p)hƥ���z���+V��~s�t�	02��h����FX(gŗ[��Ġ�Z����Ɇ���F�(+�H������I���/��e;JԘ�V}T�q{���(��e�g~\BO�6����(:�n�k6��e���99��}��.���Ҥ�%��[1�jo8 s�	�����f�ry-t'=P�H0����H��9u�,��IH��F��tcN�?j����*�������S��-��'�����3x~~~���у�(�8��0���z��;p�k)����D%}y�����}\}���T��E���h��#:�A��r�����UN��[R�}�x{�=���,,~N�@
�S�iwZX"�?][��$�u���ꕘ���u{�y��{��|N���X����qm}��Y7+r�UQ��QjX8�՘��{���5;6�`\�B#�`��T9$]�O��Q�LB�ԩ�T]x01>�vR@����UyI��P��O���o�
.�k�P4�}�E�eW��̬���77����wO��UG���h-�oW��X%�L��!P����{�5�^w庻%{;=���|}MF��7WLJ���:cW�|X�8����w�糪���]r���;��6�Ѽl)"o���,.Vy��P�z� I�2Q�E|aJ��rh�jGW�A�&q��.ǈ%��T�P��.�|x�g=%������^ڒ����lQ� O��m���%P҄,����||�XG�w8����<��\[��۲4-f��<���@�>��c��Ѷ�C#*t��$�O�w�6��]��K�ђ�s~�fW;q)3��>�C�Y�����A-�Ǜ�S��>V����j�9���
#N����&�d�n_�7��6|�$��;��*ka<�/� �g�D���ڏb�\�/`u�v>�O�15�����k��;v%� �c���{d�d�9���c�_H��6Qp�\���p��kx>X���5G�k4Nm�P`�E�Tt8�^��O|���ީE-,:<gHB�'5��Q$I�I��6&��O{��ׁK;0��$�ޒ��!�;�(�^kZ����Ky�Z��N�jhOn���J\�G0�!O5�����y!��������E�ꀢwS���&�o�>̓�17�l�_�[�](�
�"_�ʢ>��cϊ�C��À!�	zy��8c{\�"Y�,���#"����o���}�֒��+t%��H��o�4(��?K~G
��-@�?��rG�Z����P4=�'��ܰ ��û���`��Kp&�2Z�T����X*��-v����=-��
���g�'������䨰lה�)]�MN�K�"��A[�{��.�|����4C����b���%JTY[[j�>��S-�Z[�>V�b�18�=w6QA	,`?:�f�֯pm���#�+�.�FO7�Y����T�V��O����r�l���Ӱ��2�$l��.Շng�]|�z\�W�2K��?1=�[�BK���������:�quq�c6���ʨ��IByyC�wq���z@�wp�/ZIi��N���:���.SUE��Q?w��5:��\�����;Hh8:܃�HPsE	�o����]���_]}���I(��*J%��5P�ꕾ�:kk��JsZL�l��y�4WS,N��66p	��
MO�y�L�� ˶x��~=:�5:ܴ��h�vw�
��u��W�X�T��V����u@�W)��/=k��N�����TR:虓�P�i9������|�/�ˠ}�7�Ι��U`�1�&�����b�h{B����Q論�_��=q5�����Gj���*V�;e��ȹ��Ζ��dkZQx�oҴg����M�>������+� k�v��њ0cK����*�x������ǆ��{wq��w��s��4�ͥN��pxe��w8�k?������@�{ۓ	g4˻`�s(Ԇ@sҘ�\����l�>`0Z1x��������b]i��۴^�'����it�jV��\�rs`��\�Bu���m�	mL��f*��=7���[5s��]۵����i��������.q��)�ˎz(<��`h���P��O�o�s��'Iʰ�����w�ؽ���x@�ۤ�O�>ͷ\���wc ��2ld��?��S�˖�1 �?��W|��j�|h�m��^>.NʊU��W�0�v�ua�p���X忨�A�U��^c%�[��&�߅z1���xJ��9Ƹ�y�����RCS̴���V �߷����2��k�� e�tW���MgU�~�!Ei%��E���A��[���A�[$�F����F����=���χ��쳯k���{�;߫,�2����H۝5��7Z��Y�VF7��^�k���+�B��x҆O�R���LWr����IG���;,�Ŝ(�?,�Ṉ��~ޖbtr�}��󇏱��=�
{�ҲC y�Y���a�Kt�[��@?O^>$��x��\��V�����7���=ϳ���*�W@|H��zz'Wm��4��P������܌��|�Pd:a~�]v��M�VI��$���^s�i�X"58��xzz� M�	�����=�v�=��n?~�����C���q��/=�K_O����hr�s��}�B������U���59攢򭖓7��mc�f�m4L^j�-����j�jJ�8o}=1� ��wv6�g��c��G��|�e]��SD1H��y��V�H/x�bDc��t]ʿ3i5��vC���&T�y�C��5N �)��QI
��C���DY����@�o3ޥi�$�/^���4����z1@��V2���jb���i���������i�/��ތִ��̧�s��ܾJ��#,
�I��n�9�����2 ]ѿ�Ж�߈����G.��x&�j������ROk���6ZVx�#�=� 7�:�&�*Z���)U���R��Lmd�]9ڢϑ��d�X?�z�e5��-����	��E�iY�z�����s��q�>ŬvY722G���k�+ú����:F�:�pd��p|����Aj;,���m�ڇ.g5�Jļ&K��0���v��H���V@5��T�J%B�"u������golile%'���ϥp�7��s���=��iY��8����#�p:���L"_�=C���s�^Q_�.�;~D�!�|LY���n��U�&�
�a�1��6��!]�ߙ/]'��hS�����������_Dy�5P`�j`����N�8X�UM�z"�{U�5�p�,8�.I�L��_���߿��q�Ve�EO�O�KT��&W��������x��'%�����K&���	�o��D��%k�>8v3@�pU�l��d�
L�LGߏsJ�k���<c��R���z�4����l����k�=O˟��.u��|�8|l_ڈӯ�bp����J����ݿ[�ؙ��ݥg��"+tm��k�m��A3��]l3��~.�����~~v�S,���~�8u�;\O�j��X?�	W�5$���o��S���~�V�����ݲ�m�2B���d.56iG�m�\e<�D/ � ?@v��
���K��g�E���R��i�}p���0}�7/�O�g�N�$���5�����Q���H��ʩ����_� |�]"NQ@�1�!y7�n�ka߀7�KN;��1-�G8Gd����!��罓���,�����\��X�br�#��!�N1�h��\�m��q'��&�A����g. ��LF2b%�%3_�F{�F��a�����v&� �V�tU���I��F�fy��6z�L���(���og��lZ��AC��0C��0�+�ZN�~�s�¬s=�_w��pR֕�d>S�t���nS�����}��`����4Q� vN�6\��.��"$VւcU	ls~�^��Ĩ�l�F����	�����C���y�s�?c��v�߯=����,+��s޴�<4~��N��B���iF������+S슊}���1�gנ�� e�UWg?���.r؎�-��������aݏ�$��wD�{z�+�:�+��d	���G����p�`�"ȼ���P���ʭ��䎳���AhX�o���kŻ:7�(��I�<H8��	�@;��w�`D�	y�i�Z�F2{ڤ�tv�O�Q��o��p3�Ou4c�w����1h��m%�k���������㜇�LbD�eC�����ȶ�b���XIp���������9Ek�߂Q%�����u�1V�}�����A�">Ԋ��]�l�G"�Ӡ� ~)�myo�9+P�~�!��Z�̴�n�X?~Nz�O��_�֥�S��ʡ�����+��7�|�ꑙ�rƌ�]�ٮ��}���߃�{qN��Jr��T�^Z�Bw^T�N/A}�L��:/��X{��0�q�;�����������
2���:����T�ɬ�J�\z�0E����w��\]�a1�E,�C�62���Svk����d/�7i!��B���ʎ�<k5.}�?t;6��<�m���SL��5 ����;�:�G&��W�G�j�G`#����|��U��{^��TB��0)���&k�����mz$�N�Z�I�0hm�����AE��5�8x{�@�֝},Ϡ�R@�Kr����^���������I��sJ,��NayAԝ��Bqz2	?�� ɯ�B���e�t�ڿm�34Oɢ�P)q�Ęg]�0����u�ߧF��9��Wn�i��?��и���>֗�\���v�ױ1�������[��wd��ԟ�_~���s^"�ܷ�:an����{߸��K%:4̜kxo>�f�*S��t�g���1�(��b>�鿚*C�0sٺ.dG�丠]H�С{{�QXh��v����i�y���*�6����MC~��=�/B����.3�o8����&�c��2L�ֿ�Dd�6�`�4!+���jk� ������mqp�XG���*��}i�d�Bɑ���ς�����_c�h���dwW�-���Ps����e�|���'���P'��jV�>�'�6�C9}[��4$�1�9p,Aԫ��{7"�-�]4�I�Ƽ�B-��@��+8-2�����l�|Rd*�H��֥�L@u�á�#3�Mgݖ���_��T�JĦ���¢:��l��4�i]6~Ѻ:�����˟k޽�ʣ�8K�%~�}��;��Ct�|����#�VY�VxT��Uf�e-3ֿ`{)��2�#n�؆X�WV��5�>|�\�-=�0bՀ�ҞAQ�A�9�7ϧ�(�2���d�I���J���L��ǈ�<���l+?�QQ5���5JV���RS�aJ��{���VZ���[};ˠ-�b:c镊&���z,�0���\��ǣ�є�sYh��֛�����_����c䨬������R�>���۝벗�?h3�F���[+SŞ����rh���	��a�)H���I)x/��L���2�"?�A-6n��m��A���T	�2����Q�	��vދ�@�}���l�B�+7�w::+g[�չ��{k��i ��+�DC}�f��V�-��۫Ӏ1�|*?*!��sa��FP���3��U&�����`��&%e�mGr��[�m[+w���2����!��G�>k�t!$١H�����J��k�q��>,�W{ONk<<:zlD2�_�ONz<���Q�Eg�l�JsO�[MÎL%b��	�߰����b}WE�6�y��_ف#�� c�k7�qm�=���I�\�tG�[�����\l�����ȱ���f�V�S����!gக�Q[���)uЪ.��2f��9_�#i�^ tJ:LQ�_�z~�z�'-�=���vQ�a�xRXR^���	����shR�)�'kJ�Zs��l[�[�V]�B�1益q��f��Y���c'�.B�qK�q�����@�~��!��DEE��}^}
R>3�yCX��j �V$�;62|[�}�1^�N/C�dVOZn�;Z���lT�I�R�~�?௩YA=� ֨;b�T�΋:��V;$��a���x�j�c���k���p ��<A^�S0zCO���ο h�:�@�Fq懚�H򞪗7Q(���S�������T^j�>����D;�̊���b��0��Jl�������]><���ׯuUK�D��Aĝxhp��ߪ! tԉ}�+߻Rj��j0&�Zl��;]!��5���m��^�L?2���}rv�:U��3�Ώ?�t9�!2�Z��(\����c�Y7�uJ|�)�$cha��)n[�I@}�"9x�����4�}J���Ҳw� i�DD|�󞙆a�'%!q�A��Q/�G�1�sko�.�ϋ�v�C_��O��]H�tSUQ���nd�Sz/gm�Ĵ^�sl5������.'��塢$,�N�K���\rg�3��^ȝS���Qm�&[�$s7����7��p�8����JKqj�����I��b��󬵋T�l׋�n��7�^��%Ϭ7%��ht�Rʕg{{�|��|bb���s&*>�.N�b}���#Y81F�D��3<�)+�K4k\�ݴd��cK��-��ap��@%���Gy�� ������m@5����Z����-Ό�"��~�Y��c7D���ZG�x�W;c���ks%�ԖhE������D��"oCV���#y�V���C�B����a@��C(�CD$1\�c'Aȶ%7yu�'Χx$n�6��f��OF757˫��
�6�U��w���n�cm�u�v����-�J>�ɶ��[���蟲���s���C��H{��;���)�K�7��f�ұ��@-\j���a������D���p�����[����
*��ʸ��@�+rr}��t�b��z���Z�X��Y:��>�q�k���_����ҫ�fC!�'�ɯ��LfZ#��1q("Ex��� �tw~�Ŕtc` �4�T���o:cd=�9�Ix-������7�Lx���o众"�Lx��gT.wVt���i�o4�^f�����2�fY>�5Qri����O)3"aI�����!2�K��4��O�!9',�`�ۘ�B;>~(����W�Z��X��g�:����N�+=��	_('����u�_�r�����*�q0��j�N�l���L[M¸�Xdx!�W��i��X����1�xZD�T�}ڔt�����Z�a��['�#"zt9a�1����wO����_��������<`hQ��*q!�	�P�uz���A�	���(��W2��˱�DJ�9Jbz�6A6�.��7A�|i/�SK��$�/VV!M=��ڦ8��[��聳8��/�s�4nwW��f��A�X�l�GVm���<G�UC�`��"�1J䎜`��^������E������s�%r��݃�c������}*A����y��ᱵW�匛���8�=���M��[4�bB��O�f�v�ȸ��X����=LB���;�"E�<���M��Q��2��3K��,"Da���ת�p��.�����1�f}���TC�>:�uu9��s����2}������սo�0�#BEO�A��_/�
e๸�ʗ��S�a�ɜ�O8�VGA������X~������_��e��yWKF���a^�j��i����>��d�݇2An�&��6&/U�����7b��$�x�(�B]v։�tE&�z܄a��є%�fk��8P����M�{{/�S��z2%����u�mݙZ��9>��������!^�/�tGh$�;���W(nK:����4��cf���Ϩhu�����Zs�w߼����We&�$u9�{�~?��?�y�;(RvͻQ&���Ġ*��B2���T� ׼~R����CjF��DRa�1�����<� �C����.�v>�eOF�l��9rˤZ����1�eETux;������m}��[�y"��e,�j\4��HR�Ϙ3UV˕������7����FF*��?��,Ty��eX�6�ݹ���r�x�-^h���EK]��	{g�4�Xa��@
��`����g9��HG��\�рئ����w��CO �c����&��?���جY�t=�W&�m�����)Lm��\���2��^��Cȓ��w���BB �#C�m_�NLA|Iu�YmXK��z��e��o�[E���$%��0J#[�=�ga���z]_�:�N��S�K!�B��a3���MI(����o���}�����3�G�d%2�S���.9�/�T~Y$�$a�3x��HVL���Ցjn|���������ֽC3��҇�t9�LTP�4���J9'�:\��] ^��p�U�\�h)u��,�����5�"Gw��Y�cs��,y�W���SD�(�BW'��|�v�uǋ/&�}W &}_3=I��3ܖ���؃6�fe���V�Lk��_�@�a��Y�Ư致ȉ��������kyE���^�S�3a��>lz|�5Ж���]�������^̓fc����Ek�'��� ��G["��@�C�|����_kr�&aP��Eo�ŷc�q�[��;i���>46�H���RsW�<aէ\H��4��R���5��ūF����˹����끶���N20�>���s�����KA
�0���7�f_�`�	�z�Y����O
�?w�6 ��q� �~��}F��� 7�k�����Ŕ���Zc�~Ԝ�f[_z��tjH@8�]uo����V5����m���́~��y�&������w7TbOL�*y]x�=�'��SVl�U���ܸG��Q�I�,Y!]F�e\T��m8	���S呈/��^9�9[�1'��)A�Q�qDs���~p{���b�, ���RiȠ���؈:�=�3'��U���'�y���'|nO��r��7��,	yZk����ڟ���1�$;P��������~������"��PB��c^R)�إ�J0G��̰�5��x~�=�Z��+P���?�t���������K1%��Y���f[ķ�Kp{\����o�����7�4��y�H��^[h��\[uINX�w'���kC�ܩ�8Y����;�f>\V�wg_�F���)-�J�+Æ����iR�Kݟrn�~u�2/�������rg�L�k2ѳ�v��4�]�����������v7i�f���=�+Q�F�ë`�38�N�͠�r�e_��nM��\\\��7b�U� v�w�8�<5��zx�{wC	���2'�-�Q����o|M�r�s:"{�����M�v~CCCe�y�s�L� 1?��2l|����i���L���������A��2�����2��4�k��/����a,�F�����̣/���)c���]��^>M�t��Mܶ8�*���v�&=#���_w� 8bg5C&dR��������z8<�k��� �(n�hwo/gL�����8�o ��z�#����b[YY�06�͵�ѻ.�cS��=rZ�SY?��^	��&k4�\�斾��������H[��YC�@8j��=������:
f��s���U$/T@���lU%$L��Ю�&�%w�S	���a}�~BO�S�Тk��b�5gв~n`�Jab:���V��lsNG���ѯ��y<i
G��t��@�I#�4JxTh��+v�gg�+�KI�(���QS�^ۃZ����@!I�b�h������f}��3�1#iD�����\�:��8\�pBZ:�,V�d�v�����ڑ�}����2���Җ���t�O7��w��鶻6L�8�A�A���;�],`�~ΐJ��Pt����������i����^v �)f�y��(� �;��F�UL�ٷ^3����}o���	�(V��4wtT6�8aV�.��,���v��������Z��\Z�{e'���L*p�K��T4��(��b�������ƖS�� ��B���W��A�YBrZ~��Ď<{���)Vl�{�~���a���D�"�+m�s��n�@;��%��%?}��x�čLZ���I����&!^�L����O�XΧ���D������M#�/�
�IC��3~$�P��|��� K"��m�3ڶe6�8��[FȒ.�Mn�~�vsw���;�s9��O#�U0A.�c\Rw�/�!i�#�7�=���i�pp���Z@Kd ��4��4��gzi!�bg��u�9୞>�f*�˳q���U����mq@��q��	��?�fe)8KxKgQ�3k���鼃#})��	��-`���m]v�̤�d&}h^wy烑�ߔ�Y�Pa&I�23�-����wjl�)u��L����D������c�f��m�О��,�=M��47}!������=�=/'�������M�ƅ�Z��D+}�r�e�gq��
G�٨5��:��a-ψ>-nd(R$�|xI����=�Y?k�1�\27[��8P��_�����h�}�(;nB*� !���N�lh[c��O�U�q�I\-N^�V m#�DU�>�UD8۟�q��0�w�8���2J�����
�$�/���<�7s�6����N
�jJ�WNl-ez*.��y?l=��F�i�=�7Gtv���<�tWc�ت��--z���,yF)C�2�Ӂ����͊�@�$1?����A-`x!oѲ����8	��/jf�)�w�g���p!֞����ڡ>d��� 	*=
�}�!w��0x���:�_����+G��lEx��~M����egaꐉ��p<h������+�	ny%�n�0��w����l��Չ�[��q�
%ыϓ��+��J+I7�E�"�e9n��h*�o���>���e��f�����3��*F&��7�X��0mƴ"C%OD�"&	�'(Q�`�,�mN�ۭE�ׂ��ܹT� k=��ç��&^�`c�ڋ�Z�r�K�H�h��Z�1�RY���eR�!�3��k��v��j1˅�R����%/��)����6��Y�b�=��K���W�y��؜���$@n�;��iŇß��KoL�_��ˊ�?����7ܚ)HIKS�Ho>�BWS�^����쿇/N�'�<:}i�5W�~w�������]E �x��$+o⺝�F�Qpr͙��(�=��T��&�`������P#���uĞ=��d�1�����No������v�[��ZUX�~h�������k�� Ik����f��<�Т��9�k�����Z���t-	�dgA*��㬮4[z�� Ő�f.��k'g<���,�V}:$��B:yp&oǧ�V������VZ�h�8y=~��/qSաW����k��H-97��2vSʪ����{�v����CCٕ&	����SN ����k�,���l��WF?����1�N��Y���e��a�b"�)��O�Ɨo���������)���;	LH�1�+��A������BЎ}��b'�v]�>B�u�),�xI���l����㻻�oT�W'��э��yx�����f�J�h/}*�ׁ�����ɥ=�P�%�4��@LH��	��F�S2k�-o#1a�@1md���� q��OY�vF�_B
'@:�W"7�+���a����W��]O�ܞYܿ����z�ក�'>��;���!#�d�ћ(v`��X����%��!�Q-=������S�B7F���b_P	�`������&�x)T�����Q�QU�6��/�7�\^֎#��Z���h�\�=�1'q����.�<}A��s���;{D@U��:��əv��o����a<��i���S1]˯��H �X����+���KƊ�qc�I�Je�u��Z37=#�x���k�P����R�z�Ȥ%�Q�f����yᡛR���!G#��T4w��tD�?�������.o����/Þ�}�x�ě�&��{]E�a�Xt[fr:�Dq��eUf���.�����C"r݃��V���u�Qn��鴄�.����.�AZ���q�9� �i z�Oj����$�.YI'e�ǋ��ӝ_-�ɗ��}��	�l�Pd�}"/8�u|a�в�dZ���r<q'���n-S�z�'�����e۝k�~�ʹ][�������뉬�a;/��ƍΠ�PI;w��>ǭ��12c�q��J�^9,I��y�c;hׁF��OLW�����L�\���)sa��-��E
���]��7@�JY�ښ۰� <�1y�c�K�0�H <��h���t�7B��7U��n�Ϩ�@����i��0��g��N�>F��~�8��O=����I΁XnY ��.��\>κ�\�M�I�.��CM�e$8���g�=�"�7[bo�U���� �\�@k9��%�Ñ+�[6�&�{3Ҝ)�@�֎���`�����;}30���{x�sܨ��ҠQt�jta��&����cO:±'3���%���@O�s􆧐�p0��Oj���yX��F>��&c��'������E�0n!p,��+�qx����ȫ�D��\׭q����ߒ��-���ȱ�tp3:Q��o�!N���Z�Q�o�Z��Zp.Կ&�S�J��*�A����e��b����H^�r��Q3�8.S��A	Kb��?��y<��{�\W�D򒢓�h���g�' {�v+���=�ITa�����Q��&::А�뜂�2����O�+���z�Y'��Ǎ��G%�P̿�&�����2�u>�����{_��fs�'�ڮ�^�KT���?�ta��ׄBe��MD��%sJ�2���߶�ʖ��7�	ATJqqBC}�b�
{�BI_k��،�W�%�F���D���IO4na��7��9�Ҟ5�t�Q+.����"�W	!}#�gz0]A�X~䧉�`2���� �泀b�]E��qg�E�;��3K����P�l�%1G�n|u��)Y�>���B�-����{P�8��������Z{�n�VV��.�dJ1T�'�8(=�i�|Ϸ�cN48��CG�H�!*
�z,�u��L�u=!�����*�b��'��ɑ�]�.�&����*3�(�i�A%s{t�����uW�P�;�_��$
�HeM|��J2�TQ �?���ԕ�}��!��?�~�6�Ϸ5��x"���ɬ��!�if.Ш���I�����
?	˹�u�����`��t�Χ�Oy�c$uI�F76�@�oM����%Z���}��U�$44xҚ�(�Ç���zߝ��÷��`��LY^��ȳW��=|K���V�L�jFvw)������?.������+�������s�g��Xh��4�7�ōr9�� q���p�d�* Vh��kZ������Ϧ�y�P��76�ttj^�� U�6��a4�x~h��A�3)'��X�<	/c3�q���3�t둇�u��Mb�5\����X�6?�$*($47�+�9k����=w��6v��գduBB*����s_����7�G\�ZO�����z^7;�(�um]��7N�ַȔ�j�I�~w��!���~k<\��LR�j��F�O������'X�[`<U�1�8<G2�Ϩ�F���J	��
�]�5*	p�WKOW�R)���gԉu���6�hi��T�˕�����Ɇ�@oP@S���8�f&��8�Y
n�d������
}p�b����|̪~\��^0���$Y���cϕ0�����c�#M�Ӥ�E����`��Czq��������žag�����	|�g��s0�^�v�l�7����p$^���
�,9#<nJ��}i�a"}���0��ރOpٖ�L:�2T���	����h3��U��$kG\B�a \�{ X%�G6��mz�s�(@p<�|�X�; #�_z�����������i���H��ԭ-��<M��0.7�����FwLt���tt�e���JwkJ���m8���<�e��iK�����P����r=RB܎=�Ƃ�-C�ĻR
�C##,SNm}�'�[H�����/���%�xӸ�3e
-R�\V�:.�D�3*\U��B7aG�I/��\�h�8�0گ ^��aN�v�4(��qA\T�S�=�V�i�( P\��:�{_m>J����_��������Q��o皽n�y����o/�a�..S��KA
ϗ�I-0r�h �����~=Ka߿ĜB ��#�~�ׇ�.x�-�N�� �^�9�Ns�+&9��>�)/ %����.US���Z�xFt'Z{�/�Ʒ�)Q~\��z��XX{pl[?c���\Xw��dw$�~5�Tщ$�:F�w׻-����`��	À����qF~/���W).�P�c{������H	7���M,���!����f��]���P*�+/�����\8@/��m||�RR�c��vw��j0�((��<:��^ȴ�l���k����\Au�Ѣ�B�l~��A�e��]�ǐ(�ӏ\t�v��	�x���6k��$g(�VNZ��Q�v�X��s���<���1GϪ q\V\@�,�>���Q <�[!�����Jhn�`�B.z��h�D�d����: iI���~�/͍߅�X�v���6��;	t���M>)�տ�8�Q�)fG�8�ȝ���	7L��L����Y֥:L�$�f�jTd��ΪC�@2ɘr^A5>J	��5�&��|x�c�K=x�%h�ˎ��kGK����>��m����V�+}E'��[�{��.^�� �Z�?���)�����s�|pĹ�/�:�om������l|�BăD��t�N�勍�(�g�'����J2��0�F}�2��+�[��T�BȪ.�s�����0e���� y��~�4��%��i{/[EP��� %���6mq�.iDmGF>��0%^�2,gn�#������8E�`��ꚃ���Йw�4�̒m���T4�ޕ��++�BY������9����	�`�p�<�{���N�́�/��D��^�_ܑ7�s����Cʷ�ť�;�p]#I
��9��a����Ŀ��l�#D�Q�9�4K����&�Ƕ�r<�r�S��?!��{�{+?g�v���Q���E�~��Y�����R�"S@��('I�f��ﭽt3Y	�p1�C8dV���ez�6��o�E֎�<���0%��-z�*�[�N�]�d��^�.��f����u� ���r�����U�ڧ=�3!����zb��Ei:������U�L/,tV�z#� M��LA�-�]D/|Z��A���>�-�#3a���kw�CL�f[s5X��o��y�*K� }�͍��a�]'�����%�/޼�"CS�Y\��h���+���Γ�o�\]��\��wS5x@ 0圯�Lu�&�=�}+M��{p�X�%�p}C�vF�e�_Z�柗5Lӂ�7���U?Bڰ��� ���mIr��~J�������m(-��
��L�PZx)#�k�Ee�������nc�e޴��o|U Ot�/���'��N&lqNLL�Q����:uW��hc4��������i$�~�=\��v]~;��?tʃ'
�VA�@�����V�܆�l*��V:m�����$�]\����6�ŋW���>IR2�n�!]�^ihJZZ�Ėzhy��BJJ���)g�_~t�@O�Aoqz5�79H�H�n\@c��Ln;��[h�Q��B��N���6���A|����-�FX���d�g�^�����ǹ���@%F�B�O������i��N����;����WCC��	��f��2M<�|M:��)*gOo/�5��������^��{zF<��im�V+T\�	2��:�/�<��2����x���LgOV��aj��i���j��1/~�[xw���M��#�yFF*��}���i���y����X���~P硇� ϣΗ_����nȗ���Q9ݐ�����P*C���=#Ԝᖺ�b(��:� ti�rMٮ�y!�����w�ru�GA�%��݄�c �F��ͻ�º��� 
k��X~QE�}�˰'�I�\��¡�i*�J
�U5c?á�5*?�� T=KN�J����}N1O����ϟ�?,�ߟ����
^__�F����*-]-���5�M���z��jЈy��DsU�����+�������"L����6C;IC����m����5�PpGDX���(I�ۺ��%H6�3�,933��by�|������#t}�H�%�*K�y���`F�D� h�hTH�:�G�K4��ꭄi���5�4?�* �T�Lh^��0��[�ҥR��t��S�?6>zB �9Q�T?e��>@�GXn߬���G���ԫ�LpK䪘r
ss�BkcLz�^��c�E�W�U�W}��*�r��J�W*O���V�}_sxU���󦠚����	Um��@lg�)Q�i\֍�g�T�w�ݍ�/
�ۚ��G�ݬ��bG����j�A�h�W����#����~[n����d��#gf�S]�QrI f��M�ɧc�Q(��13�4���s&�M��0�پ������y��C�C������S�m��@(ɼm��Ӊ�rR������E�����h}�+�z�T��m����[H{��;���P������N?��_-�l�4!�e��t��>��q��U��ZGM���(qQ�V�H�`�_#)��!.M������x�[=|G��5�����uP? p���m�����v*}��a�L��"��w�>�� �C}�ɿ������DaKۥ�=r��t�W0���-{q��=^������kwᣟ�����������L��4�Ob/�6i����ml�Y|[}}aC(-A�Q�>3�9�&��OK��9�Xl^DNK�5�E����1;��k]&U堏_�ؽLt9�7�~��/uMp ��[�C%ȭd��]]���6Q9�~�����:'ЯAиD9��9S���� r�+yg��K�"����R��` ٛ�Y��`Λ�����o^�������3�s����V�>����|&�-�b[J��w�3�˗4���oj<�eDD���V��
���L0�T��'>=?�(%�YU55�2��YYY���$�9��b�rt��5�뺫ղ�(��C�ss��*ɼ�3��h�lC���[3N�e��m1Z�XR�����,m�Ķ�6�A��������8��˛�ƥ�>��$�`l�BB�8�⍥5�I��G9�Q6m�;]��Ћ'h��B���0�������ojg��K���y��n�0]V #�x�����<�j��l��A �=y�3�ѭ�Շ���ɷv�ߖ��hs���٤�����㪟�jl`���u���*;�=z�@���C���:g���FJ`����ŵ���8J����i1ql��-�פ���ؽP�?��m|��##�wԑ�	���������8^݊N�E�94���e1�58�7�G���o�y7j>IL��b��8���x'��g��!8Kz�[�����x4[�e|J� � 
fDO�D1Zp���^ ^��<���Я�?H�bv�1~_o���s�l�XiN�C8\h �\��!�k��hz�TL��v�㚆��X���1�ml�||��C��K+E�zi�*�	���t�>|�M�Љ�ؒ��b#�b[��qȸ�ԃ	R��#Y;?]�Ϭ���9���[�|S8�&_W>��S��o�wOހ��L�����ו��i뮦�l����DE�3��_V>K��Ƈ��e����%({su������t����(�r�2�����o�Zl��cFk��e�Fe2�Q����ݡ/���ޙ��6|�yi_��X�@J��6np� �1�!��0���w��J'�7?����FU�<�������;�����7oG�f&��'Q�n,�����܉��-�3�l#�,vv����32l���h�b�p��ٓʆZ54��e;��N�c���* t���YX��SD0@2w�U��"� �G�h�1 ]������\¸[��w����1�,���/�)�%�d��c��z
Y�J��͇�yK0���2v뭦h��
Z��la�%ȧ2����d�����@�lQ�ޕ}�Ճ��c�6�o?��\��]p$���\;�0��sj%f��gQ�䵵�]NM�ii+f���92��pdOw�Og&E��"BB±%n�.��Υ��Ƶ��~22z3�0���RԠk�@tSX�־�>1'E���/4j�e�I��D�)��w� �ƛ􍩫O�"_��1�ی�V"±��!ׯ�����z��£b|!�&�[�⯰P�o�'�v	�7Ϟ|o�̩��<?��v8����o�WA��c����&���a^���g��̦@��*�`�=R�~�Ƞ"��nC�������*|F^Z��D�B%�ϧ3�6��a��Sų�aq��PPRb�hw��]�������q/�Ȅ4���ޢ{�㰼*J ��77�/��+K��EKH�`��ԣ���>���_͇,����⢐\�$���̬:^P�|=�r�
���\�w:(<]Ōn����@���y��b7�;����L��2��t���䲶���-	��:���У���2������O�J^����ؘ��*�̳ܥ'�`=�r֓�M{U�ӟ$͐8�s�4�&��}��f�<�����	~���S�nA����qK, �g������ $�"�b.���3r�6��5�"Sh)�Q���x���&/�a�!͐�o�R�Mr����K��Z� 픬N���c���K�Ӆ�q���xC���g<"����̥�ޒ�[��S�9�s��,S�D�1>�2	}o¡� .�%G��{~9�r�n�3�hl���U�D�V�������E�$�-QC��H i�
?�4��4�Ӡ+K]�(ח�ڪ�'�崯Y�ig+��h��`���^�E�=sbUus�ȣ�:i�a�0�xv�ܞ$g�ɵ���fa��";{�:.Z{��9��4�Rє��Qe���%$�&\�;���~��^�s�o���8��&������Y���lL9�/y2�����!��
o�
n�����[��/�p�|���V��r}�ґ�Hʾ��hn�u���Wc׾��1�%}+9Z:r����⚠f����tvP�2yc� �k�'i��;f\�P�MZ�h��}��n�({o�A����vTK|�7]v���u�uB��u`���k}*ьP06AHLo`i� m�m�7��C�� ��3�2��Նy�^CfT�z���ң���wtFn��[��&���D,��4�'atfI1��u�QQ?a�_Z�I]$�n�%%$DBBZr		X�DJ@�KZbAJ�;�[Z���<�{�(�ߙ����\3�]W�E_�f��|���ȶD�\ ����n��]�n��Q�v��I���R���!��d������^8��cWQ��ǚ�2sxA����3�E�v��H�m�9+h
E�1i8m"�9v��		؞�Ab��;X��ڕ�CH���3�y�C� ӪB�c|<O����1���ߚ�c̴p�w�}Yo�JC�`j˙�c����1����y��L&�QaJϚ�p/��1���e�z���=}0��3'v�e��m/����R��ba��%��]���&��A��G%7��BE)\ ���ippmK��ԩW��#���ݨ�/w�w%(��}��$&z�Cu�d�{c�!E(�OZ�QK�(!&��a���c�<�oW9�$RTUk_6��̆�kTr�k)K^E+�?�9)����DT?E�*���vo|����R\�E�h̶wm�OZ� �D�Ҙ�;�r�D�!zC�	N��&�mrqޤq����[IK���Ӆv�|�&��As���p�
j�`��9��Հ�7��t�h��[���G�\R�9KMrJ?0찭(�0?���.��;�M ����;<��r&<��)����x�s��G�cy����{��N"�W�=�>CNL$O2c\"���Ӭw-�I:M�W�~�������H7��c���y=1�P���ƾ�g_��gT���d�>O�W�I�߱�O	X�9�� f���>��� �Uv�Pٚq���xWUc#��*���oݞ/_�v��������֯��J@�5�s���<��7o�r��EAFI AAHXX��tK��/�{��c�����'����N�>g{I��1e-�9��JKD]*C��<ٷw�Ҩ]?�|v�]&4��/�q)��%��F���D�Ndg_��Q�B(�͸v湔c��l�V �.,0�n�%�p��ؤO>SP�ǲ2�.��!��+e�� i(5777���ulfi9�~~P�}'����2L���M${�g����(��T.w�����
A�
�Y�v�_�N9���ۀ��۪�~m�"���Q�YO�S��8���k�q8��m<�zG�D�t{�2J&4��D����{���N�6�@ ds�}�B�ψ�♒��1!E{�>���P& ��)�2����Q���Ȯ�%+���4��r�6-�%�1��y?ŉ�2_�޲����h]�)/�X����8�n��(�7�	�wj��5�YJgfga���2�^߳�x@���R	�=��P^U�&�P��H	.]T��k�f����Ƨ`���'Kt�1�`�_�r�m^2d��ߋjW���Pr��w���o��nR�J��.�Z�0���l�F'�;i��Q�K�(�Z*��D���|,$j9􀗊�a�:WF��H�>&��QfJ�#I��H��F��咲�LN�	�4uC��K���%�3y���=c/���pv�5��Jv����@*0�����+�^�l����r�6�N�I���")Ca��/�&��l�p�;Gi�P�W�ء��ѧWZE��5�-l����V�?	�d�7:*�:��n�Z,}L'
`��~AшuRr�YQ�yΕ�$�4����aGk�x�Yb�<�6FsQ���L$��2US0��a���3�Ӕ]��;�|J���ҵ�11�6��ٞ�uU�:/?/���hD#t!��P鿻�[[v�Ҡ'z,��o��t�$V�u��j<�i5�hm�Í��}�ȧ��1�a�]�����C�E��S�����wp��ơ��.H��[yK�Bm_��@mc���mFA�G�ԣ���S��4.X��9��;\��/(e���k�|�~����$����m?�&������K++˷p߮�G����	X���߁����K'����^�Z�'���������%����&��h-�.��~��3�fŶ������E	�y��Ml�`YDI��0�"�I���=�c4��C ��Y��YrE�h�F����w���衪�ji�K
=HՈ���U���.Ԅ��E���Ⱥ-� �e���R�/[		:�~��b�A�h�}��y�Qe���e�Q�`�ޠA	jgJA� �6�3kM����p­��4E'R�&���������bP-OtD��z�̩q�V�\��17Q>�ΐ�_֔�]m�<򩴁�e����+�P��'>������A�U-c�goZ� L������ww}p�d`!�[f,}��G�"Zj���da=�e�K.�/VɅ
]��o545K��ZF��"�e��R��Jn��&|Z�$QkV2)�*�q
D m����DA�".����HH�Q_��5~���QC�u1�q�Ä�9�禦�Kt���U�P����v�gtyyZ�T�ޟ��百~�j�Pw�Au�9����R�`b�������S��L.��B4q[%!����[C�ެ�DV������a�� ������V��a�gZ�ӛ��wH�y{�����Eӷ���q�'Hě��C�-_�k���1z�T�3W
��!XwzS�eC��'Wwp�A�B���Ώ�ص,�媃��zlO>2I����U��W����H"��@Y�Pv�G.xsx� �&�e��qe����C��V��b��4�v2U��$6��fX�ǲ���G�j��S�}2FrF�������|�&��f�4�����]��$�{n���B$��b()�xDד�G�_&�5`�x�� MD0?�D�Pc]r������-�����±7�<���[Z3� �u����{=�����1�S3�,�E�N�"N"u��h�q�Jѡ�\8:x/�F�1>N~�2�T��Di��������d�O(8𿎅���!Q2����{;mÀ��'���-a��ꊞ̒��48�yg1�ț�B�G�}(Ѯ bMJ����Ev�Y�ŢuA$#��/����]����&eT�1x�ٷ�C��u���ͩ~2��sϹB<�윃�߄��������"�i����~�<<mX5�p���p1�N������St�!/��J�ҡ�y�B�ĵN������q��ׯ��ЛƀY(�gs%9茹���}���(�rI	[B�E��||��hA,V;��x����Ϧ�zy��I���5� �-��\Ӷ�A�_!��"d����<�HT+��I?%$�@����L7�@9�v�H-�8F�7+�0�
HJ�q"�Ǣ#r#���[�K�r��wα��[u���xR~��Y|�
��/��4^9;+�~�f+�U���ϒ���MX>�5������D��)�B�whg־gӿ��j����!�Z4���PoD  �.�%�.������㵷�P��9燤���倮��T����8������+�� �.���nynn����6x��*Lr��4���q�C��=��Ȕ�G�/$�+����pp��Eޣ�a�N�ϩ��ٸ*����~̐��"��=�it-�� [b�n�ǙP��es�3��A�[1���y�� ��n*�|I���\zx�=�7��sŊȧ�q�k�M/G�r�1AP��	p�؀��#�f��lC�|��&�g��cJ��kAI�Rܜam�k���t��+��췹��mx���y���H�����Ŭ	4����I+���ti����uw�^AUg�f�Ɔ�������*%���z���)&�<$y��;��a5Ů�i"`��6�p�۷�9&�߼y,8�}x���R����`�V�)@�{���q=�A�9����1~�Cf��3Kp?�lk�t���5���ݴt���ca��g�N��EK�D{�gr�4�Pw�A�L�)�M��D����7��5,>*d��9C$��� �\b�i9�P4��)�!???zgǝ��{Sn.9��#�����dƥvV����m��шU��	����v"���񼘥���T�V ��e�l>:q�X����������8;NU=�v����_z@8��H��B�
u<3C�!���)Sh��w���~�
�	����P5z�?�lY��~{�4�>�a'K��� e �ɩ)&g�啟Ɏ�s/�p�`1
�˷�9+H8:�T�����4���(̴�2�\��bm i]�{$a�GW��}p
��q����3D]�C�o�@�G�����H,�ǯ��sQ
kݱ�N������[�5��"�ìպE��[dq'|�A� ���N��-h�ꄾS�&��$;f{�O�����x��K<��:�~��	��"ɉ}_z�$�� d�@��L�R�����������@Xp�P�wꤪ"_� ��ީ��ʭ�ܡ���R����%)��u���� ��*�#w0��
m`P2 I�5�.d+./�sQ[�k(Zt�b'�m���f >&3�j��x���(��x�j��U��ü����0�qt��$A�ĹR�G �${�4WR}�Έ�gC-T?^����˺�p�|B;٨�vV��Le���>�z����Q�)��&v�����(�'�q�+�ٶ��߻ s��\)>	*�9���Ҿy
�#qO5�fgu�N/�@�2����h�JH��ZT2^!{fgi{�}p���!�pi���A� t���'��	��ǣ/�gR�@,���4Qמ��,7(����`	dc��W��x�,������6e��e$N/>��A�Y��g�B}���]N��
��;Ƹ�^�oǗ�?�[���\%Ʋ�O��y'��a*Ùm�FMNE�<������C��U�&�rƿ��T�(2PY�
�%�~��'�Y�5M={J'����'tx�Y�t~(���1�K��a���!M(�����ɿm�슺:�A�����yh	�h�J�}��E�@g�wS"��q2��1�~�������w�Vm��5:�<��wOMLA��:����}}�f����ڏ�1���QHzz_�`���)^%��-�}-�Gm{OcUa�<:�m~���ڿ-�_l���c�J�L�]�]���0��a�����͹��J�����_��y�?j�F3Kc���ҝ����=̿~���� �L���������ӽ���k��;���I0�f)9���=�P�B42�صG����u¡K�ّe%�,Mu}�u�\y�uC5 �����~D�mM�:`>�/��C2dga%'�h��C�h�T����H�5QL��Ԋ�3�,fh&�kFhH�Q�����|�`�JՔ"	aYB�!���e�NGO�(3�3��H��X���Ã����,�I/u(�H↕���L��;��Z<<W-@�u�o� #j>���q:َ�ۋ�s6�����ϙ�����{6u)�J�b��S/�<i�{"ԗ�2ד�gO�qN!3F�"�gͽ���H�A?�G���z������n�����X���7�f��;CI`��R$!&�}�#��5���,���|����ÿ}A��k��BܠB_K�]J�>���|�Ƅ��+�0����Ƣtܥc/��N���EO�HJJ"7p��=�&T7�0�� `V �Y���ȍ<�o��x������:ߠӜ����F�T�F֐u��Q�г���^
���B��+ߕ��~����6�����%��b�D�O��?<�:n��b_%�����,�da��4����A�2�?�D;�!�"�zN��l���w���e`����!��sX�ݺET�75eLYO]���j�ϩ��C�iF�r�y��Ą�ë*�� rRO�%�q��0���S�D�^^�G/�n�_�\"'�:��Ѻ�Ǒ�W�j��a�Z��c�_��r��Tw�74��چ���e 暰����E��0Gs󜃩���ة�Ci\��ӑ(�D)�q�Ũw�@�����=�;}�vƺ�/�#��LY=G�D;�G^w�տ��zT�2�E��^�Y=@�RlA�X�9m��Bv��mܴ6��^����G�΀�����zc;�_9�}�w�� R��Lsy3?�o���z���2��"����G���{�7�U��G��e�����GJ���7��˦�W�/O~��T<�������53�.�3�ݽ�?7�1�V;i`d�owo|2L�|�&ܮ�gX�5��aYM���]7������*-7� |���Mئ6�κ���Y�� ���������u;�a��n<�鹈0$����$��(#���yP,*&�ے�O$� �OD\\{Tm�VГ��!2&�n��f�)Υ8{e0�G���1��9���U�`]/���*4�Di��B��(=v_����DuX25�-�}~?�w.�*_�t�|���ҿ�^�dT�@[�4�â{#��bLp�0�#ͅ:F�6�2��v�,�@��t�w	�k�HS��_��*���v3�%���r���	fk{;!11���J�j2�e��a-)��<uH�����u�}��ʦY�L��Q>8rG�9�����go5ED��쐅"���So[W�܅$nm.��ٸ����4��w!3�Au�����.i����,:h�khK��z�� ��d��g�Tl���c�^����D������Z�.�A�7*���٩|aC����,3'�j	.��� ��O�SD��0�=E�^GS��=�G���eф�oOt��\��1�>����Ժ���6>>�/�)�x��o�S"���D�����q���G��_�����&&�n�F��NN���T����P�a���
���˓���j�C���J5�i]^F*i
�<֚�H��z+���<~t�\,d	~85�rU�[E�c�I#:�a\ҕ�^���w�S��"��n2���\�H_K.x����Ѯ�꘩uܿ�9x�9ã�1+��j��S|6o�ϲ�]N,��#�6������j5V�hooOQ����sk�TPޟ�rs�'��s���� Ǩ��&T[~t��[�w��[��;��N��4I&1���D�����TUUU�r�T���WL&���h�p2���^)�T����{~e���cCm���^��p�X��ؽc���Be}CP��Av,"U�Ґp�Q��'������j���6��C�Vv��d��f�Ys;�"���q��۹o|�ds�<�Tߥ���M�����6����\�y�9#6��u3�J_�i4�m՜٩�C�t�	\^C(�`z�l"RRq�D����;
���HC���%M�36rr�E%��� @����vya#�PZVF���3;��9�s��LU Cze����X�-l�v:������4�L�j��շj#�N�L�����k��2��X;Kxs0�m�]XmU�8������0�'� p����ё��津�/�f���yI{�qs�~�"���7"�ƾ�fe�t���w���s�@��8�8D�E����ͮ���!�-��$M=NHDt���٨fEM�����Tt��}��	�>'�XQ��N���2��@lni�`��M}p}�rE�g���h7;?��jJg�,2*Jy�1��T�z	�^ѝ� �Xni&S&h�*��^J��O ���J�&����\���r���#7��|Ȍ��w�����`��W�j������4ў���U.?��qV���f���r�O�3��^��g�F�����-�yo��E�j�2�|���Y�����뫢-�O�1G��0��xJ�4�]C�9�~^*�55š�q�4����!�8�\u�cz��N�s��@�pZ�� Z[Ǩp�Ow�1e@s�o��k���oY�-���0-7��ָeR䟷�O��lR��}���տ��j�#8a{|痥���z�21��������U	���/��X�D��"��1�� El��-\�B�����p[S1Z����:����M��DDj�%��p��(�*��X�_�tu)ߥ's��I��:���[2Sf\ƒ1@������Y������\�#@M//ԇg�^0f����9dM��xT_|�hf�9'����,�K�p�jX�ƀ�����h�5�tD p��V�ɟ�6ǲK}y�Z��튴P�=�\
�_�|����8N�ԌI�
Z	����}'P���O�p<����RDտ�l�s�_=�9��s�����ί�_��u'Ya��c�I�Kc�@��f�5�@�(��x0��@n(���E٢
�t�ڟ�Ϸ����-�m���PZ|�2f�^A���H�DH�\-�
}�T���o�){�sc�=�(S��mtV�@�YEAA�|�z��S�k�ȶPw!%֥��Ԗ?��^�F�X
�JH���
�!���rk�:�OL|�HR��ud���+2�y���Ge���&'��hL$��E�x��%ڊ�xE_� =�Ϸ��Iwpa��dnnn%��瑸8^b��be�8ii�QMǋ3#��h��xO^mb�����7�P�q"x�{!3���b��ͱc��2<Y���մ���ӻ��Z "����p��_� ž��-���}�֌,*��G��Qn����j#�u��ȕXy4�:�08��9�BL��#q7���)�@mt��zBh���89V��E�P�6�[�4g�kޡ����U�z�v\����%��j�7ul�ʇ�{�:NN�5K���_\x/��o7V�Q��#ub��Qb��e`�X_O*��ulfcs�q�i��ti�2�䕵���������d������3C�Q2yP�O����Ԃ[���s�٩;�*�0�G��������-�;dƜ��bn�d9 v�pg;���n��e�6R7�r}�'M�Z��"�VqIު�A|pi �X�ծ%dsj󌎮��c�TAO0��\��5��w��Y�n�$2���m��>\�-R9��s8U,�3�5x���lh�:�O��HJJ�E��Λ�N�MM5�Z�GA��J��r�m�}�������-,`��ᬭ��F�˝��.�ONO�TA�~��upV����-�y�a����=�+d�P c [�|�a��꺲�6��R�:C�$$����#��C	�� �OH޾v5���Y�Q��sE��ﯭ&�g���V(t������vS�0�(�f$ԌpPr.*+�~Ґ�s�����;9Ik�#E��~��
�S�"]�]ABd+��g�sk��)h����[��)J�aSS/l��5�fjˆ�(�����iiiI�u8_301=�D@c�He�������S�G�X���Y\�~J�Pg/��oQ�,ꖌ���u�R
��N[aDd&t^PAJUX6��(�� ��a-@>p�_{C���$�)�C� �����t��n��&�Ǻ�����	*���b���ʵ,�K�[Ā�lC^���=wuq!7.��Td�*�88�y)��f�����f�-l���!�n!�伀����o/�yh,-'��&dJ�������mG�T11�Q5G::���}�O2��!AXR�#06���	�O�x�H�_�EQ����Z�NVl�����]���u}C6��hQ�aD�tC�
ACk(KSk�-XN��P�X%8����ǖ��ƕ%D)d��ʶ
|�2�痒"�),`��E>n���&M6��y�!wWm����=T٨߽����(ё}�C��z����^��5��w,����F��^�
��s����j.
�J��D�٥�f�=&���!{���h�4�`��^���#V��.\��H�h��dB 2�V�'l)�i='���sm�� �5HK�4�@.oe`���m�o肧9��r�R��3�qK6�mŖL�;�����I�r�<˶Q�t���F�����*79HyUU���嘝��F�A�'��Wԥ��i�`9}kK�_E���$D3K��|gbb��$�;H�⑈"66��_�پ���"6ddd�}���� :7�)�	�diPto�+����<��2��;�J�
�Z�!����zC;5$/������~4�}��?�/KCK/��;_�u𔑬0��U����5���(�����{F@$u'5������#��86�sGl>��7����qz.X�W5�B�vxH�tA��à�Ya&i_���t�7���5�l6�yÓ�<�v�z�0ӆ���:���ۻ@��P/! @��8L./f�u;��ʂ��Φ)4���������mRfd���:p߭�^;<|�V�b������\��O���������� upʌuf�yVC��[�5
�#J��(ɍW>o���~!�<<�) Y�<���S{ֈ�����W'�2�P�K�w@ɺ������Gk��2..�YJ���Dj(�>!aw3P�&��^�.#L_Зڜ	"�����GrS�O,�D���H�J���x��-7��#�;7==�S����P���uC:��=Bxt.�%qɽRD@�{VzG�3���n�U�����0���?;���ǘ��PĴ�;�k�{"��_�=�P�걨,��<e�B��H*p�#��0�&7ϧ''c|���k)����И�w�����閉��-��H(ѝ��j�*O�9�l���sC}��Y>ŝ��2�P� ��Eo�X��,�w�Ar\	Ǩ��n�P��n�����#�{'�q�i
x�"�kw���Po9Ц�;w�p�C�h3�(��}����ZL۽="p��>�u��ֹt�Q���o�[X���=6�]���X�[vYC�usL��L#Ξ���<I�;A<�<�Ȋ��A.-�K�C���L��Ծ/r�1���lz_�����ϟ���>T��K�7z��qH|����"ןZ��JJ��U ��JHg��}V6�����֩{�S@m����{[�l�!�lP��PQ1sV�ꈀg�z��gB��Tb�a݈�n�����Qc��S(f��8���RH� ��%��G�zL4� ��篁� �J�<�;���좦�ݷ���]�Aev)�CC����</�����W���'''9(V����O,U�ʝ�"�W�ܖ((�Ѹ�:=gaa�?��:6��sZ�zX1ݝ�{��o����Q�YQ� ����Y�4�B-@�.���rP��OF��L�E{2��+�	B:�. ����2��6f��L��z=�>I��,I�~��=8a #�ũ,�}fu��Qir񰶾��ݻ����+.w�?��o���:��G��Ȉo'�.�a�d�%�T� ��T�`kKg\�+^����)E���ghXL�g"mȐhHw��7o����w��[��LMɖ�>${'���U"*�x�����K��9<:��)���m;+���(��)i��p�����(��M�f�>ًv�xs���H�!��`f�`F�E��\U��>�--v4obz,���w�I�����Ñc������p���{�(J�c��G���-}C�[\m�Z��f��H-�[I�"�gf�il�>V��uϰ�Bs�33X�RsS�!Ob����gi�N\\��c��b8:���ݔ=����͹5�6O-�8$���/�cьw/������<�KNa{X�-��8�s%h �Z���E*b�>�b-h�R�W�*�fd+�g�H���n���G���H��������|t��!��5L4�B���dRVT�W�KZ<��a1�4� Ղ��<��@R-��b��(�g�|��</�fo_̯������o�wx���7���Ŝ��}� {���K�ȧP�a�H���A������]02�
��˶�R� ~Ä���9.���F�d<�q�) ~�;�DJ>"t��lc�G�Y�o������1�@�
������?I�T		������{����mݷZi������f���	��p��
!!!�z(Ԇ�~~��o��G8J��4����q���D�%<����L*f�r�8������&�����v�5��iL�y��W�)�F^b@|����z�7HMҩ��W�Z;<�j�`�%~s]��{���Jc������.��c4BG�ȿE�k_*Xw�J2.6Is|�k�؋<�3-��̎.�]ў��v�����.>����ohBh�k�[Y�<%FtE��3��{�CJg��Ԃ���o��ǫ�+�؟�y�AtW �F����M|^ޙ��SS7��#��Ǿ��� v#3����Kߖ#���2��^&�%����^�2k�>!��`r�Y2����i�������[U$92X%�\�j
ME@���80�kWHX��W&��kݽ�¼��_ī�d��Ū��B"Y$Ϊ���d8��AE?�'�X��"�,�~��goo�4�#��),	�����M��}��<o��Ѕ�/i_��YL�����.3iQ��z6xǨ���?��-5ukx�d�XNN��'Hp>=l�ސvp �,xm���>(��e��f��d8�PYu���c�6�x�:R��y7}��±E ���������נ�5k�ڋ�ZE�p�=���Q�,��8���p���1U�YJ͌�L����w3�PbW�����k��«ޕ�\�h&����O�&�K����0b/t��o�QeiCYƮr��j��;��d���}�&��u��7�^�iq�o���,�)���_N������g�E_��W�b�$�I��ژ��m���&S��|I�uX��l���� \YˬB���]r�!7<�D��ǊL��(T�~��[��Ɛ�ɵ��(�&���S�J�nn����o��>�{�:-���U~{�ny�^������m�XTT���/��Sy4:���Ξi*�=,�^<�:/���'�H�������6��ϮAv;��?�0ߨ�.go�yV4V�|%��x����}q1��-A��@����bח��ß��,h�J����뇷���kƏ�a8@��2H~�(U蓪[�-0�=�H��!�������Œj�-52��Q�`��[��Xpz��F��v�6Y�
�6�ф��,[O�g���i��B%^����-�N��wBd����X��y�<�wW�� {V��nDV麘m�q�5nM�Ϧ-Z�$����s�<⑨V�6O�%9jr&P�&ED�7.�VWq�"��G�gml�@m���ojo����b�:�FB����ԁ>{��'����o�*�(m�K4!�q���d�+ό��>�7�~��9f�^Y�P�?g1`�Xg�% ���߲5TL�-s�9�E*��rx�Z�LTJ��7���%:ߙ��%J�}y�`q��u�kSS2&�|?�l������
J�ͽӥ��5�z
`���`�:6>5, Zξ<���PN"��(�g��Y╹6ä�C����&P�\�&�,�'&&-��#3;�
�G�rF8^_�O�V����^��=�X֥k�dC5|@5��g�EPU`�~�p����6�~���D��m-����F����j	/�DK�Y�kd�l��QV�gy��T�*w����Y�~-g��Li'(�E��U�Ը6<�ss���������U�w�
/dM٫�5�M+�/�?z�.�t������3j �]E����^�N[���d���!��\�.������&�+22��a�V��"־o��'>�a��D�<`M���cA�&?�I�-���jH�Iy��A1��0��,)��mSH��J�/���<b��Ukb�(<���~��̷�w�xw���`9:l���1hWFmʡs:05���׵e6tlll�&R�D ��[�H�Dr���V���F�����ӄ�.���Mhg��PR��?L�e#���Pj����{�j�e-�b��V�������3��1��'�
9���=���\����A��[PDw�4�$���ݼu~��i��my>��͙1�~),/SoH�.h���tf��� S�
��s���b�(יl4��$%T�Ы9�Ǹ�@���G�x`fַ�C:��Wmk�½4����S��|�K��/g������!�X6s����L�
C���Iy��naӢu�	���p����ŰB�~n��PH��dU�g�5&[����?�2jy����6V� �_S�9�&��&Jt�v��Hb���C�f����V�C�>j����p��"��/҅sD�޻kY'�19LH)_�}������bJ;\�]"g���-��j�]���!KYYni���]d*n���c�(�w�����-˿}���nm��K��E ���Rq�y���}j*=��{}P��] ����Ĳ��û�s<6Nf����[��E��-Ȟ�e����R&�H�%�}���>̀ ���c�N�޻���[Yy�ߦF"�@$���1^Q���wf{l��zy�Z�	�N��2cj�~�%�r��Llu..~Cذa��=@�:CE�M���ٸuJ���[y�!�`��+�|^NN����aY��Þ�cçD-�V��w�� �}(렙@Y����Z�ų����u�v"��u��->�gu���
dj?�ɉ����r��9ƞ���~���[T$���zà�(��S_��tsy�n�7D��q����o9�����T�>����Pr@���X1ȆN�E��0���M�PyJ���_��p������/�ܭ�P����IrR/c;��09$c*�&��w���)�Ԗ�('%>ж������{�������\��:F��[�r7�$�P��o�/���O��9 W\̝2�y�U�Q;�x�j�nP:J�IH,�`��/T=^�wp��uμJt�D��
�������{<R-$j��*�*����,�*b��N�B�������HYh3z ֐��)�ƵϤ h5�����A��Ik�Q����e0�3���(�""8$�I���1�����I���O&������s��힟/="
���}�����d��'��&��2�3G�f�0����s;�ԉ�"
2�4�ƀ���Tt�K0����1S�1qҍ�=��r�Łv)���O>����&��66V���C�e�nP7gޕb^�	�'���J���IDF�fs83ֿ�x�&�7d�W���~3Y᧞�=��n�('}S�f�h�	7<�Ƭۈ��H�P�gx�c�Y}_�j֜]�(����cA2"pp}%��͔12����
ä���d{q����HT"]*���[N���w@r����1st���[���NJ��㶵���w�(�O�A�:?��U6N� ��|Tc�S zǈ�|�J�!Y�zidA�[9����.�:��i����C���!a� ��b���^���=k�nQ{������J�s
Yḵ����8Vm93�P��{���"�s�wN]���)I����������6I�x������*�r)���&���ܜQ�����ty�j�`m�#����9��/}��NO�+�]��/q��7,/��v!�v?��Ս�%���vpP�����\@�x/
�Q쳖�z��*�Ez�* ��YX�F�d�ۀg�E#-,0<,�030w����a�,!�}\I�4ᵶz�Ū�`�Vʉ������bh$�О�
�_Y�42������+�q&�i(����_Mv�9(�F����mU��}Ͱ���ۃ�G���V(m�ti��� P��!h\�:IojlD:]0~!E���:n�N�a�����I������8�z�A���>��#�������c�%ķ�����_�m]�}����p�;!�f�#S�u`:f	�����$�Ps'������د��F~b�a|�-��Qm5[j)/�p㖿�Hc4`Y3�1���F�iio6d�~����M!��l�-��s�}9���c3́%Aei�Q������5Z�a�ݯ�㥩*���S��SSߪB���24�G�r_�[jk���I�dƠ��"2��1���{���n�'��|�Y�MSG��jo==6@J���Sc�M��7f:���MG)�B�v��a�Z�K���׺�z�q)X�`�`�1�-[6��o���=�Z�+ s3Z\�rKOO�_2eF_Ǿ�;��G���O�.�"��Ǌ�a�,�s���*[ ;��j���|��4uv���D���4�q01$�O��xđ0+oi�r�%�|vky�b�����sZ�:����}����KY^lH|�6��&&��`�FCTl,��g�����YC���zC]�$�y�Q���l�����-��H�u���`U�����+�����o�4"��6@�������k@��$M�}.�����]=�z���𜵵G�=�R��2��Q��B��[ e_XJ�bAcctoo5`qqE璌�"�����G�u�<O����HP��d�.���g�mlp�rßqS.�_qy��p��l��ݻw��-
u�k蘍��oP����۰�����L���I���F��� ��1������CX9�~�xP6�B9tSJ��i��rI&�l�6Ǣ��>�4>��O@MQ�AsRs�u���8�8�s3O�
�{�=������Z����w�� [�ҴGɮb���t8��_�<���C�����~�nm�e���z���Xq��@[�A�'50@4`ř��ϳ}���%���C����v�]�2,H�mo;y5r�남��9�ԝ��sQ��iV��'#�R�"�*����.��X��i-�AFjI?�z�o�ߙ����
l�J
w���5c�e��>�7��n B�Ʋ*Ԑ��U�{�J��/��{����BB��Ռl�%i�*�)zn���}�
�~]���ORj��(՜.Ob�L��}�^�]JpggHRJ�.��5�B;*���6"��p���9������U^���S�r��(��	4�"I��k�q�!q����bs~Y����)�B�6�xꀥ��C�u}`Q�'�m�0;�-� 8��]&�[�S��P�x�nR�{��:�� d�Ø���)n�ܸrK�0�o���ss�6s����;�s����C��h�W��0Y�QbvvQ��ႉ��k)iiHd���=�&}_?AB,;�"��8|�l�[ظ|��J D���|������-���9#uG��ffO^h5�;(
5��^�W�����Ĥ�P�N�k۳j5Rp���z?����;�� �6P.�s���5�-��8e�}����xJ?�ǁB��#�6�g\�q�!"b?+ ������S��x@����%/}n�M}a�9<��9���`�6���~X"3�iJ<�|D���������I��	K���읚𑍎���j�sߵ8�]]�Rɭ���X�]\\|���a ���$�넪��S��z��/(�jY��|��C�`s�����&؛E�����=A�D�*��}�"���ރf�v��%�:|����Q��QQ>��0 %��t��Hw�,��! )Hwww����,�%%�������+ҝ>s��s~���⸰3s�ꚙ���*��8�&�y��{�y��s\\O�6�������1����j�����e����0�x}�����*I�۞uNd�ሇ�w��W]�[���E�|�+Ra��G�iL����-�.S�1���:��8��+��:��������K�3����"/���+��}���^qo�~|��X�}NsɝڵYՈMz�mN�K�m�����tW�B���@H�c%��"n߾psY�qޙ�$GF��C���`��]n�wv���7@��
��Z�7jǿ�Dx���ׯoQO�-��[��� �R
�����1�p'L����ZZX��O/��r��5= �J|!�7�팋��+��_�� >~=�K�K]O�ymȞ�Z=��E~I��e���Q�7��ygg�s�7�888�E�q��u��}9��_��dC@D��*-M�<��0� X&�zC��jO�e�80��i2�����H�߮�#Uw)2�{b91V�c	��^ ՟rQ��*������Η_HT�Z�6�;��ݝӼo�;�v����o^w����PQ9a����(
�}wP1�T&�
+*j9n:,2� �RsfR|�
�W�O~��3鼕<�`i���`���KY���Ip����c��������Ze�����I/�V�z��WdB<�,�6��(̛�b�w
�����cE�	��1AЇ����:le�p�����TRq����F��跉ec�;�F�1��������o�b���Љ��m�f�D���Y�����ֹA��(����yN�|�53q�e>�͈�s:��iЋ�x�'������	WW������A���G�D�L`#Ƹ�(t�@x��S"�uV�+�����1��H��j�&�@F)Ϟ]��*�B�I�%;O=�H� �c�H�Nc3�|?x#>�75����	+�
�d!|�ǂ�����?���;R��r�E����,��g9x�hV~��002����5R�lU���2�C������� �C�:��ŷ�[�t��I�С"�\n>�`d����@Nl\��~=0��������70z���	�ۓڕ�/���mm��{Pcٿ�����&��\Rbj������6��G�b�� X;����m^dވ�y�ų%Z��cu#�d��x��v�M��������^���m�s���d�kJH��3Ux&��,{�~�=�����rdك�痡�@[�T@ۛ�.;j��9������趋}@��q���WH���ncj���t���"��vh-+k���-e*#��а�����?�XY|
�h�t~�� 
�"�����l�b1��"Ɨ6���f��m��%�\�U�ŵ�4HY��������u�5�t6a+��o�j��b�;����ȝB�X����'< C^��N�§������p�^����w������W��7	
B�t�<��w�~��_G����̜ǭrh.d������$b�#(�:��ũ�3������!�����:T�(rپzl�����؈T�U�MF���`GEv�����冷iS�s>z<ݥ���v�×�6����=Iu��do��K����h��P��y���hu�`0o*�kn"Z��Ǚ/���	������'ѹ�|v�wT[,�*%���5�"� ry
��>�(3 '&2m]]��p�vMLp�D6n}�R��k+zя=��r��xe"?-5u7`�����mͣE4j-����6�ijn��E�^	�U(��96�NL.`.Ҹs*!�c>ξ_�@H�-ͿΥ�rs������%555�D���k�{���]w�=�i��B�0FX�>D���f��hb�ͅzyLR�l�=���Y��p�'ė���Η�|�Cߵ��>�����Ed�ںF���Y�{Δ�,3�)����#�wAM����Z�Р���^��ii�z��������mA�I�I?���}��n�~F;�8�ba!�/���{�ϯ��x��v_�+�nb9��GD/�w�,~i��X;8(�N�hTUW{�����&�x�����|YȽ�w~?AP�%r�rE����б%�"1�ھ|���] *�1kZgD���~,OE�0�}�l��C�g����~V���=���&��N��hK�LhK�5�<��.u:��KD�HS��)�"��oW]�����4;�dI�|�R7U���z�֔�:$��dm���ǏX+��f�<��~���ܒ�e@ 9y���
 C�X�������_����� 4�y��dNd���u����{�۔���s?�-�A�����Ò��yv���������v���cz��O��fr���f����^K��k���)��2������$���p�Õ��4�IW^���W�	&	��7��g6$��­���]'��m*3${���//C斗�Bca�����>����Eo�l�P�|q�ւ5���:J, D�R��w]�u����ggPg�чJm��������8���)�ôFl$$��ղ�ˡ�Q"uMM�elXᅅ,�ĉ��}+}�C-�HA�qS��qHk���Ņev�� Y�3�bVNL��⼕Y�3+|�?��~52ӫȷ�{k�L��lJ���8Ą������_=I�x����0a[��.U�{3������\���-����PfH�H@SK���f|O�Fsy�h�FUMG��v�(������w2�|Y�!}�O<=�
�KQ����@꣓f�&"&~jn��Ǝ+MEU��w�d�$edꌴ��avT��@g��߀o(*%�|y 2F'FKCV������IDH�Ch�+�=����𹶨g�b���.Y��3��}��q�?M��|�u[�y>Ҋ����N��<�(���	����e�������,@4�
X��	
�:���ǣ"g�[������K�����XU�0Hs�'����x�,oim=�w۬s!�����'�/?� ���_��.��1��%�y�%)yiy_�e��aY5'������a+��:w�Wll,do�9Ҳbt�>�R� /���G�����/��L��$JJ˼���A�gV׮-�=��-��^�.����~�&�� k��K����7�r2q',���[F�'8&~�_V��[^�C�dk �|���e�Lg1���;�Gw)��v��"��9���==#��nWyHп�I��f?6����H*����)_&�������#��O��?AY�:���+~֘�vD�݊��O(�����)CCFĦ�'q�	�ܻ뉰\M�9o}����.�������)I��x\�n���];�(j#����U�R����Q,狭d���ֳ�������s�C���;��v˥F��8Cq���	:���DuWv��;ᨯM*0o/C⡧w��?��Ȅ�T]�U�	l�z��%��'���\\\���%UkDe�{��&�0ɩm @�#�ĩ�<JK>궎��i���S_��s���S�hδ��1�F��2+���dm��PVc�t�l^>���<	��C�È՛j����ن?*�����{p�-�9=�Gؚ�v��e��++lm��G"�YUĞ�Ƈ�6?�
u=:$a��
#�ĭV8�B�ry�C)$0�龮���`�����V;k}�o̪�����w9�R������lh�i 2i�ث{��*F�/.f��� S�P�
�w�y�V��b�[��������H4���.�y�H/$�3}+���k�30].����Ε�����נ]����{����z�8X����l`���tTҜ���3�b����%?���@��f)Xb����? �#���yh֪s����$��=э�[��~�`	dO����q���'�d1���Q"�=/�~����d�a���uT>�1��	 �9������:�Ur��;qp|l��	��--�^�f#�����[�hSp!˄�7�'�.|��hl:"X��fb��P���Z��&Gk����(�� Sf���
��-���g��d�!!1��1!~�����R��u�W��֞��1S�얠�t�M���d��M�Y�p$��Ry�#�"��j6�P;wF;"N�Q�&���`��.楫&�遊�m�#'#�9IB��fǖ��[��#�/!��QmR�=_�ɕ8<��R2��M%�Ð�lEmdf��n�9��#� �%L�/�!�ZŠ�7���e���$�Q��a��ddf�%  �������{����=_�I���I�x/�����8��3o�æL,6����+���
1YY��v��<y�����.��u�g�=v/���KXh('�ꪛ�fm������W{�#�mZ��阙'N ^�^0���o+�>A�p�q�/�62�Xh���WM��R;��:ڶ�Y�n����NM��@����Tѭג�,�~��Ti�}!z�`p}{-���9Osi��Xz�?Yii�{wщ��0S>�&5�D�ļ�"��?P�W�8ݥV�r�g=?<<4>��ZBp"�G�B(`d� $q�_9�@|z�I�v]�E�ynz�I����؜���ٜ�+��k�}
�!���Ǚ�0/0����m��6����`%���qP� #�B���4��� �0�<�	Bb�=�©��o���Q�0-�4�����>��7��M�ŉ/;����1���mϬ ��WI���o2>�q�K��ɪD[�o��������d}����݌�JLL,i�@���'޵}�#�Y�������������zK|覫�����Eж��d'|%���)&\���dA�U�'�83a	;r5��Iʇ��Ȑ��1���lП*��rH�橵+�xP�bc���-��ٯ_�y����wŷ���>7�61<���h=�J�������� �dȨ�ػ�3���?� �>��Y�~�CL/�a�$N�|�i7V���GE��SS�����#�ohj�C��Q2cA��J\�Ѯ��']Y���w"��L��eX��=*E����/��*%��͝�����˗���|����-,��#����^1�mE�>�"��@|Q{h���#@�>h���.)-+�7��|����0o4bO�y__��49S�t�&(����
2'������QT}�� G�_���eI�������J��o��۫���.1>\nmͰ��mE;���;=]���!}�)�1{vХ2�k��~���pC�����O�:�}_On��V�'H@Q�jAs��9t��B��Ԉ�O���_���������"��>^��a��_����e��z�
oi�v�R�rM�VM0��*�kYOwoo��svZ��:����9A����#g��r�VV�,�?�Rc�Gs&(��`T��?��J�Лiq��tO��}�����Vi�y͆m��-t��Z��PR2v�z^��k?{F|��DDB� N���+�� =}���7�,����o�Y��Mo�R�~_��_׻�~��8�`�!/�z����OS���2��<5�3��8��z�$�ܰR��9{i��Ü�2�a�gK����d�6��Z�Q�Q�UGp+�#$Kޞ�.�e�Ff!Q�zr�A�����j����1/��S��ՕQ+_&fv��NXNe�8��$u����#�Y�P5���^����>�<Ɂ.n4sQ�,1�rRXC��:�cbrA���^�Cvp`��;9_&��9P�}��;y�Ԅ/���,�#5�w?8<���p����%���~]ږ�_?�h�IB�`b��e��i5=�'�
O��k6rݫ��翺��5ƌ�49?�｜<��^$"���$�Ǐ_]�Al~w��Z��-B�1|� G>��>�&\����^�'�6h������Z_�*o�/#�7�����0VU�D ��O���,��S|d�ӗ�-��w�EA �PRQy���l���+���Z�ww=�[%2�G`��@���$�#�͆��{�1f�jv����σ� f���l��	��8h~�������W���5`他B��I��O��i�����!����=��L���(��v�Ŕ�/ŃMe�_�.	�JW_����:.ٔ�
�wk���׊�S�JEEȇ���u�u?��ؑ��.�{�K�/��"�&!'�;z�X:e9�j�����
��+<�IAaa�*������i11�*I�a/��-�ϭ��;��t�ﭜ���t��j�s*WCg��*C��x��X���Fv�����XV�16��[o�_]�4��Q���Ȓ:����_o�q���-�utxx�EL�y��[ޡ��۶���ᘥ�/ֽnv���P�w����5������^��2w:��H�4����(zt��A*#����iq�>yW��n���%���/!�����P��v��3_���jW�S�|k{RGmʷ���OA�tR���d�UU�� O�Y��_�nRi�?$b��ikߌ'��g�V��辽L��MD�O��N��qS9����U�[���k�f�پi.��y��<3�Wq&O��\ڷBo�UL���[<8B'��s��-Б#o��X<̶n�t;˻����FG
0z*��k���X8ן�����0a���Ne�iAp���i�g�k�uz?�\�D����z���Ȓ;s�X~������h)������[N7�	!�2�3��ٔG��u�K��+5��۴_"�����|q��'Yn#cq��h���9�&�<��۶,�r�_��`Z�c��e}��~oo{�o]c�g��Ǥ�'�09�-��_�XA����;��q�����C�����.C������#�i�_�n$§h	q�x��N�Y�C��ε�U
�5�-&�C��o%fd��+���95t�,���C��NEm/�>���}��ݺӆㇶ	�`Fj�ɺ��8�Z;Z:|캖�,��܁U���T�Z:�K�1tOmO�GJ�^ּ�v�6ō,��5:\�g7�;�T�/�e�++��]`t)*SssV�k��X�}���Ԅ;��	�4�T^^^Ō���II^�*��-c��"@��ו�M��,0d�3���42d)T��vy��F��)?��S.8���8�v�iX
�|u�m�ǚ�ƭ��C�*�-πmQ���p=�u���}��N�}���l�X�߿��<��yI���Q`������pcjB\�㭠�B�I�+�Ծ(���ۆ�&����ɐ�}�'㵡Q�����SW�%/��;����umE��m��^8�8Lͅ��(q�mk����N�.��4���ɉ���Ӗ��[�LII�۷�i
�x�^�gO�L�M�;���7]$�w{%�GPay�v�S���F���I02��@O�.�X�Q�#E�[m���r��\OuUA�����Ɗ��������4ˁ�U*/���bk=�]�sPz6��io/Q�:���R����8;�#"Y�_�6T'W�E�?$Ŷzpr4��p��ZTzv����un��G�v�򜁞!$�$�"st����3�4)b�#��XI>��&�����=�dqi���������P�{(Ԉ���Ü�5%fR��~��$Ԧڋ���{,$9�s⯢'7V��aK�_ZKfƟ�9ã,LpP�Z��\��Ɯ����&/ػ����B��OW��n�UVpwK�&�a�ݽ{7�R��%Tij�ǃL��1�Lx��+MIONL�&��|I�-�v^n۾�:��Q,'z:ha��2K�S_(�sm�%]4b��Ҵ�����\�@�s!us3�������J�&� ��ޖBG{K9k}��VAߊ��x2�8���>�S��!1��XS>'�}+W���\;�
ޏm5d�{���(z�1�9� 
���@�<gG��e�9��L�8�%��$��#�k5ߓ+6�aJ�[:<���		z�& +Re�� {�W虘4H�X:9��L�{��RUe�y��-�Ք�����\��d�,��l6wv�����H8f'���wp꒻@��Pe��@YdH��)M����|�(��J<
���(�0�ş���*LJV��jr�uVzw L[��o���
(�Qm�m⢃���l�]�e�ӝ(��n>p<4�ʻ���N��C8r}j�>�Aqn���a��g�՛�@�� ���%w���pVn����1������n利�?M���+�sU�PF�9�df�M)4��S�J���ȽŴ%6d� >�y���y�V#C8�.�%`�ݥ�&vf��ꠧ�LFkA;q��������MϠ1�n����3l+�\��-!yj�cx`�ɒt$�����DCs�� ������
ۼ�VRߊ`�Vn~�J)�=��z �''|��P��'�zm.���އ�'r	�$�k��/Eғ�i��|��Ԛ5@M�s��Y�i��=[lZ����(�_���㝜�N���i�Q��^c9�8�>X�9Ig�j�uQ4yP�$
j�ZX������z�$�yz��p<�o7�X�����+��kE����Bs��S����\+o��#�Ѕ������gdİ������軷� G$��Vu��x���d3���4�6%&����B��oL��$B��!��R�:az� L`�l�q�L�8��gr|�a"����B�	}����or���Ń�^��E%Q>UJ�2gء�]+9�C�����!���OdI��^��������B�q�x~�S�����]g���9W��W�Č3 vAdr�9�~�(CX2 ��[�x��9��0_`�:�J(mT�Alָ���xr?�gkce�)W���Q���n��Ut��ɟ-���$���p�Z�_C�w ~-8{���ϥ8W��7�(�Zh]�5h��s��u�6L�����ʍo�6���^QR�ԭ�����W�r��L���$ʏ)*")�|���911T:�v��n>mǈ!AO�1`��oN������H$^ٯ�DLJJʝ��L����X9�`*���-.�[�q���a��`�m��i�
�c�?�*����/��D����6�ʰ���qF]]��#�W�|t$�oФؘw�Vr�HijI���v�{K��O9h�����6�&K�k��o_�npa�d�I4��j.���y�)�AoR]�Ph�݃^BيY�g�������=�S^.���&.���(S��{�u�l�w޵�E}z�F��ٲ�k�N텳�����Z�w7��,�7��$Y\$nT%�3�����	rG��wg:ն�����ǹ���5^R�2`T���ٿ˹�Gq�.\d�W/������,��Y'	����(�����|��f#���($�+z��I'���=c��|����s0��	nE����1�C� t��ȓ����r%�@���E��qKܜLK\���C�y**a�����U��/nmz�>,�Cz���k���Y[_�w�x� ����15qJ���5 ]7���O��.�껺bT)B��Nl.Ϻ�E�HYY�t(���;/Vk�c]�K�3�.��:��M�[,(�?��p���[h�9�HT)22���e``�r݆��?��+>wp� z}X����iq�^}ش��h^� �×� )�j��s���X�X���"�]74r����m�T�=X"���ź�O�����m�g�������C,x�k�\��$����Ms�h�ۂ���t��ܰ�[c�PL9<�65?ˌpL��b��o�	#╿�ʹ�a��E?;��)�,;Ҟ����2 `���#t	6�XUB�r�|���e�v�h���JQ���Z/��+��
A2J�����,�{� A�!_k�աuw����T�C�_b**�^I�$�����m��a��E}�D��ׇ�R��8P��pvu���C�5`�4P"y�'�+��A2�?<%�iI����Y��Q'h^�7�<��gfEX����C8׽�2}>ޡ��ʑj�Z'�ӑ�]��v!
m��f��^V9�����F��M_��{/���� R�lRbE0�\���R��^$ҵy��N��67���罽��L
��ϻ������뻏�b��W��B��N�sv>�z��-�5��vQ��ܹz�C�׮��"黦&�)wz��%��Y�@�)렐��8�
�>A�LgX�$~���~�s�}ޤ�ö�~���/o��U�s�r����T�#֒�l�JTc�	�����'�*��k�J|.����G����Ax~I�n�m�׽��u���OU��@���3���t��u]�G�<ԝu�Ŗ�{�;b�p)ǭ���ۢ�Ti:3���� �����]r��+���xxT�C�s4�Ss$�K(�8A�ڳgĜ3{0T��S�v���))�KF����N;<In/� �9h�(~��ߠ%FdA�\'GM(g��|/0��	�Y�5�7�f����n�����Y�)eQ�.����+ƪ7\�ZZpl��We�a�)���� ri��|!���h���/�����T&y�v�z!�O���&ݟ`������32�U_�Sg�;�cc�X�I��x���P��E�����mY��$������3*�5���`��J<��T�W�� G�Ǳ�h�_�n;!ȌYҍ���tTJ���D׎t�UNn4��ކ߭��
���ӹ�y��;������o�h����ᑥ����P�B*;�(�����n\o%֡ #|V`��t�=rӗw�9�i�V$8�yT'�YJ>�יN3
��&���\z���؍���\�5��X�Y���V��(�܈���̥%�q�">6iO�EjkZxE�}�q�L��P�ߢC�5M ��L���-s�	��<M��4cJ���˧�T�=?=�ssݵW�n�ߜ���E��n�<���[�k0��a���^�4+P\��jhz�Ʊ)��R5vG��PϽ�s|T��[�����vy�Q�Y����;�+~�)Cs&��7�g?/q���N�O6l�<�̚�3hmmc�s`�Ά���X� �L�S�G&œ��o�ί}Y��I.������\p��"����ܦ�
.�vh2��`��=�$�D��}͠rV��B���� G�HD�ƞl^�7��
Z���������@�v��'u_6~If���u�M���Ǔ0�=�dk�?AFGd��qm��������"�ڥ�5r ��ÛLهa�**$d�C��V4,_>�]��p�=��-��lNY(+�-	�֝���6f|6e�����;G�|�{��٧���?�~�ntӷH���ō�l��O�,���)u���M&�%ni��$#$ͳ�b*O�[9^����v3!�B�:~�g^d0B�~���ntX'p%�MJֹ��W$z�$�w.��l���$��� ��@��I�Xr��u�L����i�����X櫻D��.�\�Y<`�Bt������.v/����Y
w+�J�}��jK��X��������hv��E}%��2�|*l���Y�1��ϯ]nj���b�u!�ܑ�ud����:1L�����.w[@ظQ��&��#E6���������3z���=� %�i3C�%f�x\n���b n?�/s0�����~��#k�C�+͋Py ��M�X5ĳt)�/����.��g,y�h�5�/�TV����9J�~-���J%
o`�ja�H��J��2��%߷�ɒ���>��o�����*ྥ�s7���)���c?��h)�,ʺ),1�f�3i@NS���o��-�/n��*���}dJ�F&ff�P�&���F��4���z]�Xk������g����v�q�l��߿k��;�%�^�q��CvlR���B��O��*&���UZ+����ţ��Q�j�2��2�u���@�3����Vp��Yy�"�`��}�]���)V7�ѻx��\�]����7�Z��*�P�X{x�0��]�I�W�B��W��-��CMY
(�_��茸W�a��� �0��ܵqȒ���m(�v���F���d��<^9	��9��Q�8�v���RҤ�wM����b�����㋶�Q���;�7�}
���=Ʋ��y�j��������4�A���{` ��\�����x4p���hϖ�'u�V�0--�,��»öךLƹ`�"�����y�:]QP~�V�P����p�l�X��l�a�=�*y�C��>um��Ζ�C7.��m)��7
T�N8�cI�9�n�_i@�!s����\�k��m.
��Xx2�@�k�I��U�O+�ٽ��X�cmӕ��5��o}s�og��Fw����R�C��#u��*�[�������C�]���B�#��֓�%��RN�^Z��я���Ε��x��qNw����>��UW�|0�=)�/xc�ơZ���ܵ�b6��\'h3��I�k�!$�����V^��~��
c�������j��Q>��M�И����cn"���a�Rd��✌B��
��Up�jR}��E%��Q%��ݠY���h򾿌霬R��p��}
e�0
����Q�L���%(���^{�_(�$ƈO���r���7 �g��`g� ���;��l��	�z���><�߂-Mm�D�և�NIyyħOr�s_)<��qQ>~��C��s��K��Ӌ���˼���au\w�$��� D�vs���8g����b{�D�!x߁�z��q�u���sr|>c�|���0�2 ��ԕ3V��:�ȿ������D�,�I+�n��Y��q�bہ�9>�;w�|_�7}��J�4����Uw	���(������R)JQ&_ �K�D�&ZN������2��h�P|\���	����g�2�� �����|
��_a1�͋�9�cu~���Ô���tR�=� �ߺ#�2��;҂2R���ߧ�V���f<�r>q� ���"� O��ռ=���lg	c�u^e���x��q����K�(E��XAPh�mw��o^G���.��\ܫw�fܳ�1x��G���������lpmN�"ҡ��U{af�������/��4�*^��q��K� _����5/�w@� ���`E` ���f���z �/3 -��4RB�����'論��7����v�Ɗi0f�uD|�{#����L�R��S����~on��x����2''����3�X�"'�dnb�=Z�u���\Hjh���ၗP!%%%�u�8���<����rU�4Zn�y�2WT�������P�����1'�Bnw��U�/�P��]���wA��|����:K�w��YYo ��6��/��mKY3.x

�\F�w���>��K����v�s+$m6�WR�l�A����ÈF����EP�(g�ZSdʷ��,~��3Ǧ'��F\����B@�?��<� HJ��F�돕]R8����&RL��Ǐ��4���USP�M���� �
=���F(&%����Ħo]þ�g�==��T�%��G{J�O͇>5�/ېZy:�0��[�n�ZZE���6qxH���r>�����"�g�6$��ʒ#+.�Ύ.p�>"��
Q���N��xk�}�f|;��(�d�����f|m�[`�3�?��%�GքMu~{�  
P�'��Ts�7.Ed���{�#�hZ��L�X�Dd>P)�E(`��#�H�gc��|���)��3�_��	��Wt�Zt�q\�I�bt�m����W�57���)l�U*�ck���d�!�zR["(�?���t��Y���7"9���~10��A���6�ε�ol���u��.Ri��+��_ �r����E�6�K⦣��ra�z����:*�wӍ�	Pŏ����:��;g�{����qH�t��\k,�_��q��a����'C�I�ꔷ�����ɖ�����#���s59I�x�r���c&��c�ǒa�'����L��	�vG�5w	f���[�X��?���@��X	�c�'�N���5�c_һ�̿]P�:��Ԅ�(�`o�u���1���A�M���d�˰ 
C�6egu�1		Hbے�vd®��� m�mw�y��1��JA��ً|��U��;���g��je+7���Fʙ�)�9>���(�u
egWW������?<�o4��t`�3Ԫ
Ş	�m�G>������z����B���ҭ<�a:��c�{0l���'V,rG>�黑w��0Nɿ�V����sJ[�Pr˻�6ƌt+�R�Ԅ����Bw7}o�e�z��[`R �m���M��e{�0	#x.r�^���*�O�O�d60���XPrz�"��J��X?��j���¨�������܂��0��@�֯.�`�P��ɚ�Yɖ˺���� z�,���#̑��Y�4��թQ��T�E��Ǐ?|ot�\�^Y)���U�շ~��8v�/��*�?��*EH��_�SJ����p.\�� W����z�5�N���fM�B��TOȅy�����*^{X�0�*>�+\!w4 )u�.���2d�J��IkY��8]��[��a����9������:_"+V�Z��/��O^/~���F&&�?���S�rk�*��L���VMa2 ���l���W���{�Ϻ|:B�c� ��F��EG��܈ݭ��?Fڋ�RC\l������3[2�OL|4u`1<�uj�e�/N��w(�E��Ӧ<�q��`Gw����͔�3�]r�I-���F���-�j�E:�IH��7.�82E]��_��V�"��*��]�9��qǞ�C�}@�tTY��Wj��qQ��U8�7�j	�a*!OW cj��<����|�aƗyi5�B���SU*/vBԏca������� 2lԄs��P������\��"}��H�--�m��J�;g%�d&��z���RV<[8NB�4f�q3VE���fd>"�X�YoLL���]��,���g��ơ��y?O��<�v�8���⨾��=����BO{�z����b9+V�fi�>7���cô6�-�H9)��(��ˮu��	6BOO,������7��`f�?ִ2�\�R8�`�a%�S����z��A��>'�M��.�G@?\F�d����)=�r�Ț�GJZ���M�|��cJ�}����ɐ#ױ��w�\�7���Y�sؤ(A p�ж�x�ח������S�eu�+}��p��LǊ�u�=�%�J\1�"���e�"wp����@<���נMbݳ���+�Ş$"��u����59U��"K�hm.�u|���?�yp����Oѿ�ĝs�#�M��䶅"��5kkS>q>�A��z�=v�Q7TǦэC�!��PC������i����:�60S��Hg���&7
QVd��u�M?����\#*]�������e��G�ܨ�y�qF�V8�W"�J2�����m<ϙ�A������P�xlL���nN��ߝ���KYQB��`0�ϕ�j�Rh�3̝Dh��O�GSc�T�im?�8p������S>���"qu�W��KAW������4X����611Ah]?}C������#���q:�$��>H�'�)�l���'�q��o�]b�n��W)V�S�9� ��-�CFo�z<�׿&X�����ǔNb9FFF��v����`Ry��C++YhS�4�xpejSP��P���C�g�����PgD1��i�_�P6��e���8n'��9����A�8���Pצ/�{k�y�^���o_<�]�.�0Ƹ9�����
�S��cɺ<W��C/}��s�ڤ/�`i���hjiM/^b���~������%�.Q6&� $�XrO�/Kz��Ǚ�ȧ�S�pf�{�-q�P!��j���Ȳ"�Z��u�j9�2�q��Gtx��F��ň�Y��k^Vx0���n$Ϲ���0ie��J�����o����7�Dn��r�D~� ��Z�~�!E�"u3j�P؂�$���,��}rl�ϝ���sQRW��I� 3�x��lh
	qwCJp�V�#1@���a�@5���M6����kfƫ�֍��P�k�LQ( ᥽�!'�V2`�T#�Bp1�o�i̥����gBw6e���(=C�;��B{���Y��!!	�|
� M���M���Ǿ��,�8D0ӈ�&���52��(Ħ��O��]MM�V����A��V ��^svI��T>yv)��W�[�Ī��ƣ�9)����]ϔ���KƏ�� O)�>+{/f�mDh�$�YiSh{���>̹�̐$Tt�]mh�0��]��z�֯C�X%bYx?���o[��XRh'Ij�u+��x�aִhv���V���:P
BY��܂"��ɗָGOw��J��w^fx�G��Ϋ���g��vL���d��jYV�Rr����.p⸩逾��x]+���+N���l�s��r�pffF(o����Dي���X��;K��d� ``����K z�j6���U�F�(Hu=����<�"�����DZ�M�Y��<�ҵh���_)=1g���5Xq�L����b��0'�pF��������=h�u���%�ܤ !j��B�sleEJ�a}[���{�Ն7.CG"�; ���i�O�ho`���-�
E~"�	�[�����Z�|80%SSS�Dh����0�r�C{�H�����Z�x�_��'�Gސ����fU��ǀ}J��A��
.?�<b�1���ڇavӿq8��ЦXyZS�*���<oT]]��|2����/9�l���'?55Z��H�7������:f��F�����1�+1Lo��}92���������/�&n�IuF��p�o[���sb[��wޒ
no3qފ��K.�=�_��L��@ܥ�"����Rwr*� F�M���N���͕�C	Tht��9εtv��`ro=���ؘ��x����67g��3%¿{M�F����Ni���#6i��4��]~�˅ʀ��C�Μ� 5�D���Z����]������Y��u4ڎ�<@�ͤ��X��O��m��&& F�6T�̏�,�_���
'K���l FJ�J��m��[����!nD�������`��4(1h�	����S�pm���U�^�"& 1kkg1i�eKK���ץ���%����G�o�_��KDz�t+�T��*T%���Fd��3f$�N���=�G@@�n���=?���4 �&%9�\b��ƚג�����2õ����E�Z�0U�yV���#�
"N)7/��0i��2iiup����g�###�{�ȐǦC���bD@����(m`��bt��Ban�!
ms��bA_�豢(W�T���Utz�x���� ?W���x�~=�W��Y�F�����DT㼏�:��^��8>c<ܿ�a&L 귅r�LH�m(D9�n��F;6?V+�"J�,�ԏ�Ӹ
�fMS���hPRʧ��v"��Ԯ�5���X(��;
���\g/"���!@=l�Tm��,8@�4�~qd�����o�E �)�ou$�4��>-�{r��=���7���K�D$�5L`Rq a��Л��+�[��.X�5+''�kkv�6*�w�	� �x�_�<��}���gƒ ��c���'P�.���������}�ǉ�l'd�	yKƱ7���!;��{dfd��!;�^!N�N:���N�w��/}�����8�D�����㺯��19u����t�OO١���C_�,��ÿ��_�Q7������]�E�&m�F�[��Ũ r�/�ˋ�Z|,9�>gĿ�-�e�4�W�,x>ӟ7��lh|dV��A�m�la�d��7�'�D˃'�Z�dR���><�
$ �8jNDR���gk!�{ 
s��� ��
� �ݖ��6*�&?*��;3�n��.���"���V���B��7�t���T;ǡ�<ΠG���>��^�U��k-Df���w}/HD�'G��u�+���[_::.�t*��XYY�����[������G��,>#G��I|ެ�`vv�)Y�D����,jƴ� <���S���[�B��A*�Ss���;Q�{|q�%������G�\Q=������_�>�Hߩs���V�,��'x��f�3�u��Y��N-��،�y�VV�"�痟��Ӵy(;SUj&ydV��o�z���z��2&���2S� B�W+}��Sj�Nɫ����[}������i :��V�b�9#|�hK�ɢ8�ͭo�g�ҫ҂種�6�?�F�ڱ�]����"�W��l聙�L8�TU p��J])�64�����}5�>ԉR2�WK����߿/�8����L��yt��1�#(II��b97�\; �|���R��ɣ��{8�~�-��c��c	��3j��?�n���zn��4�'�=��<1���Jw:�>���~/��u���F:�%.p�M��X���6y�\7�Y�"��ņɨ�O����Uj���@�%i�]��Ij����LU��z�U������l��i�:�r��Kp�J�L�L���#e��/e������̥����E؏m) ���m2����'�8Z*u�Ļ���s��;i�P;�X���q��^_T��X��:L$iկ]Rvf���1$z�O�v��\~-�:9
���7��(ɱ��T0����w�8T�6��uͣ��˽Ġ&�ET9�����p��wehhg�u�[�wS��?�i�W��&�1�4K^��T��.s����HA�� ����v^:��u���v_Q#q^�`�R5���ܺeZg�]����A�NB��[���-��]��F�Q\�t�?-�lUW����M.��g2���_r�q�-e�ܭ`j/�k@�}�[EE��B?���N'~ GߺN����aݩ��]���ގ��n�rt]��SR�n���Y�?n���Ya�-a<pl�j�<���~� -�=�z�)p�,�<����ܹ�x/_�
�ͰT��~�2ުNZ9,��:]������M��;�t��A�\��Rǋc��3E��f�J)�P�A�?4��+�^j=�rA0k����"��Hw����r��
 �����סR�b��}�ʵ�U�Zet!��6D#b����4�XaY7�� h�[~R5 Ғ�+��gۤC;�_7J�����.�"��Fn��|�j�e��k\?�w� ���݊QW�|f ?[<�#�r��fQ���sM{i�$*К��+��q��)[A(�l�h�e�mp��Ղ�����
��_T	$�N��kԶצ������~�$����w�/����@�R�<�F���o$7ɡ^���#�ݹ��gN��g�+��x��]�h	H�Mh�޽�Bp�ɠm"Z�xԿ�BC ,���)�ٜ��a�*Nq��-��ޭ��>�>�@�D͢��$®���i�8� �2�klk�o���¤�+�.A��g�!��N�{�<M���(4Ӂ�?8Q����5�:0�*�S]�
�ϥۅ�vq{�����9�?-d��S}��r]8��I5 w6>�3q�k���sS��\��V��5�4utD���
9J�Z{x�-��n��k'"L��w�<�&\�U�bc R�M��;>��V�u޶O��t$���81�������*J4�4S��I���z���T��բc"��xi�k�W*���ꛘ�I�G�hX��'�2�=%����Q+uZEϭK�Y� �(~�jZv'����$�~�4Z	H"�jc�g��Tq/����1Q��O����Fv�P��o�X�x$7�,S2���Nς'g��w3�gO��?��wiR�����̧�m�=�e}���ݭ.>�K�}J]P�1e���j��n+R���f@}s�Ñ����b�h�������B^�d�<[鄋Y�x�=++%h���"z#�i����S�kO}�S�+��-2av��ٌ����U��LC���ƀ�|�_~��r#^ͮ~z�Ni/�0G!�>(J'���1��8W&
G5���)��ʱSCb��u��U^[K7�).�Jj��- _{��j���rpx!&e0��^��t�˝����C�����W���^ٖ�Y�2��C��YB�)H���h�n�i�8�����)��� ��{���:I�mq),Q.5X��ؘė893�,-wx�tB�� ��K��-e4dLu"?~XX��s��k~����trA#f��+���@�gty��}��F�ۻ)��Pé)���kJ�{5�zz�WV�	��ou���; ���H0����s��k2;�o�o\�9�QR�v�/1ʱ���d�U�	D	���<�ڵt����S:6
�R'���3���C8����[�uG� K���A,�60����(S+����,(��W�їՂ��N�7L��&�<@�5����g����ʃ�)�d��W���v������~��B~���jI���T@:m�G	<h���9*A�O?�oKY\�� ��b�Φ��� =������)�Ù6I�����wD�@���/H�J�^��as�Ȼ�au*A�6�Hŏ;r�w��e���-�+��:Fg������ϴ�����:�����n���Sf/pwK���du7��8�~E�,�%��Q�WW��Y�l���r�W��6ͽ�,�J%�DA�Q=�L�؉ّ�=�3�7Fr�'��a)�p�tZ�EQ$��굎 �����>햀�*��u���"0K�|05�<en�fG�*E�5q���D��^�;��/_��P�>+���m��u�aa���*`�}�ݿ��ktZ�Ŀ9��Gn�������<�7�(�>6��N�	����㱫o���î���^�*̍Ԁ'��9�窕��Kݜ!G��_�;�7��-"B����<:!+Z�F������z��s}��u�G�b��B���2Q	�h|��� ��.aP+�+�C>��V�k�+>_5�t��G!�f_������=$v��j_���-Kr,�R�XS��=,�jo�� �A��+Nt����m�%�K����Z���#�e�����W��}}��u�<{������"Ɩ�����v4� �9	�CCT���:!�߼����x��|6��"z��M����r����\���o;�`Z[���U���u-w�5u�СZ������Q�zu\L����ddG���u�@��|���R���
�j�D�5��g�91{k�/�al�b��U��=�\���[�ɿ`�=dV��cX�K:lO���Z�ë�\ę��yJF-F���c�J��KgQ�r�޽���|���"@���ڦ�U.��������>˗�|󩿜�\��Ȫ�$�(NN֔TK�I�������gF��94�S�,���*tp��aH� Óa��f%S����D���� � �z����T�>R�yc�H%P��2�x��ԥ<�GKKW�L�o΅UO����=|8zmٯ}���~���>����"5�>iT$?�=;�Ɨhk`�s3M#��荋�\_�߄g���w!���8�yQW�1@x
f�K%кs�H�M�,�L��0B�@���ƾz4���]V"[-������ZN��?��W��ϱ7��/v��Y�5]uB0�G�%uk��}����J#~�g�zb�P-�h�gVuf�Wu�˝����W��]-K�z���קD��Qi�U�*^��2MQwq�{�Y8��7	 Ua��)�Y���q�:ec��4y�xC����2�.�Wsg�o��p�w��<}ޢ����}_��~�]M/���ߗ�9 �;}����V���0B�Xڶ���Ȫ��%�Fuq�.#�ި:$�h�ͭ%��rm�v@���2h�BO.�Ǹ[cZ�J���c�+J��,���R4��z�x���Z�U���ܘ��Zgs�s��y���@,�����^�`�kT�7��*X#]�BK��5?��!��y�^�<��;��66�=�"9c����6�S�/�,xڣWˁ_Q@Y[XA��E�H�q�6��O�/�K���%&�k'
�� T�<}���}ꎺ��ܳԄ쩤�ī>��ծ���Sbb$/D�S\,W��s +-��C���tx�{q���0����B]]}Fp�ݥ�\�����A�����6%ԏ���5?�fs���ޣ��r��N�S�����slJN��+)+�c���S��7E�1ˡ�ë����pͳ�r糞�W����Z92{)��*��|�3k�4����NnI��*-Ӈ6A|�2�x���C�w�9t4 x��^�ZK�L�ۊ�n���BOu��x���cƝ>���K�j�&[$��9�g�$6@6r��_��R,R�/�)ȟu����I�-���r�!b�\����v9$4��u8��YK��x:�w����?�rc�������跡㝳r��=�d��LӞO.=�Tz������f�C�E7�����bDa�,��I2!E�yy�Zֳ�$���]����ZZ6�*D�Ti�)DpZn�M�Ն4���>[��g�35%%z�bE���_�D��X �/�.?����Oul�wG����V�b˴�Qg-^R2 a{���0�7x>����P�%8�]�.�}�TI�H�F��HFfze7H��JG����QL���7*��)x�6w���S)��h�Cn��4��u��/:w��ۖ~����,qz?|6�	"�/���:�?�"�9X�uָjo�j mjn����H=<T/�{�"89|��X���\�`N?&'�66o�^�����{rv���MC�etq�:4���8j*j������kJfU�t��d�+vv$����Q0�>7���)j�T���z��r8�'�=NX~@�ⳋ��C&�:ʥD�:՘Ca��e�ߞ����c
}33�@+{���S��찺��tߔ�u��O1]��I��0{/��Ƽ���ΰ���e�_c����'R�8�P��j���洬�&	�Q�`"H�ݯl`��~�A�t�����|,�N�9��r����
������_c.Rlu�/��JӪQQ�}K���{�'���$�����
_P�h��a�ro��}�>���N�CF|�B�� C��{���_�����{�DgM�J��jo�Y�i)|�R�������gi�"� �S�� ����~�פS.R.�8�nϗ�;}�pR�ډ]� �6��2��ӷ�}�"ovy[��e˃�lT0�I�UvAǎ6{3nx���meQ@���z|u�
$��C\���59#�\��V���v4��o���t~�XX*O�fu?x&֦�T �u����q��{U����5�	GZ1
v��Z������{?�[O�Z�O�Ԋ��WY�xO?�?K|��+�����쩼%��Ҥ:���L��Pvvvܛ�_�$����|�stp�����X;�4���&��SbB�bAsݕc�:H��%J��O�V /��S£�|Άhh��ܩ��Q�`��}A�&1�;�S�� ��n�{q�)֫����W���Gn��Ԯ�,�*
���<:!���&5���Ȣ"w�kL*�n?��l�'kN��b���	P+r��}���+G���T8iX|u���C����0^�W�mQ�ńK����Wj�K��_�S0(8{��;A������z�e?S�!���	�H�mmꗗH���xa��k�
$����a�O�S�n�G�ЖC�42�����
����vw;�Fo� SI{��Y*hȈ���4L$��s��6�����^?�ɯG�CC�nn�d���8F��� df�»��6��TӢ	h��3����WW|�V�M�2�h�
�0G�g�}v��7@�H�f8�ƒXu����5&�����~��0��pM������:�P�o8j�$_R�Z�ď�ٽ[߷C�>4����uCq�Ȣ�f��4?������P�ӷ&��4��� FKWs��~M� ��Q�$��ǔ�=�����w�3�Rq����(V}��������e�ݖ�DW7�����+���%��^�Q^p�u����� -b���`(҈�K0� S�q�b.��V<4^�m�5s����ݒ/B���R�܀7�}W|����f|��r'�8%��[�Q�xj��_���䚟����U7u+�����1V0���%zJ[z���Ŭ�������%���72V�R�1/�恊��h��*�X���{����7���ei-!�4x@`�0&��qSpg<�X�m���l_^^��:��)�m��Z�f�2� ��!�פJuA-��įr14���q� )A��'"�駏�X#j�f�[Yyx�\���������<�^{~�ͣ��^W�Y�Dy�O??;�6����H���WV���]��i.HO�������C�nğ�[ѿ��ܪn��#,ybb���x��� D��ښ�A�=]{F�D��A澎	��}2��~�S�4�d:<!��G߄×έwoO���QwZqTU)c?�L��J�kF�/����Vl���u��[�isb^�W[ٙ��tQ���xd����wԻ�c�~�-�SQ�W�4�^�yP�~|i�,�d����Ç��$�z�a��}?W�s��@�����������COKC�.8�(�����r;I2��G5����+i�_���СB��M�3��1�jC�-��T|�����<c��ub���hۆ��Yw���U8;\W���}BPv����>����O/cX�gi]�e%�r�
��TІ���_19��şs��EE����9:�����ܭӕ�Jc�0�ㄑsӐ�'Y����
"`^?���Z3�P��q�uڬ||���d���}�������B��~|�d�R�Y����K����)4ӹ0[�u��cʝ��rB�~�ܿM�&����ӈ>}{]��jGH�X��~<g���$N����p̱L�"^h\(r��.�>>�V��}����޿��i��  �Q"�������~!h'�E颔���? L'&|18�����K.ͽ*�H���m�3Ĕ��p+<?����Z|����͢J��8�4(^&��XI�'���n	�ɉ֫��e�v�HI��yJ]�j�9ƞ�^ljZLӀU��ivy�W��|���nbbr�5'��֯�L��a"��Vj����
|k �ۏaC�J�ll�����J��K��;�d*���Sr�
�|df]:�d:�t[Ƅ(^M��S�Q~Ƌ�%��x�3�K�_�d��Ƿ�?9eeK%���k�[ZOR$���ʮ`�z����ܣ�q�}��F mўA�*rZC��0$ �}S�t��=.��ĠN��5�O
X��W��ńI�=���7��i�ԃ���d<���3い ���w(ܸw�{�k������'Ζ��J%O�_?��e���P���N��'�Ǧ ���;���s��)�5Ga���*%��_��&�n�o]����@����Ss%~O�Þ`����0�5�`����}������*y�Z@Aǝ�z$\��h�hƞ�����H�\cˆ�ʵY�����=�f.�10�2==�h������h#�;������s�� W2ȉ ��gŌ�U��FʱӄP��3�����?N��{b8����h����"��:\���'���K���ޣ�ɡf� ��DS�
�T�L�8�˾������ʉ*��Z�ZUZzzay�8όh��aUX8{�C@h�\�/�KX��d�y��֡,�//��V
U`����k�ȽR�Oy,^W|\MD]gU4?Z ��ш���0?�B������!
�|�O�?�3����s����j[, ��,w�uTK��~T:�.,D:D��>��{3��x[WWW���]�Hp����+yw;M�MX���M�6�!v��������5�Gɴ�Z$0�Yv�j[��/V$2�G������ou+�Lk���
c:�`���wØŦ0���}�߹��R'�s9��y�dnJ,��a��fya�@����O�l`�H��w�:4���o���jL��d;�}tp�>�lf�L���MW;B�!&�=�٧��$&|�@�{�*ll<�Я�4���7Wwq��.p1u�����4vh�h��#x����R0�����?��i�:;_r�>���;>~atp��*Ū�B���/+�,����,��\�Ƅ>.�T�:7���y��E�g��J:������^*j�����V�d�ĳ"��8�4��ğb�w7�������1|�ňpwI*qx0��H4��mӅHfJݴ�h&�[�_��bۆR���7T:!ae�MM��GG��~���SY?��B"��]NE�	Q� kz�g{yn�x�)��uV�:�YYE
�����'_�$�'����o������J�0KQC��S��'�ŭ�'~WcS���K��q��r�Bu���x�:?02��7l[G��'P�`�=��&��ER`0�ջ�H#22���MS�;8;O��z6/�&cK�%r�˙׿����i���̅,���!R�4��� }K;���`�h����
�\� *mr�� �?�������J��!��r1 o�ӷܴ���_G�
8�o�u-|���KsB�D�	�ҹu��_��ς9Ec�d������b��jL�;O.��N?I���y����?=����n �]��r��$�g��g��z��Bv5jz�m��G�$��]�4��+�͋�z	�i�?r���7*������N/� ��T�ٹ��������z=����ٻW�|Y���#�	��O�5�x�c��3H�!�;B�v]�Qa����~�r�tx�K���}�:߸�E�np��3���iR�q�� J0Z�+o{�|.��35�O�SO�������22qn�Q-v@�:2I��i�����s��s����~�����Ch�=%�Wl��Ӿ������}���2=�?�u(�>1��k0�%L�O����;  ��z��F�P���j�����C�8�XHq{�>���3��qtU��Y8��+��+�A'��	��켼.m|WK�,yKJK��>Y�B�ዟ{�\� ��$�Ǎ-������7N	L��[�6K�`�;�Q��f2�6`	ع���v����A����t��a�/Hٱ��D=$ҧ�:�5���wP�8���̫�;�����|llF-Q���ǝ��C_��������6�.$OF����OQ,�u\����'�j�ܱKKW�mm�r��smv��2?H�w�t]�ʛ/�F�6�DC����?�z�iIu���"��Y(����/Q[��5��n���?ݔ/�H,qsbMg���u��Qৼ��-�(�ߥ���%7Imxq�{u]W��"T�������6�4uݧR!��Ζ�-saD:���/_��N����y�Ŀ��=4�S��|{��[X�Rb�/���C�����A�|'S��#���Pg�W�-mZ�U��AKO$�5s2�V7�-d�Ȁ��2��j�����32<�I������E^���!��HN<�;ې���)ڤ�d�e*3)ָz����1�dQ���00���:��Pewh�B�Y@�r1QP�2�e746&:!KKUt�3�+a(Nt�ǘ�V��a�,
D4�(���r01��5@�]Q���G�`zh�������%vY|0�{�-��r�EE��p�%���0��B?{Aף;O����W3ݪ�j�'tr?��z�5���F<�"t�ϫq"X7�4�
��o���K�.�z{I$�@��k���i�qT�k�d�������.�,�̼2��#]�?��3Y�ך,��I�}�[�3�����ۆ��βm�R2���MH;lu��Ӗ
y,_���8��U@��̀��@�Zu�������H��/�n}n�3Z�{��-G��Ӳ�xJ���Nx�Ë�����R��Pq4�~.'YnQ���넣�Qʽ}-ҟ�i�v�W�{H�#�����S�9e�h�VE�7����!]4��WjUW�]���mc���Ã.w]g�"��|дF�ږ���$"�,M8��S5�/|����s�������,����������_��B��@N���]����RJ�U�m(^�.`���~��߷�/_88 ����=�G�6�:
}�Ԧ_��-��e��I��&$'���5�_��BZ/��H�ۦKG� ��Wp����������� =$ٷ�N'��%���.0]�I�_�NOp�0�S��`X~�2�K/Thhͤ�B)��:����S��3�}1��t��vK���(�R�e�#��_[@m�~Ӯh��\����nE��+��/��Tܻ�?g+F��������N�t:����g��\(��/_h)b\�O�:>�ڡ����V`_�C�3��k?��o��ND���q�;<�ֱ�F��ڞ+�irF��z��ˬ��E�cL~)�y��	\���d@Viy`��p��=<E�b���j�}-<��e�o�/X� ���Z�E�fK�y7�p�j2��@H��
��>�rQ��>R�#��� �J�����`]�d]�U����m�*�+22n0��:�Ak�E��,�t~c����;kp0`�)�ŗ�" �hk�Jd8��2�zZ:e䦡V���Ȱ���0��+߲�<��S��w��P	��� Hem���/?������cY�Ŋ��o
Z����$t�,�,��YF\�m�I�A#�	�F�N��@?��*~�9ְ�Q�ӊ����K�:oi��]e�9��إ�zYFzK?~ժ��P��T����OO��+]ⷋ��F׵! n�rI�����M��M� �B�xjE��?������yp�uj7�blo�~��A�K2��	�̶�fW���cCS����L5�:����D��P�(E��c�:�y Ю�+ a�%>�M7�����>p��oi�ll쮭�#��$�		>���>��uK�Q�k�[�����/Q��7;e��l�V��D(WU�-
3��n��p�ĕ8�/ٿ��{���/6u�yU(�a�G��կ{X���?+��2�=�yT�;%�s�g�������Q�l�h���y��4�2&��u G���O{y����]y|�ͣ[�z`lx�8bi��SvV��ux8uY��#}曚������ͳ(;����ƿc����}yy�d�l�dS*+���n�����@�9��}�:Q�bu4���:���YC����`�(&�cWC��~u�A�����9��_<v��g�*קIV[�n%�򮑢_H�f��ߍ�u�R'2`z�k�M�}�LBU�
p�R���|� i^�(}��|�`θ�8m2�+2@nTF��2V�9%>��f�[u�a���Jm��?~0�'��@�鍩�E�{�_����{�H���-�x�d�ɩ�^��k�r�� �����q2�n�Q���NP�3Q���=���\������u-��
�n�g���O@PS�q\TA"lA����|(]��ӭh2k��Yt�	#G�󁙝�M�7�1y��Փ�w�Ybs��H@X]�8�7��Լ�[,��{6��U<ֻ�ݿ�Iq"�:}�$b��0H�k�;���G������};6�F��n^/���Y���ZY�r�S�wii�&/���ŅYT�)�0�rɓ.ZJ���F� 
(��.�߆�g+����f?�j����jɓ����6�͗�A�[t�
�u4ԿM6��Q�?:z�Ё�"p�0�:�Ѝ?��� O�"2�("Wb�~qd��˖���+D�ȧ;\�/N�8̭��1<�͍�]�-�x7c�z�<���%�L��
�:��$k$_���.Lx�$��| -��u�s�
KH��V������m��WdW����y��\Q��M&a���8J�M�l�E�;P���j['��;���O� R|}Gw�j���1���<ׂ�X�H�+�ǬhU`B�hT7��c7��χ���PH����:.����W���Ī�����869ۉTM��j�[Ȳu��<�V9��5��`�S�.[�n�-�������(@�F:���&=��¶K��tqpɢ3
��)��c����Vu�'�889e���r�>��
��� ���2"A`aQ�8Q�eD� f�k�c`|������e}�r����%�I�0:��A��&0�|�2J���zrk�^<{c���@�P�����
��I�i���[�Ӝ0E�]�x��7�*ol���H���:E4e��0�IG���+A9 ���o���b�����`ۀ;piN��P:/׀�
m���O�?�p.��R#���B��ľ��*�xW)�T E�4Ҫ.�	�]�Ks3%�B�x�M�װ�S��!5a�P�J���Q�p'T2 忬����;M>�'I�_����FSS���j��Ys�/v9 *��S<�?��	K�k�����;�Z��|�q���J:H\�#:��U��d@b� F��ʮ��T�U܂5*?~	͇�sB��;�P�tNq�]�N��n����Pͳ_���D"��`Fj�d� �ƅ�^NA��T <ew<[-^�T���ڹTB^��P�.b
? ?��q_���˃(1�j��S��r�:P�AA����`99��pn�T�[����_>��i7�_��7�ɮ�����[�����x?�`q���'����g͵�p��A|����T� Y�,]^���_����v��?n#�9hP�7y~�����i�Akc���|>
>�1��N��Z�Գ?�0�~:�\�?~���:�rr'�l���!`�s��voTq4��.~�;�npv�e���~���W`ң�C7�\&�2��l�k�_m����|;�R�� ��e���9E�S�P@����xx���Pß?#,�_��\�rܑ. ��A���^.�e8ޟ�yu�v�	���g�Q�lEm�4��o��BL�JN"����(��T7qW;��L��*.֔�/���+m)�(���ON�3����y�-�,�l�~D��* �UW��ҭx�2��ޛ�=�q7(~mT���ƏaC�Նjh����#����=�s���י.`��y�#Α�$�������}�!�v)B<��>Z 166��C&�3�Ō�ny��s���T�`xQ!�%��sO��Gǵ՞ѳ�A��[�]�@���9ܟ�����D�+q�a*�A�yM���%�l�/o,P;�rfJ���
�����B�Թ�u��a�� #X�]���6�-�g��QGy�|���c��J�Ұ�!��Yں�7gm��S�C{{~㨇#*QQ�������c������NDO�'����g�׬��C',�?�n@������^[��$�[��]�����"wi�rN����"j=��~�����nF��^�#w��e�S�Z�9]����}��Ҧܺx)�_6B���=Ju� ࢋ��q�]�B�r)w*�Y\�������5q��-.m���-w�cS�%����Z�x,į��^���LG����(
�s� �!�!d��j�h��&"#WYyӆ���B�v5��36w+�Ɇ��l�˔��K�|Q��6J@�(���/G#�;ǝ��)�e@2:�A����	rb0h�u|��=�WD�Fi����	��}hΤz����:�/q#��bJ�:df��U�t��	��Ŗi�٧LA]~!�2�W�f��}#��w*a���.��>E���L��(`f���.�	@�����V�Ւ��a����s@n����#�`��)-t��v�+yfff�9,5�F#�u�������߹߿.��vgee%�'�DC���´,�I2�8<ԓ�����vφ�5 .�G�Ã�r�s9Kܿv(�B�k��_�
�\>�6hAL���Vi�uǱfhQ�}V�i���P����Z|<��C�� u�H�F���MK��zz�b����]�ȒH�G����`��
],`w�p�r�H�x�ٷH
�{@���ׇ�4��}�|�<��d���\�P*_\��[渀]�w�ýϵ��{(,34u{����r�Ç�(u�ȥ�+X.hOf�cF�n
s��8#c�{������g�SR<��&���X<�`��nf���QۆK�Eѷ�uZA�҅A*�,Aio_	�RA*B�/����1�F���#e�s�%�+��m�
V	�Ԕ�uM����Y"A��x��0�31��5&�K�Ԫ�T��]_T�7�%(`_���5������$��JRZ:���M�S���������ͯLOߚ$U'�� 
�9	(����l���d�;	��~���vV�uJ���`B<;{&fu5����:s��\�O����C���l���E�/?^�+�Ʃ$v�VCok���Hrt�V�6�w \�q,t�Pv'-Y�_�}6�?��"��Kwɨ��8��g�	���аn����V}@�~�S�H� qy��p�kg��˃��`[�J��wyu�M��7�|�\^�r�u��P0��R��H��+�ϝ̥
wc#�k!{s���d��!���_�ږ>� ꥒ�jS�񃆴z�S��4�*���}�h�d�j�3g�J�$�����5?���z��K���.S�I�74A��j���_:��t�*U��g����n�����s0�G�l�����I��LD;��Y�x�M�����_���'�&�/Dr�.L�BL���i���ݒ�Ḧ8���IEI�Y�����[�7+$?��]���
'������m]s�|h�Ii�
@�, xcbx�ŀ}𠠸X�3M�����r������ /S�s��Z:�i(��ԡ�%�z��vz�h�@�n��s��	�rR�8A��@��ܢ�K��tt��#$�d�k*��˯��zBo�� K��'��������ᓱ�͏�>�Ք�?�pzfU�p�j��gF+�{N��5�s���+M�>�"�!|*��-�}���t���Q~�! �}��Ŷ��s��-�������x�����17�K\���ǌ���{c�9���1Tض����
 ����\�ڶ�v ���G��T�a�yaϪ��uɉ֤9ޅ�E7�.h�ŋ��Y�k�^��d�iEmUG-_�a�ܿ 8xi�6	��' r�xH7R@''eB�b� ��!��n�],��_�v	W�ԡE7�����=-�y�'�?DOׯ�x"�B2��V�,T�X�,��ӻƼL/�a�SҐK�y��ʷ�Mj �����	��d�rs�krz�)}��ٙ�Wg5��=^�W�U��
:��)����<M;�l���7���������Ҳ;��A�P��_Kl�?HU���s���`
"*��h�ZD�;�����B���o�y6LN�W0�>��4YZ1�EC�V������μ�T�.�[?���� ���ڠR5 �㮥���E�����^���>�r؍ ��>��ù��*�����v��q��:����RRj�s�1�|p��x����n���saooR;8@��.%`w�W�'�Z�,wҲ9��c���e:D.��m|}g}���Qg#�+!�n"?�q������U#ߍ��0���Sq5����?թ���v�yo�iUU��F�����Ֆ�,�rn��f{3�z\��,�<
�o�b畩'ں��� UlӒ���@~��Q�eo	A]TBr�A'*6UNf>���"m��HT��9xz���ei��~6�sH�Q��..䮮,`�Qm��]G�ބ��g)�e��U��x$Ze��<��"��ٖտ��:^sњ�Jg�_��8��:z�����>��{�z�����Z�-�c�4���+��y����	���,�LH�����ɿ��e���/?�I[��@�HgIҐq�*b%ž� ����nD�T`/���h��"W5�r�% %�NI�8�/��|l������H�x *�2[Iֆ���{3�~^�>����ȸ�#�SG�s�ŷ ,����ڒ�V�_����Z�X�p�7`'gB��TC�����l�������Vuvqc빀�[d3?�w뛚F�� Q6@������@�oj�st�$U�ht�����a�����7�@ܼ�_�8盤�Wיbm:���]i�R���R'��&"�0�gb���E�\BC~Q����H��@����g�����4�����;�����h^z�`tٝ.��+UU��c%Vu���=�>�V6�$� yn�t¶dw����/f��=%Q �����۹�o�zl՘���K(��{!�
���d����c���B���ݵ�;�nA=m,��T{%|3���/��P�j�~�Lv��݌G�}��r�1�x��P\�.��B�0T�L�'XF<�����N��p�j�p�=jѴN���'A�s��iu���n�^�I��r�[�����8�b��Z(0H��ބ��.x>��9j��Gk���E1�Z��بH��#�u��m�����A����.�bUd#1K]��b:���N�ͩ4�T?��=������FH�+ ��ۛ��{�|�Db��g�H!%<oG߭p����ݐ�������v9)M۬����}�^��eil��wVV��9���v�!hr*��,��'�3�8�0Q~��-�x��o����{�yM,�pm��K�J��N�7i-,Ĕ��=s瞧"���˖i���U ���f�S�,l�1��r�P�OF#�[(�GG��U����jsѐ��_<̿NK;շ�mc�p��1ć�bx��`��UFǂ_�'��[����0�����
�-=��_���tSZ	ݓ�ut��|yQ�����1Zn�ST?x,t�/�V?$_�``�8��Y���&�����Qq����
fhq���J��c��O��:~V��G���hR�tX��ة<ՑXċ*� 2B��!莅���! �/L��-,D�����*6��x�~!ۆ��&V�8���m0�F�D�'T�8�J#}>��f�@gX"�*-w���hhC��v��?<T7��Rb����w���J�֭� �bX���A�����b@��b*Wāg� �`)���PV�L������bz8c��۶A�����k�(OJ*5�8㩣7��/=X4�����V\����M��A��U��a� ���S�Ҫ�1��ٜ���_���s>J`x��� �Ȉ��Óv�C7�t����!X���.>/F�����%<����	��������I �� ʰp땄2��"'��ϟa�̔�m���9��B22qYYƏ���\���ڡ�K�eV�jA�<<����#���2;?~0y�=���o������ˍ�(`��a�,��$����D3��������=7���0�FH��R�g��,R�X��2��F�N\[�6�ilϥ���6p�Q(� ���\bR��g�G���8����N�J�_��{�>sf>�x��>�IT[9tt�>Y��Lm��S~�2W�>E˴�x<�$�Ѐ�H�_>�@���a�Cm��M���|6bnP1��_�F�qc��i�4������3���{�P�}	ٷ�$�dߍ5��dI�}��}��3B!��&��i��������������?Ǚ�o	s?��~^�{�{��F9�a�H���u2�n�zuȝ�����U��!r����{���O��/E�mks�7R18��+9fO��wփ�3G�}8�'v�Ν���V��r�ߤ��0-�2��*l�C��DO�������v������y��,��Q !{@�~.��g�yb:#l��~N�����м<��*sL���Je@g�7(#B�d�z�2���m)A����R��$.�P"45?�<i_IA�R� �
��~$"�\艡Ӟ�g���g�8�6b�F+��svv>n`�R(�����x~��fF~`�����6���J��M��55*d=��/�F�D^�����s���J�X���߶>�x������.�P��6.��2���Vю�Aq�#�F��t�����$~�e���,z^a���� �;4���`�̀��E��y3Q���+> ���4��NN&r�������P��.CZvq�ؠ���m��t�f�	W��FQtϸo��.ҭ6��ܙ�(l�.��0Ct	����4_G~�OYOD�)��AL�?(�&���C;}������㬷��ʚ}��{Rg���*��|����%XN莬��s����!~� ��Z��';l��7�5�9���5l��Jx��C�5F�):��J����?�\�����nDP�Y�3o7P$�e&63�HquG��
=���*U�(�.cx����k΢�a��_�$+G/��zR�d鬙�[�5``�M�\�ɕJ�W�����2Sd]�6�r���8b	�ե�8	8I�zJ&�zQX��Ǫ��t.@�Ӯ�\�y�W)V�4��������_V%�kl�R+z�w_Z[;�YM�[)j	N����O�l��q��������u��(t8\��ICE�址�?G��x	� ��l�C���Tc@̭e��}К�Tf$���q2'	ȣ�Ww���,"��2o�^��U3@AxiՇI���bH,�p�ͦ_�Y���N�S��G�����k/*[�P�va�a٨?~Yt�r���QHP��+^�	'�a񣄸e.q� ?����8Ջ|�*1��P����S�κ=�:w� ���h׮1�9?���CF1������0��+Ɛn�*+���M�(0���<���/��X�Kр�U���<��f֥?m��-��)&��� �hI�*or0��2C^4����M���q҅*W�|�!��ƫc��J�'*z)"L��$�dAZ��r�z�x�W�h�kKB{�-����,B8���ip���G� �dέ�v�@�cn^�q����ߍM��T�Ѥ��|��F�H[*�L��ϗ�Ӗ��wrm̅��nI1j��>��{�Ui����iu�<e	<
(����qޛ`�t�3�0"`V�֨�[*ՆH���ۼ����v���?oA���X��K���hdT��s:R�Y�m5��^���Q;�HP�&�e����&����(O�,:���I�����|l����Aލ^	�pF��+�-��|�7S\�hre��'����&>��=�b�a�o|���fl�)��#8�̭ˇ{��KK�7���x,��������c 9������#w�)����\/��0�M��o왛����;����L���S}ڝ bQk�8
�*�V��Sy���&�ه:�%���cs��N�"8�����@�WZ�aϔ=��q������rne��r_���mf��,���JW��٨d�
�����+���r��_�=�]W���p�_��H���E�m�O���͸w����i��͍���5;�Qndj�(�ļ�g���9?�u���d�y��W�B�������[&������H�P)KS�u|,(�E��n��ŝ��Tq#�(���T�Y�g��˖�J�~�Pv�+v���&�28Iڀ�����������1>Q2���I��lF�vg�e�g��/��C���& (]?A�bۯY��(����9<ޠ�V�B�}
�PA�H^c��M?�/�.�}z}ʨa����U�?G!�O��r|[�������J�����x��B0L�>ց��O7��~}Ɗ�=M������*����k�V��I¬eB��L
O�d�g��j����f�&fW�L�0��V��|Iq���]�C2�3<��щ�F���I�?z�_f��=U�����F��Gls?�{ʍ��|�:1�[_��|:��?�&K&���f��$�sa����ki���AU��l�}@̬ll��	!k>�..=���"o{z��x���eX}9�n4����ا��NK���b<^<?�y�!\�Il�|��5Qze�[Nɰ������F�V~��GG+���xI��ˋw��:�_i�7\U��M�d���2����3R��6��:����n��b�Q\���2����<3ޘ=�R=��,n�UO��9�~����% ���

]�G�G4�7$���1+|�ӝO����ϡ�n��?X^]MG�r�s�Tg��^eX��鍻���Dn2�_Xș���� EEDF0O9��vv.;4�>IF�B��wxb�L�� ��  �'����F)hg��,�.mX�z!��I�4N���_*ֻV���L�ĸ4��%�Y�����~�O��{-%>�d7qB �n�n����̔G����yw�rM��Q�H��*��ȝ�*�'Ԓ��{�N������';���߼����ki-|K7SX�9,-���5�qz�f���j��L����ןk|����,��#^��6UcA�U�{p��������8_�bI��x�q����Ĭ'{!E�:BO���h������X�;ifh�T�^P���r-@�`R�0@�����P� 
E��A�:*`W�f݈�����������q14L�~��K�v�mr�����@5k�A���k�L���U�?{��O�\��ӧO�i�:�7�^W�E``*��о��q0��7���5��G^�R4��]~���<M��=�v*���|�.�n$�p[����ёn©5�8�֭[��ƝD����<��<��YYY�r���c�P�uq9Ǟ�_�d R1N�H������CA]�цx����8��gN��/�S0!�OL��N�
֑��#O�����֠Ő�S����ư�z���Iɨk���k><y��/�$u+2g=Z��M\���߶�c���w��)�w%S�u*r�iK�/��]S�u��4���pټ�Qh<[k�l}�����8®;i��2M��~�4rdD��,	\�hN�ʰ
:����C pN`�hI��vt�C�	^W&��hGt]L�Ҽ�~��gda��0��x0����ٸ'Z�S}���^f����z����D�Ѥ���K)>�.(����㮆����
���T����م��c�i@��	d��[�7��~5l������)��-
�01k��'<�Ȉ�i�W�K�Ҋ���O
-Ԕ������XԒ'�n���O G���Rl�g $4,�O�@�_����_�*�#` Ύ�4�#W5���[[%�R���U��
*T�fv�%�_��/w����{��� >Ç1v#��Im7h�[�J���%ǯ����PV��]ҫ��[[[s��cO罂.���5�?1311�m� ��p�� @eKKO�����Z2�(A;�S�ƈ�Z�w��m[�v���NQuړ+�/u`�/�B*�k���8��㓗:��4�'�����-��!/ߤ��(M
����z�㔥�FX�o7�T3��@�_Ph�'s�%�!�om��Dc�@�C��ǫCv���a�{��`p��f-�CI))���M��Xz���p�v�rr�"�K�P7x�����p}/��5�����A|S�",��W�Kn�r5����)�r#��������`f7-q!`'i�LAwx a:k��o��C�i��L��l����z��S�pT_�����0>9��,n�߃V��2��S��3�=�f6by�M�o�ђ��MW��U�B���F����w&7L-,���
й��4{�w����t��YnKQ)q����ܦ��@}�ucB�-4�i�E�z�����CQ�^O�A)��	�ؼ��$5ogIiZ�~���J�*$$�t��U�cwwR����Ζ����ww��p�}����c���12q.�uΣUXT�Ġ]@F$����as�T�F�W�H�)��:	~2�B� �'��i\".�+���ٓ+�n{w#8�o���MO&$�*2�L�W���n>�!�[Vl${B[�<�U�|Z�5BQmH�DYg4���Y5���(�&ի�0}eѼ�m���C�rq�̀NP�%eȁ����In�\𰴱����b�r%zw\)w𽥯/##����իm��m--Q z7��P�FFʠ�������/-1 ����1� �A	��V��3�P}����� q_{�xf|\L�* �@6���ai�y�s@�}�3�W�3�$G�+�=�����9�	v�'>-2��eF�D^�.)?{b�K�R���~Y�U����JMtag'i�zkϲ� � 
I�"��� 	!(��d��N���̔���OL\�7�F/m�m�.}�O�I�FI��3���񀬜����PY��r��-���
iS3t���������������SV)��A�i߿ߖ���I"6�d�D-[9����Q��[�u7i,�������mb AP
ޑ�� A��5��/(p�����U��qe����/{����PFb1���s?á�3��逪?B3�ܚ�q���E�@΀a��� �dSK,ȭ�ͨA�YB�I���N�JI
0�~�.�q���4D����l�.��7��GC�5�构�zɏ.o=�>@����R�	~��s7���_�9�i ��Q�6�Wid�\����нw|R��:ghk�$0��@&=T^Mhj�$1s�f` � %Hv|��WfN�o�:��qc�8P��O*�\*��%<1�zh�-��K/((���摲������O
JJװ��l{���X�����P��M_6���o~V�H����B�9t��N tѹ��R��,^�z��Eo P E���׫�dA �ܞ�j�0��C�S�����q�ěb���2{�A ��L
���>uj��;L�l�n���?ܪ�����N@w%�h{�%l.֔�"���Qc:������TT\��X�U�	���m���<�e�fw%�I������JL�c (��M�@�ʿsA�=����婱�@����(���V�M---�zx����� %�Qkj�6��)����۶��U?��d��ٌ4�yAS7�ɑ◕7g�j��Ah��]����X_w������EՈu*l�%��efC<}�"�����:��w���Ia�DYY�/PlX�����/����*�檝澜\2���|���e._���Ù����@�\�Y*�TV�f��{-GLx��c�/f�_�ǵ�߉A�[[�X[D-�:������	ڧk�[�N.5[����屛�+w��x���[^��Z_ y`@��;6�"�9���P��X�i�����޹�^�Δ[:��ikO?�C�2������3a��U?�*�,�r���܆�Ā�M��ųC,J�T���л����}�����_�R��J�)�G]�N#�'q~��G\�<���ee�j�Q���@فcR*�y?1qh����4;��q���91��S!���Ԙ���j屷dd�US�y�/�d�;4&4�[��� ���=pۮ��d�x,p�X{����OBg'S����+#�������	,VA4��ZV�|��bMq5H6��D)VSKC|��,ѭ�4��u��'{��I��.�%L�֚<ƨCo=��E8�����gD�Jc+'�)�^�6���T�繆B�\(׮��ރW��ȃ�TF�LS��� +�T(�m��q���˓1 ���V1e5Y�x�)���Y�����,	�q�:͑��+)!��%}��<?ur�����Ⱦkn�A,A�7���keee4��������P�4\aec�9�ǣ_uYȎW@���P�ںW�}�����v_�v�$���1o[ZF0�z�Ӭ�GG� -�т�u�ϣ޾>I�X�Aw<���&gc��� ��(����?�(Y�Ir�l�ԟ H	���NQ��bQ�wɑ��٧�|�ɒz�p,7@<Cΐ|�w)�S5�TT�:����/�˃~�z��I9���À����A>WU]��6'&�+�3M>]=������ ,[Z�c���׳��>�
�W�.|�����	��|�DG� �
���nI�;H���Y�
ޱ� �k4����oq�D5������/��lF��7n����y��;�oT{�T�;:"��weUS��ۜ�g����յؤZ�Y�l?�����5D�Ԕ3�z�z44I�Z^�Q.����hdUu3O{���7t�	�Uڳӱ���q�����33����9����Ch�i��[eƜD9Q����V�E߼٢١j��J �m�v!�>�����?}X02S+Y�1���w�)(���=�1�����/.�WQQ���g�$�;h�������ttt 7z?}��A%�	i�c��\�ʾ^b$� $��n�}�10���b����Fbe�}��:�%*] 5@
_��d���oX'�'�~?G�b���֖���G�9����&&`OeN� ������L}�ߏ@�3_Dw��앍�N�´�C�`�>/���s&
'�(��+|�/��~�����>i�J	G�zhJg� @�Fi��ç}^�L�n[���:B�:��4��Όb�I11����z�£�r�vP?���������/z����˗���oyv"��e��H��-�����ݟ��8�U5���W������=E%�l�?xfׯ_oJ,	�FYY[�U30L�' ����ٹT
�Z��k�Yu��9IEwVY>}JVf/���%�ܛ�����Y�����4N66oJ�����nY`hN��'�t�z���<{"Q,�?�R���,�"�,���25͗���E�hej\%��z$���'�G9/5L��J���Z\g���$?/�|"�2�tc��Ia6&L�7B��n��}i����)iz�H!���$��o�K��_��/�p����8�:"�t'J�K-=�?�ɒ	D����{��/Ez��g��-7����9ڟ�f()��蟞fO��qE=N�<��GX;��MM��v���;u��
{�������T���]ts���ѭP��v��\�E�֭���a��l�&�{	ż���
+���&��{D�9�nf�y�k�s�en�,L�E��3�S���s�b��{Xl�,pY��Ҥs��.m��)!A�}�
p�غO\��h�;�M��Õ�� �;��+��Y��L 9��u@t˔P�����ם	�8� &$��>R��s|=|DB���R8���cMMMnVJ����
�����6��n�޽S5�ˉ>6<E��5А�Xd�����������7=�GX�ˎ�U��3�*��²�.�|���
)�;E%$�m<>՗�tuI����G�(�0�b[*�x��,��8ċQ��T�$e��fg�H�p�^�a��a+�74��PIR���2e������g��
Nj�K.	�*֠�t�N����1^�)/ϝ&�h� ���ŻȒ���+��󶈳v�ۊ�r��y��˗z?��Xs4/���Ϸ6\������-�mv����ۤ�laЀ;�\.�п�'^V�TXR2Fg�%A���������,�O�;�
=ۧ�G�w~}TЙ�W�qw,����#B�[8�M��8汱1�ZO.��K�����|����Ǟ��E�@a11���vO�&��Ǳ�����p8��A"SCm���	�H�*�~�S�)�@���ރ��f����D���+N����q���w�`��U�w�N~��f���gY�Wp��>B�B?锉��Gwg��̠�S^��<)��~�hӉ��09H�_�6��uv�N)�����<�<��k2�٨���K�A)dN�k'Y�� u�`oY�����x�_��l��1�H]������Q������|�DP֭��������e�iS�n��574$��<��jo�����e�Y1sXz�W�	S�Mm$5�T4�BЬ��RH7pV;S=6���'{p=��q��(���b�C�u�D�g'��I�Ɨ�i���?����^�K���<�0� �c�u:��& '��T�4��i�����EyʏV�I��<��
��v&y���/mA��w��}� �QH�ڻ�-�'��S�~���\J��}��	�̈�ժ�"�AG �k�K�q����4y��[=}��8��]���(�}m�����]�ٍF�����x����A���_º��$��RЌ��`h�D���� ��O�pI����$^�*��R[x1�7z5=2V��v�O�f��<�8D��������K�dsц'��4��>�u��[�w����쪪{~���J������V�r�!��v*��Q0�P��7�F-�O�%V��L�����~/H6fXի�śW�
&66hrds��ʇ���QP��67'BW�9t��̸�O���V�3��N�4�56�WU��cJ
���o��I���ww�+�	v	
",)�n�ޘ����&��� x��)��?�K����ۺ�ip^������������ʺ'm58�[�]6��k��P.�!`]b���D�z'��b^6��,o Q���A	N�$127�s�Ӣst���F��'=~Z�aX=^�n�/�����[-k�������D�\i�\!��:���&%kS�����&ʲE���R��3�p_��&7�F�������?�:͕�2zvv.�V ��UnII�V�Z�:\~��N���"9)������a�/,���	���{������ҫ�kl4��J������lp#U�$͘��mr�C�лP��A>���6���"�cx��Z�OkclH��{�\�deto��`}kկ-h�C]7���9yvu5=c���=3*`ht�{��� <���QB١1�Hp���'�<7�j�NT�{���M�a��Lh"x7P<<�3���в�X`�"�6�S����U�WQ9#�5�c��8)�aHD�v��3}@�1��
�e�J��ױ�#>��!׳��f-�g�h L��XW�_�s�β��ols����̱�v��q߷o	k;a�/0�hy®k�.G:j\\��o\��>�1$b��uo����3gPU�l��?DyvPv�}o�%S��ۮC�yW�4��Yݛ�ݘ��ȝ��X�����i([|��|�d��e��@,(I�߻�']���/EK�$���� �_0f�Lɔ󵇎8����e��-I�<�m8�"�J����L�ͮEG.z�wWwL�
!�_����ʘ�}����i����_$�HS�
	).����xK7������ʼ��yt8F�7���S&�ir�v���7  ��i0���z��B���W�R��)P��r��'t�̅�x?� ��-�w�V���8�����!V��3r�r�k�@
�'.��0��b���0���DDl��1k>��2e8f�+8Q�Z�w���n� f&��߅�M�(=���(��$"��b���IS֎_T�~Y)`!�UK����O����}�f�Ď���b�2Q��p�	��a��k�ݶ�A�u�OwyL@2���EQ�4��>@?��|�ዏWOJ1��%�ݘ����C8�fi �<���_I,O���Ɉ�?�
���3��|�+�ZΆ�����W�>)����
=^���0<�NT/��k/��9B�΍:��o�C�¨���@���!�Q�Pj]�,����D`0?���2�弲�ȝ\q���q�����@
�lT2@8w��]����ZtWJ�h<HK�⥞POE `$���^�ٴ�NL@�6����F)�֜��8���67�'Ǭ�VJ��[�Db�ЌR�|�<�����ӹ�,����7��F[#z��;���I<����`�������N
���kjn��z"�AM<(2H��9 յ�f�~㓋�e���wZtg�/�ҫ6ܜO��s��[���?��O�VA�I5��B:��򼴽ssz��d�M��8yt����G�#:��b�/��???���V��k�|��;��no��P`J�=uu��n��"dɣ���X���}�+��X�O6�+U_�}�����$$*ob�	sMq����k3B"��1���]��PW�Z�re��h�F�_ �.�C�`����f��?>����+��������)0��w�=g�.|6%a-��m0�v62	���!dʺ�8�Ā�9�zZ�/��*�ck�d2��҅�?|�J�+b�t�ɥ)L~1]�&����V^^�S��_�6KUz�����_/�	�s��l������u>��7:�9�Q�a:��⩁^>h�ԇ�^�d𗾷�"�o{[����/�m�/(���Z i$��݈�g`�a�ꪣ��J`��ǋ/8��YՕ����6�6�P�>��ݧd�Y��i����ĉ�@Uox��5�sz@���Eb(�3(��N�e:��k�5�}|������� w�D�)K��gd��Y�Xc�����NO
��K��|��ȸ-�=z����c	����-�T�f�w,VY({��6bD\��u��֏����%z�ּ4��ڵb����������<�`z`趯��w&�	 x�!���z�py@��Y�9�T4�wz�2�t�ui��\,nG��E��⫍�~G��~���j�)5�̳S�̄��ϸ����f�߂gO���1R�O�b?��'B�䪁�i^�{{A-�+M�%3dӀ�I���=x���}��xeۭ_����a��_�7��$��cd\�$�r�LCe����@\�\sH��e���ݶ���;q�܃t��5�4G�"���P�jC((`�t��^gN����n���T�A��ȟ�m��ίc��y�ɍ�#d���ji��w����=!o;:"�x�3Po[[�u��J�S�@�n���?=��w��I2v�ı�zF�;�0a'Х'����JJ3u�=��M��>��@Մn�d�P6��v�&mƶ��?�����˹[��>E�IV��_l��]�?��o�M5���hB!%����Gy�j�.�[��s�MN�8"�~��;�n��G�>�!�I-nτnu>�ݵ<�� ���|i�]��~G{�}}}�;- ���n�,]-	�۽u�(�:9�	�ek2��e�=�p�v����#`GF����O0�kB�P�ݙӫ�9�;����B,ڧ���+[�k�K_K�T�¯B�Y�0���M�c,ޛ���ZA1k����Tv��#��~��aPe�r�0�u�_ۛz;����5o���}����& �k�����Ǉm?�΍���i1�1WU�=PĖ�RP4�m ׍B/E��N���d�zU) �6�7��J	�O��z��~,$���ݗ�&��r�O��C0w�-�N�~��аKA��ݛ;���=O���s](�l&x�vk-22���S�o!tqf˻f���� �.��Q$��uu68��$��"Z�I8�H�}"�M k7�n�8 �Ȍ����	�A7y?|�4՝�d�H�ts�c���M?a)�T���� ����]0�?�N���C ��D��C#s��h�z��9�����S�q\4z)DN�<������ez�q]�l]�i �*���__$NJI���V�MaB4����ؘ?8�L�x]r����ɚJ��1��Z�gI]c_�8���v�{Fed�R�"���Ԍ�2QW�3f���8�����а�yrF�|����I����yYHy�y�A��+��;�Nn���}q�ps��&	������7J����L�~<�/r�b��U�Qss�Ǯ�T��S҈��:w鐣_�b;"Z�<1Ֆ�+I����J	}�_B�onK�l`މ��H�����ye�*%�>y��h�O�'K�'��]<���iexj>'hvY�n�h�<u�'@дw��K�0^CC��~����>�S�?�/WUU�w��-��{�N��,�� �T�����Љ�����/���d� F�2.�}�qnƞ�܁"�u6��a[ޯszS�d����:����`�x7��z�0
����^Ͳ�9�����@��v#�\HD|�@��vs{;� �	�kqqqv' �&_dd��;��Ufi����n0O��[܏�>~�ذ����d��.M�0J��o2O��d�*����_5J5�[̢�Ǫ� �+M���ݻ�U�u���J��&�>�Xizv��g;vJ�3�8nݪ�b�($D��J�yZG{�T�8�z�y�-��?��QLw�.A�쪲�%�0����4�\�9*U;��b
���"��B�њ�b�A�q��^��Z�G_74��$�jKL��R�71��M
8��B�� ��Y�M��������F=���괅��1��i�dj�뺻S�D�Km��Z�Q�\Q��đ\đ
�Z����\�}�3�`R]|���>�Y���h:v-������F<b�R�n��}���gX6
�~����;HA-|���Tm�?c�qh�R��
������W^������E@�I]Y�˛g��9���UU���_�ih�T+��uT�Z����O��,,��i�A�=d���Ƃ��o��{��j��� yz�}����D�"Wc |0��
��������������w8��������3+/�F�.Բ��zS��s���#J��%#Cf��"����Wm*��y�v���3A�.ǹ8�5���貆�)�X��ܱɰ�rۿ�|HT�Q�M����
��������!���MX�k, ^y�M�/�L�����`l�\����v�E��.{Ab�k>_��/���0����%>�Bݤ��uv������"/�
 �FԀ:y�#G��v'A���"����s?�}���Q��*Wc��u�YN�WK���R����xQQa���d2�ځl&�T&��P�<�k�{9��򧒅#�|���k���Pκ�2L}`p��0��B= (�P����Z������M����*9��-�ƵQ�
>�k����MQf�ܱ����u��d��'i����iw�`��J���b3W����iAa��.cy#�UJ��5�^��P���x�˴�H [��KXBDE�ތ�<�J�$d�ݧKmFj�N e����,�A�('�������_)�<	��!U���w����~nKe$�����Yc X�h%���7iO�U�E�%��-W|��r�.���#�`I�#y����g~�{{Cg��ꥱ)P�}�.B�c׀whh*Ѣ��z�)%��?r�0�ڲ#�'*@����)����0�
��p��E�p�ף�����ax�(��P�1�NA�aU��)̸o�����׺��h}|}[^�:w�����d��[��2�M�:#/�+Sѳ�4�d��=׸���:ć�C�5$����gO�&>R�]E���e=���[��f���8x�a����P�3
=�E��G�ȑ-S�5��hR�7��ӝAQ䫟H"�M�I��7��\�G��z�nPQ�ç�d�i&z�mc/�3>&rK�ӲE����y��X>����)ӄts���D��u�sH�߯-������v�8� �:W���W�.��j�ta�K�oe���0 �  o)'1Y�fFV5_�s�?�y����og5�u������!!=M.���9H���'���l�eݎ��<k���U�3�	3��\�����w�$B�Te��c9N��~|Zsi:!0p����9)����N��x{��2�ǫ�����_��d��! � )B���@���/������3�Q�V�m��q�!a��5QkiM8 3�\_��ˁ���"�LM#x�c��==3���.&��|���(|����]g��r�9�]��Z7�
�S���/�6a�N�Τ��LO���1r��.�\�%�z��L��fl ��wl,F��5]�>3x�M��rWUM
�%y��Sg�W�����d�O��:���	c���E@q�T�in���K��&�~��?~��k (�Om%��sˊ'�^b��u�	��{	,��?IvL�G+���pn�������a:V�����K�<��5��.�X1����Kj�s��]���󚚙�f�+^? #C;ό������?�z���L�����J���2���͒����E~v<*Q) !�	�#�h����utX=�֟p��iuˡ5@ii�G�>>	H$�EZ��Ť�Ěm4K㪓ӛM�5�m��ý=q��}�l����T�������o��v�Bv:��Na�P�:�xŴ�[u�;���3W�EP�_����pJ��~�9��X�Fw"��藍a�Ǭ���&�Ĥ�����%�?'�Tֶ�ce��I��^ON��{�av{[�����'���5�Ӯ�ڒz���	$��h=��M͍p����������2����ne��]�vr�ů�Z�v�~�,��w?����q�*'D�K`�mm�̸�si�YL[��ͽJ���̻#<BN����`	�
?Wpf��D��|P~��N�a"��-��n�V@'��5��[7!��ϳڝ������4���J{f@� �ـ.D���j�&g��n����&VU��,�F�g��ݴ����0.�r�xH"\rm��[m�d�y�a�G�����C-��q���ݑ��7���YXx�.{X�źZ|X�wq��E�#_�n������/�_G�����U�ۀ�~`�(��.��蜎���1Κ��4���x*�T�:]Ġ6������<�,k�kq���$��P�l	q��OB�e�|JnFh儓��k���4{���VJv||\��mk�3@����WV�A�?ceZZ��m�ԎCk���B���W�]O=@Y���t�1>)��uHt�R�_b,z�.�L�C|�r)�����9����gɄz*���8y�x�W;V�P/G@X8y�~��c��rJ�<?������2��n7���d;c�2)�H����@|.�W	��#��\�۾�t�4�D�:ĕ���;m��}�a�b܏�Ird�%SQȘ�1r��(8���Iw)0!�P\�9���e궡�5*��9''#ּi._u��z�y��P6�~HDY��\Dv��3s�_�Y]M�4M��
;�?�P�V���M	F�]�*��g�խ^��1׶��5A�������8Ug���I�ŷM5浳;8�b�|5I��~�?��Sp;�c��_���^j��K�F�Ts<�6|�܌Zd�v^����o��3���:�n�e� ���HЋ��"I_ 9'g"%k`�{p \|.��r�Z:�g8�Vˈ���ρ4�=�Z�Q�/$>>9�b��v�]�	N�02�	H��������,g!�1�� ��\�%�i �T�ù���^M��SS#Ħ��#��\���-9��A�2��5ZM#�cE���/����� �Kb�8�69ф��+�nL���GF٨d�? �*ȇ�XC�|ӏ01�GJ������I����b�<3	Pf�����|�--�ͺ}l����N�-��G��VU�
������F��+&��ԙr뙶����s�*
���3q��Pc,;�NcQ����㖧�5�Hd����M-��k�����Tb�kMo����i�	�i)s=Z��:�]W�ެ�e�C#����k��Ϲ9B������+"��E�Tо7�y規U�ZFOO��A^U��:Uu���(��<N���MR��`����_��¬��?!_�~�lV���n�����1�����؅�X�s����L�?���+�7E��O����?�GN��7g5�X%BSq#Z�����p�o��Hn琋$F���|B�;
i��2��qNG��:x���!v�.�ʤJJ׀.��Q<%ԛ��E�x|�|��N�H�%��Ӧ���%EH��T���Ta11 S�7�Ą�n�X>}z�ڰ�����+���>�3N�uMM��ޜ�Ԧ��(o����l����-�}6�a��';����j	P1Z[[�e��70�b�f3g��v��:9҈Ny����?I2]1@�X����L�?���������9K]�gH��Ot����Ψ!@Fn�x"���A?M�����q�f���'Ͻ��|lcC��x�/�������m����)�ay�Ӄ��6��H��/+ �֫�R�IV!rt�m�"�F�
~Se�	���.Tڽ� yI��om�/8�zn�]E��C�����(o*��;k�9;���@>��G8)��hh��w��[V�]�����Q��HUV"�k��`�U�O������iNU"yZ��Q�Dpr���CVIf>;0h5U�V�~g�i��K�K\�}�[3��]����m��i�-c��Eؓ�LQF��f��oQ;����AJ��Aj�|�߿�xN������"ŉ1)�m4(�[Ԓ3��Cx��8H�����
'q��g-�	���OAV��Ul�pE�ab�5�K�,[�48%���و���H==�N$@!S�,\�M	?�~>^?��n�Euiv��?g`@w��~/:�8�+uU��d�V�4��D>u�	�o^F�LM5�7A!!l�X�~��ۮ��Gk����s���# ��P��bY4�����Smp��g��4yU��]Oy*������(f]�{m5����ed����2-����u�z6*N�:�.��t��p^3�Q�n�^�3����.7VS[��{@vS!�45��W��}��,��)����o7 �9�z	��,,ϖ#�����[ҡ]Q��U��_��f��b\@6���*�F&���⒓���Y�#8��H|�}����������˰��/�zQg�'� �b±�ҕ񂢢P��[�ǌ@�f��w�7'ɇ��~�6x,�T�F�&���n�z��<��	 �+f=��5H}7O���y�R���Yuq���ܖ�ְ[pp�Cc���8K*�'ɩ\�/-��tY�q������7Ƈ�>h��s1�ӈ�l"�(H��R|��{�󳡶k�)�3ѕ��-���_i�bƁu	6�o����Ʈ�o�VlUlnݹݰ�������������T7�$}�KS.�;�q����S`4�˒�C-�ZZ[�zzdѺ�OM���g��3�D/y���������@:`��]�޵�����|�������M�?D���x�>|$�;��r(�������M��7���B��	�Ma��Б�����5I���ֻ�l�-E��[�t�-����Io �G+���?���KM���0����r�bx���Ðh���8�OK���JԿ:������^��D��ΑDx=��%�$� ?9��W�E^^���H��,�U�D\]��I���XZL���l���P����<x��EQ���8���v$�5���c˞��G{�D	�Bs�̌��$��t���Cg-:�'�����$�w�������1��(�@<$,��S�4:�H��O��'v�V�=sB/��p���,�p��L� N��#k>@E�h��j���sH޳�wN��D+�R��	A@P�.���Bж�5���?�a���r�hZZ[�a��mTU�荥��3��V���&q���sgr��~��7��\�K�X#33�cV�E{��]c��U�*�b͚�O._:t���@��������}��f��2{h�ÿ���Xk|��<��z�t�ʁ)O�s��EV6*n��<A����W7O�AQ�-�����gc�܌U.�@������/�"t��"�|M�Hq���	t�����;�����U���{%$I�$3\3#��M���2CٲB!d%d�nH>�n�^)ܐ������;���sΧ�_���1������Q���5�!�ӿDI�k��(�<�u�l%{dR�@�k wv��e�,�y�|�Gmln�9K��#���ё?�9��V�G�.J$�;#�����N �U��	 50�x�93oؿ�Y^S��1����O�9������ݜG�P�z�V�CxK����%؞�-����Ѿ�cI��II���'��� �8}t�r��Aj
����p �g�cZ�A�J���봵�',�%"ۏ2���4:6��4�?h�w���!���U��+��:�*|��o�d�~z�|wbU �};$9�t6n��������O�Ngo��N�����E��M�������&�r��d4Wrӯ;)���n	�R�Q(m�;��ڴ�K{�a瑱<�g~�*+,�>!�u�.|���0�b�`��B��C�m�dzd�`j�<��9�om��w3;�xbbW��]f��T����g�i�J|��)�B�L�@��1���8�'ov�l nq�4�g/85�B��Me_�R?�9.���7�i�fp�Ε}���<�mNW���-2�Q?1��n�)��������w�y�� ]m^^^R3�\��H���0���>��`�}u%���ekP�!�R�Ӗx���|��o�$l?a�� ���m"{?
�ݤ.7`���+W�"/�XqՇr
t@�qS�n���,�7z��2�5���*�3�  M���u�G�z=$��g��vg�Hv���c�a� ��O�<���T"22!����ܾ[( �0��g���֯���D.[��ȷ�W��buea ���a.bktG8��ݽ�A�
�@���1jd��6MmJ��{����hpe���dʒN�C���Ы�b�F:ѫዪ9fyvF�Ȭi�ɷ�	 ��֭���Ȝ�)�??�<������uq�u�����m?�^�����G�W$��~�=�v�UM�*�#--e��v�����~�_,Sc����,K{]�E��nD7
u]����;�I2v��%�eNO����� &x|\8�P�vv����I,rqwl���E*?9�6Y�� 0TS��Ҹ<�&S��I�Ɠ 0r�sH�gyJfv���,�e#����;&��X��eȠ7��agdp~�r,1$,�Z�W�߀!��WU�kϬ��:�I�Sn�؂�4����ME�$��Z�|dZ��rK�~wãQ ��$�yZ��������\TX2�.�X�:/���I �8ھ��G��W&�N�:/.5+���v�oo�H�\zK�^J�y��h~B�ϟ?5q�{��dh���K�o���������aQn!U�4B+���_=�+��U=����9����EHkF�*�ٞr��\��KO��1���_ݏ>�SnS �v��\�0J�R��"E*�o?H**x��������?�E5��S��!�M~�#�$;3���g�����L�6� �������ָ�g�8�ƆG'�?��0̦��k�F�7:��i̡OCBdt����U�SX�����N=9
KWu���P�e��m��P΍��%�w��׌����:�~K�LI����g������x��y&Ck�yt�}�0ir��Se�׺��Uޫ�	b,��w�1{�����nJ��k8��J�}�k�gC�5�﫾S��k����H��p�W�[�(�F�������~�� U���!��۪��J�Փ���x�v�c��s�l������Lul�g ���N֌`+ߌ,�;;w��D=ԽLɕ������j#ɦJ���_���m{%,��޺��8�	|b�j�9��^F�l0b����|�y0��H�V"�-]�N=t�t<�� �^�-]�P��T��,Sߥ�kM���F�ǯQ����=�Γ���D�mZ�R�L�z�J�RZ
��/LDq����}*�ぶh�������9���N��m���/@�T�We����"/������@N(����Ҳ���>��l��y��X=���tɓ�x� �'�))���8� �{�G��4��q���l[�A��)y��̾��A�ZW>�XH���EA�$/���R-��X툚�1�����l��l� ������s�f�0�L2��� "�K�4_G�P�;:׌ � ���T�{z/�����n��_��֮=��i5>`5_�{q���g١�Hp���ל�V�76{�����ɞ$yf^9ՌT*�<k)�ci����ǓZ�9M,���^/9���x7�@`C�fc� )ҙmiiɜ�>f�c�e9Q���؂��/	�gh"�����D5�qZ�&7O�q_Oxl-aS��k���f ����oO/��{s���$����� �<�T��mdnęH����BNv	�
�?�����}�j�N�404l�ￒ<��v߼{�	,��R��*��;���1Tw��B��W5��O����c��,�o��u)n�z�:s�F��^�{cN�ڄ�����u�@�F� �2s�K�LW��d���*�9;XI. �*�1��/�W� �m-�<n��%4���H[˦)^5�r�w�ܚ�����(�fg?�M���!N�1�/���v �>���B^����d}&߽�$������6ֲ�u��:5G��� �n�%e\�+�"P�y��vوt��/\-��*�0�6��Izzy}�wwD4�R�%:��RRR�<}A�F��L�g'�y�c��4��Ȝ-�P��q�<>h�
w^�y�_�;_��]Mu�`�����uk�YRz�4�\V�"�������S!�W�2{T��ru:{zȁƎ�Oĸ��wς P�����_���G֢�����'��gs��Ą���	������y>�Oy�>�lV9�aLxc�SG��u��mEE��~�����(t����#c�|7�{��	� �JC�#�����}ԉn�/�JA��DN�����JI4�W(����c��A�OO����ڱ�L�)�'
�ؔ�g�`���jӧ�T5��x,�PW�aLŲXǊ�m4]��uD�9� p��[�٦������Y�l�ҿ�* 4�A^A�:.51m\���T��O�)�V��YZz���z�-�Nك�}���[4X,6��LJj��S�����扷��6;w���83�I)�Ǔ Z�[Qt.rGc9F �輦�HA�J��n���B���/"d��+!JR5����ࠟEȜ�e���)�ˋ������H����#5�m��LL:eY΄�A�zIf��&��2~���������k��*S����CBv�����6�o���A�N���N$ob�Ջ�����������j�'�����s���<d��X��s7���S0�E_2L��^�}��GF����w���u��^�xWT8Hh�L�+�ã�����F�~��D�r\�o�6�t�b�D��٢'�����w+(��|�^�G��~�X$��a{|�G��*ێ�ﶴ[���p�<W�2�D8zE���� ]�a���婀�`��b�>
���*�V�Y\������\�o�r�����x��w����NMq{=g}���#%>ʧGBAAQ{#�V���s�t���ŋ_7L��i;W0��?{n��|䴜(�������2]{{/c�x�*��s���C�/Gy�A����%�Jj��3f�ra�ü3�Cn���V�sTT�Ѩ���4K#�q����l�P��e�e���1��s�F���U��9F��ϻ�xn�\��|@-$�vB5~����}x C�a����b�,,��e��m�KR�(�*���646~X\�!�m�c�䔽l�5gZjc�㫏}�r߻Շ����y��x�O�"�Q��H�'�]�ep�x`�k
9��������������U���y<�4��Ī�1��Ҧ�,�I7&�J ���}+��s�ė���Ռ��4�[�� �v�[���d��9i�̹&ɋ�|��TȻ�s�K���b���R*X���265%��?Kw��ʊ6G m����o烠kD����y7��y�#R�is�o`v�ɼ?�a�a��a�<�I|��L����8��r��)@f �j�'4�%���+�����o@?D5#ǲz�Roƕ.JI�ț̬x������<S�`��D�w���5.�9�z9ǜ.�l���r�8RIpf�B�������������N�����	�~��͸��ѿ��UUc�>_c+�ȴ���;�-
5}���EϷ�4o�WWF��>���<�H�[���uO�I��n8К��h��SBʿh��o�9�v�5h��?>M��/���?�\<�p���/�k���m����d}5C������k�^s!F�$����0+�T�'�}.]�|�E�~q�g�̟���h:�@ٰ�*���5_�(cQ�f���d!Q��8MM+����C��^��E�q��&���5fw�\n	һz{�*�Y9yx�]k}�������zڅ��ׁ�Y�����+%��9q���A:g��e���e��Z�W�a��b隠��E�W~�YK"=A�_� �s)���e���nRbG �[8��)4�]�9 �x׏��F�TR�ޓ�^��QCJ��T_$/��6²			�{x�#m�d�\Q���������U���/�C���]H;�ݩ�##S��*��-�B��>8_߆�=��66���ؼ�j�yyr�K=��ov���9^��9Q��=�_��i����ν)�Du*U��"� CT�U�2E��J(���E��2�ْ9���=�-s�N��b{j��i��H�B�
nn����+f�sK����4װ����#�����-�QQ�߽���e[�ջ���S�k.�����T�enl�tv��Q�� ��:��-��8`~���͜�������y7�������%���A��6��*�=+e�W�0�6�Ry���e��>�>=�8����0��kb���[�QiЖ�Z��6*EF���}����C���PG�;nnoj�&=
V=S.��1�z�Ї��{�ccn��Ky�"��eqӝ��?c���� ��=�8�B�[���i�zԽ�݌vـ�G8\����g/��H��殦�Ȣ�x�.G)��˽��֚���yԁVA�r��el�6K@M]�DĮ��[�8�u���9�Z�����]M�]�2fBY	���Kӕ��nm�9�ėX}�}�:��af3���U���8�2���j�VH;D�zg�1$�I���A���ʥ�OF/��ܢQҡ�@#����i��(�4�M�9^�4H/��Q7[�X]$�!U�n��gLĢ$n��ܹ&ԝ� ��t�jgz�[��ϟ�yIxU�\w���my���^ǶࠐPwnR��[O���_��PPs�̝s��������9�i1"%1g ��P��m*8�#�a���gyKԇ?�:^��;Ҳ�(�i-�(�pK��z�� ��Ksi̓���C�F>aR�����|�P+�O|ӯ��1 y.����j4�hT*.���{B�# $�><��C7;��~�B6��=<2H$wN�>��#�?���J��5:4��G�E
��C��E�� ��I�����4�R)))EI�{��d����\$D�h���������=��=�ǫ��x|sBj1%��ZhmP�"L�G�)��N��./<$��]{��t��C֡T_�>�B���K��Zt��������YH���:�"=犟5�Nh�Z(�����@�{{G�oߦ�@s�Qf���r	��9�
h�z5C����3 )e󍅭��(���σ����c��4�5���k;��X,�V�M�>EH��m��͹n�&D�����G���q��7�ϥP@��AyO��H�h�9֌l-5�)ր`��}���7�;8��2u��RV٩��KbL�=�)!-=9q�\�����p�~�4����e�|(M�k� �e�\,1�>>���Q,����$3B-��}TY��_\��A���ҕ+�[��-w�غ���H k����6J�4����7#*#ceGM�_o_��kv�Q��5NR�R��=�\��a!UK v�����Q6���� S.����{�I�	;qV�*�����*OD7�SB٣�A�M��M�����V��#��7��s�\�_��p�^5d��X�\�Ƹ66$�)���Q��h���ZB�z���z$���A���QFbSW[��d��IͻZ��ݵ5aaaP8�G��_���S���$�����[?9&B�>�o��=����<==���Qዽ�e�]{�t����������:t��L�u�q���#:�����1'��G��>�}�B�j�n�	��� �=�3R����a ������υ�U�n͹K:��d�y6|�u�h-J��R���xb�sm�,��KW|��%�}�*0p�Y��e����@�r��0J����c��}�s�gg���~/�olz���
{�T1t�E�[+g���C_��L�v�V����w/+�˥�h_��������4J��5��*��������w�ZB�<f��;���X��!mTH�>�^�k.���(��������7�7-w�@5��ǿ���#>Rn@���@�H(gB&��"OV��4@�ic������.;i~AW��º$f�>���A.߾�b�����Z�k����NH�G/�H֌�,.���ArK��ؘ|e����> Q�f���>s�o�(j�C�TyW��s�Ld�:a1�S6���R z��￮m�������^H5�%��B����
z���c-��-'�r7;��G�o�Uv��	7�����*�ں:7�lĿᗝ�*l/�-���)�᝴ް	��˷�2��>�zP�|�� �l�	@y�X��}�Gi��KK���"TU��!m�ޥ�p��4ܡ��m�d�{�Id�����Ş1-�!R��~����$9�}-|�:@���a��c�aM!�s�^*]�Wn��Z�R)�����#@O�L��a)�Ť�qx�_�,Ss�Q�zʅx~��`F�؛�n��=U�?���<��E����o�\����y&��Ũ*�
?.���N���������+Fy*���c�y/�Ȧ��Yq�[[�E��Ѫ�÷����U�I��u��P� ����s����ES�����9U�'�M:��.����٤4�zђ��u[+��G��v��� ���fz�Z ���T��@yK_Ň�4YQ�F���]Z�=Bf���~-��op}x�<ћ)SӘ�rp�A$~��x"T?|��43cFP�W)���X��da���7er33��"dܾ[~�ڽ`�>-����f?R6����L�ES?���ݾP�c�oO�����c�㬻$R�5��ܳ!&$DF�;���B���泞��mmr|��bY�AWFK�*(f
�>��=�ҟ��.,��i�Z��)�A<�\�$�$�+A��~�G�(�DA�4�:�J"��k';�@�0��R��TFF7���$���]�"<GW=��;���2�F%^k�M�̻�#|s�<2�$���oi
y*���'��h�H��yb`4C6����b�H�Nii��@n��ܿfQ���}x�A��F��{Ș���T�}�3'KJJ��~! �M�����]<7�B!ޫh"x�� 
aD\\]����r:�y�������<T��=�n���	�S=�Κ�G&��p9��U�u�#���7�brk�*U�#�%���~���X�������X�[�5���|�ds��n��p���t�xr�?,zZ�۳tYۛ'^�ʠ�:/elf�;�D��R�Xy��aN�&&ӿӦ�r�=c|�gq֍��W��'�z�
�o`��D�x���(��GB��J���8��oR�OI��!�82�2��!�k7<����9ɩ'�	]����Ty��z@}�$}^s��k�y��컦��W9��7 ֢v��=  ��[��J:ߩ4�EɎ�(��ۄ ��]	Cs�R*R�Nf5���0����sp�Ё� +{�-�Ħ:s�θchHVe t[�%�[��}J?}DL� 	Fy�-F��4�$RL-��>*�ы��1q���jtRAq#@����ne	���z�,�Y�BiJU�C���p�����1�v�� ����O�Ɛ��~v�f�L���eh������y����s6�ڟ*3�`h﷥Sg��t=U"�*f�.X|���oF5��h��=+1n�s��*_bx�L�C��"�$�Cx�\�b$8i",�	"sd��l''�9c��ûl�!N\��~Gq������8IZ��~�=�m���%�Ɏ�v��=�VW���W��vV��lXqqw�X��W��>|�G19Y(�]J��ec�r"��KH�W��b�P4{��y�Ч��Q.��T��3
E�,i=��'�� � k�E�(�򬌅�<��lA�*º����)�����Q^��Ł�f��e]YFrĞ�|�)��n�43����#3�����uY���%�Y�
&''��peh�L��F�r��ǐ�Ώ���,.CD\".)s��4�3�U�xe������3��	���'!wh-��Z�+�e�h�.�$�\
�@�īv�&��)axg�4��T����O���q}��q�g{/������3e��>��^;;�tE�̛7®�'C-��1ǋ�$�b/æK�v�hѓH��<� ��:�$s�*E�������'��^F�?�a��:l�ӊ���v��z�#�s��q��R�����ݷ�Rl2�����{�	kB��Pc+�|�T�0DɃ�^	Vlo�������b����7��P�'����k�E;�O��{r�o��4G�Z^PS�ݩ�w��o��:O��5Uoj.544�\���I��l���n��HV?��ə3���"�CG�!"&6v{5��^��M)ᶏ�:h	6y�T�C��͆��B��~{�߮����>��k~s�9����ȧI��5��hWuu�X��߿g�G�[�]Y�.t����M�Q��1r�q/���ĺ���׳F��L,zZh � ����9�a@kԉ�y�睏n�v�EEӻˁ!6�v�Dw��!����,^��_�
"O���:�X�]T$!#3%>�҇���)�cP��.�8D����Fˬ�r� �%ؔ�3�!ӓ��R���Gꅖ�Z�<�<���C��4�R���w�������M���\�m���B�^M��r�q��jN�@�����ͷK|à%��7d"�SX���	�?�`��3r��ǖ6��� c��-1-�	,q�>$�2���;�H� �}U�\>5��P,���pF3f~���	���pUk�� �r�x��p�U�u���G׸yKyK	����?Vy����T#�����8�3���i�9W�T;Kvzgg����$���hŷ�q��?Kcw��.��V��͜�E��.6ʷh�!:��`��M*b̔�P��"��2ҩ��pv���a򡜞^` R����������'�w�^�9O��i8x�7w�T��9��{�/=Z睟Fq���>n�����2���=;���ަ��C��g������L�W��|��������(�&?����ɮۓ��T��4���%��n���8��-����E�Va���?�{b,<R��<�]������&T��� il�Hz����[;:�rtVO/7��?D��L�λ��_�[�5�����sx�>O�P;%��n�����v�(O<)�wN��Y�D�|��T�'
�,T��\�G��&)5]>��A�g4+�%N��S�A�٢]�)�'8���Z�΁������wD9cNV�~] � ﲽQB��qj��y+(����	�:�C����}�� i�gC�K+k.�Zh�I.C�V �o���H#e������888��{��E��/zά㮸H��>J��95uĭ��J6���f"���O�������)�S��-:�B��������lP���q�Jf�Sǵ<�y�����O�Vb��z�Id�b�h�A���|
l�>�MX#ˉl���U�(-�xd��/�=��7�.�Ą"ύ����A4H4s����hí�Hv�j%��7�t�������O��{���5�z����` uδ]��;���;0_���&�g�z-����%~�Y��q%����TĖ�ϻ�f��>y��٠�/���z��}ґ��V;�����r̵�����������Q@@�C�"�y��BUTē���_g̱5CK"i`�44tϟ}о��ۻubL�c�pZ��aO�q�B�E��/o"ۓ��Q�9q�Χ!�V�N꘿!��ʊN/�<
#bI���LN�) t3�.���8��Ku@6�5�#C�u"�=}�/��!Js���S��{@z��y�A�K��a���i⯬�!��H5`5dB�zV	��,�_��	2���</���ےC�=��Dx\���c�9+����˾&��m]]�����ѯx-.v�"^���u��f6
~�N$2~6H���~0I���Z���yņ�?�H-,I}�IIdΞ��Ӧ�bO����<�_�/���� �x�ÙF��V6��I��Gয়:\��G�i����tTU�Q�Sj�.OMj~�Pe$!)�j�VBi#�\��vQ,���\��tsg�fcD���)���>�6�`y	�{��h�LT�[]��Őc�f3*>��δ�(�w=��^J��	�u�މ&�X_����s��ǃe-��ς�cd���TB�l-*>�Դljm�ս.Rv�H0�~�y���!w�X��sN׿iaF�d��
%On�N�x�\e����L��|�KW`�*S�a�l�B�г8���Sǿ��c��5�V�IR/�H=O��3t�Q<�������\Xa�������S�-n��\��B�K��IP��m� �&Щ��n�Ik��*�����fV�J\}�����/ڋ~�+@�7��Z���YO��便�����c��<vuuM,$`�1r���T��O7����q�$]S.�NN/�2s���7dd�A|ԀmwƟ��9�zI
8kA���B \j4���e�y|Ȍ���Zc����+a	�\��}>���~�T�������i�D,1��\4'�B/���}�{�����Y-/���u�H��0�Ú/�n�ꨈ�+Av�T^}���BQ����v7���y�����W[i�RI^�Y�:= 򷕫O�i?�G�5�nʠbxi4� �HIz˿���A^�#/+<L��M,tl'<�4���7�Í�!T�1��'??�MTÆ&�����P������b��CflU}�Վȷ쾡G�}��_�`6��Ў)�m�L��dP�l0�땫�����Ӧ9��`"�;�"�֢O��k
+��j0$�<O"��!��S�޾�s�ϖ̴����7}1�����?��NI�7�<&{��W�Ξ���>���d�tl��\�ׅ.\��?��r��Q�ԉ� uP�~vF���fcN���h�j@ �ܧ���0����؉c��n�~�7@��MJ=��t�9opm:'�yXn��SݹS��z��YGW��:���g\y��;�R����	�D\Kq1.��s�$I���S典jl�����%��0� ���n��R��k�w��m�`U�`s�3�	��~�3��ٯ�x���G/���&����vv�/��z�n�0~���m͈��RH���Ej`h�;���,"����R�.y�;�������5�Ҷ6��C	�4Jհ�{�����$(xk�GH*\�l����ec��W�b�����FZ�Jj���ʚYX8E��>�z��x�-2h&^�8Gb4FP��
����.շ�HQ��l�>���"��x�-��a���?G��k!a��*=,�oo�HM�Eu噒��^s��1w�����Inv�}J��꾪:$Y#_�i��|=r`�.�F���!�h�7.9��1�"�߬
�Q�P"�ҡ�_�UF������XGU��W�����uf�/f��?��[^�PzM�H!��އ�O[��Q�go��x�Q��2�T��t��鯤[,�r�$�>,"7���i�,ˁ��(oﯸ�_`�C^�s��WINՌ����#::4a��P���������rW��k�k=%W�qd�����\����WMmC�"r�����:�v����^���2�Ts����GAlQE�k���y�V���3�I���B���3kkt~�Y|�γ�z�1S�Oo��sʾ Zg�C��*��d��������-���M�E�*M���
�_(i�1�W�eukF���}���UK_��y�x�t�)=ނ	9�����e�0�����s#5oب4rl�]�F��p��eo�Y�]�v�%t{��j]�������l`Z.�o���-��7YW�)u�L���\������f������(hPd���Eů�P�8��Z�k��A+�ޞ�[X6s��xK`�Vvt�u�[iX=���;�]��0�u�p�Je�5�R�`�b����oC�cD=6���y��2���;���=��P�u�,7EY��~��x�����U>�o���/�5W�#�7*�k���������U	�awo�T�q�=D�+��7Ǘ�s���=y�|h�ݳ�-ON��)+-��̌�+��;��=bb.t'��ݖ��ܼZ�zQah��E�W�TJк2������Ӡ�@��K��T���ہ����:�={
�Y��17E,�xb��0U��lxg;Ǣ�Gs��QXC�3�{5Q�9�G*+{�H�M����ÖG�G�(���p���
"}�;�ǅ{{�tŞ���c�
����>��9�O����>�^K�+�����E�����nHL�`x@�&ҽ�`mxТ�����K���-�t~˔z��ݨ�w��3�W��]>��y;nu���e^:w����ΉrEZ�u��K�<�9�>	P[��ޛ����|�'ǈ�(��lq�q�2�����O� %>*'V����r�E?��Zv�
A�񴂲OȨ���u�]�7��S��햮�]��]Ѱ9�!D)�y�i#uL�4�C����|o��	�����p��W��ǎ݇G6�Gf��<4�U=�r�)��+&"��O����4;�l�H�D���BĴ���ciW�i���׉
�x����������g�w��ߟ|���E8�y�*��e��b��mQ|���nT�2u�/N-�8��DV/e��AV'���"�\}(He?�0?��U/��h��{{{!���*�_�h��~��? �X�s�����4���!W�����K,��o���dc4����]�o�s��l����mFDs��+����{�p����e�
�������FZ�x�>Ř��V��$Z���0I���Hѕtr��o�-D캦�<O� Wf,<{�l�:���KQ�2����kT:�ݳ�yx;��q���<���v��5�ޗ���=6C9�C��"o�p�Ցa����i/�}��Ἳ��NfO��P�`Zj�@��S��� l��3ٓ�|�i)t�������� Dy$�����|�)������2��	.mB��u���ۙ)t�#=����O�<F��S�64�Vz�+�/]�r�P���pJA���&Z7��G�x\����H��2~��IX�&��Gם�TѧhTI����KR�F$�n{�ܫ��&8h���j��I��H�C҈��a�P����bKs���~���F?ۑ^5���*V��uI�+r���2�K�����n�R���w5}1�O���˛g�a���/o�4z��5H9o�>~=�&���,��Px��� o��2�E�Q��G�nRo�qxyyk�X��p��EZ\�wɊg4�OM�/̎:]�����Jn+މ:��������w�Iꖁ�e�
�_�4�^o�X��n�
����`m����(��2�H&�p/얻��ȺϾܼ'0R W��x�/eV���&������?�f=��۷��aD�VUE(L5������U%�]�+8=9IDI�D<�̂vE	՟3T��)Ar�W�1x�M:z��k��M���1=n��ѱ���|P7+W��ip�����o�Uo~r/�ū"ss���i������w����_�V��m8�-,Ш��L����뚠���'&��+���yΫ��@mz�z���Ąb��ڛ����{�{�����|s�5L^~L�� NZ�f�a��]i�^J�I6NN.��nd(������|d���:� @��o��ze�+��
@Q�������:��!A�����/\�;�M#��I )Ҍ�)E��7�cE��+;��Q'�F��_�9"�m�����J� _D����u�N�E���*?j�����;�W���qJL���♖���ݠ�Τʨ�9`�����tQT������~=l���)�+^0(�&�g�:������̏��e�Q�i��c ��Ҙ�G��� 5�mn9��FY99Qx�~������:��ӛx���xc�֖�Q�Y�B�?��#KKO����)���u���m(�#�R��}/}	ZEW0`yZj��īu�3��6��ܱ�u{?��!5|;�n6x�����vM�v��5������=ы�?.rTs�$�W�c_Ot����)��il���T���]]�^ƾ��"�;�w� ���nD����ؕ�Ţ�kj�aD2K��e�p�U��i;��:���gM���Ź$-��$�Jku�⩺^��3�$1��Bl�?��z���d*$$��^��(���hۢX�*� 6�;g@���s�u-�_�V�2R�Rg|��W����߳MB��I��I��S��ȝ;��)�ߊ�v�L�)@w���E1�wm�I�b¸��͚fW+�t���
Q�Ǐ����)���O$�4��#9�3d���Kg�#z��
{5����G����DPQ�Sh�0�	#��ߵʄ����%�j�D� ���2����s�N�~�`0����$}�.]���U��z���t�[�9m�\$��p�����L,�?UԿ���X�ۂz�;_{U�
�GR��`�k�.{���]q[�!૷���}ۋI��J�N�Y�S!d��v*111��@�%�w��}ԥK���w��R��� f���W�kk�HP[�{��rpU~�����D�����'we�;�z�4�N��F ��g��$�D�@�-�ȁF�*���+�6"W��s�ĄM@t{n\�_|N[�+/.����Dn��H�%��Fw������m�?�ϑ
!n �z_���fN����e|�E��&��#��X�(ص
h�aV����Ǧ\��rb8����8���ъ����0OS���&��!����ܡ���`҇�j/J�؆��>7+I�:�����ss�Oό$ugSFK[���u<H�M����Ύ9-�CJ}�m,Q�,ӡ=��u�+�%D��p��(�_��k�T#w�c��?�b�� �i�3֯������c���y��꾖�>/+��o!������S;;�

�E4�\�|�"s��<�c���%�ʅ��J�����:�/����L?WOb2�m�3ر�x���~�mK'�B.�W�������r^[���o�����D���XkÎ�i��ץ;>MOKKc��3-��Q�m�ec���k�����y�k��F7ve��A5Ci�&X%�k-u��H��.iEE���N6�8�UK@��ܰ}m�{$��I~��󼻅��1ᔦ�N��G���Z
�8�<N���P1���/�Z[#.��	��TXݞ\ߙ\��>�V�ks��)����Wo`���J���Dk[ݿs�_^��u��l;I�fH�~u�~����P��}�]���.J���g�J��� ϞR}���'��\a��)�-�<��Oy]��/F|�ȝu�JH����/���tt}79@���Ni��`(;A�;�����V���|����"�O�i?[&�raF�@L$�W��!����h�-�?b_=�q�exD��ۂ���(�F��]�M�[�IE%+M�ڙ��3ݢx���X���\<�y��<�FĂ����W���y�Ju4��}E�_�9��i�c�ַ}�"��%�,�H���ʝ��e�̹�|�c��^�Z���Ž�IT�\;2E����w�D��ӳ��"�X����!
�	W����T�B�`@0�~J�YG� t���Q{~
'.�&Ǚ��r��w]]]��7�s����_"]�z	/zץ�$[0V��9؉�L��n�~��ѣwp���]Ԭ.�}��=�]T �$$>�\������*�|>�#��`�x���)��ڱ��ص��BLV�����d]i������Ab��臃��XIM� ��h������3֞�gdM/]�ߗ���С4�vF6������q\V��mU{�'��������I�'��t��3�7�cPZ؉0��N�c��#e�&Dp\]/h����� ��5��:�g~^�%�m�N���'��R cᑟ���m\��A��,����+��Ñ[$��CDi,�ߥ9���x7<�	�`z�+(����_��,ͧY�t��������w��.Pdɲ�lr�NM�$��pwo0��u��{��A�&���Ib�-��AY�-�	�p���v�~�f���Jm|���xE�C�3����g@t'#H����Av�8�At�.�7u����<Q����^T#t�Xms���0��u����u���v����*nv�&:%�raEZ���XX"��=�42��8z]A�rԳ��^��Z�gh�[|�.p��_��֍̒���y��#�!�����.o{�n����S�Jr�1�<8hFl-0'ӻ+%!&�}��e�g���:�$ȩ��ܾbm8Ψ�j�h��r�EE#����=��"���,"&v�� ���O��{=A�R�ib?��_�H��YA�����{�1v;o�G�Ȇ���I��e������f�{y��;�op�f���2���� �B6�^�s�~ّ��7��<e�����)-�	9���W�V�TBT�p�2���M��%�����nu�x��}@hη���>�����rn�}C�2xl�(���P���?t�r���pM�I��a0�	�)�w~���ș�r*��I	�+�RS.��G�%�Ƚ��c����_�x`�X��;��4䮫<mW<�5�[|�h��F:Eѝ������/j��
[��O,w��H	��*%vv��6j�s�S{uC؆�Y�<S�ck��f�y�~�5|���Φ�<��^�3S��>xŮ\�-/���+�Qr6��/\���a����`8vM6�siI�@�k�M:����&�鰥�%?�p������8�[qY��r[�Vg��x��'�U��ʫ����m�;�-6-� OZ9��:D!�
\o�ȢӶF���3�;/��g�J��Cdx^�8J���"WzO�UfP�m^C����[[��(�5����s�d"��G5� %��(��R|���ff�k ��j���<�H�u�xOvw��a4�X(�GT��_@ɛ7C�ẂIo�֩��J{�^g=l2Ev}�Rz��t��)~~T�P���t��]̌	߉�U��"O�W�l�;(�|��WO/(�u5�s���s2�P�V2�7e1�X��1�{�+��%<2��!]<7.���fy�	&���QdG�h����˛�"�����s�\�	�����;`j�N*0�ȃ׸t�^�ڎG�1#�/�=�+�cs!(rS���3����yDY��ڬ�"8&������S�j�Ґ<�;<Lb,�R�cTYZ
D�⇶6+3s���wl�pT�ֳw���q,��IVK V��.�ۻ���18;�?\j-���m�dvfIɩ��$ǈ��rs}HYF(8R��1(w�'*1!b�NW�����<��-!���}�(�FӋ��!����"B�g�H6��1����=�0(�XN9��9GxԐ���nU�Rd�ϩ���J���(,��b	]�CFA�)���� �m�����!"|�J���I?�A��0�	�H4o��-=r��Ŀ5GF���!F&
�"�範w�x�P����Ҿ��\�|>�Pط_�fz�7��5ց��[����%N{�'�u��}�x՘�c�z�S�]0�{��G�TBQ����ɭ>d��t�1̾Ѻ�a��)�@YTdi5�Tڵ��~|"��0ӶL"k��Tǵں:e�$?����O ,����zx,����RBe'�HI��PJv�ΖU��3��
!{e\��I2.�2B�&�����|����qw��q����|�q�gˁ�\s���3ˮ"��ñ�/�w\�WN=4�[�w���R<��'�Ali�-q��4L����3����|6����w@TN���9?��� ܌����y0>dN�����F��&���FZR�j��j�`YV�f��;��F�N#K���f͆ƞ�ж���r|��m��^��_��2X��C��/,�X��z.���=q�k���^��� �voHepӷ��3�x�ȃ�PLg ��Q,�P���Ґ�vp�L,IbO��~qdL,�KS��&�J��}��e�A٣:LE^���9�M Q_����m��
5�?x��="�#d��BYp=�+Z�`4���PUZ���v�A4���!�Ǉ��>��cR�jV�{2ȫz���?�T�K�d󹗭2w��i�m.���z>{���K�P#�=4o���c��?~-`��y▴x��%-���������U�pk׺QP���b\�4�4�̓�At��nq�$�>�͕�f �i��&�`j������!b|@��N��F h!�$�.U^^�`���[C���!k8�l���%'�O��[�΋a�m���m���Ӿ"oem����76���W�F#x�F\=_�����w����t���;w�u&��/���v�K�w[T��e31E���E���j�|.*J���-J_�y��I��T�)5������EZUu�O-id[_�j)�U�3�N|}|�l�o����qV�:55uNSK��er+s
��j:5^w����ъ�H(�;����� ���Z�K���|�P-0=��HNª�ȍu�z���5��G˩Y�þ�ö���>�y��A�UY�����J,L��!R���E�ww)���l�������MK%u�F�!򞨻i�����JDee����ʜ��`�N{[1H�'���������n�5��[��0�ڃ4��Kn���=y�����6��>�	!!�@u�����i�����t/�3o�s�}�8Y��<{�J(�%��Ը�*7Z��[]9���\��~	D199�S��	Q�y���R��v!S��U*�9�
�ZR|�'Z�WV��T5�3Bڅ�b(�op�BCK+��r�P�ZUٝ�D"QRZ���W܈JW�1��rN�QdM�!��pCs�-�"�����$���dX��"TZ����B����������K-��e�@��2U�8�REȗ�j���q�w��ՠx�&�@�Խ���%��W>��^���.��q�W"�����S-ky))uuyEEC//�荏��ے��<uby��+�HZ� ���8�|�SP�0��~94T��f��=�<O��{�m����	Uh��J�G�Q2��)(��3Y�er~%�ć̜�;��"�Y���:F�~��[.N�W~���r�nٶ$d����pF������Y~&|����|>>�s7�̧�q�*.��$	�K0특gm���u9���?M;d(�6�u
0_C��eSE����}6�o7얦L�
�x��iS��
��@SWiJ�����\v��^��sp<�N���U���j�?�P~��ia��+O��-��25�����&�yq�U��\&�B	S<m��^����[6�B(MN*m���]8����F�tӃ�����K2�$��������c�g�$^��*�ѧ� �xmz���̪)���sN����ww�L��]��DDD�5�\WTf�F����cU��p);��$�p@p�����N�y��h!a��ؘ�	��VWC��h�=���h /��.p���1��:���
��^��ӎ�vT����4�?ͥK6ږ4w}�AF(9ٞ#���'���������k<"���J��쑗�ކ��a�ݙ�;�� ������S���l�va����s���_��U�kb��˵M���|��t�+'v=̵-���8�M�\�)���I;'�o��>-�a�J{eZ�����)i�2'��}d%���}����I��Hq�X�ֳw@w�.M��$s�t��Ȋ����QQ��$'add�g&'���O�Mk�f�T���{YR�W�5wF�-@���TqqqāV�7T+�I�_o�y G봺#������$��'�sJ�T��a�F��-P�w#GG|4��>)�Is��^�11~�����1ί2�)\���ʊ�Ҥ��?���V6n:��(7���<dg/�{���'o�%��5�!��Tʻ|Zr�6��앹>�� .	��+���L�}��z���7X<l��8�%%B ]V������~%�lX��C����Ńmg7~�,���kHE_�xꜝ:p�}_�uO�C���$��_"{5��	1����ȷ|o�^ ����"����T����Ez		��R��|�����^��an�]:)�H���l�3r�we�{m�����Q�VB����nq��A��m*���|/{zh�;��j���C4���'^^'pUL*f��nz�9F����Ĭ3ŝЖɦ�=����555� r&%��.�J{��+�Tc3t\�*�ML�,jci��,�c�{�3�\�o��ɮ�q}�fWÌ�����g�e$㘽F�=���va �w+�����ݼ���l�Z�т��?�W'�[��8�WT1�!�Ȱ����`��d�9����nk�׊���C{���OC��`���L��ߐϒI1ʂ���Rk풙�N����v��z�e��zz4�y�苈����~W++�Ț�Kڲ<�	�]��Y$���5
.ęV���*8�3�߱lu�k&?-idH�'Z�ᄺ�5�����;����ыp�"΂��}vj�7�ODw����~���iE�lZ^I�	���3)K��ic'�5mkI.��ܶ=�)�=�g"���v}=���я>�vN��K߀͵4����B#L*,=�B��R&��R���ǋ�~���Y�_��,���[W�h�u^��Cd����0�QX	P�.Jq�?��F�%����t\�����������L`�]f-��T��l4Eh+���)��cS��Nlmo���|	i�P0���܌���Z�C�༕�O���wR��`���X"�e5)f�e�_ߚ�_��M�	)+;Gt�Ѹ�6g���X��pUƫ7������eh�/�dO@Q4�$�U�@`,�0�g�{�Ė�(u��߿V��b�DZq<Ԉ*p��Ar���8E�����Ld���g|��տ�o:L�SR�R�?9mh����y��ѳ4�ŵ
�X��5�����������É���(���I9���c�gY��}�*��*B:�8��\Ƨ���H�F���!i�̺�Rb���P�|`�a9�
��DK�2�簢��%K4%*��A	��L&��hå􋗵T���6��qC�� � ,�L�
��J������+�}|RL�1���R�������� �k&���Ȉ���mP�ᛢ�F�*�h� 	�~G���5<�o�zƓyh*2���+n6%�(�v��Os"�:����{ɼ=���k����&����wn�@�O�E@�����3F�vF~$Qz��Y�C��u���4a0�_>q$E�E��##�^bʿ[�fp��j���uo9�a�����~*yy��<69�V���!�m�\��ː�N�r��)�cp�
�2硺���a�H􋱅�0�b	��3Ǉ�,�c�ojQ�_a���UP`Y�8������$f?}ͣ�ܿo��[�%����%�>3c^k쟻�
$�0a5q���e��.i�N�f�Ezp�B�|��	�]r�O�=:�$?57S2E/C�rq�B{>G�B�����e wIEE@]�a4�rU����kK�m|��DғQ���-��U�B���>�h��K�։�E��P��''f�IO��FB8%дϘ����Al�M8%��v��X�3��׃�������-���*�gs��/��%��5LL���p��p��T$���ߗQYdi2��:4tb�2눣�H=$��MW"0�����i5�X�,��ȶ�:��M�_J
���R櫙6�5#o��K뱄w:���G�������)��኏��yn}�k-ųW��3���W{�Ï6_K� |�����Y4&ni:<�,�"ě�5���j�@9U�g�O�S��S� �ύ��E�����Jd]�G��ѝ���>��k �fg�(�Wf����;�YJ��U���1S�Ǝ�b}��)�����)���]��X�P�;��T��B<���Tʏ��������6q� ��q_�3�'w����"���������6��"o��V�3���O������s���ع��𞖍�9M�<a�������&�"	�-���|��������H3�G2.����-��<�И񆔪�)�����-�m���x���y�mN$�gς:%�e��p�/Ҝ�Rcޫ�b��u:&������¸�ۧ
پ#�b�l��--�	<D6x��.E^(((�Pp�pc}��J���o����L�N~_����e�<�?0���;#�Z7OO�p#F��8'�$>�������M��A-~���uH����{�Pc����.&PE��9�����`ck+�:,���hd�YpQ�A��5p����&#M�������V!e_���YV����r�C		:�p��d���K i�093OS[�y�����B�̵=�Ĝ+�����*~6Zŋ����W�/e��y���)��t¥�qN�j!H�"|��r�DW�E�Eed�t)��4��I�8S$RY�M�-��&��B#�Y���:n�I�����;YP{1��zD+?���%F�9�pڱ�i"�<���@RjT gW�~��c:�{V�%��?�2v�U�+wŘmf��o������n�{,K�WW�<"C��ea�gf]��07/��8��j� p�&p��vYv�B�z�"��ee����f)U��^�8+�}�`}}����`}��S���n�"&Z%�#������rװ��J��݈{M�]�����}9�ސ'��E�7[׏P/Wʞ����9h�d����2uOh���,שHk''Wfe��rM�GGmm/lz��_�=�{�-i�TR�i"At;3e�EEnU����_5�KQ���w�;��_J�zQפ��MO
C,�k�Ȃ<���m��_&+r7<�Yc���^~':8/�M� A�o߹���� ��UfrR���d�$��q�l`��HZv��U�Z�8FO�hp$��u�c0�պ6ض�翋���"�F�̲R|���Fl������!�pr�c�:���5�Wȉ�����*�yuD��_��1GV�tum���j^��X����O�gCv���kR�lF�^<{��(�s� ���������zv��6)�� ;��6p��xa����l�O^JJJ�V��D�a���;���`�y.�������i�Mtܫ��Nf�������)>�vj�܊G=�� )0Αw��UU��&&�ߌTES)T��+!�C�����*-��jT��#�<L�*���)�Hez��� �<å���p�������N�R�g�E6�W�<HrrǟXXk �X*+�f���Rm���R���u/�2��tI��+�=�� �6����|a�&�71�+�!��KM?�����=��xz�u6���'1����tƏ׋�/Ʌn�Fp�.F�������C�D���%%ꁕ�e���ihh^��o�Պ{(|������ERXz&y�W_�"�����������%)�x9��Kr�QPϨ�i�3�扅�Ɋ�����5�ɯ�(��~��$INGNp^H��#&!���}��i6����DF..���g�(��S<'~wZ�����<���7O����4���+,�������T���3�&t@kt��.����1��M�M�N{����7�$δ�J�N�x��85?�.А��SKs�_����"��of��QSS��HX3k!��+$h���4�_o�ޏk<����<�3���<�	�R���!F^^�ف�4*h���m
��:�.�DHJ��%$������?Ń�D �c�^YAe�̵��&�4���r���5�E!Z�m��)�e����n���aLk����Y��[�3��ӧK(=6K�������kP�/����L~R���V�&���-�sr�*�0�k��t��N���(D]o��P&򛚺
z��I	^��r>��I�`3~�C�c0Nը���*��f�+}/�\�
��Y쑻���HAZ�3����j�BӃ3��(X�+<�gi!�z��Ċl�Q���u�ѥa����Su�JO��+J�#��m�r�8��j���� ґ]�Z��R�����������'�x#�]^�+��69>0 �IOjlmݲ%a���(�96&�cn�;M1�,{f++�%'���B���:_K�p^SV�3H/|�u|���xŞ�N��V�y��M���[L�L��Q�y4�EE���s���cb��y�6:�;�����}|��?p0s����X�&�J����=�lj�N�۷�9[�~�
而,���L�0��[�Bݼ>fO�&�<��J�V.���Y>�n��	/�=�r�)s���:�Oc#��oss<з��6Ų�N���fv����kA|��ڨ�ff����­������C��xD���M��jt���8_���P��nz )���?��w�ɓ:'ffhw�OQ"��>������,H��3���'�,P���,�g�cۦ>���=T�rt0�{���,@���iʐPă�\�JII���M���"���E}$�dʧT7��"���b�s��|E��g��D�C�k$n�9���a��S˘&�����)�7٤�Y����{{�)\��o%Ì���R���=ill�����\��6	�C��	�q�rDF2�-(%m��[Ȁb�=ST\�Z~�n��Y�%!a(�Zy�B���R����;	u6z��n��@��X9$�n2�����^�z�(R��3�*mx��(��\��?ҙ�oXm#8c�Z�l*�	Z9���f/�H�B߇���q��ȭ �����L��
B�R �J�L��ՠ2��ui����ћ��<���������z�:��I���٨#-�t�0��{-vB��/�B_�v\��'o�_���O������F�*�P��%�v�N_	D�� *�l���*�O���/����9�5�4Zt��;�{�VR�,��lZ\�`x��x�FQ���s��*�r�O��t\�5)!Ư�(������<�:�p*����Uف��?t(z�[P��.�O�-���R��`�vBa$n���6͸��v���+/͌������[g�Lx	>��y��FA�����k�����rvKNⶕ�������zI�&AV#w�S�����CK�s��H��",/Y�@#�a���ڃ�s�� ,�Z@X0��>Y ���B�)1Y��"V�;���w K%3�Og����w�_��q7�; =H����1�/8�wY��`z�E��|�J�t��8�=����n�11UG��݇ ��=�����~�0߆c��#�m��uL�z\�q�(��"�P� �olj��0��+)+�J%32��T��(����-V�`j�[卋=��4�.5�Ԥ�tC�Vh�TU݀�{#�|�uйL��e��Op���E��B�c�d��^Bn=�*�`@�����g|��'*6m깭�����> 9Mg"�_@%ي�d`��`�F���3�?������IW��Hj=z҂�D�p!K���
D�\."g��j`@��ޗov�f��~�>��T���%��JRg�.�U*��͕K(�?f�9�{b��@z06����M�.��K��O�Ѕ^E·P��A�AZ��4���8w.fe�_e�A�J� 2��Йc�7N]�y�� ���U�<i���nbHP���%��|��C�؊��y�!	�_�F�pM�i�aŭ�w�^(��#�?ۆf�s	$�6�'��A�,��/��-�Q�p�9-(8� #U�e�������oz��=�f��7a�_K_������?QXߐqcm�^M���Io�Z�p/��$��]R�� xV���w����>c�6�AM�5�bi���FE��40��Zx�	).�|0����ܜ:�o�^�_j�=����c������׌�����9
�x�~�
K��{11�̔����g"M���(���Ln�9�Mc�~Kg�<&��Wc����������{)��B����OMx�e-LpuC�8 H�:e}9�|��Y��}� ��!����W��}��P���s�"��+�U�E���
.�K��)����_�6,Z8[����_���U �&��[�5���GVS�o5���/��n���x)���;'g˴C��������o�QxX�e���������,�����b� g^^��	`�I%�~������,�_��sml�d�eO�cض�\n����w!]ݩ.D�~��I�q�:�L4�^��n���H&]^'Z5I�1?R ;���4 ױo��֊�.'Ϭ���G�]���b�{����ͤ[C���n�B>Ͱ��r'�z���G�H0��&+�΢�x���٨_�eC޾=�I�.�磕��]k��|����ܵ���f�-`+߱�X�_++����Ty�M����6ge��lnz0 ���b��Â��=FE!'"��ڤ���<����TŃiPc�,��롕�pʑC�����!3
Z	6��^��Ky���&d�O[G\�s:^{N��a�lY��@�^�"+?Y�*�F�]SF��o��Uy�(�Q�H���o������^M�n�S2,�����w�l�9�n�k���ײ��w�";��ؤ�B���]��5	|Ԋ�G�}���e��.CV!�%�x��#�<���%���b�nP*�d$-;��c�����bg� ��׷�������C������:cp�z�<�����Fl�C������!,*�C�҂�	B;��`��)+�I�_�g<�z�_W58��Ç�k���w��jZ�n氞���<j�����OP�e����E�����h��p��m�$�H��-1~�������n����Ai�r����E��.��ۯ���sd�m���c���������H@^�`�MP���W3�K�:Ս\�S$�S��SPxc��h�
0P�Q�c��;�!òq�ab ���	��h�ar�������>��b�:#)a��p�c����e�,�ۮ�����''��E�(��;&���#�z��:�d%X�
����8�٧�'9ȉ���/Ȟb��]Uf��qQ�SyCHpT���
�Wk�G��u��ō+�!��u�Qnb�/p���#�A{��4���)�������<99��О�(D�-�s,�FR���+�x�����>�A<w�Aĝ]�,+��q&�2(�X�6��-��.^��x���:^43��%ӯ�]��:3C�l\��g��E�[��N�Җ�9;��)�����ÇLADp�mN�e�����%(�y۸cH0,V�h���M[n�բv�a{+��g{���שiii�"r�Oq��_�@���|hll3?�؈���f�����ψ�l9�F��������������/�yT;�t��EE,�����O�-�B^J�Q.> ������gx�3�J�����}����
��.Xw4fiB�bJih=��z�2���h�O���nBa��o4��?�a��Ɏ9�r/�{���/���z�!߀KKE��v��/���ǧ�	�RHT�iƅɃ��wf�Z{��ub]���xO��QZ�Hx���z��m���5���
��vřI��˽σə.R}J�oB�"�O�59����f���x�Y��*�1]�r�HBB��K���*�b}��i��i]e�jӨw�Q�K�^��O#s��w���U�:��yǆFqr���(�G��%��lB����hV'�$j�0!A+<�qUkѬ����嫸���Ĕ�����f����JW��򔒞2,u|||�>}�[���,]N߄�>����d(ѓq�7b��}}=<��95����~���ͽ�Fu�d��ޭ�t{����G_�-<n���̲�?��8�חUe�m:���XUUPX�I�{be$,<���7�3�x7�`�G�2�_�\���B0>
�C���$
%
W|Դ�q|t���VA^���#'�ؿi0��CXD�ҎM����^[�M}�e9mtd���Zr׫�~��[��ܹCKC��{t��UX��ܯ_�Ϟ]4-��&Z|ŀ�$��������@.��4���]�|y�,�ԤG=wk��*>��Ϡc�$--o
���*�^?y��cs����nAX觭�[�����Og��w�ccMk�<g�+��8���XZO�Pf7�F�P�K��4_�i�/ڞF����0��lȷק	��989y�\�$��Z�֭2ڋ�M󲲮Z��pRX�qg���n��[2�������ٳ�j��h5���x�吿677���,�udb����j>�� �7;�Q��N��p��o o�jaaa���IS��6>A�\��H�������HZF⦲_B�:*��N`������)mos�H_��:;����/��1��@����� 2{��˃����.v���I����D����d̠1�Ztt��<�4�	���������)#P�%��
:�J� �BCm.�='�Vx8:�7������ѨD��!n�;KLOkkM���򴆆���\o�e����u_]Aޥ	�0_X��ţ�>S��3M�0��.������P�������z۾V��(��J�O(�D����{�g�x4s�s��b-��g�߳�$zAp��qB����=j{�>�����L��D-��jt��pr��-~�x�r!�38������������Jm�_�n�*�ȘL\�7M�ѯ�(������m�<�e%��0A�fMNR��E�KaW�n���>\���_�H��L�:�B�s(��Pn�Z�I���tQ+��M��柩_�Z�M��t�k����on~aUWi��:kni�*-D"G ʐc�;�ijJ��ۣm�tG����prv9�D8�������?��>EH��V�F��2K���*�f�^ΨsO�wNI�d��J�u��Z|<�;����)hp3�[P���ټ�[衡�	b�=���h�O��iR�^�=�
��	v+mMty�w����ei���g�f����bi����z��oB3`>n�����`�%6�ʍ���@0��d���P>�C�ml���6Qh����v��-�҂�������[)ii7�;f�Gl������_5Sq��m�]�{���%��ޛu�==ʘ�iY�D-	&n�Z넆���?��-��p_������P�[y:
F6L{�*O���sh��`ajǽ�L�v�P>%%E�� �����^����d�~��O+g�����8�郛/�'J0e��݅�?��ƣ;�~7�1�+���}Q�=�C��jt|��k�{�������3с_�<�����͵���'%��[�m3��y�oݔd�ʏh����G*(�ڑ-+s�c��?��t=,��g�:��A�B��ɚ ������^��:�P[��z���Z�v�+;55W�����c&n�LQ�� J��Л���3�$2����Պ�1X,�Ma���W5M˴@���@�6��~*��ө�h�x���D��bʪ�KR�Y���z'��	H��s�M6^����֖��\!{Am|L����������O�蒐�X����_��o���D�gQj�j�� N��M�[�S�c�8�`|��ring��?��ݿ���L5� �53{���M�a���k[_5r|9BQ��E�X9tq񣃃����.Rny��c\�]7�N�Q�gR[�yW�lY�������#P���ng��\���v>�)����+U�f��
Ϟ%d�8�f����޾=0?�����'Կj�LUG�u�������������-�9�c��}$���O��.�v{�!�K��/loG�G�c���
��+�-]\[Z��sPٔ74�ttt0�L���+�ݏ���?^u�hnP�T�,�����B:!�j��R��������
妧�� �]3rMR��|b��[S�a^K�kk�o��&-�������4mu/��SM��u�
e�{�Y�\�A�;�GE"ˬ��VE���Tء�.����< �,a�蛿���7sww>7�����:��|�}t􎶦�0o�ewwwEC��z'B���\�^.I!i��[d�N|��ޞܮWj�7�,Ĩ�9@�����^�6��ֽ��<t[����p�*u���[Y8����_��>7q�"�ry\��1��=F�<���O�b0��yk�g�t����*J��ܤ������>Yl�v�7Gu�����r�1�CV��1˞$���_�W&�3��w�����.]Rzwʧ�����*��Ν�b�s|�Ƿ��L�=9]otO�����?%J;�x4<�ZpY�Ҝ����uGh�ڏ�o��ߛ�
��e���ki�g����8��N�=޹�QZ^���:��~�]/����u��FHHI͝�����@�۾4+��誷����j
G|9�>��t��x�#
�4��d#�9�V���ް;���:�34�xL�6�o``	��U���|�<����f~U�#�Z�̯!chǅ��������݇U��N���e���l�pq�tT 	��j��WA�m.��tu��n~#�l����]����30�|1�N�9��a/`�@�A�g���ٹu���k��;;9��֮��>B�{�vk�t��M���P�S�9�T����eQ�:>O�{ob�UD/�蘒��6�j4+��L����/-+�=3�;h}O8ݛ&0ci�&[�~~nN�w-�	ZYT� ��v]����*D�<K������#�<�JC�mv��ӲoO���z9y���=��oz��-�����mm-}}#�n����R��޿%�Փ�Eu�w\0Ԏ՝b��v�h��f����W�����e,��~�>7��d5�L��8�#p ��D��N��~c��v�����>>`
E`Y��� &��E�UU�vv�C2��H:J��6�+�*�Ch���:�����EE6�</e���h�e��:���������w�3��i_��˙zv�p4�o���v����o~��d��!ꕝ}M+N��륿<�������<@�aw7ak�e�'���X�i.��J�d�'��}��T�Yj�����.k�YC[��z��_<�� ���xl�4��II���ISB�,>z$}���Tέ�'��^Pp
�H�>y9���ޜe�c���]u�dT-*�urO�LOgsrq�(?�/���f����Y"ş߿���p���tvv������x�V��/^������8[.;�![�>Ꚃ���v��"�[.�����\7���̀��uO��2""��-ncG6b���C���,�b��� ½�ի�����F.��B[u�<c�lml�XG����`J�_��I�2�!����݆��[$[��-���w����f�W���[����/���{���D@P���4��~Q]�Ս�'tttFۜ(�|		����uH�FD��9�O�������*��>3��c��oΤ�{�)�q���Tv�KK� m�F��D��2F6�^�g#g��<�=�Q`�*}N0����ښ����z�O�}S��/�VP�od�آd��ַu�{��z�mQ�6�B���Z~2��QM�; X����e?8��zz{u676����M��:��!V�����6 ���?���`�L���W2+�Kl�\l\t[�����`c-��~~Ǩ$�u�A#C�̎W�Y�����nL�j){��&x
���;����E.�mP�k1z�b���4�lԡir�U1cg^�	�l�6s�����������z�uʔ���ط��ֽv�f�I�n߮A�ʋ��z733�?��=�s�{���@
��� ��)����b�HW5g/r|m��t���O����:Eʔ�8���*|W�6HDŞ��������?}q9���&*���C�c}�%�ݷ�&bZ6���s����#����s�0ߜo:wLT����Y�^���2ۘ�2+Pc3�[�)c�}S���l|R�[y>������N�
����m��v����:5࠻���l�N
Ed!k)9�Bv>>E�����ʷ������z�t1������(�!Dun��fB_�w������b�R��ۗ扻���W_�<��N(�յ�?4��=G�V)�M����7'"b��L�3���|*�y{�u�,-E��n-�p��X�������:e����ߝ�FGF�4ٽ�|��^TП�Eu}؊�M���Q���iW�ieH3Z�����Cչ�i�c<�Nnb4??�Az[ |��M~@	� �[������ŧC[3��-χ��G��1::���j�V����nj*k���5�0��11�4GD�]��G��Ć"�Y�%h;��{]}31+����?��������4�i�Bh닻>��nm݋9���ɛ�ϩ�[��f��#�ml��lwhk�\�Q��d��h��Лԡ޻��"oІ�J�{���,������9y{�_����,�l�:��8Hp?��^oqii�1��b`45��@?�S��}�^���	/j��6��p2�����M�+���BU��Y���«S0�;���Hl�1O�Y͵&�Cu�$���
��ؤk����Z�qi;������|h�
7�V
�Ā%@|8ڪ�P`Ѱ�}�ַ�>[�:g��}����ʬuz�6Om����3���K�D���n���N�KIK=}6?d?}svvU���l5�`�I3�>�
�ʚ���/���:,�>�1�t�����B�:�pkfx�=x��iu#�nm���:^��pB�u�0�hbR������sxk��ϝP�B�����υt=S�8�߆�W�WG���Ū������Δ̞|%��J"�T����x���v����.ӭ�QA���[�@ ��c�w_D􍜤��{`��xs?"��k8���\���d�a|�5���s���X��  ��,O�!~��G��M�d=Ī���`S����}�R�m�,Fn�g��x9���SO�)��f>�t��4�ql]�kae����s&�J��0����
Ň7�{�5�7RM���.JK���v?7z%A[Q"b�=�$SU�o��K�?�r�l{���.��H�/���N*���W�F���x?�8#*���8F�&.nl`E�y���뷧��{���Ò��������G�0�-,`�MdJ�i��Qzw�A��aPH�����K�>�/_jI��ha�ﲮf�>���33#�}fB��*��W�÷�o������q�	���;�f�>.��M).���Ǝ�x��0 ����j��a�&�|Mv���>��*��OPK=����c�ӂ~%TV
����G̗��=*�L��Tp�CX���9�ow��O�[��ȚJ�	��z9D]~>pr�����fJL�@&_���1��P�{^�q�(��w_O�J���_�<����&�sa|yj�0�W�Q��a�ٚ����J�?�@�WkiG^r��VXK�ﻶp�h���1��UP��]�S�o<�0l��<�:t,+`S��׍r��Y��`Oԏ��d�6�$�!��sX��iqp5o��Ȑ�]j�v�dis�$`�K�4�t����eͼ�M�qw��侙uo���-bճg��^������p�I"�90H��Ν�tAa ��ը�*�|�IO2�%�ѱ���}0�K�Shl��@?/�����֝e�,F��������{ݍ>:*G��� ����[^4=�P��U���d%z��5��@/TBˠ �����%)L�d��M�lt� =���w�2?�̈&$1VƩRX+,�a��<6E߶{�h�
GG�ӚnN�|�`��`�H�F�(F�����J���o/;9�����a]��7W�#�������JC��W�C��D�����_��%��=f����D�M��>���:F\�r����]� 7�\�v���r���sЫ�;��*�#����y��U�UU���"???�63�lYK˛�c(K�����?|��ԣi扄���=VTU��ؠqw�o��~:�-c��b����6�������!��k+�4�h3�|7�M�C����,����5��l��C���I���J��ɼ�|k�}0�6N%L���i��\����L���P����7���ia���Ðe t�����-�O�(/P�8p�6,�t����[�D)Q}���*��ޤ�3n�>�]]7.E��yg(��ڒ6��uV$�����U:��z��lPx��כ �Q��Հ/���c���O-|�v�4~�݉�a����N�W_��!�ܹ����?v��)�M͂7�Y��1��R�:%�~�S�}˴î-��PK�qW}��B�p��nS:�� �=8���%`yP�{�d�� �vb���X���{Ga���$��d��ՈG2KY����h�Q�ȯ����uQ��؎�0�l�c;L�[>R����=ZM���|�L{�=��յ�����x>���&I���f"�����vgwR��I���曒YV+XVA�Ap�F��SB���G�q�5��z~I���뜺L��À��1G�%000__�3MDOo��-��w{zEEs'>����p,BZ_���3OL{�T3��5%�J��!�����:��E>{y_��`H\G[5�>"Q��h�{��!/�l��w�n��}\�嚱���k8e�Z��Ύ���忥�+�U"���

0��q���zv��(:J#��c?o%"}��[����>�`Et����u=+^�����1_jO��D_O��LF
7~A��}�'��fDDFV��+O;�t͡&�i T�r��LӉ��V�gCv�pՉ3��+�펙u_�^�<��W٭��T�T�J�7qŨ��)_^P�����L����<)׷��M��R�\�������)' ,`�^��&�T�N���B��8�1nK���,ů�Cs!Qp�a�K���Q�6gL 
���VA8��g7}�����Ľ�:�5�bdp��-;*n�ɶ��ib�}o��P�q��|���`����W�*��>2��8�~�E�a�q�+�+�ݣ�_�����7m�w�Y�O����A���I�iy*BuFpxlL��Q{��MV��d䅔�T��Tm8����R&3J-��N���VaD�@WwwEU��2���:{�{��8q˄�~�}� ���G|���^lb%C׬���a=�y��I�++���B$�H������<�g0��R����h���uT�|����FZ��b۷����E�0?V����r�no[$���SH�ˊ�����s6tZ������x�K��>>��='}��

nn7�b�Ġ�����������[
뗉^U���6O�X�cŮP�����Z�_�
�ۜl'��v����7�~�!��:K�I�"�!KsF�7t��..9��=q�G>Պ߿A;]�&u�E�Ҳ�����g�Oy�^���0����zA�t�t�}�����L�?
5��AJZZ�f�%2�� ��j��e�7ݳ��)وL�߆����΄W�=�����8+++�X���`����G+77	d'������)C�?++�����M�,E��~̓�V�.���o`���U��u�^�Q7p���������Q�k浇˾�/e����Xp�	��P *M�M���>��^��[lS�SBO"��	���L��3�O�:aa������:---�	T��~��g�&�9� �'�q�-*Z�y( ��O�o�R-'!%������f��8�c�4����c:>y�A�G�����e�
a"T�!ST��G������A]==s�]S�~p����{{{��" ���2@��;�\`����:vj��ҡ�pq=�ڜ����Bo+?{�c�P���q��9$L.W�Ȝ�g�Y���Wou�������Ւ--��(Ym�e!��,c��F����졲�J�&T���(d�R�&&��3s?��������ݯs���z/׹�G^O���sD���9��E�.�*�O�3\�V��j��Մ���历_�UQ���K���+��V��������ˎ,{���_=��E�/�QTT_YY��Rl�Pﳼ�jv)x?����D1�~�/�W*Y\<���7%����22�~�2����4����'Ѿ
���0�&��9�2�߅���-3M���]z�)�]V{3'�{{꫰��-Y�9��ⶀJ��K�.��R鶰��r�2 T�^��	}���k���� 9>����a�O]ll����A���ꔕy%�����_��[�{���Xp� ,��t�S�2y�-���,��]ua���}�m�����r�b<��B�{��Tx�W�_�q))))��w�}Ꝭ�m`�+W��}9^SS����C�g�����|~{;*+����|����?:%�+vra����T!#&JO��������
H��
�ujW�*]�P��+�Y2�p�.}~^9����73���0�qQ�"��ߔ��|�/E,���'���c���=����A7;�+m�I����"��::��{S��K���k:�(^��+���U��4|��S�@���:�;^7�����p��>qږim�{Ğs�Xj�aƥ����ɫ��I����Kbmdd�Y��`��������hЮ<�oh�������5O������?bt]�,LP����q��k�+�]�2	��rͣ= u�!���ӝ��,i�M������
�v��y�i��޸Z��ձ5�HH��-.$�z�3o	*�E X���.�������Ӄ�怷�#T(�**Y��K��꒢�֙��vZ��� QN�������}��?�޶�6���ގ�Ћw���KAA��ӳ�/��MLL��[���q��2��銊�#C�N���nh��\"��{�fq��1i��;-������͵SE�Q������O�������_^W�"'��[ZjUj�p�MѨ����f��yiiihK�b=$Q��H��
�DM3s�?�72!c���'��2ԗ��@|���OmҸ�066l�5%���f�Bw���e+���5qў|g&= µ5�?XKѡP(��5�o�!�����ymx�p��l$�Ç�FG�8��GG/�$ܸ���V�d�z��ŧ ��b��*�"�Κ;��;Y$r�n�s��#�����z��ŋw��U׉%�u�%z�&|���;32�]3��6�[d��CX#��D$H�۷o���.�+�,����;Z��(P�wv��Z�5���ɯ_� jÂ_�|��5�p�۷m�&Qs�*��<73CJ�=��4�ɨ�S}�߭}!))�� �o�Q�}��1�Sh�o�^�ݽ������Ҿ``o'?�3�a	��?��e��l-v0]���|�Ȧ��@x
N(�!��v�`X������
>![�}=:%���nm}xK��L&������L�=�������	���Nb8����Ƈ���3�Vig��qx������,0�

�CC�0Ň���A����E?C�.�з��|�&s&�����D�=B1��4{��s�LDf9X?:�<�/��h��t��@j�0�,�iei_��終ώ�<���Ó'������M�|��u��09�ap��	Ԣ<��87�����G�\R�UQ]]ޔ�'��hk;�Yk=V��NGG��ԛ�R8�����@�������� �[s�G!�Ү�@F�FrF���!��x��7T���ҩ_� �=L��!z����V��I�^Z2xQPV�>�U8.s�n�ؾ��0�ea��O��+�k��]�|ܺ�r��M�ߥ��Ӱ���w��"�t۸O���M��C�2��
�k���(ͨ:������V��`p�"�_Ł�{�Aw]��vq��}.q��e/�`��,oHw�X�M �f���1v}HU�zWV2�lٲc���	��))�9D�bEE�#5�K}��Ve��Ь_@J���ˬ}n�"-b��vf)R��)5F�W�Ė𻜪�T�t����__Z^���Br�Qi��c�kA�����h��

K>k�R���atj!#�4q��!9ע��J�By,�|�=��x�&
����Ԕ�W��J���J���[��S^GmB���h�]����Ꙓ��{���©���:��~������������쑻��`R�{Ǩ���@��S�ڟ���li���R::n��t`�c�� �Tq����]���&k�Vʘô��ZYY1nsb�h�/�#��`>'k��+"ӿ���o�){[Ў�!<TH�s�����)W\W���n,�ݘW�=�V=H@��S2,��	� �<�L1���AKED�uu�u�����q2)D[V��O/L��t6����EG�J�j����{D�^��KJv�)w�L�0�4j3O޵�*��Y(S�{��;:���ז������6�6�B`��jk�z�vlD}*���#�-
Y�f�=C?@����uk� �\+�L��C4;�U�6`_���65|���!�w
��Q1w8��{(D�b�L�T���[�0LQv�� |�!e��5c6��t�4�5���yy=Q��Hyd�<�߭T^����7���5s��^p��|��D��kW<�:���p��UL��O��~����穽;7�C�D"m�\��J�E����d�ě��~z��L�4�ş�����ǌ�|�߈�SZ��yә ��Tb����@S��]�9�W�Rk��WU/0��4鉠pɕ�G�w�|�j��/��:(0���̚�qg�g��g�m7�a��X�%�5ƵĞ�ޔ�?i��&󨝡Lˏ�y�v�)�@r������5Sy*������<<�?���}�f�/��Z�����ξ.��;�@�?T���n������y
f�/�eW������g�m��K�C�>.++C���С����������ʸ��6%���d�t����P���jo=$�h���=F��X%_��1Q=~&����a�������k�d�`.6U�^d���ݎ�svt<������TESS��ݷX���+`bll���+e<K��ikw@J��\��G�@vddCj�+�Ϡ�g�Ev1�t^�"��j�ݨ.�Շׯ�AG��=MJ�(GT'�����>���s	�		����$n���`�+�3X^^���7\H8^�����,wQ��@�#:W����ݭ�<�;��\^�����ޓYz���J[�K].��B�Đ��/J5�L6i�.7O_����K8���Ŀ>;/"�J-a�A�}�Bz�ϴ����Ctt��W�u����=�A bl��ӂ!�]��@>�U���!A����)������1�}6{LZ:�'�i�a˵Hc/���B@x���g��<�e�W�d�V�}�n����_�E��ߌ�p���FAnL��!?�=1���$:.�#��^�{К[,�}bb�Drr2D<�$�fvv���t��HN��ڝ�||�R2ݻg�� |;6�t��7�fm�XF�쬀�nW������� X�o��c2j^qB=�sq��<Wa����������r��q[*jj�XXtoڙ�^�	G��%�%v�"�������>H�������+���5��MMi�~ yq8��dgg����±b�.jycc!�H|�.�D��{�d]˗P�@
**�4y��s��^f�F����J�v�i�s�U��Ó7Ng.8�SVV�+F`ejzA��%e�0��b�d���-,-�&&�d��/���H���� |,l
{�C����	��wM��?���tO���6E�]��	c����O����V����O$��~k(-z�[÷�e�	�y;��o7uD�[�=b��fV�<�'P�B�Y�Q8��������������ń��/ttt|����.&{��,.���xT�~(�}G��}!�*G�Z;���)*�d7>a��oĕ��E���̻*?��P%G2[� �-ZP1��}t��E�I�A�D�-�Ʌ���#������d�=�aO\�aXX��̔O�^��ȫ���^	����;�NM�*�`�r�n�gd譴&$����)"MAV9Y~�� ��_��"-�����\�<�ڂ�a)hz��)�LFG���SDFN��sDD�ĸ�qEg�V�թ�隁 >}����w��<o<�������z�������6sPt\���$��X�剠=��L��_�jt�>Ä�K�;s�L���d�,lXEʃ���E6��uu����M�#�[�����L }J#^���8�rkhA�ð�N� �z?[�q���

f����5��o�?�:�se�kj�b)O)�I'����$�jӹ����J�[���D-��>)��7�#����t��&?F�ۭ��r�9����W;���q�������,r� �9����skFx��I���/��5,M�
���LO����ֿ�Y������� 9Y٧���)���T [*՛_@@4�!�p��T:rĜڥ�诗�)!?r���VVBo��F uAt v~f���E|�^MZ��3>o2��8	wx�P�腀�]؇^t��$���l��5��8�dť��@||��ܻ�x��w�2����h�����ݳ��J���[�5�z''ol��0K��|t���jˆ���ٌ�ޚ���#;���1�SS��q��ZG�3�**v����nn����̨D:�Y?�ևd����0��\-D��]�#�f��\K����XU%rcC��$.G_Qe��	�_����m}��5^n��E�xo6���G�Ch���z���Գ�M���::;�_<M����7JԬAz�ZAa[jZZ)�D�ڜ;������heȆ�mш�+��C�.��m���fF� �k��'������ͨ��sX�7�5�y���߾��vC���O,�0ͼ��:L��\�q?7�!�H��������6��:��5��J$t��W�ъA���F�r���o�v9�����J$&0n_IU��ř�!�'���LH[�D�XI�|ӦR�Tb�{yUU����jH�e4���*�tJ��qb|�
��WS.n�=59�T���9C+$��� |��a?�`
0 �D$�[u�-�2���P��Ӎ�Oʹ2ܷ�	�korj٥	8�~�bOb�^�����N��j��G��J>�%�����ڇ�w�UgeYC��ޝx:]C{����nU�n,<Y4��'x��llc���,,�@�>!MHެ�����r� ���͑�ԓ����岪�� �@�����n���Z�;I�]td��1��ە��8��i�����埓�Ew���3WH�_?F��)z
�~��������G��
��/xB�u�n̿�w޿m!�W�����)馼/@/���ܕꔚ��A7�+\ve�Z��C$yAډ�cJq;l$��3%*=G73�;��"� �	�jɐ��)�����#��tB�����l��]s?kj�	d� �A�W�N��,`��D�@�E����Vk��p�"���I�7T�WL��?U[��t�����=����'�v=��u�|��>`�9�H+{�z��^G����Js�4Nt�څcF�>�z�x@�3@����h���!y��v�����o ^Ss���QAQq:t�y�y���
��:~nYi.|`&d�E��BC1���J7{{cF7u�8��b�yA$\��G����,�6���Y^F@���<r:���(s	�����5)��,҇������Nn�k����2���V`H!e`�w�И
}7a��1�f�Sp##6VV=�O� ����|��,++nh���c@fQr��T��׮�G��i+�?��{V����i�t]���Jim��ٹ������7�9!~�RߠB6�ÚC��sO>޸��Ѧ���������z�({㶤{k�Xo:�6��7$��ܢ2�A����{O��$��-a9X�BJ��h;R:GwA�0������P3I3�x��rN�;��gf�7]g:A��`r���]J���_2\co�599�d$V�����Oo=_6��p�v�����/I�\޾��ƙo�jPaֳ��M��>pxG���d�\��1;��Х��ߜ�XN��\�066�;l\;XRY�bĹ֪�S���=wA*����W��oE�*3�}����r��4�$50#�o�Ĥ�z�/9 �c^�`Z�	ߙ�zQW�<�����RJII�0E�&���H����V�-z�O��L݀4ٱ6tt�j\����۠rf`�Zh~avP����K�pkg1�D<���~��ZQT���%���gYJ#�ޱ%Ŏ�o�j+rC�.n}��ME6lx���{�S�AV	�]-'�uSN��Oт�F��ԏ�)%d{�6t�a�	v���L%����'��)��C���r㢽�������s�4���KP��2�y��qE8���DF�Ȭ��^���w��?�V@r<P��`�*~c(��N���]�P�Ha���Z��ZG�i���u��l_[	�eb�0�D��c|ㅖ�E����Ś�L�
,�ȹ�Y Ƛ�"����p���q�s�"�g��!��cW���P��d-kC ҿgOk�D���������~~��IZ�Yu,`�v[�,1F������2�6�u�̟Ǖܻ��:��B\�Br��I�G��ϮW:�2�󖽽D8,,�Z�F!���׸n��+�i쁥�-�(Q��� }ĭ�4] �[���z�V�%w�Rː�Z��l\*����kᓱ��g����96�|�%����ŏ6X<�E���l�/�]-+sY��Z>oh�*O[φ���kR������ʪ����=�X32.���+�M��*ͫ�2+ޓΆI�ɤ����L�� Za��W�����f�10�P^�P���s�E�U����ʔ�e~!���a�Ɯ�!���k��9g���̔��5Ct�(��Ҹ ���[Nf��=_��Í�6]Q�"���#UC�huMv%e��(�Q��-���Y�w>*�B����Srs�C͢N^�:�?VfY�g6cX�����=7w����Ϳ��F�
�K���ۂE��rso�������77�k��L��1����L)��]�h��7�C��o�ml�7����O��p���9�fiQb����v�.ګ�`"�h7�}�&�&z����75S��<:�a����>�7[�����|�5Kˍ���Z�m�S>�.2� 5t7ĻU�������\f��K:v�chu\P@�}MC@>���׶��dz�����0�+����+gV	��0�W�mҸC��Nx��]�^�����.��^&�u�Ndۍ��b�8�@t/;*"� B@����i��g�b�=u�w2P�N�Wl�tK�\YQ[���DY'�S�rqp8c�v0 SR��v���&��gx���Rj;=6M��6�`��1#�0�q&j�F�rei4�Ce�C���(����Ak*�̦�Q�_�}��Z��C���6+���bî��%?�h���>+L�ܔO!i��Aw�s T�8��X)���_Dݚ��n��N���3S�!���:�hr�mr^���O2��͘6�,��~�X�y;Gkk5���3V�.Mt����z`�>f`�s���X7)}�^�	�4 =����P��)9T��gJ��U���֞�!�S��t	UCh�e�n*����E&���u���3ƝƋ����E}�a�j
ƶFi�߭�������V�f�Я;7`φ^I������wz�T�o���?�5_<�o��E/G&hΦE���G0�C��ֹ��e`^y�2K��":��q5�����\��:5�n�5�@��1/�wc�rr��_��q6���]+==R���{�ď[n��NMJJN����h�^=��<��2Ǳ������C{��q�}2�m�r-���ʦ���T٫�cHe�m�+w�k�0��#0���7n�)J���3�*���;8�F-"Ħs���r/o����hȭ��.����~N[w<���>a�6��)io��I2*%�C-�#4��w����l��j�@ ���-&{j{޳�[�qnra��bߘ|真��C�J�1�ƛOi!��7���F]\\D�q�W�)us�ҞI��;[��p-z��0�C}�D����IY@�����M疖�����8�2S���r��i��=��8�D }�T�פ U������;ZVV��\��se�:�A`����<�>�M�V$�-������"_*���}B�@Ƭ@�!�vG�$j:ySo�~j��q���ő��+�l��.��HOTe���+ �c�����aG���u�a%��u}����믕�S��B�DE7��I�'��.]
�pJ��A��r��$v��W�SqII�t~����/3@�[8�S |��0\�M��*|�n�J�cY���.�`�ii� �_^~�Xp�ā�5V]�ڰj����uto}�|y��[TjG��TZmm�>��U	,��ELh"aLV.�@29aD~�bX�`�b �]�6��e�:��P��y��ϕ0�@�ܜ��񮾚�ӻ�m�ҧ��{񌾝g76 �p�ڥ.s���;�ZfV�a����lR^^�����b��d�9C0��kj.��RK�K=��i�ZQ�����WKU�.��E��/$��LT��/��~"+�B��Z@/�8��[�JKKKM}K��㓟�^5���9�^�m���O����v���U��S폱G��ۻ��sF]S���4�4ݹ�.�Q(F2Zt��Op�%)�Xi��kf[й�v�E	�@�Rף�����ܫ�Y�C�=�u�N�1�
�K�4�AG.4-'�!�zN�88��?�dK�~Jȇ\\�Q�o��`���3>|�&n�����s"CxLsi�Do���`��E'ｉ�}�d;���|����	���J;�'�!*QG�l��������Հ���Fy�S;�uܧm� Ϙ�u�4��= R&��{�%�WF����&)ɫ������e韸��S�v��U���ң��. ��<��3p�x��5] �\�|�6��D�iiy�؅�mQ��wv��u�$��qT�K��A�q�%���?��y���08G�(SwZ믤����!@|���b1T�;?P3N��K��9��1��S܊C�xMmu�����
��q,J�5J��6��Ӛ��q��;q7�hGSN�r��&\��'���4��^&1ݵظ�v�y67#��r&�{�P�m����ڔ7u�u����l1Ցv�����C�.������1~�/�:$�*<�FY��d��k����g�v���>|���,V��<G���7�5& i�j��8�-�}��ݘ�Bc_����iŝ,������ݗT�}�0$����^<�Z�x �8Chp�0(Ez�9�,�h+�ZLzH,�fo���Z���;WVyP�����v`��#���R ��VK6]���w�0��u.�q���� 	oC`�{�f�$!������<���twOO"D��l'Q���c,��!��`[a�9�.���:�1ݘy�dB����&$���RrM7G\>�-��]�g���}��f�����x^�S�X�*���=lڷ�������d���ʚ�/$`BL� ��>��J��,1+>_av��l��זa�'S�?9 "�q�\�`�fk�A�z�Y��,/
�1��q��;�����UU/�	
���h<��4����6W�A�'|��]�D��`�7R�b��&h����x�L[n���g���j���]}�"�����*@7�����>���4��:�Jd7��n������
ћkl�젛z�Tk���i!۶�����K���;�x�U
��M�$����7.%��(J�C\�i�Fu�����c��%���܍nd�d��-���d�[�G�Ú�HOc�Ʉ1�R�>��jm�ҴB�	���Xp"�ԧ�Wt��r��Ҧ�A�����E=�E����9�d��������r|���$/���ri\0iH��{;��o������C4��<�Ǹ(gf�\����2��w��V�Q��
khr�6n� @J���k`���r'AX�@��I�9?�O�YZz)R|�w���Gx)Xt�'������(�$��E^�%"���[�U��9��[t+��F33c�:U�[潉}���ht϶5o�M�clB��4��_Z���}����kB�oO���O�-|�p�����y��l�{���}��@�6_�5rP�w"�5���99cl:֛���~Ϙo^�.o�T|�}J}R9-����g�R��G�:yԨ3M�XE^���s*��ey���l��s�M�=P�2(�/f�8H��ĭ�%��	0^� ����:���;��ew��˩����&��5�8h\��6#W������VC����La%�kgJn�+}hb��D���C332�<�'�~i�)��c�*e��(��=��X�^p�m��q�۱���5�� H+���>
W��V�O�������N&��}m�0|������4d��n`C�1����Ae.���q�2s:=�$ȭ�o�B�3�!r��3�w�A�,-R��Mpe��=�o�9���3ss���'�85ni�a
l�2��K�d��h�({[t����Ύ���E�@���^W�1�5������
�Y�by��rG;W��+$= �ܢ�XƩ��y�YX�x��죀zL&��U��͗_p����?�щ󀇰��q�\��<���������sv_h�t��>���,lP�q�D�S��8$���+���N��>x�;��A�AW{�]s��e����T���d��J�ߡ9��:�q�
�v|�����ƻ�A��S����6��Yw�:�ͦ���^  ڊ
|q�����׏291q�Ҏ����637'uJΊ�L}����F��ٿG�CW;� ��
�gE��P�V(���Wң���v@���	fffIN��كt!PV&���y{�-����2��`�
�3!��4z���!t%�r쟋IŶ2�5m�k˵�3�d~Y����yW�h������ҟ�h��F�sC3o�V��d4��5=�\�%Zsgٙ6���<O7|^��$�\�\F�(�d������d��Ø��O���~�T���}�f����Fx�};�����nP�D�@�M!v��s���/�kγ.��q�;��E�!��4��4�.�(���w9��'�Pҝ����#�s��<�:PL\�H,�A��L�o!��)ߺ�X��1����'g$�6�����M�g�%�wSb�'�~�V��o��
�u8�����lsj}�����G&�=��<A��-7G��`�ڗg(l^��.� .yqCa+}�y��q{�ν��ۿ-3$t�������A݌ǀ �V�;�K�ݭ~P�#��b~����w��_��,/��qQ�b�M2������<Ig^�Zp�`��lN2KZ�n�[�¤wf][��9��ZO��x�B=Qx�����q'��΀�hH���	P�Y����(�����Z-K������������;�*w%��TZ��m�u]�P��-�R��4�����i�����չc�k�ux~|]z�p�9p��۰����II���~y�����x#�5�e�v��qp#' �ε�*��`=<,\ȿu�2h�L'^���<um�^⋧� z���;b(�\��Xb(���?������S~�oqG�kٟ���:�+�˕�h�4��t�!�gȜ:�JYWCײ7�c��!t����D�8��uj���N�� �v���n�7�H�*;�U�0�� )ɮu�t�8	�_eG�bz%���S����㲣�N��|�B�b5e�ŏ�0���r�; jb����n��ә��Fe��
DY+6�ymϜ��	9���f�q`sD�I�u��AjzzO*�ȏG�`?~�����h���,J\P�Q4ں?�b;��&k	 kq��e�Ly,�Er���_	\��2)s�o2�����������_K�#�9�#�K���p���S���j$�<�y�:|�*���9KP��� �h���vU��׮ᓚkC�Q�?���J t������1�W.r]�^i�!B��oD$�ġC�\��Ls�T�n��U�e���� ��fN��E�V^�j�D��~�5V���&�����oZM4c����+A��>��)*Y����Ό&��0�X�V# A��|w�3�%@��Ж37��Iڂ�3o�֞�����y��Y�k�-�ί�P}rle�3O5|	����u���9끭,J� 8}}u���9G��(4.��!Ϥe�(7����?���J��Z��芠����:{����0�A`7�؉��B�Vu���H�Ufe��հ\��24s�;�xv�j�������o�)M�� \��]e.D�Y���,�Nf�iiğ?on����s:;��Ԕ�+�ڿ��x��������]��S�//�s���rϟ]�$��ӕ�����rU���	�4�ي�G��--��X��be����z�w�����o�fΧc�J��@�x /�$v:R�
�-l^��Ҡ{�b"v�!3�����o�����mm=��$6lW-YU*�Lh��ts�� �5`(�8㤩9��Z���@�}��� 
�Ʒ�A��!���wa�-�4�WwG�����]��g�7�Vڟgi�����!������!3C�!�ˡM]sb�^;�o17f�m���(�5Ue��V����V�n.�v@޼>�!}U�J�[Tw����G�Ywh�����4GF$yB�V����C9�aa� ���X�ΑN�^k���F��+�L+]��-���<���T��F�.�h ��|��>ey��1�ԑ#;���5U�3-K��cϵHߒރ��A���Y�'���++-�H�C���3M�C��ۏ̪�qO�����
a����m�7^݁Ef"SYE�y�B�O��i��ο/�X��5�?��c�wÚ�-58�Z�B��E�t��`Q�
�vʗ���N��fo�\{����ǆb�! $���D1��,�.r@a��A��d�|�zUI�[�Z����^����1���[�{�K�5�������]���A0=����f�W��J�3�I��ip�-�]�.���d�RZ�R��j���FQ��k���u��ČP��T%K����z��\�DS�h�-�ٛk1??w��Ѵۊ�>��AyT*���M����S�����<5N��e6�y�w��ø��'OF�+�^��b?
�K�I9}}�I���=��/H�w���a�Af�"A���JlWzcB�1�D5�|�0m���(c�gc��
�]��.̟�����Sc�ĳJ���F�)tE��5����|m_�z�k�.Ձ�#{.�zVVZ}����2)Z�M:��؆�'��|)/��[sdRY���9H�U�h��uX��\�B�(�s֫=r^�@�Hs���0����_��α5퍤->��/4��){���s��c���x��C��Z�#4����Z��'��)�*��sd4�]� M �ǋ��X?"��'5p��.�������.�[$퇒ILw��X��U���Z�\�\W���0^�J�_<"�D�fr3ƾ,�̢�����]����� �{ᅬjӣ������������11)~�)���v[d�S@��|�pXj,������V�6��Ufwth��C�N���N�����U98(#���a���6^6t%��c�&
��$wvv�&/�i��>8��ЛkJ��&{�f  ���n������Ǭ�h�����ކF��Y	�Rf0e5�^���J=�����Hk�ng\r������my�M�'����B_"���B���J�⇗/Q�i�p�Z,�FC����Ds� M�U�C��0��$�������VW?��R7��W����Ӄ����M;c� �%��i�5�m��ݞ������p������a����Ԇ�����@�y#~<n;��񀌡��b�R?���M��I��8ŸS�l�J�cP�]ӓ��(k����[ɹ���^�@}�~��L�<2��.�%v[��ac�+���s�ݺm��D]G�J7��ס��C�bMJ��^�2�	��������5�e�����d\�y���(=?$"�g�9Y9��TD����}<_���W��r�J3I�j�ݭ��A�'''W��i��{�T�UMi��*G�`��n�����4�Y������ik�	��._

���u@�������m��\~NMi�����d��<q��tq�f��A�jN��n�uJ�z����� ��O�����7N
Ƞ�Zs�x�~;WsI��yq�����>�)��r���������v%	�ր*	\����M���֞�Y�Q==��"}	��r�'3���J�nd�4}�jC��q��0<�f"�D�A���m\��rǿD��� 99vv2)g�H�rg�$�Ҷ>ał�`q��z�P�Y?�+(tO:-�⣭�&مď�y3I��d#�D�c-�^)������l+Ã��}�ωce��vn����]�o�����t�����n]T!��Ҹh�9��kg�~��6~V M~���N�[<���c�0�����h��e�����(u3�(��������������([�ͨfT���Ie�[������R�m���l����!��n �ԅZ��*�F��!��\ߢ�������g�a.E@CӤ�>S��xJ��Q��nk�5�"��]z*��QQ�wƶ���V����?ɸ�q�6��u��[�P��8} Q<��Hգyx�;������j7F�Fe�#G� H�
�v�~"���J���Ξ��
�>�����f\5N�;�0�Q��V��W�{�A���Y�BY}�\��ˢ�����g�y�W�ä$c�NP��Dp���[�0�̏��ԋ%��"�
�7`��ϲa՛Z�Qsr2
9��p��P�A���;(�9�h7��[���~�n�Z�1�]���^av�_P���X��/�6T��.4srw�\�;B�3'�3@���y`��- U{z���ڭ�뎁PI�y�)����\P��c��3��RJ��J�g�^$!�D�ؓ�iugD>~���dT$*Ǥ�+�5���=���b<�qnrtTz�Fߺo-6cg�����10A�R�U\"5 �k
>�/���p�����$�M��\{�p�am����P!���/�xoo�}̷T���
�5`$�L����7��C�w�2D�ls��)��Vq#�!!�>
���_jY�{/K�ڙ*6΅	߰z���<�j��61x�Z�㌧֍�ي�Sb��޾��V��d�TԄ���֩M�b�������\��h�.|uǺ�L�κ}u&{�y�����[Ǵ�`C'��PG��c2���2Vӟ��$�ס��}�P��lǙ�q�u�E�c�zn2V����ܱc���IvʁMB�E=>>>�
���:.��q#�a�gM�=֪=�����o�B&t0]Gj��^��0��*�U������/0������!�lSB0D���$�!�
�	��CV/K�U>��r��ZL�st�Io�Q���C��ds@DE���N4���|D�1�5��߆��`���
5۴�<�����k�M-A��Q��A��a��:%E�֮;� Fǹ#�z_<�TrZ�w����e#�>�����l�㲓���7Q(j�zg;����(��7��C�X�	���1�����Nv#�n���7�rF���^��"مn��h��B!�r)�\?���������\�Ʒ[�^C���m]7L�,�Gd������� x����8v�C�9\�k�����	����ǐ�Z����9�碷v��q�l�֣u� �y��Um3�)��b 0��-U�U�4�G���p��ZV�@$�H��� f��Oy�|[�X؃�.=��}�m:������.0{l�.�˥������c���d�36�:�1�-]R���b�Je�`�z܌�`k6��7N�)��^�э�������Oh��� i�:c�Z5: �k�4N[�)�W`0*"c��L��˗*\�4ow`�k�)+�����s���}zB��I����	w�y��|^N��7R��o��,k� ��U�tqq�a2	�Vh\�p������}������m�D|}����R��.^�0��n.nn���v��u��i?S^�8�G<����w�R'�_`:s��a~~����?`eE�<��UD�"�" ��OP|�����69vv͉.�aQ:�蛘\���F�ȃ�2K�S�����%jLd������C�0���s�r&�@f[:+`�w�f�=��;7��9m(��|Tʨ8c�W�x�~.�4�s�[� 7�~���>���?|Bt*.�8�U��' ���/7�
�㕠��7J̋�ኚ��A80̥�	�:�②,��4�[Xs��<3�~7���>W��B� ͝;�t��88-����+�p\�e#�g�B��Aki�F��㘃=s�7�QbQ	i������Dͱ�y�[ֳ�8�At���KF�K�Ҳ�=r$[���M���~��k<�F��1*q�2��c�n��ݳ uԙ�[��w�:�`g�I[Gg�'��%X�(�O��W�i���M-ޝ� �Xt�W��K�����WP]܄�c@x �#qפ<�����]W�p�Q���cF!@���5�.| @"Q�T.ϘY].-��X�'�,q���1�5�T�]�anF�;��_�f��Q�Qz&)�w&n����&��kzl��[�8��w෕3M������3���06�ç��f�K�b�B�B���P|�N���Rƅ��۝
`��v������ �=�	��:��j|c��߃.,^e�OP|����Y�&��M�S�!�.��H�B� ��>sB�ݎ�(m�?}c�%D�M��B/?K�5�}B�(2+΅�;�|j`�~x�qqٝ���u��!�f@��e�/���þp�;@�g0�-���4��/�[\�#4��x)�XѨ�؀�~�|�q)bz���ʹJ~����Sx�u�-ҟ�Y0]u��KK��\{y!Hbb茰����Ў̡�!�I��n(���#���B����'��`�:J�ŚW��}�0���9���#Gv�%��s�?A	/<$������qvsS��&�r��o�f`�T=�L�?s��0�1x�b��~�Z`%�������hJ�K)��v��5]����u?��(@��.?�,ݽ���!P,�Δ\Ђ�7��@'2��SÇz
����	T�� �~�����[�\��k��'���X,�?Q�"Y�L8�7 �p���Vp�LD3��f��>9<�9�;��4W��#�L)�Qƕ��1�j��-�k���4s��#���L�2�����֌"*c#
�q#�$X�Qy��q�0;
��55�M\�,��q�����M��L�������;{5�D1����ʨ�	���H$�!�TNO��X�2�����oYZ`YJ��E�k���qS,Q�x�tB��=...�bX�vZ�)�%	Bo-hƑ��ҫ]^t�gU��k��\�/���A���HT��\��\qu�Z���a>�J��I�.p牡X�ҕ�ݔ��o9�RYyq�ѷ�k�H@�_&A�+H�$�eV
-,r�;�"�i0Op����� .�����s,K� :�f;�E�<��II�PNٕ��I��WĆc!@kڒ}.��=^�8��y<�x��Q]�\�E��dŏ>[�/n$_�;���b���K�z��z���Gd=d�_3�&�
�eR�>�@������`�ް'��?���B�Ƭ�2�X�����ፆ>ˌ�����յj��u��kԧ�

�¨4��q��	��^���p$�r��<���~�J�!���r��IT�ރ���OF;�ŸЌ�b�*������Nˤ��d.I+��c���U/��f�3�2s	�ڨ�Ь���"�8ϛ����{��@~M�֩+r`� 3BQjFR�Ad+�0����2��`�?R�=�-���V� "X,777:����GT�7�x���h�,�p�ϕ|�quA/K�P�.�Ԣ���QQ:�_���K�&]�|��n�W����=X���$�1�ƘC��Ы�F�p�y�� �.��E��9fm����B����yfI�b�U0,Z$�=_OT,S�10�,�p} �_=gUE48�Mx�~�Pnn6\V_<ѫ3����P�v�p���G�C��!!F��S8�@/�CȰ��-�NT��zL���1�`fON���$������XA��_8d������u	���y��f�9�]#S��v���_e�!ͼ���0��N�8u y��w�j��CѸ��r>�D|�E%&�}zFy&]A��Ȳt���K�ܸ�`x��K_��2p�jlKKH�s7��ǻ���^9[���cm(└�aP:��C��E�.��Z[�����������j�����&�P�o��t:'�ꤨ,�RT
5!kG!Ր4��![�]�%ˉP�J��,�ݠ��11֡���`01��~����_�N�>��<�}_�u]�������ۗ�((8�δw,4=�.��=��$�\|y{g�e����a�O���0c{�%�x�,F�Ըs$��E���R�l��W�Q����r��������O-��|�����zi��\�ḟϟZ�{A�˵J�.���ik������s���@E�n@gS�t�`t�@!X� ����Ǜ�C�y��⪗[�)�feC�-S�j܏홥.}=5�D�rd�:�͛����_7�;R�)���%u��Ⱦ�~����pW����R�"�<sl�`{:�M�����WV<O7 r+�vt;�̨p�|r{AW���V~��SSץe���־P=>,���ޞ�5<-���-OR](�f6-���۷����	�R_�1{�X��7��_nJ5^�>�Ӯ���J��<�3�+������<#�evzl7��@W�69�G���70p:F������e����Z��h�����1����rr�룭ee'�O���SPg�ٯ��

f����������w��XwQWA����|�FK�6�%=���B�F9�Q���{�[�,#�Y]�o@ա ��=~���D�/>���V�����]R"�����$�v�;,~�|�Xh��3t���6��i�'A�fG�g�K������sↂ٪<I�%QI��Q���V<�����Cm�4�\t�� �[��i���R�tH MW�WB���5�C�j��.|ln֌m�.r���8jh$^����ء���ľ}�RS>����S�G�e�L&�������)
�*X�'��w��f��)Hצ���j�������4N�c9�[��xI�!4���b��,L;��u�ķ+�/�?z�YN�۳����pp���VffG�u�Msc[�t1GG��%e=�����a�U�p�&�m�̭Z��õȘP)�:���9))	��?�,[����(�R-���fJ7.q�r��9ʸ��vv����m���1�����^[���Zt}�����pެ
eؚl+(�SW_�~8[�O~�������v�e������Z�~[qu��އ����K3�ns��?�u��b(���Ņ1���hsf雛��,f�v0����g!�j�"�k���###���ή�.��t����IMYy�C�_}s�����a:���	K������ݾ��a�_�md�#ި��Yd�Ht���8��_9���Y�y4m�T�~�&��J��x����(����w�;$�������=���[B�ޟ6����騘��`��zT}��61.�W�CrHV8q.׽��ͷ�\���=�`�-i��9X�dޢ2�A�|!��(A�R���Ɓ��Wx5p���npf�N�pi�:1��?�z��4�[;<�YO���E��Ix��xD`���S�p��kGr��|�2|�x�Kk��77��n�*���5����NjN��P�/�	�<�4&������u_�^��.6��w�[YXD���wvG75e߽���K��^S`ЕV��a_�����z�����l���@ʰ���6-]*<�@�-�y����� �>�6��|�H�R��iK˘��8��	(�2���٬�q5�[�'--���"s*��|���e�Q���[;?_�����G�~�C����P�Z��yʱOK?'c�Ύ�e��4�طhƔ��o���R��Pz�c�$��Q�W�� bup�a���2�C�5Y�)r.���崲��
boedd<c�=�5���7�v�Z�А:&,�Mv,���~HRrr����Ǐ���-NmF���h�[�Q�=���r����Cb`���!�)���4��@�q������RY�
�M�n�%8h�n|�eB��sϘ\�����p�.�f|2�tjV������m/Y)�>��g_������cr���K��_O^{�89��oK3�M��܌��6�t{����T�E�����X��|in8�l-�"k������D�zW�3���
7�#!w�،gg�ڶm۬���{u%kQ���R��y�����Z	�?�lYDӂZ��Eg��H�����^����|]6�hhd��=��T��\_U��Ko�Z[�����w��e֣tg�,��|ƹ4�|�e۞"�����ߠ�V�雖�qȉM� �0�:�N$PW8 ��h�L,��ޕ�{�Ïa��:0�f�!R���Ac���Xܥ�
ڭqNDЇE�gV��F�@�ViQ�W	���0���t5.tuN?�JN��@�XC��Y���^׎��2,]������V3�����d��'IrǏo70�� ���[M�R8�����l��ƺ<L�-�WU��P��)��			��+6s��D�IL�%����;�E�=(&��N���>���dCqS/s�����J�?c��sP����֣T:;������������hY���Ϫ����0���Z1ˢ"##o@�y�єS�{rt˖-��L�SU�]^��8���XUmWvJ$q�Hsw��w����2,�Ѕ3�_�t�a�yF�7��7pc�r}���l�zuXfff�
D{zzt���_8�X\�rNw����Q�|=S�z�� �d�d)>R���5���֜V�����k�S���ựE�J�<��*O`��cTaٳ�P�x%�V<�9?�s�+�[B��P��c�j��$�ÞL�8����2:5�B�l��V��k��Uה:KO��?dv�����`�[	^���E��;37�M|���g��[��p/Ǡ�6�������+պ_��2�s�#��e�G@�rG��a�.�AQz�;�A�,c�˩��=J�o[���=Z�һ�t�@�inn��X�RQ^��0s�<�Pl.-���
�D��ϗ��G^^�ܒ�B�
��7|�S.Ek����ˢ����������I&�)�^��aw�SL�Qi	)��C�Wܥ������j.�	��#��
��a�{��ֲ�5n�w���=5���^ӟr�'ME�\�"8}AJ�Q��=E�gr.Ͼ���7�{Esz�L�˾�	�~�1��|���|�C�A�N���ȗ���zs7O\7fT��MO_f�A��sK�烊�V�����Oɖ<Z>H)��TMQ�H�25L���p�L�� ������ĪP�+~s�`ƫ+�g^vwuE�R�lk��R*�� ��B��w*A�����$�5���.�>��� �v��s���e9i)K�`�ҍR�08k�2�������-�3����TmV)+�B/0�, �Ɖ� ����rn��l�0�Eƪ�I&��!���/��N}?�O�9�L���V�4���)a�2*T��*�Lf�����C>��kв���]̡Ξ�)�㣇ɉħ�q�'M�iqd��xƩ��L�j�Rǧy�������.?��fm�*�F�W��p�,�~Y��,#�J]_�\nt4��֒rPjh]�2��΢l&���1xi�f%�(h��w�GHY�T�>�x����2x�\ӂ�2f����n�5���ӟ�j�/.yr���T"IoY%��T��\lU���k�rD�a�N瞺Ky[����Њ����2G�S��p��[@V���cJ�-�B�-{K܃����"�A��}�`��՗`�"������9��p����|�����ԪR߾��O��b~wѽ2�g�ީϕ�+�y��uW�*rN���jf���ܣf��@7�|h�2�:�m��Յ�*��Xڂ�k���,��#�RO�H<��*�k���9_:F�O�3��)�s*����=kI���*(آ���أx�����W	A�QI>�����L��osCc�즞=ل���3�VG�7��I#�=��;�TD�2���!ђv�����XC����/�L�s �a����\���(����s�jn�w������@b��`]$sr���I�#���6�/<�COZ��X��z�������e��B[�;�@�2G�=K�2�[��K�SaÚ� �~J%���a�c�lq���C���ma) w��5���<��p(3�e����=v@k�"�Ƈ����82$Z�h��	m��e���-[Z�1��L]�H$Yؿ[�(����˟kn2����j\�A�����c���LA�F��m/���'��Ř]����D��s�'m4���z7X3���a���[AnچZNY󷵎�C���y��Է3_
������-b^�=YM����y�:{�!_��b���ӜRN�mW\Y������f`8G���2g�e���=	0����9%�)�O��LHS�T.����fw�ݐ����m����q��-� �GOY�,�ฟ��HV_6�b��N撓���e�Db���@�<v?�����{��i @>"1H�XD���qֱ�̭������C�f���e�\)0�K2���_�4$�I�W�xE��ѹ�)�֛B�ۘ �M�����nT3�͸�����2�K��?����-G4��b�`�SNqUK*w)�v�dh�ق�T���6��C�u����*`#X�DhEn��E5��O���aҞ9kP�Tql���bs!V�v��L��f_�	ij�0�|��d�j����* ��N�����6u� Z�^�U
�ۜ�rg��ԡ�%�'�	�8�Gų�����&���.` K����H.���TR*9�[p��MLMá3�b��R�u��@���$~��N֧�ݽ��a��o;��]4s ����zCS���qw���<���v��_N3c%@_뾸�,�OD��b��<d�%|�Z�):T�v�p��<�߼\��B��>7����j�CP��{��� "q��Gԡ�������O�×b ��_G��Hj禞h<r�b��5W��7jj�3)� YasT�n'���[ ��T�$�7�H�J�`o)[N����2(=:�C��T �o�t�|�_vhµ�m��r�zL�_�It�����2YdL���kC\#&�l��9�lOm�*L����^ ��dr��@�6��nr�I]�a#��TJ�\̣���M�l���kn��v��}�O`?�n4�.Z�C�|�i���+���>th��� =���[���mFSa��m��b�ZEg\������"�*���� �F*�ڷo�$�t���ڛ|��7�d��������<"'7ݩvwQS9/��i�&H���7o>CH3�K笡s�|���Oc�\��ي�x�߈�n��SZ^�G��On;�I$��B�e��{`�}u@��+k����֣z�ia���-_�0�����D��8Gr0,�e�,NB�ի仱�z�1�:�?:::PrZ�*�҇o���;xh5 �Q,)K�c��y$�K��y��α����H �|���;i��=�֎8�<�u�\�>~7��r�:@a��Ī�Lt)<�+�x���~� -<E��� �R������byH�f�}��Y�|�C��I�xQ��Y�J���4�+�,i$����S
K���S�W��oa�⊣�j(�&#騸=���O+�6z�2�wbJJ$�!Ã�:`�� �H`۾�-����хpD	����1+�4�M�N���2O����u��g�`v!�.��).��ۚ,�>�>�`��򱱱�|7�V�$#K Gndr$Q���s7��b�r��x��i]*�Je7]I��E�x�w�I}�Wz�r:15�#)�M]�������13wF��p`=Г��3�i�R2J�1S�¿�Bר����3���B�u����y�o�P5'L⫂"��m���]�,��@]���0����چQȭ��m&�v���!U�!I�f��`%1ϛ�� �E,�wמ�c��WeK7�\{:vba��v �yq;{ج���?�li��c9�u'� ��7B�c�I=���Y�dO��������z��\s���I�Oʻ��?Z�K��(74����k��T�Qn>�}�Br�aXL6C�����|
&�3��s��;3��u�}2P���q":=��v�Q^V��KKK}���,g�H~>�Wu}b{�v�Um
zڷ�	= ���~łf�녮}ŉ�Q�[;L����Id�ʞ&�9?rNe��ɮ��zG ત$�)8�F.�K��R�LAO����3��h�ݦ���#ebH`�����"����8z��K��:���z�G{V&a��	XCG���3ؑ��Z�.�.�4˱�è+��0��M��������v..j���ٓ/K�MU�}S5�[1_���+�W�#����%K�C;OD֘�#���m��0P��]���!��a�D�m��;�`�ı^8�T�¼,B�}=��T䕖����S;�r����

_����\�F�x�� �Db��-�h��ύ�&�/�{*��O'w��+�Qp�+��ܽkT'�!t6�57߆a�?�n�	zMM����)+<��s%��zx���{�0d�=���Ѹ�M�!QM:�+H�Z�����H�=B�l�ɧ���C1��Q3��*�>;Zjll�C��~��JA3�$�U�B�E��o�儭�#Z����x>_��aAg��+��5�<��c###K��T6�
iа�U�b���#����_}���s�OvO��)���>����)��Q��xC����B�PŹ��ԎLIS ���y�>���i��D	�P��/����t���Z�2b u.�mx+���Yl��ɰ����9��C�o{��.��
I��j��kj���<�Z�WQx2%\,�cm��h́���Ka]�jʽ��� 6}A���0�O�ݠ���UZ��[�B��=ox����vQd���� �W"P��h3�9@�%=�T�#����0C>���Ta�|�d��^j�M}�r���Y�9�899a��Ә��F�1�X
��`�,��,08j�e���PV*n	E�5;kh^��� ��U"�j�权�i�f�!;�)����d!TH_P3���<o[D ��r�-�F�FTH6泲��f�� �~�x�)d9h���9i���M-նe�ݓ�0c�9%�C[�b��~z<�9�3$��G����+��J�*��{XB����"<�hg����7��p�֜��yR�2"�,�� �u� |�`��y����j���g$�%LF�����3��T�RUZBf�U���l@^�����?�^2w���$tK]������T��5�������(Rهr��S���f��$�J|s�^�jtv '
º�x=�I���"�Vh���|~llj:�t[���X,�6=V�Óo8)�^8zKN��s�$u*��1�xE�:$�G}�A�nBЏy�ׯ_o6ʵ�ʗ����#������̊1��caX�"K���̈�4���n�=vl�}Kjtfff�A�I֞bW���X4��c�[#r7 \C�V\�,A��XZ�,��Lj��
Z덠��ĭ��{���8:2���y�b&�8�r��_ϣ�t�� C��ya��Q����6|�y�Z��h�ژ�J�j�E�@X!Ơ�<&�~��VӜ|*Vc����V�^� �Q�YN�·cV&O^�P��~�s���IY4�?[؊��h_��v|�'ߍ�,:-�m�oIݐ8ӴY?:�20 ���fC�7��ֆo��+e�`��ڮ'+y)M����T�
����/n�S�x�x��	u�s�E7��+�o�)sH���!�����9tfu~�C�����$x�fc����jV|�ba��M���5����I7��9�4�� s:I���C�S�rH�N�ޖ��o߾��"K}E�\^�>Q$t�v��f���b�(�~-���;]}A+e���0��KE��*r�:��y/�]}J���R�2��6k(����������L���R���v������dȰ���w��[�l��z���R�.E��)���o6,���a9,��7��B$@���S�uN�eW�5Fqq[Щ��W����� #�\�<����^��ȅ_�Nf�*�z&����8j߬�ډO�*Bf )}c���˧T���`�4����XaKٱe�"���J�����8�R���oR������;�p�	��)�mԕ�L|͗����M��������n�p1���-F��s�[w=���([x�5�O'F">>~�s&��B�2���5��F����GPS��AW|��C�&[�Ғ��1�� ��QdmAA:�U35��4�`�Mi�v!�`�m�t:=̙����B�oN�W���A6��5P2��W��7��ʨ�8�J)	�7��qO48I�?T�6�Ec�hcc����G4��XDh�UB'�h+�3��ERw%FW�?# :p��e��
l���VM��;dGd���i\���"�����BM�!��<�ui�4�s5���H茀'p3���j@;��$�_44��y<L���cͻ�I�<ͫ��]zْ� �D:ج��n���P�����<#�V�L��y�V���q��?ʓ��v���]Ͳ x;x��bL:O�4�=��Q��crr�3tS�n߮E��$h�Tx�q��?���ؒ(>�	�HRH/o2�c~��@v�T�4oA���H\'���^	��!�]H����CbKx��4x�si� �N� & ���W��6� Fwz�����ox!�&F�!�BO;�8��: mU��7Qh=Fʖ��H&#�����P�Ԍt������1�W���V�$���|��s(YX���ί"cf*��5t/h7:x���E䅈�16�.#�S���A-̙^J�>���Lf9%�=Üa袣��>�45Q*�(:�g/QW��0q _��M(P[`�1�����
7�hr'�Zy1ncq�}���N�u�OCCZ@�� '9����^�ɕR�Ţ���5��+S�'�ƁS-�4��ҭ�b��9���IJ�7_Ns ��_����.�Bi׉e̡�)֪���f�y�&���^�L�@(�̃�e#[��P�fr��	��"y b�k�f�_��eY����嘬��
�Z�4N%�������M�����m��vq�CZ�7z�,��I ԠS��Lt�-f'qH�*�ů%ڕ��~���UC;��G;�z���9�rj@�rf_8�= �f�G���A�Xc�<𨁽��ކɛ�/l֋��ފ�f�?��&gp�ig+�\9P:1hah�5;�=��a�#"kdFŇ<u6���J���&S�SBvb����/�XRv$%�,��ma����5@O��������\4̥��Kۙ�T3h��9]]o��E!o�d�-���"J�W����8����s��nʽǏK0�@#/��S(mIc��)�=M�7<��;��M���>��mz��P��?JI�RZ=�����h�H�N%7~=e���J]�UR��ۮ�V|Sq�3�T -C]�_s/��`�����o~K��ޮ�d��F�2y��b�*_ϛ@TNp��T|g���t��>0�a��ѶPK4F����O�@�%P˩�u��ϼ�Yӳ��~j��fP�~#h�5O)�A�T���n����i��}�YUt\\,��S��U-6D^���Q�8�9l�'�zQ�����h��0����l�/�a���|��R!�E:w�k�I�$���p���K��ߨ�	^�[����"�^t�O��nQ�:�B�A�!��+A:��)�Q�a��&;Í}���%��Qp�����&�B��;w_Z�0p#�7h���1���[$P?zb�$�X��k��5��e�sO�˥�2�`wQ_;O0������GS(�a<�t=ЍX�ޖ�b��c`e�)
<2�c�s�}�����Хu���o�ai�2Yq3��n�T�k���x_9��ߑ��]�Yn
� ܔtceF��w�=���M�͵��HZ��1�_��"]�V��KA��"P��,�^u����T����p.�*��$�S��St߽O2���K(�| ����u�@�I�����r�ѫS���HA�V��~zQ���C�Gmm�������^}�x-�8'��\�A{���z��۠�pG^���K�7�>|�l|����q�X�k�pE���*7w��5��&���d)�7�P�P��*�P1�M|����Fݘ��XR��j�z��9x�L��H�m�͈��sH�E�֠�"?5A.�r���̲�O^����04����c�S=E�x/p�D"t��vO���)�^�x��?��!څ�����wM$) K�q���ec&�����!��E^5;�����ҫ����?�t��B�o�������]�x�)2%��/64 ���3e|�	���A�����z1ϛ�GC�����##.=��G�����/b\{y�,?�`�\�,ggϰ���@����՗24׶��~K�s3���c�-��Ik�=XU����JMЬ3�B뻌���8��P�v�-w��<��]	�Ç)�Og�^8$�.�t�-�Q(*.��G��-����L�R�(NC���Z{{}9=I�����A;v�D����������s�J�/_�~�����h�J8��)?� ���������@��X'�W{������]��H]��`*�`�w;g���ƌ�/꿬����I��m�蔾������ݻ���-BL-p������X;5u�իW�����6u��F�Tȁ��pHe���
��D�B4��j�p����P�H瞲��ȪJ7���%��_�-/-�$�3E��"�* ̹��\geŶ�2S	t;���`l��7Ͻs�s�:Q5�q��-@��K��X�bYK���9vnmoo m?+˹�9�K�ڍ��bK�� V��s2V!1yD&�c�>�k]�N��5�x���ɬX�R^1�Z�F�������Zu�Q:3�	���^�~��T�nW!ڐ
�\���'�G6˹	��+�Zs3jg~�����[����+�͘܅�n<g61�6ta	��$����ccو�����.SB�p�!����:�ؐG ����h�L�S�W�����ܻwr+�30қ�lش3g��Q�o��H���B�~�7��hȏ@g��gdr�uO����h�kE�Q�+&t/���##�%~l�a�-X��e�*��6 ϰi3�Νhra�N����Wхc�>%wz�3�{�-�D`��jM�A�D��!�=�GBSD�%ٻI
�5��#����U�%��ڧ�*��]��#� I��� �%��Ӽ֧�A&i������Wβ���Y�>6�8�T�wuإ�s��?�l����>�D���ߛ�9��׎<a�Q��M�_����p;����۽��?;�(⢏�,ge�rTC�d�2�� ��*��꛷�p���sO/{~?���?"|��X4z3�ہ�
����m>3����?_�ϊ�yV��ܝ
.W����ꔃ)���:K���!e��Ȱ�Txw��^8̏ѹ�H�� &�<��c��D�B��I�J����Q@@��H)w�������X�EC��Œow��P��!�RjJ98[�n�Δ���П;�a���s�8~�:]��f�I�"�8�NH��ҝvr���BX^���� ֣����
�C�������j�E�tg~�G;ٞ62㐸$�������6H�v#]�82�)#�5Ac����Չꛎ���zE#���`4�"��(�`~��{I3��L�����~�ey.�{������-��7�m�\rڄ<).�G{Z�M�t#�k2�O�������eLUnWK�R]i�����MU�$ü��v��BS�ΝIݝ�S�᷿ߕstu�SpQ	&s2�]�^��s]z2�x�9sje�A��=���Mr�M�IB��M������
�.|�r�K}`+�S	=c��b^{�\����>|J�8tW$�GsP���Fv��z؍�]>�6�ٱ�ŧy1p�S3���K\�'.	�L��+GZ�ǣ�omTA���@�u+4͆�k�?�4Ìv	Y��j�/6 %���-#��|���J�}��V#l��R"����wd��[�{z�tzΔJ�b���
��{+H���c�9������^'�\��ܾ��QϤ,7�aC�]2w�N�';��/>B�Z�E�h_�N�w`Wa��NN+R��������E�'~ExSY���D8�� ���V���3�6ю�I)\�2��UA��?i{����	�m���6�^`��o��In�n��Qx���uQ�:��D����F�k��Đ�נ媓(tSe�'P���t��y/3��ր&@�(�;�_>��/�rrr"֗|��رa�����W�̋��{�tKWBRR�c�O���{n���9����V��PwO�U��;7�;�r^me�����ߏk�/�<��`����$�#|x�tc�u|<g���N��d�MJ�AȞ�	@-GN�����)� �pa�2t�_�^��"��'�,C��r�c��r���P���1UN)����u�^���\]�b?��("��]�hq4�B1���V��)�|V/p1��7�qP��Ι(~/��3��G��&�!frYJ5gn
d�;�6$��#�--U&$G�T���ff�f��K�B�EEF�U�l��~Kkt^�z��"��a�ֳ�i��Җ�4c%�Y.|���3ߧ(����Q�/}2��F;��:�\��
7z)��q�v]���?f���ţm���q��X\?������t��'�Vm��5l79�R��e���M��|z�&z��)��+����>S3/�1�Y�?&��R����gc�����,/X'ly�����f�#`yϮ[v�&��Fi��X�f@>B=��u;"��I�CP�I&s'0*��Qo�:ۙ����:2���^B��@*\��q���O�+���pn�F�W��
q�_��閗���**&f�U��Q����z�ZJ39�K�Ts�\`N�xȹ����b'���I�����LL�@ЪƓ�����2~���H���ZVU�BȎ3x��Hj���p���<C}3�X�E���ˢ��<cI+�K��D��6������i�;���ߚH�Q��ke�u����O8
*xX���	��cޅEEOu3�D�[G@նB3���޾�i�0�6d���
��+UyP�@u�D����'K"�N�O���U�i��	.7@IE�V����O�f�|��Q������!c.��5�1h�Es����$1v���Hl�e${�F�Yvq곲,T��d^*��vU)=镏�o�N�%�V	L�d2��# ��W����Q�τ� �i�>~�W:�����3�1�Q"�2W}���h.��Q:����ë?�%KiM��u/[����-[�Eƞ+�"E0�*W����B%��3Ϯ�KoIN���g(��t����?x���t�N\H$�m�Y8�Zdg5��q�\�^6=�_����XwL�C%Oǜ�s�rsp�Y�b?�8d	=QZx0���)���j8��/�~q�Ι���͢p���(�#k����W�*�Pt��v)��0>��Z�^�r,Bn��=(��=�_Rx����&��_1q
Ӊ	��T7Z��aip*q�t$���rv�0�砂}>�lX�����?.Y-.�H����z�'�B�	���Urhׯ��i�t�A�l�`Gw�?�꯶��I���V��'C*~я�Ȩ����?�qk�>�c���ۓ���l�5�D����������H�j���-��S�5�Y|�|�)�1�/�ʸ���o$���!��l�J�Y�_��M:WEW3���58yV4�X�q��������@4��3`O�`�׀P������� �
:12�-��5�:ѕ����)K]�;�k��!7_�ۤ-��k�˗uLx��U��u�^�;��ļ���d�)9v�=~�0�i��/_2퍝��M���g#x��(��4tc��f�u�F񈴽mD�v�gm�[Q��}��7���`�s�5(�LG89�?5��U��N������acɢ��k�[2]�i��PU�|G؆2"k?�,s\\��/���j)�Y��B���9����P�#U8����G���J7h���#��1 1�n�Ю�H%�Ĥ���!���ѡ7�dj�<p��J�Z;�s�qo��tb���i��_Me�/���e�ݔ�D��������+�h�Q"��T�i"I�IY^��_Ey�:3`��xD���T`NpU�ڑ9�[���̘虱�)T"�#a��k}�[b%�2<���{���`hVX��?|	��-�kO�&S�{�;S���~Vԍ�QMh�BT�̠8�X�g�G7��vVcmFj,i8 L�3p�	{�x~fpvq/n�ߤ�Z�z@HH��K�{���#3� ͏��k�{N�bA��S:mxbq�An1ɻ��)�αTV�.}�xU�*�l;��^�{�	�Z�ݱ�H�|䖛Q��Z��*���;��y�LJ�a|p�X�cEs��L�i�9�Q�֓�>�֚�}F�wtgH�[�!&ּ:s[�s+�_A����n�O	����Pȭ�d�����~��ʅ�OG�;�L��A�ڙ�`���_j|o^T\|Q�6�a��W�H���o�2����ATO!��5rg�)1�/?L��ib���z��k-�9��Kh>�	��&��Q��w���P��#���Yo���W�������RVl����Vh�X-�4���q�+ב��A��N/g-�mpz�5>]9r�>�F��i�M6PSxI����a��y��DED~�E2�s�a��Nc=�~�		<RWٲR3R%>���d���\�MD+ʾ�u2��$j暛�knް+x�%?Y�!1�����6;�q��c���w�T�gDl"
:��9KNMg�+4p.B<ƑiM���ͥ2w��UL��?Q8t#�_����*����6���!�����U�u����z�Դ�y�pAI��ݝb1s��Y{#W�4*�	�zjiXƏ�� l���)��e��az�˯��*8;��$m}XA�0�����*2)�!-�$.eF��q���L-|���wo�h�Y���%��A����&��\�]��í���t>1_���_^�ˍLL�������Pfo���/!&ځ&���D�����(1*��f���ڕЂK�x�U��G��3�q��o�	Pu02�ӗ�B���G����DFOs3s,,342�h���\�P�q;v{t��ه�j����]~HNh�+������^��G��`0��E��G*)��绰8�k�j�o����vI������qP�'�����䐩&D�e���37��By�L��@��ԙB�B{ky�����]��0�"qkB��[/3X�]�-T1����m�**���?�)B�m�l ⫟Q@no'�:��y^���rv�(Y���"���h�o���05�r<A|$ݨ�T����4������2���Y�mA�\z{��D�Aߏ��d���ޮ}����R��n�7U@C��� p��Z<��GF[5'3���k9@���L�R��Wa�������5g�N�����u�۪�6��gƚ�
FNW�&C��|[||l�V���L�np�G.y�V*�d _��Hx�g[ak�p:C��UNь�;!��/vrқ�_ p��8��`%T=�{u.xI�7�͕�͠CSf�V(�*�
�I��;��@~5)�V��ΌWg�Ţ�;"�;6�1�P}����P�3�o�}�^6I�1 �,��p�T�m�޼��Ј��� ψ���͔s{+9
u?Pl��L��8k��&.D���z3Q�w�3���j�3��N���64�scn�������j�Uq@v�U"c.-n�FX����+���}k}$�+�q`�\]�ſ��q��)ux�dT���}�D&�x*��+�w��^"{�����"���$�y1���)�e��|,�5C��l� ��_�{Ї==Y��x[ۈՇ)���z��|���#0F��٨6<P�ۗa��J�-`6�ҭc$BbH�YC�9��VV��o�wc�x,�,������O�9N�G.��m�꜇��G�ޫ|��� ~�� ��]�~�����7���k��������Ti�s�b�E��	��g�����H|h��IM��j��+��#�mޠ^���&��sb��+V��$"�R�uw}�O��X��+wwu�{��+��ۥ�H�~��.�]ۏZ���99�ҍ��s'�t�:�XR�|Bn�H�?(�f{{�����aJ4X��\�m�Y����Y�T�򾧟�֔j@�
é�Y�u®ً�ń������Qr~�����	n��Dl8s
�ܔ�EF���X%�f$����͹W�ޣu �촥Д �r,�P��!���^SKsprhs���9�JV�	���E��/�w��|��o�>�����	ݼ��§͋W�8�$��k>���!�]DJkw����z�a�۫�˦�M>h�?B$��6S8�	�TyV��G	��ߗ*�����J��o�`�zD�5��@���zb(�+φ=�}������G][�T�{�uM��N�@!{�F�׍a��99�����z_�^�g�rή���qx��K;ِ?z��emܥ�yU`hha$891�;�7T������"u�b�Sл4��mV��@/�%tE�[��]Z;B(��^�����_Gw�Ә��������e<��.U?ې[�靀2�ҳ��$m��,��p�o@��q\g,�U�q����l��,�e�]���ЃR���ǯ��?8c�$�Tq�_yU|6b��K���4"&�S<d��s']��9I��{a�mxA��u(��t�3�IVu�Wb�/Mm8c �dw6���/[��A�o�\����1i8$vZ	���T�r�[��j�,h�|Y!ˏ��Mꄡŷ(�N��L6�J��/�T���s*G�Q;@0 @Kj��o%��x@�Yz�	�����}-lu�]b�Ui�[��Gaq�w�H����љ�%�lH8ʶ�OrPJ�p��x	�6�|�:�4��8�!��zkڧJIq�:�r��'TT�q����f�a0��ݏ��8۫{u�lv�2��i/Oz,=�������T���Ф{|�%�z� �j���nVk�cն_��~&�ދ����l��W�[ �)���4�1��V��6��Y��)�k�r���3��-"��|R_����aa~,�7)�	�Ώ��m�I��#��v��I.p�ĉ�]�S@��kmZ!��?g��ӹ���^F��,����]��uRJ*&��(?K/i\�3H�#��M�u�_�EK�ZG�p�HÞ��Ƭ�Lf��s���B8��_x�NH(lSpo��0���o��be�!������Ew��֛fi�O><�\�J(�㶷�z��.��+��8�!Cdu�.��&��ۮ�G%�=�m>6+}4�B��.��R{�C��
�:�$G�/8�dw���&���~a��^���]���\�ȝ�j[�7��Y�O\��@�/f?���lk��m��}�3y1m4�SH�X�Ԡ�ڮ ����MQ�����+.��3��:�A�I�[�W��>�󭤆~���3T]G��Y/\��]�w��^s:����iOq��Ch���^���w��O�4�S:��x�k�~l�?�
T�'4
�>�|�Y��7-�!��q��\�8ipN����Us�m�c&��ܺ ccc�!!zt�;S��na6��-N�7���3(�U��>g�jao��1>�����r!�fuɟ..�U^=�k�/�s����|���G\6�?����W��ЇuC�#R��G|�-	��S.�/�*��Sl,\���1\�d���"&O��>�F>����[�5���ĕ������==���$�;�4�7}K�k�^�P�NP�)�b���$~�n�͐C��}Ƞnۓ��o m��|��jϭ��#k��gf��XK�г���|稤5Xy���'��kg��6�9�E|��*�#�:}�(5���U�YG��W3��+��nޚ�˝�!p���1z��
#��jj" a���S�f$O�̩����$�Z��&B?ޖL�>��6�Ρ1��<��k>�J���E�2h�p�@�1��� ��'���mU.�e�Y�A��ۛ*���J7��$@m���DCcm��>K[]\�q-��p)� Mv��B#�0VCY��j���S�Q��5�lIrv�H�K7�ןݾ�G*'�-~㙣H���\���z�:>�f�Gn,*[-�����z�K�YR�j>U���y0��t̷+Lp���?6o��ٮ�uUQ�܎���MiG�!�1u��ſ%��Vt|�x/��6��ݕ[��,XGE<李EO�E����/���_T�S�'[��������?��b��j��i����꼫]���WK��,�z�tds�O���ѥ%J�y��lՐ��9�I�<�R<��\WG/�8�z������Yͥ��&�EUà]��^'F�����T4��6i`�@�y��NO��w��.�{dš��>���&/�����"
�����o^�cX���;���&6����\IA��q�O}�%�CW��<��O�i�-��t���͐���2��B����;����7��VPGA��ڈ`T�`1"��A�����Ju�t+̈!��!E�AJ$JҤ�B��|?����u��de�˓g�g��>{�s��O�r8C]]ʮ�bRB�깡��ῒxju}	Q�y�v��b8f�������g�����Bj'�'`�ď�4*o�J�z�Y� ��k>����\���w�i�VVT�}m�_�Կ��������N���H���zK��dݘq�?������̄=~^���O&R�@Җ�	�Z���4��5*�m?d��`!�)��<xw����A�Zn9�Wk�rKl\N��ݵ�%s��T�U� �ݒ7O�'�x�Q(R��!~	��6[q��R���~������ ��q��m@�F%b�C��"�>y�x�n�ҫ�tl2��ϙ�� FN���i���,~T��U��e������ߞz����Q�8��E|Ɖ:x8�" �h��:�I4����X�UV?���b��ҡ��X����g�r�������g�M�i"6��6�a��7�G�S>�>Žc�P�w�ι��r�+�/���pE�����C�����+��8شc%�Ĥ�Aȋ��f�M ��S�+_��^�2���KQˇ�"�yp�j��Ɍ�d�({E�ZˇF���-)��C�r~Or���]v��
�+l���FVq�&��\�/�8R�;�Ԍ�p��rB�"�=�_�խ�)KWX���B�N寅t���W ��Rp~�5�(~v�ο�4�X/~�Yu1qI�'�F2��$cd@��)Z�^0h'_e��ysGҖ+�ޢWazf���q�����++��F_,N��#In8�&��}O7H��J��#��=*�ͯ����Љ�2d�������$��~��NP�DR�k/9y������[,&���$+9�K�d�xV���aYWU���7?vA���։��|�`������m��Q�J��(�%�n���Uv�Ck�i���1u��Q&�w��>�(�Y�ē=22��,�y��zE����@�az�
ӗ֌_*�N�#/+��1����=A�?�������)�F�  }�yW`5�����7c����ٸ)�p����X���������ū����7 8���,�����7ъVnٹimSp��*Bȍ��۱�G��J�g�d4w�f��f���(ﴃ��"��@ 9{[���8y��f�/v��tCQG��B���j�Ҋi�	�:�
M��ϰ�q�ħ.�Q��,��e�{��
�J��u?�L{`��-(��*�1)��ҧ\��$+�� �J��Z�5Oe�*5 �)��p�
�.�8{҈�!X�J���8��b�%���P(^��?/�]h!EC���H�UͿ��T���]�@�d����t��?��7�8��BFX�z��)����m\r��� �dL���I0w7����A�HUA�eV4u^-���!��`�Bk� ����U:6.�m ��K B�d�mB���,&�-��A�9^��;���o�1?6����
k��:��_Y(It�!K�&��@�p���d��uÃф��Θ!e��H�	�G��ς�ZQsk�����%�C��N�˻�:$ѳ����
��w��F� �� @�F�R�<N�cF������Q}�,
<��w�@�$��SE��
H�F̃n?����ߚ7�0lp���c���-	��f��,�R���/A>״��������6�����0-�M
<���]��T<L��e}��s��4����俗�� ���a0굍q����u�e����)�+��/�� ��R� �+^��U�����ߥ��
��}_���(`8��e�`� A��t{�P�����f���!"�d$�z��#P�]EV��%�9H�EUz�pӁI3h4Ȓ�f�$jf􏏏?�J�A�b�Q�F�9�uG�\��.��"��H~�։# E���ws,�-����u���w~�	,�����1���l�-埥�}si�-�m�������0�-���A�h�%�P���h��;Y��#5�֣,��\��	`!��~��G!E_>K��O:� ��ew�nGW<�'"�t��Hdu�D�p2o ��F����]�.�� >(I2(��dl��j��Au�wVՈ^�Q�m ��������ʎ�:CZ�,�ͥ���\w�3����� ����9�@/�ZrabtDjU;���8G �{��$¼�4�;w$Q��0�K�oP{>!�!k������	���Q�M_o%Q�뭴�n�+nuY�@���-���Af�VEE�n� �TE"(,N����J��f�UR��;|e��!��bEÚܵ&�$�e���D�~4 ��dF��`��&jNd��1MT�6��:�!g�e�M�Z�f䡽ԅ�~��Wf�s�%KV�^��]��ݘ���+��9�_����ƹ�Y[�;Eod�d�-��e���q!=�	��ȷ���:/|�l����Q�`���D�MV����3��W�#�fe��D�g��S�h�`�N<F26}�yz����G)��dD��[9I�U}��%%%`є�H>�#`߆�VF �2x��൲ׯC�Z���yvDYE��"b���Z1��y3*��]T��n�Jj���qR����ZW��*�b�˪u��M��s�ٷ��6P��F���WA�Zn��1�7+Q��G�Y|���B��iI���Ew8�G<�.>T||n��g�?�>������J���y����H�Y?�˺��i:q5��k5�#ȆF�ז���}_������9�\�!!�0�k����Ю�HO6���g+{خ��F[���猪�#�������{�u��K��������QUo0�A�R��ؑݻw{��@t[��N���s��3�֡��w��2��2Լ\u����p\RtY��[W��F�M� ���nj1�ܔ��w�Fg�v�Ai�~�֚�#��h�)pzF��D��Y�t{�+��k/�j$}�%(Iw�[�~&qX�{�Jl:`�]IlW�ߞ�����@��̈�.?ᅗ��<&�#������>9ɮ!6	K���pT�)@�Ź)�����@��޺×���ȵ9���d�-�qj>ӄ�ϐ̬A ZK�����g��@��?��O�#N��3��neHt����}�K���׏B���$P<ӧ�{����,Ev�m�3a_�}���z��v���98{�w+���Ht���Zc��F�S��P�(@��0jT?Y��x�$M�����I)8��0�H�آ��Z���ĥ��>�X�Q~���ē U|�<��:��G�O����>A�������}�A�}���5��3�^��-�w�<]�bʜ��RZ/+�I���=�/�jż�V�*z$�v�G9��f@Q/]E�!�_9T�:1�[��=�U�g���-�3�M���ǟ�Aj}��G�����>$���?��,e,�L�� s)����$yb$��Z۴'�������"�J+�,w/�lb˩4h<�����4�3?�����A`�Q� ���*���9�\|"����\ 	!����Q�ɸ%op�M�>�X�]�ԛ)ZZ>���6�V�ҩ��[;��1��	�gAY`�h)���ڥ&0�ϣTY����܊
ڲ���]�O?׳�cIgh��s��>�vfa��,��c��yg��"I8��>['��T�~��T�.
�T��8�I��͇e�E��u z�Y��ݐ�ġ�m���|'�
�kbd�A�tz���$X;���_��@�:���;���ӸUrx���"2�:��O>���# y]��{�
�f��\�}DMf|�&~���z,`���u9�����<j:!�5��K���9 �X$�����⑕���?������}�|z�j���\ZÈ�6�$H���g�P�qv���'^N�K�~"A��(�ϑke.;|�����C�#�������d�Ê�! ��.�����~�W�]�d��	:{�[Q_��Z���b��+U�Ϟ.6��.c�
Q��7ܬ�>r�jއ��ˉL}�g��,�7�p��*�ɀ#�[8�xH��}IFyon��M޴+�zk廍w���ξ���_�,J�BK %���섾�`�q���lɆS��YXu^�I�kL��'vd_e�1���GC��Qr&��@���o���̓�a��$&P��L���0���LNN������}V��5c����/��ڋ%�2��6���G��Րj�.x�G�c/�ս�8��0��_��8"񘌚�x��k��6QD�z�qR�����Ꚛ���oQ+�a�:[��40��6��a�>�u}i�}��`�(�\q+1I}8 #��j�NuA^��ێ���݇�?�]w�Դ���֧����Iޟ۸�d;$�2�%?n��Ã�@����;�ۻ�W�f\8�&���k�&T�1@�j�D��c���k�$�O�8�'������	C �H]#���ߍċP���D&��� [gk��m�ȈNa!ǝ�T+����h���^�٢�F���\)_�zw��:O � �jx���<�niI��OL\Zٟk#g��:E@��Ja*$�s���H��2'@�	m�-����%�Di�c.DV�y��L��f,²���X�f2��0����K�Ǐ���2�������ك�+/�?Ǧ�3��*�-H�1�,�-X�(oB��1���0v����u���`��j����kpDxxڅ�Ja��N�W��|.^�s�U��ԙ�I��dm�Z`[�����ط��U��"ӻ���']UrU�ML8��n��7ͧ�����]0��?�V�WGf��g��͝�ԒY�ل�!�����b ��D��L�K���!�n~�C�}�8�l�8�gΎ#d��ޅ# M()+�����˫}���r*nu��p�U ��z��g��Y�Y����Ӌ�)bEe�":�
uk�=$�=�Hd3~��W� ��4��P��GN�ED�NW��7�ǩ�U<	�������#���u�;�Gq�j���l8�^��n���4a�7�;�~k9I���F�h6u�pp�i]��u�y�39lƄ{�H���nؗ��"���ܟ����`�1D~��G��#q�HksI�}]��3PAX�C�ѡ굆4�ӟ1.�)�W���<�i��NN职:�*M�����3��+��.ɍ�9�w/<���S��6�U��"�����u@;}�	/�������	p&��{����]���2���[��G����bP�G���2�{[�����/3����?��ӃhSki�ㅬ�[��ܼ���>�Wk���V�?D:V�u��s���ݸ�� �V��5.�a�q�j����'�p*NL�dG`�9��0D�s#�u׌k��^�_l��Pd��UL�ƛ33a��ᣥ���3���{{��Ig��&/�zEi��]�7k����"�1õl�f7{��O#r<T�rz��ʕ�����0�z*ֶ�*�'�-BM���u�q}�����ټ�0�@�-)�LV|�a����	L�X�s����oe����4[��s����Aov�S#M{b��c����v)���:��0̞y��[\wM�$�5!\���<�QK�b *�2�%�3f��¶�f�z������bj`]�%�E�\$�n�����#�R��n1��� Ѯ���mq��9#��z �<R���V�a"�\�;_�ߔ�-	!]�j��!��ԫ�}���{��'L5��?�1���Ev��VF^8�^�2��+�\a�	C7�ٗl�cT��\Yk���6?B	�2cц|nf��["�
�u�!�c����c��M�%h���OR0����2�hJn���]sA*�﮹QT9����J�.�rF����o��B�7�n��VDTe��Yԕ�]3	\���	+���CSʠS�����g�p�Z`�k.�&�c&����>��D�s�R�ʹ�U���\x�!|J�Yr���{��"�s]3T[��{W��G��;Iv�n�-�Z0���BVe,�ZA�g��K儚��!L��U��'���l"U�Q�`�$7 /k��m��:\�Q�a\_	c��[�2��,���
��{~sl'	�NĪ|�n�$��"R���R�YفT96y�1��L��c\�O^�f`�a�{t'Zź���w�W=�B�������0"Ùb��W)����NDF:�&�Y9�{j&�8���:��j3i��O��g�h�W��:��R�Y-��T�e�
�j�Y_�5yY6�z�j�����<����h�F��Gp�uj�pMÏ�����ܑ�D�� ��hka�B�l&��b��]L����V���Ϥ`+3{G��]��-{yxhTd
Er����"\\�[��b�z&x�Ӏ��%� �d����׌���6�������P,o��Bp�7����n�ָͤ=i����X�Ǽ��1~(zt�(�SƈL��B��:��6��[�g#Xmq���DI�T��Iʈ^%�Y�}l�cH
 �񳙰�����g;�J�L�-�^"�����Ԏ]ų�=�T\G��wAQe��!O!8�
�S`��������ͷO(W�M0��Rnogg�p��t 6�'$�8w�=6� M 8�ʁ:j�ʪ44����(]F������Ʊy8�q��f�<I�-jD�&Q����俟4iT�|��~���������X*�D��W���N=&�T8��čj����Ij��$�I.�\&�Lr��2�e��$��/�.�C N�f��_&�Lr��2�e��WI
ٍ�N���;�qC�Fn���7��8�j*´��ҏ���T�?�~���������#���	.\&�Lp���gs�%S?�V!���I��<��Ҏ��Do�C�?�]r�r���'�k�Z��&�~4F�+��ѫ=��:��BM�L��4ū�P����$�0�Q��7K�:أ�-��#y����/>_�����rI�:�����j��Uc���e��UI�?U,����;�(��Q�=���÷셛=��D#,l�|a~��� PK   vOXhT���� ċ /   images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.png�|y\����Td�D�+!*ZD˴qk�J*E�B(�F��-��"d�V�j�s�!5hE�(��}�]gD��<�>�_�^��m���s��z_��u�3~�5�7od߈�`6��(��`60ƪ���/�싿��8����������7ت�s�`v�F��)�����vCQ�������/a��Z[:�_��$dcoE�a�`x0�
�u��}�R�8��w��`��&���`>�kq���x�i����-�S���q�A�rg1#u�]�u�\��ʖqѽ��D���A��뗬M�N�Wj��S�1N�0�����^a0-ⷥ�^2�;R���@�z����f����n��=S�u��x^����:v�5��+�5����;����w������;����w������< �M����R�̼��CwR_y��ح�|2��t���S���]o�[��}��C&-�Y�5�	Y|�F/	}<W�|i^u��b�ud�MK�e��W1�F�]����F�I�G������&Zꅽ��c������7����Ϳo�}����������lY���и�vKr������?���dfE-���aƪǛX�nd��z��"��&�99����]�ʎ>��4��u�8�O �d�%���	g�}��&U���x]a��{+�;;�٧xՏ������ZB�����A�ca投�B��䠏����d�������l�i
^�QHȤ�����[W����9�9�nj賍q����#I�_��Y�6l���xrR��Ӯݙ���\�/_�Ħ�:�|lB¾���FB�q%%r��~ۄ5�*����i;�)B���q`�~�*���;gF��:+�l<�'�%o�9�I�?�w$�+j)��˫�,ѺU;�_�vRU8������Z̕�~�!rMG bf(��ْen7�����^ &F��}��l���^
�ŚU����M����{���M�yWVRPPP2�9A-�s�[���4<��ʕ[����!ܚ�v�������lb��ˊ������x��e���fii�����C�{����ޘ�׷�u}xv�n��Z�iĔS���߄{ƣ��yL�Q�'L�9���\-q|���M�99G'�~�)��璛����Y6%-y�c0+� 6&C��uO��\v�zK�W��a���[k�L_���g����sRv��Ǒ<St�fF��d[h�J�l߯}Jv�OP^+5+KԺh�J�`{�����ʬh�}{��٤]&��oү[gnjʣ#�w�f(A�N��ŕe��>298##\Q�jtS}���$Q���7�|���	N�f���k�:9===���h<��uA"������o�aDј��\Y�v�
�U]�*�SSSsbb�≔C�An�U���vRڑ��k^�7ݺ�3���k:�H�WllB�ڔ�>8xnۏ?�{W���o߯Q1?\�=\<m�6���˽������^ϫݧf�^�L��@vp�4��p1���5�u%�m�B���뿼��/-�K۽����I1��$�]��WX�֐�J@���Z�;hTp+-�M\կ��r��Ü������~]�!I��0?��f���󱣃;��ACC,��������l��Us}ͳ	Q�J��`�mk�������\gF!�?77��au��[�I���%6��76oN�.?��֢e������b-��3��&'�sJ��{��p��;v�����R!ս����r�#̓㐣sRY!«
Φd����hur�����|r1�;�l���M�Qd:*��D"���rdY6g �&���^C6dQԪ�U0�h�i/�^
��]Anb�.��������?y�ĉ��Ϧ��Q��[��;^��\�Ӟ�,��_;:ǉ�w���>>"!Q�.B�+ڕ엘�H=қ�w6�t�,/X�	�}s����6Zǌw�ڔ/,--=OM�c���-����A���I�'z֐x�;�\&�KܜQ@R�.FL�Fʝ'�͇ۋ����b:R��Mi�;��)��L�� k���;'�MB��m������[@~�	FٽV�S1��Y��,�3���-	�'��j�Gf��ή��Q����RT`	l	�^�4�$i�]e@j/��~^��QQ�)�vLJFFF|I��.y~W�Ǹ��{�e��i�������335�M$J���6:]�,�4YZ�H���¿�n�E��SR���eV����T.f�}v�0�ݺ:C6��G!�Ĵn��p���Q%���uuuN��������/�Mca5�=}��o�G��~+!d7$��#��H��n��F(W��8l�d��G�V�8���.���˺֘�4����ݺZk:������Հ�q!r�,�"0����l����D����|�9MG�A_i���Q3Z�ɄP��������y=���7��[����㲑� ����Ӆ���c����m�/]�v��{�.��hW!H�g������O��:�8C�jr[a�XwM���=Z��;�vG�ef
���h�! F��-�a�� ���d5��0�!�sww�Y��ʺZ�x ��T�|-��KJJ[j/�.��h#��N8��JTfm�y�?��s�OԌ�%x6�Q�jn�'.[�TI�	�]o������ͩ'x/rߏA�-��6O�=�&�z�x��8_p����C;�ߣ��E�/���Us9V�ºH�o'��ЭoM}C��2�
m1Qd�c�b }��~�ª �	��'���-+>�����d#C[�j5)b�ޅ���e���G���V�E����mQ���7l狧v
��g�v?2b/�Ĺ�G&k�l�ׯݔ��dIOv(2!��jf����
�Ľ��h G_J��?��@ �h�Y�?�m��I�^[�{`|]�I1�ʻ��1�N^^Z���|���@E%%Y��j�^}��`q�����J �@��]8���fn�;N�'����������v��ф���1�@pnR"�6���O����z�Z	��<f��8���=�x#/���?~Fޑ�����8���f]�۠����SQ�v
s:��%E�%���tF�.\:���I��/�Ja���;[=r$ܥ��n[���n3ʱj�/�hhnN���Ɯ����oC!*~��A.��LG�[	h子2�����Q�uj1@F�!C�=���|�ܻ�.��5Y��\Z�c%�@o�:<\���	kD�<�/��ikk}'���o�!�v��% !��@)t@L`C���\��L�V~�X<�;�
V-�z�Ȇ[C.�?��4�Q��o4�p���-�Y�	6�cC3�V��M��� E��{ ��P���-¿��=�6�"�M4d-t�L,���jB��R����D�����Y�(	������$yp��+3=�<;�Oe����8�v�����Y��Gk7�!7�m�w��i6��D퀁/@�!��K�[�mpHyP��E�i��B����E�#�Kz'�nr��>���W7�?�]� >�������˓���F�f�LZڃRG��<W�~j���
2���]&�I\��^����E�x�g_L<�O����kF���k�a��?�4�z�y[��&�?��9ui��p�%'����uA;:Zͭ)K��Ϸ��C���X���NX>�P�D�:�bt�����#�~Jv�%�4�S �� �.r��^��B*��S?��!V&�|����(����2�b���kq��%�s����^q���T*?#jjj
t��O,�fVL3)�����F#��#�)�Q �Iѡ;��#a1{a�%b����J�|��q'���>���H	���Z�!R-[)_ʡG�e�����[�kܧ�X �թ-ɺ2�V��`������'e��i���=��c��f(��E(�W��sW=IZ��!x��g3�|��}^X(A϶�q����Uabj�*�(����4P��w������~Ϟ=kpeWt�?2ӭԮ��{��E��Ln�e��uD죭�(����KT�3����^:S)l�99)� �A�-�{��Π��?�í�կ��?~���Η=���CP��_�����"kFA|(��˿����dXN���m@��|j&��ʦt�8v�����r���&�?�OZ���lqn2�"��qf��r��n��v9��r�{F����wC��� F?*s'DN�z���H��_�����2L ��-RE�D ��m�	��8Pg�� �S�-�4�M�_�۾�
�7P�?V�p`rrr����"B�K��e� ��T�eg*#����l)�YR ƾ-h���U��c��xO�����uR	�8�|�KlT*�\�Fi�A,#U��@|"%&n�rυ�j�.�Ifs���qB�6��X��vC��#�X�n޼y��M�
���7W>���[%�l``@͘=fɣ�ň
Z��IW�l=A?v=0�V��?S�ɉ�
J��|TR'y��U4�jSG�JgV��ԹM�ʊ��/_��2����pE���p˳�ޮZ̈���{��1)գ��գR��FR[��r@F>I=�M�_�:ܧ���S���CC�ww��dX��WZ�Q�8�=C$\�� H9R�S�I�^i��U荌����39��s���`�d�Y]L..�����I���M9lkR�d�������(...`��)�CW��m�����{�߽��Χ�H�N�sǧ�N�0�);�:��^��V�WD�c��������!AduP����zR
Q����a���[y�z��sܫ�A�ժ�0(�I5?)�[��b�eA�X�#��G3-
>�����p&�rJ�o����%ub�$,��Uy9�=���c��׍ǚo�R���]�r�ލ��e��Ӎӭ�0^�/�+�,_7s��e���+X���NzN({2www'��5>e%X~4�d�ڵk���C���G�B�t�������r��囵tu#���x:5##��&2�nF�΃$�n�����R�	��;�ϯ�͢_([4�=�)uGT�D�5<��Y��2���=d�|��2�:�}�Qءgx۵�~�̽��h���ԟ��H�K�����⤻IZB�8y���PEP�c4 Y�N�g���i�j88�E]��9�r�I�]��e�Ϊ撩�Y������婎��ojj��ۘ�lIK�Dw�w���9�&T�,��))0��v�z�j�}͡?W!=\$���57�ܺ<�,��z����	���� �����Xj�F�F��_-����h#���'X�s�,�E֋�-��I?�#  (��Ǔ,�q�9^�֔��/$R��4� ��?6>�*=[�8��&hib�Gxx:��O���M�/�zӭU1��ꇧձ���7d����|�� �`0ã���|ڹl3�֌T����sM���#�&Ï�HK�����T�>���Jܺtqj�آ��G^Jj**��[o�z��y໧�؜r�E���x�!�������\*�XGF����u�A����6QS<�#�w�S}[H�/��YlBn̤�^2$S���B��C)��1I�d*�f-"��ɕ*�nn�<d�S;I�G�W��?��C���z׉�2٨Zl1UϏ�y�˖���HJdu��1�~�rJJ������e0}ю�j�s-�v憾��ٚ�0=���iC5�c��s�bލD��"R^Ϻ{�l�a�S�e��ZFFm�yTO~sdnU0�������0/�����}���v]ASs�y+
�<ON�O��n��0�l�}�Νb�Z9B��x�����H�#�g����S2��5�Ɋ��v?r��*��6�5��7�]m�率�(R
���I��^�"��L����##Y$ڝ�mLVOS0^4Wj-��n�M6*8���k$�7�<5Wz�D*[/�q�n�2�87Ox��S�i2�3�"DFFVs��	���N����d�#y�����kը4�H�f抗�j�f������v��z�M�T�aU8�i����2.:j�*�Q�q�}���r�s������Ʈ�m�����3�v���3�]qBT�,���u�������we�_,3��r��ܦ�ӭ�R�Q�sb\�9"���y���Hj0��jL�3�pv&�\��*aݚ`L�%^�M��Ή:�}p!�cl�K?�K��z���s��݊�á����J����P}��{0���ȸ�UR�ŷ�o���p5���T�?xP������s�[ �	2��u�̦zXdm�e]n����S{� x?�Qov!��2�|QؒD��"����A,
�I�cJvuR?@P^�o�娭0?�(.���������Q�˟�7�
O�QM�A�Ņ0���  rST�:�<̿�8����:��CWW�e��ݟ��+�;�N�ZGRx��E!I���f1�����8��Dq"!����[~�U�$lb'�@�G����d�E�����6R������pȆ�|n=]BWH%�T�3�i������c�+_~�B6z�T�Unn��p����!2B���7m"z<�����s����!������{8��B����qo�06����ʹ_3:������'r�Xt���39��������*���,����o8:�؟8~�833��ww+���1oxsO�03��(�K�����'����E�s�.�aY�DJ���0v���q���R�Xk:���E��
����Z�0���>��uuu!O�x���C�^~����CA�]��@0�c�Ν;�&���{<�<D�@�7g�̰�9b�ޠ��q����!��͂����Ό�����h���w�bcy�N=���4�y0h�|�8a/�&�]a�:g�N�g�Йhkk��r�좙�,������i�����A�a|��a�����5�[g~?�OmvCfLsYqA�;s���G>;q�����]߇g��DB"���%���k+t����(]�t�T���Ј��xUp�m�\�E�g�'6������.��/�X==�Wyyʎ�ӟ{ݿ���d;� )���l-f�>+�����7����&1��l����x䞟g'�$2��0*��߆ey./��zz��%:�EǸپ�������,-���{aK�"M<f?��Q>��+IL����\�_SIM��s��21I3&���	�5�k0�]�}��Μ��l�UU	�g����($QV�V���rc�D���e"� ���C~ʒ��9�����)�&9En㘟��>?U	����8�:Ɇ}��Ri��Rdew��.�ˈU��n��e`����R�0_	����x"ɴ?�|��W/�����D���?��������uH�x3�\�qDD�����d ��$��pH�Kٍ^����ۇK歁1I��ޯ�v],K�}��+W|��� ��4���R����"��=��T�/�c��JKw�,u�tR��x�= lX����:�S���qpp@���o���!������C������B��0>u���OK�`����g����CȻo[{l6646Vf��{H��<�����{xc�	gE�K`u�_z�B�i���� �:!�Q����W`�3�ی���K	�pهG��A�K����yB��dŞǸ�?׊CA8��:��y�����If�ux-==0��X?�Ą�}��c�g��j9���K����(���"��Pd �J�7ݺ�-_:ܧ� ����i��J�����1���QA�)��֛}yuUԼ*�yZ��u����I[D���=d<M`�Qu�c[�w�;85�q�d�{���YH:Y�c)���y�� �m��D�:�aT\��U�vr�%%�ggg�}�l�����L[_�˗��)$EԄn�gI3sUm#�]���,�H�H��,]�Ƣv�d�A���	�b<
5��.����a�v_�kQM���H�ud����,�Ůĥk���B�� cCCN4����CYכ��J�Q���eܨA��K����Z�UZ�|�tqq1�(qGN��c!�p��˾��E産C��* ������C��������<OM�X��rnG�M{��--QMM����

(�!���i����Ec���5z�4J~rʹ�͒:|$�{㓔���N�с#xo\z�!�6�
T��9�5���0��7nެ)�+�N�%o����EJ���XOm����]<��QP.��^9���խe��5ݱ%%r�܊�u�����:�RN��'��2p���+KaBa)�%�\�����p봸�=�B�� �����cW�C�Ҝ�e��l�P��"i�o?�������/I�����,��T�<".�X�p�һp���*U'�Դ�ۉ�B���כ�oF��	%]�H`>~���F��k�ޥK���^�I�̴���Q�%e�uأ�*J],��2�����~u��q�Z�_#��X�Yu�Ȣ@R�}��C�/@�qF�:Ec�k�׈|G=I����G�Xl�y�:2:wZ�Y�*�Cð9�PL�٨g���"��|��B�!�Y1��u2vB����lVgz^�?�'X�9HX,:nϏ�Rvo�tyz9��u:zqF]&w,���|"�uzz:��ӷ;,�3/ف�4
aꋥ��X7���"/��?�`��� �mY��I�F�ʻ�ө�%XHgz1��3C<�z=�������M�/n[#��%�$"n��j�kew^�������X�#��v��8��V��WM�=J:_s���ANV�;��y���>-/.��h�B'�)�� p�t�7գn�UsK����)6LLlv�*��̘M��&;��]��		␨�
�0��aW�.Q�Y�'�6Qc%�L1R�V�ER�6��������CB�d��|с�=C&gg��z�y�������I�A;H�(���r
O�y��	�0l�u�R��:��P+P��_-~�����"ؙ���|�׾mmmZ999Z�f rv��͞�/�a��uV���)@4���.]\@�9����q���]ee7He�3�l��
�uR��������0d�h�����_��}�Ơ~-c�����7n܈����>w�-U/3x��Y��8�h��:.�#~^�ok��ez�L	.��+�7�@��E�ĹI�h+2=���tq�!����+���#��0��]J�?�vHFN�d`ˈ(��T?�4�Ƅ�ֲc�5݈-�d�3�e�"j��J5dv:���$g�"�k���X�p5�,�Z��X�:��!;��͌ҥ9h!x{ZA�C��ސ�ɫ��=hX���%j�	斏Ʈ󉘛���s,َ҉�K㨬�J��F&` �o�s	��Zbe;Y_"d���@�b�Q��0��:Z����An6
2t=O�?JC��I1�Vw+�pJn�l�BMZ���v
�M����$ J7Wo���_���O�>m#�Nʀ��	�M]`M���|��nSDqy����%J5E�2���>��@��Ȣ�=�*�]����_� ��^ֶXq�W$���n��⼁�6���ظE-�Pԉԙ��:`���[YŕBvq����i�<�6:1q�yd��h5�/�Y�<.��Њk6B3n���Y�܌��4 #�:P�hԺ��Mi�L���<�q���[�W��ᦦ��K�e5b;����~�'ʦ
�5�<8���=�AR����P���T��ػ�xzQ�o�֬d��)oɳ1�׸�;�jD��

��أcccr]�0���);˼鸹��� K?E�Lx�9�=��Y�bH��4Bg@�Y}~�����B"��ZO����w�ޤ���j {"k4n]H �Ine�,;	�� B�{ooRm���uxHˍqYwV��`�%3_��гx��FXP?�ۛ�+�%�q����e�Da��z�~t/��L���5�3��>�wtǎLL�[Z7m�LZu�1�k�5,������wd�������)bB���Q�$�~��%����LiN@���^!v@��-��ء�84�;w ��>�F�������Ɣ
:�������/�Ə��r�V2#�H�5H��m������ˋZ��[��x+��g��>e�v$=�8Ib<!�-&&-�:���у^ޖ���G�/Z�63%��R̓�!Z�k��P"{�ñ�4�i�g�S����M5�jt+@�7蜭
9���D�.y���A��ao!�L��|�F.s�D���F�!ȓ�N0VfzL�J:�����B�l`�]w�p�}S�����4�KD�����3ޯ�9F>�A�鐺�ΟgG D������Hۖ��"�qi{����܍�!��jnOv�Yt�?�)w���|"�kvv69le���������q��v ����C ���}�D��0!�v�x"� L�����cb��Y�/�yu�㶈x!>Li�y��%RY�Wx��h�'
�;��Jĥ�
�}���:�Aڣ�`faIҠ�95�2�n�4��ЗH����B��WWø_z����iS4�ĉ�q�r���u�+D��s��c�A����h�KK5<�D�^�=��z�OK�}�UIVbGC�	��r0*3�b�QY�wɲsHX�����TV�Qؕ�Sͣ��U!�]����Ͷ��~?�v���� n����d�P�̑n�g#j����2�d`SI�(��f��o�*�ink�B�r2��܂۶����,&n�M�,��Oǰ���k=���'�gGa蟀�.�vUT��&��X&u��y
<y�%yR��T����VN�}����P�1�1k%�|��46�ST�:V/��ǔA�A$j����2�QZ�&ɁFl��¾f��#�)u��i��K�;�Az6��:�*3�7�<�;�`;3���Y�s���uA(�v	��4�=8�ʾ��>Dn�
j�E)`�|���!Sh8��X����hD���
p�����g6 g�����J�(�k,֑�{�&���e#�HQ���u�� ̻0 �E*1��1��Sh}�wt 5S���q��t��]�J���cSRP��WŸ����	f�:��G�4���_鲐�?j�꓏��L��Gb�uO�\���r�M�)ӄ;D~�	5N��A:�����M��yT��ma�sLj��&�zz���Q��6G� 	4����MN;`"~ZqJ	+<^�r��x�����/���9�pw�qP��{����сO~�AjMMMX�\YSSs���ԗ{����)w*@
Tz��ڰr�R&�K֔�ԑ��fj�DĶ��3J��p��'"��l�q�`�P�|��G�^�H�d�б����ZU{������~&�J��2#���6����S	{'d���?�mi-�#��K���'V�>H23�ۨ����a��l7��DDDh�=����b�Ce1�}��0���^)�G�<fPhݼI�h6rL�Ja��xuW��.��Y"j ��x��2�6J���>)�gQ�V����r�w~�T>צ#����#i�D~���¼���x���w�O�Q�d�Mu{�+���,W�r*H>�� 3��c����
�XY���� �{
X��=�����f`���E� �@�.��$�5�]�TUo����FY��o���Q~�va,��&��<+K5G�rf�vr�{E�� Z���=n-���RSfT��g��!��j�	ʚ~�l
W�a(^ڱ
u١z� ���' �6œgQ���y+`k` ;�F_���񩪪�<��"%kc����Q
�)dط��χ�n�`ع��.��Q�8�8ر�hW���@����
�e_v�
�?�L5�vG��kg��p<b�O�W��5OhSxx�o�F��V�\���<=]Ok�
�k6�S���yFF0%˰Ə��B�^\>dH�=>�j:�q���.�	�̽�>�*�PB��ѫ�L��x��k&�L��O������Φ8�����w�i��<`�8�pSF���/y���Ѩ�J����J:�]<���,���x��×�1n�ŭZ�������A6E<Q2�j��u�O��h��J6�z݋���ݫ(�zO�/�/44�R0�����~=pP�hkadHU�`�Al��Q�*�}  5�+?~\GWm��JFb��BC�Y�.���MX���H9P
����<�XEy7n�hV��Ի��ⅈ���PH����%�S_Q��TJO���u��c�GG���2?(�ߐ�bE��-v�{B/ 2�L��'�]F�`D Ea��2S��pT�Ӕ�����X�3�J�c�~�@�0>E� �P�?<\���������I[J[ZX;��:��DT���C��@@S�%��9�`۲��Rۦ[4V
�	`p�H�VN�<ʘ��{'��c���^�խ���GU_�{::6\��H�L|]4}:������G^�.�8+7��r#�1�݉���ʼ<�D��^^�޻uF�{K�X�	/�L�?�ޏH$�IqE@n�G��!���M��	����&�o�ܼO����u���_�%��q�������$��x�Ow�����W����W�&j�VN@��WX�踞����U�c�8�>0���@�w�ct������7��9�\D��r~o4+$��kAlv�/.D	�E2�hyxx��O-����Yv�T266FZ�1�V@�9�3����&��J��L����IO��5ݔbP����7�����=��8n��-��̓���Pj��l@�Z(��쪁�ch�V������\�h���իW�5Rvya|�8��s�6� �r�Yݒeny�By E��>���V$G�]6�S6]�˽˜ঈp��21}�j�@.�N��Ać����ς���AG�a|�'�ƨ| �>�J~S.)��%��6U��ڿ���OQ�r��Uកg�cD���GI�C8P��P�/Û�/E��s�{�h��c�!v��v�#�N�b�@�no�֜@��9v�9�퓀��� )G5�3�ފ �Da��_���9swf�t�R>�'�)�R*�6���sb����

����&@Q ��8���Vn�X��(K��]@5���mG�g�q���b�{{�o��d��.���uG�ЅW��U��ܞ�,�Lj�B���Z�ῐ�?G'�ھ�\������K�X�k�`���8\%Z;�C�䂚�>�4ee����>�9�X0&$$��=cg����߁�{������î�9��2�{���k� �)W��mu���z)))�0�e0�@�����.��b�e��H��b�d*'Sѣ�O�Ao���	���򳪨���AU�njlA�˛�e\B��_R$0G�k�˱I2�ߡ��+66���VA`y�⎺��.�ꜳ��4�ѥ$t��.n�ߣ�c���:�N�����A���E+� ��S�n�r�b4����K~�3=���/�aFU�ъ��r��-���Ы���n�1�}�|�5���"��Kl>�a#�YhnnyIm |����*t�1E�'�r�x��ȆXH�����B��:thT�sB�w���K�_����
��BB��@���kx�.��R��U�:�mܺ8Љ5d˹���FFF��Þ?��7�.F�����(�FA��ϔS�v��E���U���@G0ԯ� �> ы
��7���6̼��t�ċ��g[��:��k��:Ŷ�J�Y��}���c���'��A��{��7����X	���`0��l�T�%F�P�̼�+1��r��,�T	��-,,�����A�:�42 ��뼎?��9����D��FQnq>�f%���*U�"��|��^��Hq��Rί��ji1�:������L�H�Ofz��<QX��Zzzz�ʅ�y����M���?%��m� ���x46fO�H�\�~ݰ��W/ �(�4Y�4�F?Iыq_����1R���葘E8";c�04�>�+��b��s6ғmvvivew��b�0�ʓw��#���~y	�{86�����u<	>��m����7���}jh�7�l�A�e�V)�#�}�Qt�k�&v�=8�SD04�vw5�.�ܖ�;BJjJo���)'�`����!%�ݽ���=�-��9(���!yd��X�mص#�t&����A�������#�fdϛ�麻���3�S�x�Q���/�H�dmS��wWh+ڦW��]�G6EGI�帖���	啃dr���<2Y����x�	:GV> èV�N��O�H�.3 <ѹ���Tp�'ORΙ72��+sEEE3z��~9�{<��|�$�*UYY��-�t��v�Ζ;��={v�g+qT�L*{�P_��y�a����.�O��	����vS.T��]:�A,�F�NR��qv����xI����r��1���(�u��;�v,�Dw.�����R�b����u����F�G�tK�T�~ѣծ�(��EҖ�����T�/}@Q$��m��eSZ���[� ��3H��H"�4+��.Q��7��
���@����PzKQ���1~aa	ۻ�#���ZN�m5�!��"�G;�
��tZ��_�Գ���w'̍� X/�.N�#�~/a`�N����εs~,�pٍ����j��Cg�讽����\�h�M�A��x'�1\@���	�᪞����Ћ˒���9���&Ƃ~BGP+WFD� :����o� h!R�{�-�#@� F�Q��;�y�P�Z�����D�|�AO�O׊SB��(����h<@}��8nE`li�s~�&3`�_//N+�R��m@���*��U�X�6b%�t:�%5袞��(� �#����r�Z����Zq�P��?�\2}��f9���.��_	���� ըe+����aJ� �|萐xc������G`�T`���0
��T�^�F��������o/�ɀv.G�G�d��?{I�V����ۇ+~��5$�P�<�H^����;v��>`f=��y_y��=B�� `������/z�:���9�Ά]��Մ��Jщ2���gm�	L����pr$����+��%(F�,6����Fm��@�mQ��gՌ�5�/���rFyN$���#@����]j&sg(L��%�&����Ǧ���u�?QeeT��1X���X:�Z�o�������Wj�i�{�Y�~���F[�AZ/����A�:y���C�����Qy�H�cS��y�."��}}}*����$D�������s#<��EZ�����sM�.);��:�D���υ���7I/we��w����G�~�U�c6��~<��z����6��ƛ��C�~Dg���4v�Q[{_�?�o|4�{�y��硭���S=�Mt������M8�Ǎ��$�bZ����Bx]�#��~�ć����D�v;;,�@E�;�x���{"�o3���'c|��i6��&�z��<ʽ���1D|���v�m~}���x��4mL+/�-��k�>f)B�|�� p�E�W�kʼ.?K����$�U-w�����b{'DnNE��Ћ:,�Ѧ��e�Ś҅ {�t�3 *yDA�Mt,/v����Р�ݤ�A�:��������4��*�/��K��%�i�2��өO��a�F�|9���J�Erl:�ҍ��`���:v��A�K?}�">�%����*��!�O1Nk�#�z��{��$3���[�][ڑ�O�A�loLs8�v��L�D0�4$�h@�4��9jO> �]m�����R �#-��E�Ν;MR���ӂ��0�@1����f=�]y4#�X	t�ϳ����������N)(����wov��=qx9�/��z��z��Lt���Pey:�+A1`����s�Nx<Y C�;��[`f�1�z�oo�3���[�n.]�Z�_2O���vb�K
�c���=77��z��_�}�?�؎���������7)������dքH�kld�ϵ�l��!m���Dz
lW7(8�|�1��dV
��޾ͪ{�1*B�288X�UN��X�Ɣ��'�;��Y��_i�ndccs��l1ǽ�o��.O�}������b��6��dv5[f'��2�ij6�2N��=Ϟg_�s���\�	~=�����Uv�ų=QX�@8�䙇r���ɲ�ȹ�?����SH���`fjqqvm�ŋ�5��;�|���v-??�e����� s�˗�X&i"[�]%L�o�Wx�}�I��f�~�z¥/i��p�I���/*xΔs�1�Ӓ�h�lIe4׿�z�-o*�������#���XmC�O�.RU5N���cץ4�Ь��V�Y0�Ž���n�x|zZ��A������w��}���1K���$�o��6E�>��Yv�R=}ݑ&g���q�o���F���4"�Y���N���;�g�����t�u�>ncF�ǲ���Mh_�d���Zi�N�cRJ�6����r~����hwUa�89R3KR�^��5biɣ�9;G��] �@d�B���Ǘ𷈤+<��		��z��uz���Tp@Ȳ��^$�_p�M�q�����+7��k ��q�^DH���"�W�KZ\\<���U}qq��?�h"�b`qM��`zZ��E�_��20�@�ƺ-�/�l&&n,�T�����j�AG~u��器�y*�s���z;]̰�w���XŹ$Ϲ�ꏏ�Ů3�R_K�Ù����O&���rȮF�ib��bbڈd���ߒ�T��0� A����0�q�ܚS4� 4ū�M�:Q~l֭I
� �4ИFdgA��$rt�G�BGC<u.�ᇆ��v¸p����]�9�H�8����X�5��	���8d��[��~�M�W ۀ�����&6�RFaa��/��7��/H��T��񦦦^M�8�M�~Ih�J�d����g�ݡ�Hh���a��{id��~�̅ό=f/��c��u�v��,�2���O㴍αL�%n�E�a�m���H�� ��{�f'����L1��I�s.���|� ��F��}dL���kW�f�ad���Y��q���a�4��=F7�?�d�dD����)A7;vip��1�Gn�DwTB����x
���j��2զ!�tI΍�,��&2�i�,�D���v�Y�ﱕ� �O�m��`[��ۅ�Y��YJ�=�\Br�*0�<p�|������iڶw	��z �%pΗq�mhh�K�K��Y�	@Jj zL�]�t	�a���		��tth1s���!'MLb	�,g�TPp�(7���Q
.B�LG3�u�oJ;g[@��DY��=ʯ��o2��	]n���S}=�j�;��e+%i��Ra�w��v���F����J��C��!���l�!j���:�O,�2�������۷��-����I��)�v�~�)��1��w�d2�����V/���8$Z�̛�2��x��֕I>:|��ev6��M��D���9::�&�c��I[X�8�Q���){��T�cWY�ʮ^b����� �ޕ����I1M����o�U%���y{��� �y�<~�Kέ[~���ӷ����@2�yp����7LT.����_D*�D��g.���~�g����1S<���)[���0}�����e�m�[���P��8~�̀.I����#22VT���	���132�6Gv,M}����*�㘽~�}VZ:]�+CEL0�H�qƽ��T�S�y�i!��|Ȥ��*�v�â~�d�ê�<{�ۣ�v����{�fY�@�eѭ�[d�u�s�1�,�\���ڎR�[����|��K~��xmmm����ׯ�2*�	����L���{	�a��5i�1����i���*��m��~�E��o���?iz�m�}(Z�]���CZ*#]e/���I��G2� v�DS^I�2�{�n��ӧ�B@�R�����9u
�=�Y�1ʦ�^��IH��D������Z����x�@�]iLѥZ�ʅ(	��o�w����4���^�{�QUS�>~�G�e0�V��5U,���6�i@��[�ݧvĢ�s��UP@���.h���տ��p+��!��	w�ڵ��a�%�ג@�#�d�t����2��2}?~���ƀ���`~Y�i-�)�7@�&��Wo�VE�[��J��6t@�����yрf��e~7x��5<M<��=h�{��ly+���t��� =��mbB��6��(��~&�g��
�.�=>��m��}l�s�Ƥem׿��"��pJ>ML�dp������Qq�%�����@��l�/�۰xy�v*��ZXh@!�w:;�����8����1����f�{IK�hJ��˄����z���'A�׼���OHH~�ܪ�ȷ��e�G^�d0n�Fd��.��7��l��عs I~1���ð
��{Eh�@F UW�Ux��4NG��A(��[M�X�Ƀ̄����Y^��-�J%A�U�jy��t���x�c��`��,��bbaa Ȥ-����|�P>Y�r�wö-ws �r1��3��z3��у&%�����������k8)H��Ѯ�q]�K�0�ͳ�9@�x����`��V�@����QU]@P0��+ `!���}���?��4Uo?P5���b��Y`�ɘЯ��H⹊�\�^�*��x.!!a�J���&���
�A����EkUqpȖ[�1���/z�1�"�b��?����a� �����{6��*�����}��s�U�h(��0F�p�V�\u{u��o���ÿ]�_�����?M����2,M�ѵ_�_Q��jaٜ����(0�9>�q~��zLI��_1L`DoJV�G*�T5��%��F(�'Ҝ�&���Ǯ闸�g�&��'�I"���_��6t�c��q��*?Y��+�Y{ěVYhY��q�s�˰��ΝsY�퍸��6�[o%J�HJ>oLՃt�
�G$�l��3��/$B��%���dΓ315�ĸ�7<�t��Oi1X��Y>$���V4���2�)�UG��I��ЍQO^�� AW~��.+�e��a�n@���/.��B�`�QWW����؀fF�Rwlp�x���j���d�
Y���,�b���l�C��끙'�g�<���3O������qtI��6+���~�p�Sa���{�8l��r���u2gv�����������-Tɚ�*�7ک8� �}�Qf<vd=H�4���T�#7�#� �+]�a��v�ݻwG��d؛���$ &VP"���4��*M�R�����87	_��X'Z�}�į�l���1�O��t,@��x��n�s�Nѹ@��z�h���>��$R��jH�;}�=�Nd<dy&dŉN�l�]�	�hT�.:G��a�Kc���a�g���Z��M��g�StS��Q=�w��irLW@@��M�������D3Z!;�J�Yy�U+AV���I��s������g��	��m*�A�]�e�s���X������Ů�����֛�S�>���;�ž�J�TDYCZP�d	�-�ز�Ѧ��&Y����-�#�R�PG�Ph!��?���������u�y���y��k��~fZ���<�3�kr���T��l;��o��ߏ��Ղ�������0�枚˙F�O_�U� x�V��RV�	.6/9�	>�G�IJZ�@��xɋ��o�u��3��sѬf�?a�����^!�����	׃���ij���U�x�C���9oE?y��*�0l�t��/7���Q`ᓮ{>��d}Xe^DI�a3$���dZ~�:FY�#�W�/���나P�[����4��#_r��N��S[���%-��[��%�o=�{��?m��9���ϐ$Y�G���{���;�������7�+N慞)�����)����c���p����D���GC+׮�{�ҵk0��6E+�b.b��Cs5/~$��[,d�C/v������k��}W�k����ۖ�R�:��s�������*z�}�^B�IFY(�F]?�n�rt����O.���0[�ߦJ���mlh�˺<==<W���(�꡸@�U�菋7_b~"��6�RG������$\��+��~Z�IT���I�T|����<>O$w23�s�, H0l�Ѩn�A�Ӥ�sqr�}41�:X�+6��G̷��޵.�"u���6M�z�bbu�E�n���ih,���>!���ϗ\v�065�-������}�����5;"�Xk�jr�__LMҜ.R�r�|�s#�H�<s����n[�+8�� �yp%�p��Ƒ+�J��K�#�:r��������lB�˺�;s?8����	��<��҃׭(��~,ή05���D�.�s�� 8�X�_��Xtf+>���ߴ��G�
����_��;�z��Y��	�(�G��T���F-����)��]�&:r�����p��j����@�����2w�-#��ѭ���.���5###f�����k>�_!W��K-U;��3`�~��#�_��|Ω�':8,C�

6@���E��R>�[��f�9V��Q?��adj��7L�[[gc�r��f�_�2���O��5����P�����毚���/�6��u���=���Ϫ���FjEDD�����0���NP[��� ���r�y�,�����.����b4\�|�l�3���;fo������4��l�k�wo�<GG�)��l$<���?��9�
y��@IR�������߇r'�����gՍ�����\Z�J�Pk���0��nnYR	��$6AN���~�Q�
����u;���]01Ȕ�n��D�7�WR��&=R���m����|�Eꍐ��DB
�0A1���w%�
�*{���H'B<�=<��㋄��Y� �w�}�$����;�\
Cd�Y�[X�||.4�I��d;��m�����r��Z�	)�!�eʆ �x�G��Ā�Ʋ�FT?� I��ם���1�շdZd�<8���م��ѐ���	�˚;�y�����7A��f'������/p����>����ꁘ�����J���LW8/��EQ� ���o߾v���D��4Z(���V�`�R"I�~��_�1�����Ɯ}率K��v��+�ظq��o�}؆UH�M�ɑ�\���Sʁ���:�N��C��g�8�[b�ns�˚4�`�˗{ �H�ϒ� 'w�8�|sG�]>>�$%�֯$�g���i@�?�c���Q�Q�D�qX\�����m���@3�ED�	'l�ܖiII���� 'e#G��ڙ�����GMì�~�{]�,���+���L������\}�w;�����x8N�%�dU��]���Z��3<�			Y҉A��,c���J�>;�{�)|��A«�p��R���o�[�'n�raQ�8'��K����J���V�wy�'�َ�_�*4ݻ��fZ[W�w��(�~�r�����j�A8 �8��V�	~l/<�ui���f�����/����˖�kη��x���gq��#���TY<��b�������\ s`Z����Q��`do��9�/�A�Wo]i��S��*t���*�.����gϟ�|mN �8�����1��������c��LDm���U�.:�D+�����uu��6O�)a�#����a�X��� Rx"T�
y��	ϴ�XS���6���Rk�s�yc9hm=:*i�
!�@xq�������|;����g|�㟜����#7�����Aj!��D��l���9���{���4��:��,8�1�	���zg�;Qc�?67nm�ȫ,��_��U��c�`z�azix�+/�	�t��! Bۥ��J�*�~�T0n��u�~-�ɐ����J�b�iچ@�m�sihmy�|6o���u���E���ʩ%��+�n�1[J|�
�u��*\v���_fuD�8�^��K�46�cW��:�2w�#�����;@k���"��>���;w�Z��ܧ%�B2>��7��M�W�޹��wA�elf�}���\�!�u���#vg7� >ڛ�L˵�$'!ʹU�b�*�N��� ��e�#o]�����+�:�<��'�<��8�v�|�~�j
z�%��� }��/���]����U�Dc}���oQ3���>������.��z���U]g��Y|��E[�e*H��>�Ƈ�ԑ�]�l�Q�>8	:s�|�O��I����~�q�����n򠾎�a�+XT~��'kAjj�*S�л�[��7�u.��J�һ0Ѯ0���<2�⣼�$ �h�����4�Ʋ��<R���1`㕕�w��%OX���������?K������ �/���k��z}ĭ�l��qV���;�*�Sς�j��t"Z�ќӾ�m��� �������#���J.8�������\��odt9��c˖-w��[�����!77ܠ�c&�UC^Y���葿��^齺�DR �~��-����6���L�V�A}�ͭ��*�>|�xhr�ם�,rwVx8�IQGWy������]�bϧ��q*F����QL������CA�v*Y�9�;w�v~~�jy;XS�������	��1V!�;�F����V��^\*��@Bn,��o�"�uiH��\V6��ikk�U����1ɹ�=�P�U���ǻƳ�4f,�	(���3[ݓ:�s��i��	| Jc��ywn߮V�[�:��K��O��|�X�h�Ft?Y���Ĥ4N���y�֌�#�0�S��?
0quu}~��V���Դ�H�W��W�%j"���I���o���|>�tr$;���f;�4���B�DUU�+[�$nܿ�8�H�:��pb<��H	�qrUD2�����O/�[�f)mؐ���*A�;7on��/�����9��L�������M뙳�{+d}����ǊO���+��L�򙚘�R� d������/G��a�7����(������6_Ȇ%��ԜZ2>%��r��A�����2Ѫ<^����l��n<�<���������{V�6�|���Z��Q�%������j���e%m?�;'g�}]�}�ߚ��ys)(%=7��!8���s�'h�N������l�`6�:�q/�էDd?��?Tv���ݻ�G� �W���fw�3�t2�����d}���Kw��	�?̴���?�����k���oK|�!�^�v--.Nt@�VQ�e�Ye�%"����L.,4el��d�fC.���Чh�����L�nMN��Ȫy���߿L�ulP�o�����K����3��O^M��O}�o�2��K����̋�	�&D���kK�o�4���eN��
[p-���M���A�� `���ANsi�r�<l��4ѽ��*�{����k�e�'����ۮ��ד�w�����|}Uל\\�$�qpH��'����/�w�����hbgle������'q� j�AII�w/j�� ���e`�u���6����SQQq'=R�b����7SQ�����	�5��f��~�u�4p]�9)��ش헥��ʖ��~����YS��6�7�����ϱ��2��w�j���in�HJ������`H�����$<��(���|w�K�'��_`���kͥ�0C/�x����C-�d���b���q`sCÍK��ܼ��ug����������g�i �1�!���H�Qx<���9�!c�;������`]"%׳��/^��d�	����[=����/5��B�����o����;�����2g�rI����><�����g�r�����e�VJ-�o����@��Q��c7|8(U�E�>��K��8�X[gǫ������塀�����f��m�%�ȃ��Pu5*��o�}�L`,��o=LJZ��ڊF�|�����I�5�#�!We�RZ?�>M�tUwk��Ϡ-eH�1����+R� ȃ7�⮂z��h�"A_�pA{��pE�ɹP5Øne��[r�j�����'�օ��)g�E��p���[���K6�[�]Zj0h+��u�2D���K��\��耬R�?��N.A�\ED����bbc�8�L��Ib�ǿbժZU�54�?���=�,��$�q�W��	r@�m�)ɋQQ�ǎ1ÓkTY�;�&�����}��SU֢e����0��<�4�z�W��ADt��O�̿.���,����/g>u�.�q��dWГa��OODh+�=1�"�_2���ᑃW�q�瀢� ��[���`�#4b�!i��xzz�v==�ւE�?� ϓ4�9wm���f\�;%�&O1��E�D�܌��GYoW�9 +Y��Ջ� D�Ǝ��*�����ھ8u�FU�B��̭���Ϟ=362JvnJ5s,��$���de�G��R� /Z���m�D^m����-s�	<]�k$����5ı����i��F.M߰u�E�3fy驩�)))xBə�d��9h�!��������̢��b�u,�d*b����f�҅����Up��tnTlr� ,�ML�b���ۼT��#�<n
�x~]�e�N�5k���Ӌ ��7R��b��V�~�������"b�5�IL_g'']���vo�~u��z2�H$������TTT<�L����m�S2������7y��<6+D�]��@�3ٶ�$�q7O�)��<��u��q�j�+�s�?ʆ�Ĩ����w"����EڒP�P��ލ��X|o���9E��L�H��@��,�K|���K�w��?m!߱..B�R �Eݭׯ_��z�~�
�r��I�xR������p�ӈ<E_����08�k<u��K���F��r���t9IP�=Eu���7X 
�Cʻ�?�̑�������y�Gw�cy�g������[UK'N����Ͷ	�(`Ïϟ��i1-���ҷ(t313�ο��6�Fs�q�v�2�8L�V9�+Ʌ����_�ƁO=y�y��{ZW�^%ώ���9�	a�᲻{1y zVƖ�;�h���׫W�RS��V�r8��ڮ~����������ny�֙IK�X>��6����?";v�(�4� ��d)%ʭ�8X!��̥�B��?oߚc%K0-,�R�d�
��ۜh�]^�5`��x6��$��]w��E���RJ᧊t}�y��R���u)�ғφ���������D��b�Tb}h�C���`�-���xYڠ@��Mg�ˑTކw�&�3���vH���k�e �E��;|�i@��׀)"��$��ϫ���\�� �m��'d�xpZ!rsVi����]�G�W�̲e�/�Ф�����׭���a��q�	d�O�C2K�B�°BC�<w�&a34Vœ��"&�0�Z���\,� �=�g_��f>�,�p�Y�PɮY��n�FFgH*���X�\��o���E���G�JnV6���d��ITrK~6GFFa�}�r�����!���\Z9����,,,o�d���FC`VW�\!O�u�Z"�?�\<�$%�;������H;��l"������?u�aA��b�/^p�G�A�� M7�ڌƂ40�/�W�Us
�W���<�=u{���OXy&�3eٵ5���͂(���4Enɴi�2�	��Z�����==N�t���g��Z�ǅi�I���rk F
���;�
%�>-�]Y����`�J~a�E/AY��Qܘ'g��Bۜ��X�����5�,<-Ԥ��A�T����HE�����5Y딕oi+̀���� ��I5]���+B�iw��'�1�=�.Ϻ&���hXg���g�n���y,��7�I������2�U BCZ�����nU�#�R�mʘ�MA�kq��Q>�[�K��a�S!.��򗭯mij*�b��sf�ׯoWVj��� �|������F��qk�	PGk�EN�����\�
�@s HO��L���hl������M�]k��������P,�(e�2>��C�28]�@���b��2��7�<0���rN�<���Y���>>>�(��
�!G��C<�Seպ408���g���e$��gWF�~[��P��y��ё�+��Ő��{���(=9�B�/}�a�����Ԕ!���D؀�z�,�nޢ�����o�ۏ[y���@��٦t6�����
���Bƍ8�бS�[2\_��[_�!: I��c˳n��'Z�� �1��QrO ��6,��o[��,��]��ѣ6"�����W@`�4Uǣᐴ7��W���pOv?>��Ԋ���KT�,F��E1�j(x�U<Z�Қ�|�K��v]L�z���O1�*o�8}����]o�n�0V"�'��B��W$�x� ���
[DeC��k`K+�s6F���~h�;���0bH��CLv�l�ڟA~�@n���C���zc�N�B���ooAp����ת�� �C��J\�0;���W�1�n=�=��b/<� ,fd�|���}-f�h�,���QB*oE�������lr�^p��9��ɉ��!!�DY�Ǐtď�b�t+��j�X�=� < o��X\y3�������*Տ̧�s�6 	*d��m���ԃÎ�ơ��^��Z��E���ڀ�{���OD�V>��}�ˀW>�����9ŏ���;��-����?0�pݬ=�������ON���̿}�Ύ�ܝZXh21`]|�Ӧ��w��'�����zEE�c,Ny�`�ʌ�D�km>����͛7�F�������<�ܲ A�m���[�GL��:�!'\Pa��x��$9rY��Ǐ�̥�R�]�����H���x~8�8�����	&�&��ǿ�9m�nĕk�/+�q*^W���X���?�f�Q���#,$�G[����.����ߗ���x��� �l�:M�<���6$M=!"*�
|�?G2,�.L��	~�W\��#��Sz�L~]#Q12:z1&D�f�+c����m����ݖ��P�N����e��A�x��9r�ѣGQ����7�����!��� ��'!w����|�E�����),�OXke�eKy��z&�ޯ����)a����9��^c���>^j�03�~�����Y�Z�u�l�w.ã�<�ٌؙ>��X�lYuA\�'�r�.#��$�5���������̡Y\�����ލ�g ���� /�2utrbN���2��,�
��y��
�qtt�Cv�����'zS����p�O�h=]a�!��o]'����:_C�4�P�R�v@&݀VM���۠ڐ]ɛ���ޝC���e,�N��N.9��1>����x�(��9Q.�k�B?�m窔�#�dN�W����Ct̗޺m�ggƸ�I҃�W��cR]����Y����|�6�c*��M.8._W������%KT�75>	
�?�iR��l�uy��j_㇂��
Gww���V��_�Sg�'��&����0Ǆ���fkx��y�t�O�V���{��c��_�{�Gz'>�hzz��l��,m4}�@�S:�Is���~�]q�?/�A�E�)���J��}�O�##��Iˈ��ѹ�lm�b�~�C��{_��J|���9c+Z��%�i��2�{ڃ������X����`B��TI�DV�5�u��IB�E�����x�~~�J(2���6Ѥ9a�]ݱ47]��)\��Pk #` [�[��m��X�sj�g7���&����/�����/�Z+Y|���<e������S�X�Z���H�W�<��D,}�?]��BԘM���!�ZQ���|+�b���j?�d������H�Bk9-?'�9�������A�)�i;�V9�4�g��QOu��Dk`���?�S���a��^�|)(.~; EٛNkN�`�_���A�Xק��Goc�CL����u���sm�������Z\�e�ݿ����`���X�ï;;�s�lx
N�yf���_e���Oה֯���-�
d�������� �0L"2����ã�Ѷ�X�뻡`%l�����p���*,���ӏS>@�ߢ@� eQw���i%��,�2�a���Ԛ�~���q�w�K�v``�8�A�W��SwRۑ���<��to�av}J؛��2���S�/�!�v#􌤙,�o����1�TG�J���[s��4r$�N���_�C�b�)fMg���^)P��H�'��3gμ�Kh�8ƨ2B�a"�\��q�RҤEq9 N��Thm��e!�|����Z��^S/�lw�f�9ƃ"*�`��ttt�p�\bx!۠�*��g���?c�|MP/|��G$���g#ӵ
�w�Oj�k��⍱����L��ze<���\Ƭ�E�k�A�arH���;�0�i����Jh�qQU3�=˨\8�i�$}���Y&��^"����$o�����=�j%�qH1�`o5��|�k��^�>uU�̯*e��R��1�VvEU뤞cL"e�{%�&�~�)�C8>{�g`&l ���5I�i�Dԙ��?2�'{d�w�~�p��b�rFk�l�	Z��xç������a<U(n*�o$M�+>��1�Y��E��
�������+��d2��`sxC�Ŗ�xC䎔K�Ҹ����5�.�C�N�! ̍Т�B�c�A�l$,�,��$�kAK,�Ԉ:_h�y�I	�ʒ]s�@�rӜ����+�LYմ�v�D�W7�� -U^���K���"8���tV��"N���rD����_�`w0݄�V:�o������2��;	j�`+�ǵ�+8����c�/YZ���rB��Z�K�~���lD\kK?6jR��k����+=f-�6���JX
4p�?~�������6t}7�\&��� ��y��t���U�u�����? ���*���c�W��v�^R����*��=���c�ب{��;����b.ChNl-��ݔ�j��f�y&�YTJ<�
v��݁�{��3*� ��'s/���$_Vq����O�J(��X�OIS�8�����L�̌ցt��fc�IA�"m:^6�(�ƎrbA,̚�č�uww���`�噱;v<����bߵ�)uԌu�ηč��;�_he8�"δ|f�ɋ�f����R����O,��b��F�ϬQ���O�$ު�`����w+�SZi�&("�t�g����GP6j���q�ꆏ����U�!0J��Э�:� F2�Ak@XPPwz˷��al1�3�d����{U����*�|�yl�ڋ'�}��,��̽�V�iӇ���<����P�+!� *>!!aŵZ��죔C֫��"�g���se}�,y`2ҵ�����♈繬��ò߉|�z�I[�*e0��!�ρl�����#�x��9���Ǝ��Z���%�i0i| ڕ���gdx9I��Z	E~��Z43�n%k��M��+ ^��9i�)��0���/��7Nb��0gAmijk�~�05xh�J����ʊ u�O �H�1�	=`�~��4W�:� ��Ev%{�7��f�q]k*�m@` �<�:ᒃ<d�Y�$Bn������y��'�����-^�v��j����iXrk��e��=��
�k_kA�� �mDg���Ֆ���T���Q���szPU�P̫nn7�����j�� $:se�LO,|۫�p�4Y9J���e�5�ˮ�=�t��qF�LWc=Ǿ�Rt��k�[::��	�!���	�2�s�f���zHVn�Q ؙ�r��(�<�c��=���,��		��A�,Y��bG��=?<��b=g�;�"��I+��vދg&2Ņ��LZ�>��:h���R�T�5��ʎ����9�Zq�:{oFL���Q��kK����G|[U��3����'�V�E��^o��]�yA����%��ep���~���5�"w&�xn��BEM�*++��*���++�t���>���V
[�����hG}N� �Vj�����s��s��/�z��j�ÇeQ~z3�MßBBBH�Q�aXB�(D�|���O��fDb����[?O��f�w�t)0�mϋ�V�ӊ�kxѓ���H�jg���2_H�!,"��c�e�Z[ooE�v^_�g�Y�T3�2}�:|7v��3��@^�����=�v��L~Fp�nan;��CCC�߸���p�m�ņ�Xu�׊	5y�dZ\�Q�ˀz�>4r'Y� w�0���3)���G�	�/�w���[����@��C�5,��Y����&@��z *˴�/~��y׌�v�2�:�`%4=
!�n����*B1�g�e�/Tg��B������Z�`/mpk����[�2��G�P��B �~�h~x���S$W���p��niQrĕ�����x��`;v�	�����C�3 �;���.�"���'ѠNV1�&l˱����{��9�^gpd��n�
x�	v�gcg���};��w��ࣤr�\��<U [��qq��a,�����a5u�ŦB���8����f�6�L��s���
��7��2��71�N;ԝ�?bk�Hql���X����ʈ�6��z��1'D���;�V[ j�A���ͳ�|{��`t,����l��c��y�dD!�Hp�������f�n�� �/ 
����b�NZ�n3�l�Ś���euQ�e�h��(a�� E�Xy��5̀}���P���B��c{�����'�	`�T�8$�?�c#�S\a`��5vAA�@��Ǿm��a&��1�م�J0C��K�9ۻX�c��H�ӟF���&B1
���n�ʳ��c���J'��B����GRٺhZ��:~��)�
�]�v�3R�ՙ`u�m3V�x����H9,�k��5Z�FZ,�a5���dBA6g�.��
�#Y�[�}^�q��:���r��)'!��������������h,܊�Ϝp����#Ǿ6
����� �+��mutt�F��8���
��3N�f��Ԩe�>���J6Lr�s_���M�'�Q�2W�73��P.NNl�����V���?'��m�"T^^����P�XvycE�ɪ����Su�Ũt�D�`�&^��+�Z�m�\FPo�&qU��xFб�_=ܟ6�`T����us�l��6Fm����𺀾xx÷]ha��?ݓ�̫�n���׶��`����Y�8�aI����ྰ���4[q��W���mٙ!O	[��N�FZ�v�e81�����Y��1ܻ�^��r�����S��p)l�3+���dyE�+p����w%���U��e

��p��S��l�f>l��	+�Y��R�"��:!�F�)�k���:)Ǳ���������m�j�m�J��l&"�>M��}�7


�9$H�:�P�0Ya�S�	mq�E�v&� ���h­�z�X�j�n$�H�	 v2V�D"Jjj{��5�gī���Q[��K��	�w�bo�>Lb�����`���-+�$��ͪ��zS�-�?��FivNN+๊�؁�FӚ[�v�;+ 0<8�B��=aIm��_�JN;����:��h��Q�'#D��ɐ��&&O��hT����tEEE^P$JX 9\dL;M�Kd���K���1pF+r[�#���-w�x��M<S@��j���Ә!}U@7�:8)��4�b7�(����h-� >�	����qk�oΰ;xP҇Mq`d�K�]�^y��x�����HL8�Cv]	Ђ�i�s+�A�A��@�1�n�2�<�(�ܵ�e)j�ۇZ#G�r�D�r��-"���s��It��֩�
3X�g�uWyn$	��-t�f���>�$�\8c��~�������]Re>��~+))	{�!��߀Φ#*cl��=}���6WVc�� ��zʎ��DO
;�Y�oӶ����^�0�3����\�|�5�_	5P8������#�z.��g�C*~��Q�?�O���z�G6>�j�bK����B;ʽ��j@��A���:���wz�Z�0x�౮CT�vtt�ąr�؛\�) o�'l��
���[ɗ�}��ϨU�iǣ@�{	`�
Vl�	��AV-�qr3vnę3yY��O�3�-H����w�X vU=��j�	Uە�6	��D�$N�H�՗��9�a�i\� H. �,  �)��F3�s���&̟a��֬��7ia׆-��w� ���ᪧ-v�255��&���1:�G�V�����ؘn0�������(�t�]`H���y�&Ҭ�E_�~�Ƃ��틲��oJ� �[R�b�GY�����ts�����oǦ�e"s�>+�9Q�f����23�!�J;BJL	�i��s�:��O�GV3��2��`$�r���*�p+�T�еȥB�KԚ��d����x�!�`j������!�1�
�>0,/�1��896ޫ)~�X�ts��������lق��Ţ�$S�2��=fv�����h�M� ��p��1�M=�4Y	�WX����㕭h����#��:2:px�k����o< �E�&ȭ��dLz50��72*D�W�+�H'z7�O��E!�׮i),�b���|ћ��%Nd�(�X�N;	~�_����뜕����1p���se������ p��h�އ�v����|�+\zޖ�oW<�^-��D���M�H[?��f�j0�zS�~��j�� rlu)��%,B��='����ַA���3�B�Ug����?��9����g����I4'�+	�ɣG�<����y����K�������1֘xm�w��_p��ޓ�w��h� � M�¾�I k��l�VN��� ;����	���y�=���f��MMN�+H(�ps��ϟ�c��u���h�1�1$�"���Ò�3S�C��<�b���������ua�	�cJ���t���ߐ��ERHHֻ����̹}�������3G�?oq�qf��@�1H����q}�z·�)�f�8�^i/��`:6��U���-5�6��&�/���X8ۓ6���X�ct�f1�-ja��%%�w�=ִH*����uv6B4���L:d`F=}cA��	~���$����u;��,Ì��pw◥����5�m�g���`R��NΜ�����dQ��(al�c�]��y��ͫ��g8
���� mX3~=}�t��A/y9�HU���»Ӎ�b�Ep' rs-,�����Ƈ�Z[����%��vN��~����R�2������T⹨�	�����ۃ����z�!G٨��:|��,���0e�?�5E��΀�0��\�����y��11���1�g6bbD��-����d���0B�9h�o=�D�fv�Z���X�{��(��\kjs�����䛃PY��.����w�4���=���Z������([:�}<6��>������[�Ӵ��E���b�J��oP��$��Bü�R&�+^�޽{�>}��~��݃f���۞Ţ��1_��El�η3�%�}��+��"���tɕB"�{��tV�<g�s�;� �N��7��k�}�.읁�M1�ZI�<�������V�'��1�71�#� ay�Ϫ�132��`s���^/[Z JP� �D��s��@L��K��},�o���g39���j'���q!!�3�A`pաء��u�ò�,I�!�T^\���I�Ý!���o�r��X}�֍3Ww���(�D7s"��F�����[���#���ۀ��8�h�J�G��UL�HtF:�4"D�	�� ,�e�����\YlɊ��go�6���q�ĈpZ�s0TAHÆέr�56�	Wc�p�3�Ȼ<
�kc��ao)�O>l��,��g��e[��A�l����ӊg�}	�]P�<�Ӳ� �:��e���$�6�sr����IWά�9V��<0����z���åd�}`��އ'�f⪦-�����F��J�Uf-f;;�AV��|�u�aXƙ{�S�Y����z��f��"�X�Ǽ�`V�� ��:��^��b�!���b�i6�����cSv�#B�p�<8�mH��i�賰��5׌�-Lk�J���^����Q�9����ʊ�l�Ӂv�}�V�y���$'� �ʏ��(.l�bx&Y�����Ǻ°�i�5G ���ʿ��B����`_Zƽ��2��_�V��T��hF��ꂚG��t��ޕĮd`�ب�\:�>�xrrrү/��M�t��M��z�?o�!�f]U�Ob���0��߅A�������bj�w_�r���Ǚ�̫�@� �֊��K�ut�O
X�&�m�' q�&E��ܩ��P���^s�!+{�p�ģ8X�̜���6�3����2���@'d�>�#�9՚J���{�d[�]����gk8'�1@H�!<�Z,�#�Q �i�q�/z�����ζ�h��|�x��V)\w�a�2�y�=���X��b��ꆆ�$4ҍaTJ `s�?��<�
�{1�����G����x��C��{���y̆���/px��Uk����ث��z�77fgY9Դ{��E+�[a_��(��khL>��fu�V���_�o�0�������C?��G��4J���(M�⺂�Ʒ�Ko�{��gZ����"�:ܲ�Y]�Rg/��bUY��\�Y�?�T�_�����iuLN�Ǐ� W�ip��y�)i��gx������`؛<��}M�**BxԨ��F��o�85�5�N[[��O4��*�2�C���L%�ōWg����11>��ގG����/��~��^4&�RP�9~5"�Z��&��e�Eك'�^��m� �>P��_���9rD�>�м��7/djOˁʹ�NK��W��*}�n}
V߽��׎��S㣅�z�,��h�8fH��>bӠ?�S�O�&`��zj������\o����nę3g�G��׷�RjU���l?��.-��qr/���(� G
S�_X���\�Htl
X�Ǻ����"�=w����0�;{J�n
j���x�\���
�2@Ew��ġ�/.��X�.݋0�kL����e��7o�#��<؛[��M���N��?�ǫ��yvt\���3��|�"�8��L�|��t�@xż�)�޺'s�]]��<�
;����� �h�%��rMUa��+��+���=٭ ɦ��c�;::�F�M�]���?i���V>����B���t��	���vUҏS^X�������� z����Z��[����x<�Ss�t¿� ��>p�Õ�����q?d��S���u�+�؁��+l�'���j�s�ʖ���=��I7�
��z����{R��"���>�!2Pd���HYq�⏄c�N��Q�kş�RqD<��ӧ'�Tk�4���.EW�sZ���-�>�a�� �p@"�<�# ސ���޺���,Z[qG�*�/��O�/`��?x��5��i�c/Nn-�w�0b���~��@��!���q����3 �x�u׮]A=[]�.t$�=�3hb	fb���<,��v���|@1:*��+[�x�>�l�6�
��w���^��Gz�m}
�*��@�)�t;j��w���G�Ѩ�@w��$�$��ȥ#�������@E"~v�h��=�z|�+ׯQ�Sʒ����!��ޛ����Ii�b�yĞ���,���X�k����!W������N�gO��ѽ4B�6f��d�$SO�+T*���;֩=E��[vD���Z���L�Q"�!_�x�/�Y�w���Ɨ�w�i�Q���W�~�J��C19���Q^��ٱ&͉&e���@��o�!��ʔ��e��
"�YH;��H����@K�6�\�|Y~������	։��⢢�z��ކ=�������̟,�m_�]�7'E�;�R�>�*�/�Rw(k�x��߿�G�UVV�����
o�7-=[�0����py���c��F�>H��X���hZ���ʿC��'��MX_P�R����z25�g���J��"7,9@��G��AQ[[�����x�l�hS��]��J��o�@��!P�79Ih8u�'*8�CN�ih���)����p��C��4�v&Sl���=��8nȼZ���R��7&ዀ�!��=>�)�L��J�R�y~�O�T�o��t�џ�H�xI��y9���x/�`�V��3�!M���gv<��N��U�����
��m�U!�:����j�>W��9gqK��ʹ>��˅����q������\�m�ǰ������v�������C��)��+1�$�cw/�;9k��� ��~�냶�Gھ��{3P����)�oT7�U������Z���6h<�i��%���d��ǚ~�G8���+p
^�.��3�ߪ�b�������7�zh�=\�c��={�<P=Y~��Y��q�6��2R)���D��8��Zc��>^��#bu��}���fY�C^�����{q0BK���'�C���$��}xp]zW�.NN'oo�}�ҍw���P�����mjo�������6�����/�Ic3��;wd2��3=��L.���CP�W��;&�|��X�$Q�����w�Ը��k�b�v�̡�CN�3�Ni&��
�,D%އ�L��w%)�
e���S�^<�BQM-��I���ķ�뮿z�:ܽ|���e�d��Vel��FAN�5x3GS��@�����;$�zA:}���O֓��8�*�?E�ˍ�u����7�����!������� �޾�q�\#��d�����o�I�{^�x��rM���P/e�T�,jyb}Zc�!$��9���I�l��0ܼ{�[�������h9�ʁ��G!M��V�K#��ŉ�H:'G Y����6P�zB,�|%.Ж�\�?4�J�� Y���|p���1cu���ʢ�ᇅkך=��`@��g�AOOC�_5�rr6 ��({��m���)4o�l9m1�V,I8:j����E].��6�� ���C �A 8��P����e��W^�QS���L[|�~��=E��H	��φ1u�o�2W��C���x��x���X���D�� ��� `� �@�z�Kk��d�.2QQq
�Trko�w����_���(�V�D���~�F`��͇2�T�G�ȶ���}��.��̒��6M��O��=�Ѵ���e�%v�\���4����*��M�\6x��C���ܬ.�!��{f���oޘ%������XZ�G��L�G�b��q)<�+�NMM�US�k�{�Ň� T�-�<�GZMfϺ�p�OYA�~vͱ��o��Pm~}���{�+�z*,�/����{�/��9����\sBΝ���dne���Շ m��{-7wh���,*���܍����s���ۼ�4��Ws���o{|d����c�N=R�f˅#�\��jdd4���oP��[E����o�(�K�Y>�<��ĥWw�a�2��|��d=�իW�=���M �k߆��Vbk�E����/�o`9w'E���ΫL��[S!��n�0c�F�
M��@Ugx��v�k�?C�#�t4/��\�
$-�1��l�R��6�o��b)ؽ�V�#���ۚm������
b>�}��<
7��TZ��ԇ%r||�cbb���<y\-611��M}pjN�<���(w�s�$�P?�ɛ�*
�E��Z:�a�O_�r�l�:v<JK�1�`��
lnmM{�rϋ�ϫ���e�c�z�݋NQ��o�1�؛���e��w�#�;8:�hN}�<���9�8ٗ���<��o
2�	�|�W���D��Հ6���@ �c�����哓�.������D��gVev�(��{�\|V[���RS��-��e�үk;ӛb���&�/7g�`?0�� ��'��6aϽ��։�������Z˗/OŕS�򋻤|F�MFFF�mm7���3��3���Ibu�
�ۯ ��.f��͹��#Oߺ�����,]I[��`��5��n� ������].>y�~��T枟F⇂tJ|�6��P��.��+�k����k�^9r���{i]���~�"���\Ǔ���1�>����p��E[�43���Hi|�*����A�azS�LV�%W#�+ tJJ��_zS�'D�܊�E���r��bq�;w��ǽ߾}����R?P>>�1���a�.m���x"+3h�~�n!����ڵ���^�&��� ;��/�~�d�~x�(l"u�l���#���|�R�klhx|K����C?E��B�w��7e�����ޠc��M�4j:�i� ��� ��$5?   !���нշ��~�㛚0���P��~|>"��WH ����=����u�m_�`d������X�v�<W��-�~��/�&Bb;��Fl�g�w/�;�P����~�
���δ�����ڌ�/ޙ��?8���=�M޷�/)2KypS?��s�m	.��������U��oѪ-[��V���pD�}i�1PO½�U�S,���s��X�m�֏�@/�c���K1����F��y���Jv�x�[�-Փ��ӬT�7�����v��I�}l3��G#QV���}8Nh[�9D<���((h�(�L�-֪���oT�WO���_}�o�H� wT$Q���~~�j���"~u�qm�t�~�:�F�������;��6<�����lx�U��tYi_�@l��=�reAs j*��.ޟh^�{'��'��7���q��)[�bU	��(wۗ�5�4�nQ�8qJG��W�үg��A%&��+�������C�N|�+0�Q�_Ɓ�E���������mZ*����+=9[p�U��s�<��,8	k4�۷o�cr����zn������~�"0�݆=<��9Xm�c�TC�̓T;��ي`gh�l�v��IIe�o�ؾC�2�/kI�3sW��F�/RI꼴>���!���ǏV�0�&?z��p ����f7����b�
[��j&6������
�[5��1����?�5���QҔٵ��X�ʓl�l���{��K;����%0ln��r]�0lA�_�����g��aٌ�V�֋�t�������V��~�b���/Gb�0i1�xt�RUS[��~���ڬ�l��.Q�d ����2'�kP9+l6n܈�3דU��R�˿��u_�+&"ף�-�-[���5,@�N��(�޹>a�o��5;�൴�lc�L @�S�[N�:��8�EP�!,]�Y�*�@9�X}fh��~d^v�贝*�V�2DWY	fXX�_b�u �wC����]'�2�:qH�AL�(�3�ZP�xb�I�9��<�'�*��̅!�����dSC���]� t�=&&)CA�j�\]I�~6T�z�
X��(l? �x�9��8H�*y}W����}}{d��^M
	*"mx/$V������N5s��(���C?4y�oL�hvr��ց���Y:b�[�\��0$d��k���`�.�8w.���"�]���6�f#� ��򐈄���IH��g���+h[��r;%e�cmZ��%	!��X�@���9P���.����M�m��ނ����~4*<�-U��P�ņT�X�7��t�K���R�<��kc܌;����c�;��L�nX�U�	J4�dQ� eH��"9)93�"�JIr���$�Y@�9���'����ǳ�Qf����n�[]]Mـ��p�坽�0H�jۧ�=&��휁�#@
��Dn��Y[ZBq{�a�fg�w��δ&���}���a���H_��j xm���JJ��[+P���������/
�j��fh�b�U��+�*U��?v��6����+Xmym��?){�ȵ �4���F���9����U�!]R�m'T�Wl	_
&�+U��y���N|���=�9��>���f1�kN��`�����I��W/�g"�xh#c�w�H!��]��Nyyy��i{g�'x�i1 ���]oϡ^\?_%����U�N��`��j4��U���/'�:�������`Eݰ�ź!��w��gK~��y�
���b��U�����ͥh`��]��G�_�Y@��	�`�.e 5�����x�)�B�Af|�0T@�F�nA6����r�%��� :8}4a�0b �e 6|����2�I�9N��J��E_\�������|Ϯ$/J�z?�J�� ?�J�ؔ+ @ި
<�lL����뱿(a#m���[{��{���˲���v|Y�� V����Q���}o�e������ 0C�����ǏM
��d�z����g�GPكs��)����\���E�������|	�s�y{Պ]�[���Z{z�C�v>@D��eHp_mmmD�C�����w��6�MOW|/n�ng�#���y���t~��:���2������N�@R��Pel���k��iUxG�S<�q�R�2�nDd���>yBaT��:���}y��ki;�J��cכ믣��p$�S����F��Ҟ��iMM�Ʉ �9t�]iQ���:�/����uE"���*�F��0��9#��ϟ?aC@���8��g-U�'���g��:���n�I/b@� �3�:vI�[���|�UFc!lO&�����4B ��BqدJ'=���p<�1�齄�P��~�/R���{��6*q��!���
i&��%��LNN���%�7������k�G�P0�a�|��q��)P�9|������@W3���)A%j3�S�JP6��i�N��.��8�~��;^:�y^h��~��HB�C.X1�C�i�����2��� ��ځZXc�[bN�� ���).�������Tٽ� �F�JެP>���iH�����6g(������vnT�@6C��<*ג�3�E"��4�&��I�8��N���-J �rO[;rh��Zg����g�4���^}|#�q!�8\��^LB�����#�������˗�QB�'���z��Z++,�A��&�QS�_vP!+G�vg�7� B����Y�j���=z�Cv"M�VW�?"3���}6�<�/^�B	

B�70�)������(���1�����֚o���a!hX���@Y�77�T\z���M���P�1�40�	��KJbQQBX�� ������HZ���F.VQ=���.&	
</�êCR���`�=�&�}}|!�� ����|ow�9�n>��C�*4W ,���dj��&����� !�h߉������G�,L�z�v}�B�c������[)�䴰�_��a �C,,,J��-āW�+�S&�����g�߸���5�u��cx���;������
�K��q���
,�e�r�<(����.� �x=!/������~�CgExo�t�Tո. �a�0�	@�fg}�-�30R9S @�����d��)��Wƕ;�֝$um��i���W�~�������~���>�}�"d��e!�s´���yN�����e��C���$����d	`>��ɨ�Dc���}||�߁���)*I";�0�����L�"��zDRw�.G���@5@Zα������QUh���C��/�F����oW�TÎa��Xd$!�y%�H��7��6��\����G�3�s'`{Z�K	f��N�� ��}� �z��������\u_���@���<H�ˮ��㳧�����.��uN]���� D�L]خ�اpf{m���˰�"���a2hJ�ӯU숣�DY���*���,~��^XЁ`�mt���@гk����*(�OP�����yRԢ����A��'�؈���� 
��z��8���M� /��"��PƐ�l�wmmm
�hR����I)�Q:�6	DR���,m#�XwC�}Pﰋ��zK�T���sG4����5 +o:X��a{��u OJ�����G~�ػ�N�		u�·�'�В���	,G���|��
-��_ ��l�u�����P �@̀��@J�������\t2Q�@��KT\��I�b2�,�]e��wuYW��8I�!�I
��A1,,,%���7>�R��na�Y:�F�;X�E0�`T�t�
�oÛ(���;�Q��u++Y[[kf�ק�Q����y�+ѯ3Ka/bW�.gZ�S�Q�b���Y�����,L�'�n�;:����5�����_r���q����� (]J�7l���$Vo��>���y�����I1�޵vvj^؜t����Ot���#�� �!1����$$FH@X7����v��"���'`+� *-�G���F�p���Ā�-D�����6M1b�bG d���C<��M~"��b�:;;��v@�������O�āG755��O�
 t���г��wDxxZq��z-��x��ߪ}0���>,�t���Tom�Ѩ+q&M�$������9m g �O��i������;����`�C:����|
P���|"�,������ ��_�|�����ݎc=��;�מ��\ȫ��Qg)���r������+*C/���t7d[�f����>Ϥk�X��}� ���<����]:�΅Ċ
������ِ#�'��陙�1E��X��2�q\]u���=���a_��A4Z�L�F��sڀ�Nt�1���~���<z���Ψ��En�SC灷�X�~�n(
b)B༯7���:��&\:hY�br'��L��5�yp��7�8�d�m�YW`��ɴ�

bW�8�X�Zs���x������?�u*�ב�k��<��h�R3����[0٭�BAF��&lv���l��X��.�/����ܡ���˿�P�ttTo��;�@�Ng����qη��� ��� ]
<X޻��E	�_�B��+L�@��y�K��$����%�Z �28�3S]�_�*�m�;vjdh�))� .��׌<&�@���)�vD�=��_�5B�;B%�9���<�[������~yy��Q�0�.|�lO[]�\\K��\
�+��
P��a.ܵ�Z��{?�܆|�*|�
}d:溓T,�-�AA���<��OX��RIE��크`в��R���-�&��bو�l��"��V����C²xxdπ ̰l���%���f���o�����Jc�s��?c|X��������(��cA4�ar����J����M4�ml!i��mӐ§:�ٯu���H��f�='���cR���Z���.Ow��#��:�B;~�WS������f���z��nʒM2��4G7�����%n"E��yy�d�c�Q$��� �P��}��G���������y]\]��Ђ �:?�)*�8�r?a�X��<K��fWN������g����)�<�F��*ĻթBB"�pKO!��㙙��.���ʤ�e��l�i(خ�����A���ߨԹ��Լw�>i�g��C�=|�����@�{�uw�Q:'K<G��	�/� R^��F�Pc���<�y��Y+��p��3�;)��Ϥ ���3�a���H@D�	0u�:�%ȝ��,滉7ˡɍ���Ȱ���#�BK�Pp�Ѻ@� 8�<�<�Ȟ4�frE�L�{R��p�&�@ �^������n&���%�������yy��*�n�7w.8��\������6
�j����kddT�`�v��y���a@A�7�c�VVm�M�	���o��x���7�F���~� Sw��Y�%��ж7qm��y����o�r`r{�,\����%
�V����c��2�E6[O�[m�.����?p�YH��< X��pq���A:H��O��Z�es�TX?�r a��x���A-Aף�����l'�v�w.7x"""Rޛ�@����ʀ�p��n���M�_8�R���D[�4%���L?�@)�K�$bIm1�"=M�u{g^���J�&E(��L�&�l�c���*kȘ葟v���D��@��m��F�(�%xP�r?�㼿��x�/2�	#�^|��ׯ'�6��77�	Ύؼ�~�3�m�r������骓VO��)V֎��ʬ�����Ux�a�����߁�]�'�B6q��$[-()����S�������h��,�����^���<"��o�ʌ��vX�/%9��˱3@"���tD
�ɓ�F�n�TNB7t'��P��{ L��/%�Z��ߑ^�؂������] {#��^�{X��\�Fx΍��J��f;	c0��x ��?�w��ϟ�a2|��`����yҺ��84�9#C� �I��۷W���VQ��V;r�d0� �È��[c��޸��VUa�n3]���D��I������֖@/�\4�K؆�S(�6��*�x�RC^�����D1��Pɀ83b� sss�2/ ��HA�w"�L����$@
X�F�`%�K?Xa+�J�JX�C��q��DpssC�TVV�&NM�@{x�VPP|43�^2�E���\(߀j����x�a?P�0�7��W�8�q�}��Pn��Ʀp���lⱍ�? ?�`B�\o�	!�(LI���խs��%�}/;��Xܰ4���-������\�P��b�.�FTF&n�U�
�L/��^jr��6���<z(G�A<<�_�,z�%�.3J�I�P��N �:��Ba���m&҅�ZzzV$�%sP=%%��ɶ$���p�27��U��&��0Q��x��VW����B�J0�23�@TE�`{��zmw���#� ���HK�����^CJ�+&��@�wi�ۂ��iiJ�(��D^BX8�%��˙��@�7;�S��#]jZ65X Gz��w�%��2���cv�U��M���__�g��T���6�� L�?";P��` ,���G��*�i�Gڒ�����qqp?���aA�S�ɟ�
UI��XlV�Z
q��uH����g0˫o`@H/ANL��p��=�a��#(0R�ٰ�`��T@!y��L�r����|�e'�ԫof�%����,�92b<��8���1`_t��񪦦� ����^<��Z���g�����wO�k-tc�K6����LtW�q�~eK�H!x9�%w�����&Y��nOG��Ȉ��B�H��F�l�_H>�� /�+�P��Y�P2Y��E(�(:DA%��R ��Qd`߂1*� �A(��e�q��_R�!9��!}�~���0l�
�Ɇ��ۋX��.a߳I߽o ��ȭ��=��m��-S��W��[Q|(�N�Lr�����1�(K{��Z��u����4�AQ3yI�Q�j��w�H�"yS-0Z(P9ЅK�|[���A%�>����R�wkO~٣|y�l��g���Ծ���t�`Z/�cկ=��U���������W\a�<�qp��a�����Ty�ޱ��Ur����G�b^�2���ֹ��O���^	ȸR;�} �p�W�V򨯐G�
h9�wu���,�z�,p�#�+��lTu¹8��jj	&j~o��P02oi�^R�Z��չ7t)+�G���š��Ñf�:�QYu~���n�8�]3a.v�UGZ&���������k�@����*�x
}���@\��z^*_�����4*	QϠg�c�_R�X�L�85�϶,%�!P&���R8�'��u�ЫW�Ǚ�O�h�;s&?�3)�j��֫Wc����ǘ��n�_Y"٤�:�R���#�L�HY�����\T��cv`���
�:��<J�<���ϟ&���y�h����;@O�w�;���n*��JS�qF�P?ф��c5?��?J8:z�N�4b��u����N̨�JI5���G�X^e��˧񛚚�#a1�)�8VDv~h�'x���#r��<��H��NZH�pce�`�k��ꨓ�r� cɇ�L[������� 3d��y����������Ⱥ��6:!w�e?������\�+,�[��K/�~$j�pp�<�)��
@�2�cϨ�`"�Zb@��o�9jhl7�c��>�����e'� Q��������|����2ñd.@�h#�8����<~�D�Ƿ��V�5ӧ�����ob�=��{A�*��W��^�-��VTF��gs-�K@���ʩ����Hy�<�+ѝ ��e8�E6ڀ2�����N{h|zC�-��z��Pz� E-6���3b���gu�Nǰhuwz�٠)	Ơ��dm��������:j����Ð�I���U�|!�H�kR\QÔ���M'�I�d [h�P�.��"����vz��6�!:S�Xi_�N��2Ӗ��G�����[k�����ݲ���RR)�s��?W�OHX��[hτ8e����4�����r�dUWH�U�0\(l��������F�%ÖsM�x~Zz�.3�����5��"�$�5���f�\�8w�}�a'GXXY�['��ݬ.��ṈT:�[~�I����jc�qC��n�L��,���> `���[F*�TKIiEF�]��>^~��φOL�h���D���������*�2�[��7��W�5�X�K����_�N����5�f��<� l���]4�'�F�I�g�$:�4�����xԘI��]ӚuM�Q��/�a������L����������E�Dfٞ�A���堠`k` �~Nj
����^�ee�$��5�D�z4�(*!R� ws��Hw�o��C:�fGT R���������5�X4�Р��#����Q��i�j�q֥�++,��]��/�={6������rM�U�x��XD) �����LN���:�8�$[WW�"�㍬>�X*f�v�q�T�@��n�ϟ���Y�����Pє&B�nX�}kVm���XE+Go������X���V�p�邺��*-"�?Zi���y�J��d��+�x2�%��Y���X9��c ��ڣΆ��<�@��7h���\dV���7�(bN��lh_�g3����J���G�B)����J%�~�x��������sjD��+��&�c�B�ވ�$8X�^W�Cwi{xp$�֑g��`(���AQKS'#�O��^��yTuG#Ͱ�s�"���p-M�E/_�����5��ε'�YB�x>��C���|c^v��z����?)�f�!�!�o�jo@�y�0�8�bicx��e��\� U֬d�)Փ��<�P�֪�Jߒg֘kۤ�I˦�JϾ��Q��m��Y^̗�w�����/O�Dc�[��,�na��:,�C��GS����[��o��Y�;M�^��±�*�:����;c)u1_o.�1��������QQ���%Ml��/��-TU*�~.�K{n�p��ȑ�B��.��Å����,Z�u��5�.L�nIz~�h}����f�SD�u-pu���XO���ڗ�(_����pA���L�C�]l����LU+�"l��������ѓA�_���	"��#���%��2�2Ӟ�JA�t{آ��),aT/W�,�������;��
V�b��RB����Tq�F�s��{�޺.������?e�)��b�������t!�D�1P΍�*?�r�(J�,���g�Z�=�����ɺU��F�~.�p%>�J���`o��Ʈ?E�¤%�!6�@Yg�"�jx��խ�G�f���Xg���}����Q�������	�2��J���S5���~���U�%2���^�����ʛ�hS t��*�ۖ:��*��ٓ�1m{_=�\[:"��bar-��NH�����ď���"���D�d����s&ǌ�y�t���v�66H	����c��h`�m�y|�~y��ܬ�oV('A��>=���"{���ykc�fD�Lji�A�o4�c\���kn�Tт�4���M���4xs��rx�4r�Sc���Hz���!� ��]��L�C�O�^W����b��㛥O)#��Q���9ؑ��Q&�ӓ��s�bģ/��e���"ɬ�'c��m�%�a���l��wpbS��K@�&��N�gD�)�w�k���V�z�/z2l8��R��W�M.�ķ�����'	���@Ȟ��8�a3{�9��ۋ�M��S[��-�WKǵ��y�5�_���P�Zk���VYi�*��W?1f���!��*m��3�q1*_�\;�ؒEg���X�:7�q���/
sH���9ѷ�\��6V\�p��Vʪʓ}����ˏ5�i�NIW]m>�� |��� 'N����sԃ*�$N�<�=b�;nkg��x��1�<UuY�X�V����oDӏ�dwť�pڃ?Q���Z��*�4NB��=��Qǘ��4�Tš��@���4�}��H%S�l� �l��lO&���њ��	��'~s���Ri�|���C�w�37�$�C���Td\yu�_��L����$3YGL��C���� �&g>�.�����)��&��0>�(�⸓���V����XM�+�+��0���5�&����Vg>y��o��*�[k	`�=��_����W�N�,����j��O��CT\�����Mwl�=�(���%��>��I��s&&�v�I rJ��U�e�k��hT��?�(��;���n��\���6[G4���z� I��礖[��4,�[�;������<��F�&Bi�.Gww��[~����0\!�fUŃ�7v�T>2���Y}�i��G�:�}��=�P F_bT�1��+��}]�i���,:�C��]b�����c�^�^lޑ�/�.������G���l;���4xm�6��yF6�܂1�}�@��-ik)�%/ƍ�#���O��S!\��썔\�H�Z�D�wG��/ֺ�>P����Ko��"��v����z�R�ԸH��D����%R fx�x��6ְ[,����ۢGC�xA\<���[�at@A|�EEͨ���_S�@����e2���l�ӯ����;�;>��C8\��5s3� �R�!���ܜ������_���w��}�:����SL8������Ot�D ݗS�
�^��Tϰ�2�w
�9]����T;��,P�Lc����,�BV�2����I�q�իW�o+&����b�4ClR��$�"�?G҉)�{�r��{Y�o��r�������IӘ��:�Y����Ԋ����
��1��R�@,�G �tCW����Q���)��9'�e��U��F�IQ��Mܳi�wnX��P�����T7�O��؊4{��x����qn{K�J�^��y�Å45Ӯ��:]U��Eg�@'��W�e'�l��2X�i���-杙��ۂ������9���[;N�u��}�:mM�E�"�>Tz� �����PD"���S?Z]��IN�W9E7��{nn���'U�
=�i>�J�
�����2�J�&�9�'� �J��a\o��O���y5m0�&� ��7���7JJ�p|���8P=V��^z"'��п���g�`�`%�(w���%��W�/*�",�rqQ�?��z&�ag ��ͅ��k�q)'��h�µ�f�5һ��K23��u��%[������|+�5p�{Q����7d232��v�v�/���[��)/��l�잸*�βQ��31�;�@J��\�@�5���ϬՏ�5L\]v�Y��ز�9�B ���Y��7�61���D����ۭs#(���
9��S�.���.�;@�D� ^����w��=ȱ�:$w��V������R�=���hص�Z����IY� �h7-!&-�(M�(-�(M�-��&�v�/*Pb�Ґ��C�1��^/'m��Њ{Yn9�d�����LD�R��R���/���w�%���1l��2]��'Mt9��k��n;I73�2� ��/����S�\f�x��_�]�M�������ȕ�"�l�$LS����{i��ɋ"�s�;���Ҳ��m���`0����2c�(�,� `��9���-Շ���������|�+{�ό,���9���N9$㞸t-�n�,�P]�zvv���W�	f�I���蓵��)����Ӵut
�?['�yb��hh ��5ͬMcS?����͎���K>z�S4���˞z�X���p�<�w]� ��5N���/���)�8z(��1��V�b�7YY�Q�B%��ea
�uɯ�`h�	�]�CT_��~�� ��U��Ҧ^F㫘
��h�$}��V�o���Y&����=<ܒBl�h�s������jk�^X}��C��_cA0Q�gK��{���iOZ�@���}��aɖ9�^\�p�Wc�P���QVV��	->[��(�|�gB�#����	�Og�����b7�ucгL�+�9��}�)�T<��uO�bN�sB��Xl�ᯒ��/o����1%�m!��
��;��[ȸ⧶�7]51�on=ۘ����,�Jc䳛Ӭ2����z�vR'6�34�;٘ +߂?5�h�K>n)�I���U�"�ۡ������<Hy$��]�?�b�*�V��/�Ԇ�G���4���#��/�đM���$x��x� 2+e)Dqc� `�j�� e� i��o����럞dm�g��Txm5�Y8C;�/��
�fs�Ԧ���N3]v����+�|V�К��s�<1��[W)�rv|ثG�ir��<1��~?��q���z ������'&��K�H��iӎ	tN�<���C�NJ����B�#���qx�l�:���W����Qvz��}��lE�~x7��@��d����T9�R'v��5�x�ڼ��1b��sҳ{���0�SA;��ʺ�Y���o9���0�W���ӷ���w��7�-滖{e��%&�� X��"�;���<���p�g�H�v�H?�->����.�o�ɾ��xG��RrTǫ�R��`K��8��u�YI�)F�9�ff���v��������q��,�ʴ�N�D��R�qW�y���>���r;������__H3����:V��4�ބ�~���6I�dO�-2$M�����RN��.���B�U����w����'ؓ�6���Q����zZx�w!vn�*����s4�v����fD]`���ä�s��%$o��zqf�?�o�`t�n��f�̅�5�U�.H����!=5!G�"6]g�"������o������^h�{z{~T��d�����T���l��3"�/����,�#�Wz:�Cf���+ր��k�1���/�n�,,�3*�s�ڗsm�--!���U�<R�EM��Yg3��Ɲ�Vwu�\/�#��/��B�trr�'dǮ�m�/�.R1�F�b�n^,������4�v�<����8�#��x���c-�d��k�4?\ln�Fk�q���|?��{���|�������P[�2�d�s�����Ǹ�_vu��`|%��`�b|IK9�>��`̵�k�*��TM��?.��XЇ��"���±O_T\+�c=�H:�N8���o�zSN�����\e&#�����.��(oc.C�-FT!�[k�D�Q�Cu� S�>M.6�/�Nj	*)�c�y+�fљ%)+�MW�bW�f'�'Q�S5H~0�	'm�j����=��[S������l�K���mOr��ƬV�nJ�vdA$ZH���@G���T=.k�F�K\�ƻ�d%}gV�MԖ���S:Cm5�
��n=�[��9�t�SNM�gнYgf��ga:d;B�;��%���b�=,:f��T��x��1i���/�LFE��_��~������?�}`����0 ��3�v���Ng_���ם�y�ʜ�dZ��cF�r��bP�@�����@�0��~0�g�c/���h�r�̌�t;V|�o�U�uq������A�v�zc�u�4%�P�!G#��gg��d֫��"Ͱ��g
!؉�li������+���60�k�3���gy����y��`����9|�C� z,-W���W���H�I/��`;��?:n=�3�e�h�1B��z���`NY{��6�9 *��d �`�֖� �Ǜ�h�ء_]�`vL��g)��SVL������3P�.��}
�ea�A��\�j����n��`��k�J.<m�	�6������Ϩ�؃����������'{i`�����өy����;��O��k���8�s�f��8��B�$`/[� �澜C��h��+\ݮ�y�N�Rp|�����xjwt+p���W8y��O]�S_����Qv^ǣă@���<�1sU���ypg?��Nޚ��$�6{���v�9�����u�F���xI��hifZ�]dpP�n���i�1�R��G=�:N[,���β�q�����a+绛kg���Lk����<w���<cc8[��;f��g�v�8Y�.,��(&*���j�5�!�D5J�l�_�~���﹟
㓀?.���3Łu+>L��=qJ�
Ӳ�޻�?e�QL�+��a-��әҢ烵Y���v}�4�`��F'J��K�S��*����8?O��.�������2k��̺P�D̔�P~qqZ�EUb�"�I-)^YzN9�[4�Wb(Ki¼i��}����=TVt
��b�0Q��,�?��hc��\85��c�J��M�*uވ��"��h����^����� ��#ƿ�߭��0yasA?4�"��y��Lp�1�t��|�M7@.������g��#�fL��ڴV�5��
&�/6����� ����9�՞),D��#`K~nq<��N�����=�Q��r��3�cH� ��v����f�E��0����3�e��<�nK�r���|CߤO��_)7^wI�j�T޷wޑfπ	,�9���VPP�@���]W0:QIOwBE5�t�ǯg�,��?�d������Ga�����8���������j6ݸ' !l�M�'V��J'(6z#;O i���δ���q�̀��j�P���R-g��b6)nҐ�KC(�e{Պ�7��������i���L�6K��y������)�g��f�����#'̵Fa��q��@���-�P�����a���q��ȇ���u����8�T(�f4�d�h����R�vܒ	�Ɓ'}}�v���lAR�F8K�D,���ރ EuN&�4�� ��72YN�ӳ��֜�e�)+��ĝ���l��7���1�)(�7��V�}����,jy�1{����TT˂����W3�-��9TT9��D
A憘!^c�Q]����2�`RI�����F�8�s���L��x�.��";Y�;O��X�Q����t��v���'�J3�b��ơG$�ZE ���p��E����ƫ
�pٝŦ�&�z��kٚ���{3�ן{�:��n�j0<8r��}R��K�n�4�P/�Z ��yx8�D6#����3��+d��T=d�G�2���^c����8�P�u�E l+A���z�Ų5}�C]��ʋ������C=��oő]�����2���\��xЉ�f����Mb>N��P�������e�C^�|��qB�I��StH�9_��\A:.�kR��&s��0��؀���Fk+��9"ɺ =Ҽȗ�h[iy�����je_i��l�����F{�+FH�*�9��^�iŬɎA+��$�h:x'��f++��U?�v���Ii��������I���Ur"/�r��zfM'�IM4%���e��jYҷ�e�7��q%O�Ctן���%.pCr��u��>�B�� &	�T�G��P�b�iv�����\A,�l�Ȩe�n���1o��}6�$��t8[�e����{Ϣ����Izr�\/2�"�3ѷ`�'����Zv�;{����7����W+��%	>��?7Lr�X�!V��g�.k����&Cfe�v��ۮMuK\�����Uq�������?���x�B�� a�?1�T�OL!�Uo?���MTU�lA��Y0�`)ջ��ie�o�!SV���kb�H)��Qs�D����ª���kzm�_z$+I#և��W"{����� �e<3��8z�(\�:FM����Q5fvr�����QK�tA׮ )��$�c'a㙾������B��������Ѱ���M&���{|L��I N*��n��Te��@��ʄ|\��rj�y�	��;�<�]�Q�1���ǽ��JpWۻW�$NĻ�.�,��hx��Ӑhb��HGJU�*�Kkp����g\���]8�I�"��������t����y�i�ػ�J�<��y�&�!�p�*+��BF�[a�v�xz�6���/i*��Tz_�f�307�����P'�V��63�ʳy��S�Oߓ��"����#���2���kpv�3<���3�:T�x�v�JџM/����A?À`�q#�E ��T���kjY�z������jI�t�*�>\d��
I ���o�3x��_]��B]j�-��УZͽ��ٹ���,�R���]�f�=?^�`���<���ߨ̓?e)��R�''����,��u�|���
f��.;�}�_���J�VQ
��yrFT� T���͗�X_<ͶQ�oRà*���W*�w������x
�s�&��	g�M��t����;7�!�R�g1c��n����M�F�����׾&N }r���@��i
�Z�x��N{C�'1`���Ϧ�95��Hym��<p�ј��5�/>�l�R�0�3c�)ݨ�Ȍ�<�� �`�����4 nIea�?�1`VEX�ɴKL�b=�]���t{RԴ�=�r�7��V��/�#��a�?���c�`4�����ܽ8ͦ-̶U_iS��2�&�geLo�n�g��Ee�����9�0�J�&�'B{��=y���Zf
��2q@T[�Z���lR�j���;�k�ǻ�dߗ|#s)�f���ꆪ���O'�m~��Ɠ��.k�jO�)�:��������k
�P�'�G�<V�ÿ� g���y��S��SN-SK��-�@��uD�W���5Ͷ�?��FW�r�Z��� A��c�6��H�T��Mʯ�D��a������͸���)��IQv�EH�ՙ�TpZv�����[�!��7�)O��
O��ʯ��x��u־�T���`���o&����������]�b�ȵ,V��Afw�o�!�⾮W��.]�
�aQ}���(S�EQ��) 5 � �����B�մ���

��?F;�:)y�Z�֮I�Ƽ{����&�X��ĩ� 7>�Y"�k���9L |�c�	ƣ	&�)�Ƞn�������6���n�Ɇ� ��ȴy�X��V�@�Gk5�)�L�¦7ަM}�c^�b�K�4�m��)�[���B�z�TG�Z�о65-�01�����Hi&��h�a�iB��G������Ezp98r����/9t��VL�U��������*D�Дb�9��7��=��69D�g��_��)�̀-��:n�!I���B�Cj<�p���s0#��9�.
��/7�L�}��Q�M�*�G�c1�]&(�_'*����-��{NV�o�@i�QyPN��o$��ef15����ӫ�M�k�
����s�Kmg��L����!S�4����"%�ͧ$!,I�
�I����Db�ru��=���g�w@z^0]�� J����>�c�B�+�e>?ʯqFw���[�ϖ��fژ=�� >-�G��S�W��oɓ&����K�`�NX�N���zRP���9�c�J���\���>R���;-Ast����wx('��Y�;��v��}�0A�s�ӎ=�r�FJ�S1�QO�br(<�S1��ӤR3����X�[��F�[�H�X��7�r'���n��`��.iSL���r
3%���w����	u!C��m��ÿ(4������pz��0u���gJ�F����R*�M��M�x��yk�j
q�݊��h�Ĩ�qV�����^�?Z�>��5��":��,I�2�۫�w�ϾT��A'�)H <X@�%���l/۴a,�h"l�VUt�ٰ�c:�j���5�~攐�����8>��[���V���	9�W��_C�x}lz�Z�8� /��o�U5����"���j�*��	��9�����6�j3�u���UC�mZ�B�3�?�V�9�=FwH�sڋ	��`Z]����ȣ��ڱ<�lt����i_OO+��"uo!��.��Ƀm� �K8#k��f;�{s�|j}pl�sX�JOM@��v}�
7�2�������K��c�[5�)�򌧜�]�������S!~�Ie����#8�p�sUaLLL;XY�n�x�0dYC��
uo����;T�d�m��l���k3�CL�5�����Z)���.�o�k� �T/����m���2���o��]�UqUa��T(��{.KAUV�<h)�l��E9�R�{L�:O~x����A��Y���,z�Q��[As,���O�o�
1�Ƕr���W����v�>pq>���I^���uLP�}��ѵ��������[��_��|b<9�Ҹ~bSyB����t��VF�`������,��T`���r�.��igx�4I�}�SA"���$�rg�� ��yUL����7�v�M� �����S��ՅŮ��%�D��Vc7�nKS�l:�jLCD��p�t�
�hpX�J~��Ì��C����<oG���u��A��/j��'
*|��L�E�.F�JA6��f�*�.FG�~=KA����M-�L�{�h�}��/�y'��� w��|N~ /�+ϱ��	�vn�M��	��9W��mzӴR;�U�Pf�lLJf��n���H�IT�f��0c�bBb��>f)�kS�c���,�w.�U��	9�B�:�>Z��w#̀@���b�q�E�M�J]�c��l��gչ߻�[��t�xٌx�{�M<�UK(т��1���8�2��G�$�:�Zd��Iz��T�������,�#��U*+=���)�j(���]�LH�o9�0�̰��Վb���� ��A|��A��}l�*�V@ ~w-[,��tFִ?3���U�lz�����:��:������R����$����D>���zN6A]�
�^�QIЇ(Ed�Y�aRS�i���7u�ƙ�5\\Bb��?kve<�Ol#�X&�10հ���@!{�=A߬����}>�m!��H�y8}�<�G�a���	-���熛I�^�1M�-)h��-�3�-��g�5�5�O|I#)w;l�� ��?u<��,��~Ӛno��E��]���� n�g�#�WI��������Ku�
���\Ӂ��I��i�P$I��뤠��;@,���8-ױ��iJ�v�Y..n?�:��?6lo�4�e\�=�hͭӾk�'�&JU�����6����!/�q��p���,�NG)"�<��h��������#�����jfh��Jf�l*�[!|A��� �*�wS&��>����I�x���tg���f�k��w�[h !��:��O�^�9-�$7J6�O��v�E}�Bd��hB/ƇormR�F�&9�G�<c:�ri�3p}/f�4#�� i�*j]��YX}CC�Dٳ찲L�����Z ��ʽ��Z>o}�Z���orr�i�!i��\��ߘNмD������+-�: v/�m�H��!A� �X:�{�]{QF��BO���-�u����'�U����7�RVF�PC<�o��k� ��ş����Wk���D%V�2�{ Bd�I\s��R�F(�Ó[��� ����7�L�}�nq�y<|�i(�W�i��������g\�����b�+��>u�����苫r̓{�ȵp��&��� [^f��S����:��$2��F3�r攺�����}7�R��1�G�����y���������je���a��#�8(M[dv>��s���*���1���ǘ�vw�z�L��ti	�x4*�[XNc�u3�M�h�Q�f����	��;���%�o�g+Emi��H��|���J��H��p���M8���a�G�k�C�G!
�����������~���Ht{P#����V�|F���䯑�R�|��[&����%�Y�;	6��@+X	LI�� �_�c� ��j�q�qFKrP��_���g��Y�������/M�ca'K}�����u|��u63������ݯҋ����^o~v�"{p��w�ɞ`b�$���	��Y�lyt�L�Y�d=[z#]X0"�>�S(;n���a+Ol˪��=oAp?an���Wt�+���q=�b;�Э���TT8KI���Ǳ@���3v�qU�)4��o��n�c� ;��-�\�j�\��D�8}<��d_ܴEURP��\JW{�4���U��=�9_2�RK�@���������j�����ɦ���,=m#�����m��Q �3�w5�o����<q�R����Y�.�L����*v,�����h%R�a���6����Z�E7#X�mZ���.��p��Ն<�4�ns��N�!�0�M�`Z��0^�0���M�r� Q��n�������������ox��D��R�z�B��l�'�z�8�.��ND���z`{[�hoYd��
�1�=���/��:���M��R����(
��BM�D�$�%�d�5M�B�ވ�gYBeI�d�ٲ���;������3�y{�^�ܳ<��{_��)�y*B�f���K��������F�l���IIIFj�ed��߱��ח����Htkcr���X�^=�e��.|��� ϐ��e�ofX��Lz+��x�s�b݂gF�%��;<�ڵ��*׮��H���PMM�!��(J��Wod����0����o��&k�^9�?���Pc0��{<�\g�,��W��}�Ҫy�c��j�ո	�lƑZ]�u��n��Ƙҋ������>>uib�1���� |���h.ޯ���y�V�鄔#�I��r�u�᳻4D�t�T]k3;���������Θ1���v���ҥ|k������Y���u鴤۠4n���b���%����}�z�#՚����B���� [�/u�.&&&Fmd��}nӍ�T��d�l�k��4>Z�޲�%:�bb^$'>s�v~����������T�.��/�n���ԥkH�~�������d�	6�#_i-j�di�L�~���9�PR���࣫C-�&3�dŗ��Ō����Y��1���.���\�LS?�k��K٩<�N��h��z�7�Y�h��o��M\j|m"��%7��vJğ���y��Y�ً�n�)2�;��������"^7�:������g<�F�q�)~���p&�"��'�Z\��<g�6��1�l�����J9S�n�����W6�j�Ƣ�j4�_87X�LD+���tkLOO4ۅ0��y=�Z��s���t:`�m:��t||���=I�Ul���.�����_��s����ӓ�����o���ï��ދ���w0G@�.���{L��q���W�D(��=�s���/���=���];~6��N��/w��U,�n�j�d`⯕��.�Q���r�{zD�����9Y�-vx��z6 �%~aҚ��9��RJ�� _0��|+��c��]Z1#�w����5L�Xv=zd���B���k��,�v�P�Ն���v��5�w,;l7����*7#������q�y[���=����[��ol��X�����F!�4���*�OT�;����2��ܻـɩ*ߎ~�H}ˋ�]�@\J�<��·� Y��J��wzys�ߟ�ΎU�d�<rƦ�V|��]�j���dq��i�l���u#:�����M�ͫVX�V��Nc��_�����*/`��}Q~#X}��3Y��f�l n�����w]^4�o,;�`�_��6)8�:����@�L]uL�^���/Y0�J�~����y�o�bzƇ\/>��� ����=Lo��!.�=&�-�����+拄{��Wy���H�o^�`�ӿw�8~�g���6�:���/���Zt�*>�\����*�\���:rݰe�|����c�E2�j�.	H������ᙙ�/�}g�9�M�/�t��L��,�En�2���;�&!�c�3m��@�v�O��y�s\�t2�o�a�K�2no��-g~u>RNf^�������m��y~hP��������
5^�������%���/�S�%�r��mL28��-�_S�-}`5���l��\��sms���#w,��V�[V&B��Kt�Z'd�c��@QF�Pѡ���?d:�?R���Qxd>O,+��k�[L��x�8���,y�n,�h�i�!����~�����ꐐ�f�a9�n�yќ���,K6Ez���ױ[ ���
�\�xHm�Ȼ%�

���q���vC-�w�`�9�������(��)�k�~�L��|c�{g����?�׌��Ͳ�O�j/�tx�����=T�	����F-ZC�9ӆ�>���Ek��ۜ3���-�r��\߇aןM��\G��au�G�-�7��	d�ճ�ۏ#ڿ�i`zd��ЏG�wx��άʙ�'& 	��#�k=�dr<ȱܠL[�*=ykD�,�@҈۬�����~Y)W����.r�,�낶�t��8;���ZɆ�S��^[!7�'��?7ƒ��a�V�.�g����������ٺ�+mQ�v?�8�{�;��}�ï����*�X����W+3�W�i�l`z�L�S�%wy���������7:\F�rOrΙ�Y�cY]�A��%�IF3�2�i���<#/h���������Zﶁ<.�o�s�jD���SAY1;��s��f&�����"8 �&�*�8�rGw���Rg��m>=���]�-�-O]�9�x�i�SwG��ɱ��(h��p��Z��%�xf�~Y����_ڜ�·�bW|��?�<=)��]�Z[��M�,�"�BdɫrEO��aW�>�c�� ���Y�_�.��:J>��z�
g�9����tk|�my`|���\c����-��ba�M
W(ᱶr�cꔹ�7���S4��*� ��E�N1ky������O��>������0�^S��yӛ�Lҋ"_@�zmj��D����j���_[�V&���}}�.ݬ e�쥜����?��h$.��8��*���:A��;G�\�g���K1��*�U�w�o��f,~����Cf�92�-o��;�q��R���(��e{�E#�k��*�ҕN*]��t���9���,��x���&<=/O���f�]��,;�t�jHB��G��4�>m��O��"���HZ�,�]�Ƚ���v<�5##���Tt	�e�6;5^g��\��r���x���M,9�ԝ?1�w���B��H���RR܍��Xa��8�����������{m�m}`xFZ�G]�u��,�Vqu�20)�a��fYܛ��^��,���h��{F���6(���Q��rؙgZ���DH̓C�a�]�R�t˽��Ѿ߮�վ�O��E=�y�2��1���1*��:�#%�����6E=1(�$���~��ik��3�|�@� ZO��/�[�9����չ��rS)cm�J��M������i	�1j���"����of����
���14-�Ѽ����8v&?Sݚ�n�%<�\%X:@�r��X�%K ��m~Y���q�wtW����d�/p	K�i�c�4~JX]�>(d�ޝ�5�~W(L3���9�X�dĉ-��ϲ-��:9'u��p?X���Af�
I�'I�'ܷ}��(��`Luy� ��d��a���.���~4[���aE<|������I�vF�L6�:K�9��'�@�G����/8?�d��V�&S�Y��,	K��@#�4�0'��k���u�lw�	�[��}ť.s��GF�x!��S)t	;SL�V����)3�i���g���OoD�/hL'�F�p�xk~�A̯zg"����z��3*Jp
}z)��Ѣp4|�ڋK�w��S��1؜E�����`j0k��$scQ���@i�S� [y�s�1����5Y��|����(��H@����J����g�r���鐇`�bo�Q��5G���p^c�(����h� 7!�E�022�oL�����S�?5�S½�k|���i��`	��;._Xf�WVZ����+��GWY��6�B��ɓ�z������i�o����x�8�/ϼ9�}zbH����г��@�x�1Hr*2/���O��he�X�$�� �ffJ�'����h-�(���VE_���"��^É�1#S�*����>���6Z�:�.�,gn�o�g�u�(�Ýa<x���d'��lAJa:?���%���j���_ @�+�z���'�W���gn��N�(v��$��i�O��W��9���Uֱ��׵�LRz�L�SR�����u	T�-�5�w���I-�9SLФ&��l��`��_rI�4��+K�y:w����K�kρ`\i����P���p�f۹k��:��i3���"��[���W\��H$�3^Rv�Ȗ�"����&[���V��n5�
����P����m�	f,a݈!sƟ'�`���Igf<���$�"(���{m���7���[�(�4��_�c�Hd2rt��j���6����S;� ��D�H���G�=8!�+�!���)֜��Wn���J�cĥ�<���̕��x�^UUq�^� xD��cl�����r��>�����[�)�;Z�}�m5l��x��]�:\m����|���z���H8�OE��������O��n	�~m���	r7�E��5�>&Wc�L���JR�n��rc�W���u��6�/6��С��ڨ�3�;@���#��2Ĉ�A�J�I�ٶ�6���aT�UU#����r�>�sދ�	��vt�~UQ�v�A��?���Ul�qLi��6h��[�Hv('���%�_A%	��Vy�:!��[� qT��ы�E��8�%XE8 �E�;���Ȅ�Waҿδ��;��cvf&�_�H����K����;R���V�6y�NOѵ�Zl��{�Nl@��u"ٸ��U��샲;��o��hGx7NRU��V�P�HB�]��Q��Z/��Rp��Ԏ���{r�W��㾭���Ub�B&���H�!�����_��Fw���t��!��l�)�+�rg��R�����)ہ<</�p�ۅ���o��*�L_t<���"nU���#I���w��� �(� l�����@_�~Y�y����Zp���Lk�S��Q]>���=�8��~�צ�U��ik{@&:��x�h��'�����=Z.E!�~Հ��3�[	��x� �$��0��e{����P��ޏ��'�g�5R{΢��V����8�
�=0�E�:u��X{$Q�b�^���S�!a�t���n9�k��s8�NP��lB�p"�3� 8�̔�llB��B�h_'��IZ�+�dZ�a�NB���-��h��.nt����{�����"�:�Y%�8���0�]`�/���5������{�?��)W��g�h�b�ȕ���@�h���p�u� qm�W�Q�b���;�	&�?��J1�P�+5�YMU���5���OJ�m��Tay���������m��<M{oJ^?��$��t�%�@:ݛ.eG�|u�CT[8T-��9������<�.���T~tو�3Me��:�8��G���i��`����w�m��٠�>A_����R	W���&8��Q�eM�� ��γ�u����U@9��u�ƛ_�hf�*#�����h<�	@%�*!7��-�d=������T��?�Q�6����n��qzfB\��W��D�N��"�}ޱT$���s����bBP�UK �����.35�`�dީr��w��h2����EP�?�_ߘ�W!�,�5!B9l�ξ둹��E��9�9_z�l��@}���y�C*3��Ӆ�ڇ�/�L��#]����[�NAݺڢr�=�����7�;��`��Rs=;�H�4� k�z�E�U���x&a�G4�j{~�5�==���J��?	�����q�P��\ߦs~��v�C�&%&�'�~n�*�C��S*k��uN�[iЊ���AO4����H7`cERCُ��It����o���j�����q��\��G��FiA�
��p��({�0�l�ך��@�d9�j�
fH���]b�l˥48�;�]Q�u�ŏjG�ȷ�ŏ,;?�$|湚?�y)�A� �|P���"_�7�Wy��W�@{�[1=7=���+�B_�k�l/ ��Ϳ�*<uҪ�#}��Z����R�x)��E�yL,�Dx��g #(V��h�������T����6XHc�~�S��	@j�:,���/J����E?;Ĝ��;>}S�:ؔ��+�
F��rJ��S����k�i�����m�W�_��lGF1]����o	�.eR��">�������]���� y}H�
Ņt��wKx���{�Hl��Z^�K�I�S��i����*�L��@�5�ހcV.8�&>���E���;���ہ ���*T5�	�-z�`l���Q\N�7�n�Lz�����@����,L��Y]�:M_��2�y&�b�a�b�ؤ*7��${6��X!�^��\�H�����"\+:���m��f�n�sl�L]��F�� 1-?֋��xl7A���ȳi����J^5�� ����$��U$C?�r�w�oL" ��Vޑ�C�m�Q���t��_���`��YH�AM���H['ʥ��lX&��x���Rrc�|��@�Q�m�j_I��أY���B�= ��+�w����7����e��}}�~U���F���4���l�4�@z,̰�g����H�17�R�_��U�Y],�9k�Fi���JΎ(�^����#\뎊�B&U*@�M��O��[��̄#�*|����ͱ�1f)$�}8K�J��U~�5¡1�o��^���;��;�@����_r36��ƬAA��l�e�2,1�K	2���C�%LuY�7Z� �]J(��d%ˑ�PRV���}5>�"dJ��"<#H����WD����b�W�M�&vkm�g�+�L�2�T-;��5q&���N��D3��vg�T����aP����bc���0_oU�cD��j��D�qe�v�N�2���n��/���V3�HG�����f]�v虜�,2R�g�!�'@KE/�?Z�B ،�<�&�ylT�i�t9�=�it�cEe�(�ȭ�$ mF��졄P�[5�gF�a'�Z�q��Y�ϳ�5�o_��ӥ0}�Ɂ\�1��, Zb� �dL������*�4drCqZ��w�[?"�����.���j��'ٔ�h4�����Gp�ȳ��[t���'>�g�����魮A�L����x��=�҂�1z�ǳ��{7�� T�,D$md;/2?�]��w�ژ9D�����觗��l�gtt�x������-�>'((�$���n$�ð�"�(�]���{��0߻ʂ������[�g6e���ת��&T��Q��`�8�[e	�%,�+��񾺎�hu����Hv/qP�£�|�
�C�M%��[��.���^6������Ծ������QA�!8`���?P�ʑҲ��y�Unʙ6/-/�(w��$K��G3�٨���w�v��I̔MV$ e�0�H'%�L��s!�$���%ؓP"MsZ�^�ƨ�\�G��1�"���R��BUI�V����XO%��r!�4�lݿ	'L�����_���/���d%<ܞo=8�y�+���D���񮝩�+L������Q�ǳ7��`���v{�`S�x8K����I��@��4@�r�k*�D>��|KX�fV]p?���6(� V�T�w��M�CI&� �Yv�-�,����i�.�<XS+�Q�* j�D�8�G6[�����L�"~�pZ�`f��{RSf�+N|`Ү�W߀O�(�%)k��[ۃg�6�\gF�@/B��̞n�,!|�6�����%ȱ?���Q[k���i�T���������>����� Ly�X����"�^��R���k\{ .���� ɝ4�B��&>���}⸼�/4v�DF�����QZ�5`�r�� �#�;e,�� 
��'jD֗�O��Db���*X!{�hL��bv��X�RŹB~�B��2?񐔼-1O�'Yf�B{������0�;g0q���wl`r��D��;�l?�b���Ͷ�����,vV��9��\<��r��-��R��د�qߩP��j���O���>�/�1�,Ј�M�&� )�)�ǧ���ԏ��4���j���h,P�O;�X�wy	Pu$Yu��ʿ�Q����=;F��WWO\O��y?���v�$ڦ:226V7��F�Ȁ�l7�fLd"�r�H�ҽw���m���-�6���{ ,��jv$1\�FZ���
`��Ϳ�sIX	*�8��s�˖�N0��ig�D�ς����\MT ]�nÚ�x��v�anO�����ݿ�x�>�T�X1�@��'\_2��\tצ-���Hd���h����喽_^��Lu�����͚���0\J��~�9���7��&�:g��S���3fgj|�fNA�]/��q��{�'lv,t*V&X���߿�hI�w�_��la�U�����#��6��${�f4�&dZZ	�'`�N����1l�����"�J��!E�|�5��FFۑ��'�`ɀ��Z���4jPfo����]�g����������b�5��B��5b����[R'GM�x���R����&�0�x.���h¼U�?K��^�>�E��އHzh�#_�Ep}��p�6�}�S��I�N���߭�&�������8�L��uI�a�5M��~5��9.$W�w�-�Z�t�(���4P��·���' #mu~� ��s�]�$/.Kފ���W��qS������Y1�!�8��W�v�z׀j.y�y��W�g� �n�i��Ͳ���V�x��=3{�G�ǰEZ��0��l0�jȰ2�Նr��2R_=R��������@c���f���ysm3*;�w�災%�on��*\nPF�^��]��O�" S!#��8�h���:w�bx�
i�_��]N��	��/yksrb�%�	����q��
~{Q����Q���ݐAmX�a��?~v�`�L��wF Q�}��A£���;��g��6��A�Y%��e�p�Q����k;�$a0ʢ:01��`}���b�ױ��Ó��~��@���K�$Vs���>8X��M�X�&ڋ�LOx��ȝ�O%3c�}�-��I@�S�bWFt"(�e{o"������LKpYٟt�X��T��ǋ�~�[�ل|����+����3����U��"����>V��G�K6�)H��h�q#��8���l��ɩ���*�}:�l�dD[v~f�hm�au�{�vG7���dS�b�׷N���k�P�xı��r�tjD���>��G@���˷B�^��2�F�Ǔx����+����� 7�7V�٫f�y�@�h��/!�8�;Q�}��?/�X&�6���>߬��Q�#h{���>�wWߊ7a��ގ�rTL�@@}`����4Ǔ��I��:v�=�n^@*K��*!`̸���+xӪ����b\�M��	���x�>rc����F �#E�6:	vg��DLKV* ����+:W��vI!ԏ��kWi�o9�C0<���{��BB;o�:��O&C��9�홹|��k���զ7�3��b�V4g�	�v0�(�j��OQ�ݡt�+1t3��$D����h���� ��8��)�tVhcϥK�?ho���≶nUU�p"�F��k,	+q�n�z��:��{���mb���5�f����q�Ӡ��h���������Z�����,�h��%#���l���!_/p~_b��j}�Q9ܮ����s���)�� �u����י�rX���)�����ҟ�?J�Y��0)����<3理u�I�^ml���y��^��n���'ˎ�6�3��8=��P	_�f�XrR0��$�}"%k1��42ĕ�n�	w��dA]�Jc�_�P*��3�� x����'G�8�x
�}rrC����Vt%e�
a8�r�i7�`��+�-Y��(©49:�gK�ݐ�,Xn�8���R^&�lQ��.c�<�7l�28�6�C�O���| 4
��������;��
������4)��:DM6�n��z)�A>� �#bv:��ΚQA���eE�!ޗ�AK��$�����i��B����eSު��''>����e�Lj%�?�A���:���Ew��/���Q���]����� �<rɖ&�& x��ߚ���b�;����Xa��ܛ%
sB=�,:���ju|� ��Y7�:��-�9\��#�2Y�J�o�@��$kT�����������y���7�$~�jH���&��F4�_v%`����I��`JFת��T-�਄�9I҅����!��'�m���ī�)(y4@��pV��vk����/U.��;��7��-L�s������p���C�E�W��Ԑ|��F��QDF���"�����H"�w؛�M���Xh��Q�/�?���e�t��8�F,h�����"7c2��"Kִɡ@=;����� ���@��t�4�mw=�r��1�V���d\���c$��L���dg	p��_?Y1,s4w��7ٍ�\���g�Bo�-5c�nr��΃(��i�fɺ��WTdj;��L���*����ȳ�+�3	&d�SOȷb��4�}B�j!;�]ƨd���e�,�y�2Nd3S��.�9��_�:�ʖcg�-�W�{�#6�3!6���ur3Çѷ��y���FJ�`͗k+�i��z�x(9��qW72V�n.J�}�1�#�&������g����1�p��
�i��H��¡\~ҵ'^S9#/�Ӝܯ�8���Oӿ���ʳ0w�Tl���Ti���������w-�¼����MR*w��H���y��Po���V�&�^�kK!��j�h��-���&�^��N����k��[g�E���sPb)��,�!^���A�O%������g)������!%�󀾴�����VPk�?_���I֖˹m,))i�>��,�טq״I����;���+�-U�;�OC=�t���|�O�z,�Aޓ�3�$�_��kW���S�]f��?�Ĉ�(൏�����8�\��bdo4vC��H��f���7��gR��o���7$�O��T�S��9��!�!H�ɯ��~����v�7}��p�͙V�*3@�`���8CJW$���oN��m��r�{�*����ߓ���P��<�h�� ���N"o;΅h�{�9��477�
��O���H�N�A��oM��2�ID=���/L�������`@vٮ|g"z���ޚ�wDfw��;V^��8��< �q���@���X��ޞ�����󘗒c�~_D>0b ʕ��P�O"55��q�(=nj Ge�v1��t"�Y���TV~�y	����
��X����vv)0�H��.!�Y��[�J��ّ�o޸ͻ�m��W���226
��J
`L��H-?2�-��� �$�n�F���?6��{��ڜcֿ���ݫ"��k�Y��ח���c��">�o.a�74܆����G�*^���FI�: ���I� ���)�%*z����[�zb��yLv��q)�.��sr�ڣ����D�u]��\���� ��<J齜�U���V���hs[f}�S[[[�{f�J �"�,.Xs��tP\e��5R��^7���"bsy��%��.bN��"pd��hV�����;��d����\܀�v���d4A��\�J���߂�JC�#êƜ��j��o��CKpA��I�(�����a� �u�z�߮�R$���2�,���U��oP�%8��(�.�@n(?�_lS�B6r2d����J|@?X�g�y���!:E5I/�� c��U���^5fFĻY{e���'��?7Jۯ�r�
���+�PA$��B1G�t�Z��=/�S�m/���{����jO��%��M���9�v����7�V��N[�����f�I፲�ļ�dS�ɕ+��������G��bY�njnQa��i.�B78�����O���24���8 !VSB����Q&����?���^ݭ���������G�mNڼ9�<@q&$|A�J���mYK3.���TRo�A�{Kwi�4���˕��mETVH5pV7UE�v�ӥ�¤P���T��\�Uf��nl4E��'�,��B�e�wY��L^B�f�P��+�}�w����iR4��^^�輯��<�|�B��.X�a��`sI����D��Ŭ �$���5�q�N���0�)����ɒs�yO9lώ�S���h���Yy9Pk��~qq43�n�a9Dd��?L���.3C.���ޅ^E������/���b:�ҰD�&��������骷O{�(�w���r��9�N?�}��UܫI̲� �
$8�S���`�KēiNc#��gW�~l̲ѿ��H%����)����V�U3��?����7_��M�HT��7ֽ��h��W�:��~�|-���w+.:�N��O<5�%�<�j�'(p��`�/�����,�q2Z�8S�,$u������ �I��ԯ6 �#�#�EV7{����o(=ۀvI�u�O���q� Xs�~Ă����MDN3�Ej�Z7]	b����`�����$H:�.�m�?!qC�LU�[��H��MQ˿#�nZ����'ݎ��+���e������u��7�W
�"��W-,�L򐘄]SK��ۇ;��:Y`锛F노�k���v��n���	b���ݗ����S�6x�V����O$���ĸ���W/���7,_��yq����TF��TK���M5�����R!{�x������i�O&�𦬉��㛳��E����������?-���D�����q�m˺p	`�.I�ɑ����4���O�$��o~�y	��9r���N��`5^��Ϳ�#ֿBk������G<d�dj����$�;*�M������	o��^��sϼ��-č�m�ߌxn �� }�4��l����&E�ͥ塷k���E~)ѮTE��/��F�'�m���PT���l�m=��WC?T�Q�ڞ�C�h�m)p;|�`\t�T�����aH�# l�"�%cA�w��N��K��r�|[@����Y�C:��f�L����$y��6�^.o2��JUZx�S{�����C%TU'��&�+G!��VS&MPoZ��� 
�4�{���W�w���j�i%)�m�#�����ߜ��ͣ����>��i�K{B~ۆ G�� ���`'��*�&��'��z��ojྸ��K$=�d����V�5YY@��5 |�=4L6pPI��Iqߍ2^0̮�˨��F�],�k���	U2����WJ���`�ɂA9Ř��jr�P�y]'7��wHu��^R"5��8�ZJAW.�2#��ܣ��>]����RO�-r�|���פ^L��cCN,qj�A��7200 �ٵG岓i��Q�e���l�55�G��t8��&�T,D�?!�FF��6�;�&�#�� ���*�B� B= P0 �()R���H:ե�Y��oA�bV���Ѐ��/��h*�5y-"�qy���f�������*��w�+�=�a�v33�|�7�8�bU?��n� o	�~p�V�y�\d���/8����V��g��8�R2�
��W��*5�u"�e%yCs�!�-���F'\��{�W��=�Ž��o^�jr�.��`�uC<O�wc��:(���$��W���U��9�J�#��i�Zd\g$6�8f����R "�n}�p�.Pq�BR3�B"�Xl!d%�U�[�~O��_��Dk�Ϟ�*��s�X5�Z���8Gf����UBos)�Y}``���h�w�С'�b�E.a�L�d*ں�����_7��}��K����m�l/o�$�
��!���_��˯��R��>e�{��Y�nK9���P�n���n0��0�5!��7��撥�GX�h��t痜���ז@�rO� ��ᷚ"*'��[:2�!�u�y�))�!�(�=��Bj���s�.���k+q�k���� W��D�B9ڏ��O{�G��'����ɇ�6�?�����_d� �&���wE���,)�s9(X�PbU���dvR��˹�R7���w����0@7p[�ՕS1��:IW�e���L���_�P��迅��%O � �Y��P7I`0��7��C��'�.L��� ��Y�����ߠAю�u~�e�m��M$�]���V+�{L��1�o��M�/���������I��J ��з��wp��G�ӟN��i+�c)��C1�����?
��.���n)Sb36ұ EYL�^�7��u���?}:Ff���������ƌ�wEՙ�'�Bĵ�dv�Q����0���CAU���V:뭔-�L1}��su����7�����#��d�RX��a���^���u�A�~���n�Ŀ�`�6T�C`����#����`�r"23�M
?4!�=�O�p�dē"�e+�z��'kNZҕ������m�Ů�O�\� �i#�%��J��M�_����ad/�/������,*>�$���
�-n]@�klj����o���?�n���<���c�k^����}��������{�D�/��>���0�0�<��Ҵ��<�Y`z�+*�=9���nAA��p�7-+)<�>����ĸ"�L�K_5��Q.�@��vu���+5�g���o�e��i�#e���L ����V��|� �F��Q?.��4G/IH����J�%`&ޕ�����'�%��3)���t1/��4������ȇݿJ���T?��+܅�#��Z-A��3��q		H��G�,���!�\���ᦅGA��t|w��Ne6�E�#�S�z��lFvxz�rH!R,b�n�J�H�hf7]�i��d�zۡ�1")�֟��F��`R��X-��Q�W�^i�96��<�Y:1{B�p�`�_��@ 봵�?� 2����sӹ�R��F���y�/"Т'����s��HGQRNN0z�eZL��'�����P�����wzI%�Ԭ_C����)��g�|A�ս,�p�	�|>إ����>5��6�ih�i�ȍ�Nb���n��.痳�hnn�m٤�IMJMe�|����&�O������(ĸ���V�K��<}0�h_�sG�z��Y���;�|\\d�u��;@&,W<ȢY��m��#�����9O ����C�����(=��j!*7o*荎gڔ�e�1=D�����^��[�O��-]�M�s�&TKa�[�w�$����7cy��2�A�ڙ֯4����u���~'�`�����7D@=��Ө�t0� ����P���Sdg?�d�02�H:��

�r�����rvW� �ǜ��APxT ��N0�a�y���HQM�Yvdڷ�����.W��ICCܖ�fm*�RK5��4�H��漉0b\��P.�l�/�g�� _ so�~͵��2���h!(��X|��$f٧������һ�ZSSC �"�j��>k���E��Dz�5t�K�8���z�!9i��+W};��Y���L^�3.�K��X�*��z����dɞ�lK����2�s�W���ՠ� �ǅ�Ї��%��Y��B����aoQsy�P��c������E`����|X��S�fޅ�]SM:�n�QϾ�� Ϯ*a<��H-����������@����,�i��v1{��Z��&���������OB�%V
�:�������8�i�Y��e��`J_��|��[v���|�P;��ʧ�Y��O�.��jS��UVH��]�1<p$�g�QdA�7$n|xq����}T�o5�����"	�?57���'��k��Z�B��Zʵ��"UI��|)~�Cސ�2ˢ;�=��ב����*��r8�3�s�,Al��2��$xv��-�YK�6/)!| n;y;���`SF���!y�3蹞�����FQ�o�P�Z$%'?D��c���p�#�|�[�,�i8��,�Z��C��]x0{��؛���'����8��3�2�!*+�V�H�
�wu�.��!T��A���Ch:_�|������7�C�v�X4����)o�p�ᶃ���k�"#)M�HH�2���"�V	�1��!����q��:(x��z�|k�͟�S}	���&��"�z�1p���������B�
�q%�/&������}���t?�	�v9]�Q�|7���F6���@A5Nn�O�D�_^|���}�z����+��GG;|� r/ bYA}�t���d�������>�k���B��L�������/�k-_w{I�b���l=�nC
�i��h8�VVE_䗺��qj��U��'|�ȑD���ux��XB���) �]�%��Q'�h߃"�ׅ��F��H<y!�vI��j����M����A.y�g�ΛU�s�A�[j�"O��Q��b�Ή�2���i��°�u��KTBߗ����B�?����Oɸo�Ƚ�����*�]15&�I�za���p��@\U������#�WY)U9VC*�M�!=���W0UF�Dxu}]
���C�\ޭ7ZJ��[��xIÆ@l"A�*k�B�c��M|FRe=be�&��Jo��'��J^J1���9S>�* u��X�+$}����9���J&7;�}<�����Ѳ��//��#���V��m�=ڍ ���\�eQz�c [x��~kaCe)E���j�ܢR�jx1��9�Gn�o���n�!�p��?�B�W,���D�j��o4��8�]=�?_��p��,�̄�D�dxbL�}��� r�%r7rBFi���2�YP�4\��%++x�3�b�o�k�vus�H�#���B�x�1���	YY��eDR*܉���w���:�_hΰ�GL�K:72!������o��7�4E��]�/N~�8�� ��.�_�?��z�1E�)Ù�_��{dg����ri��[%LŽ$��P�a�afH@�����X�s��"7<-y"T�����J��a6⸡��۬u,�C�A������#���O�<!))k���a�4�-0�L��T^�F$���"I��t��n��C�C��1 ��>{���|+^�Hm���,�@��Һ�V��z��߆v8<��Saɢ ��̃3*g��Y��@"l�Fi����𸝧,nuSs��G�e�I���`�,�Q���A����!����[(A�ȕX��H��Wx�Ȋ'!Qkq����;Hf]�	2 D��n~n2K����+.Pg�XЉ����T !d;
\��7��[:耾���
�G���R�9b�Z��smz����|6/����Ka���R���Y �� XX8�J��� ��ꅈy�u���}���	%�6�
�x`�Ӱ���E-Û�Z�{����;(I|��yU�N��5���i.��h�r�|9p+�'v���ֵ]L%Ԟ��3�įh41c�h TIii�PO����h�$����7ϳI��WAꕺ0�&C���>R��F��R,�9U�:i�^߿�M���g?E絿���w��#��E4yoģD!\7]�T7�-�<�(�1�=0���ȍ-(.���'�4֣ffa����������>0G�'K<`�(G-P�(���E}"Y�������V\*������.e�r��T�y�H�Ql�Ic	��V��i�(WF޻���=��Z�����[�y��H���D<iY�$kѾl�c�j�ȯ@E��?����^s��W��_�R�>�Y�eW(�J���%���d�QO;���������Oi�s�Ο��ӱ���L}dS�a��WHGd)F���+��䑂R��ʫ�FD�� �*��K;��@�8��la���hl��KUB���O%P��V��͸)x!ǻ/��4�r�"�pƦ��V��g� ��sɹ��ȕiA�W���;����R���w�.��ޢ%��Vi�.� �b3<S��')�����=^w|?�Cb�(�x��qL���4��4YZ�A-vv� ���)d}K0"
��t��i+�ۃ'�gsgQ���=��4]��+m*De�AU�T�7��e�.��р\��ٹu�h���G�F27���]��g��O|k�v��a~�[`�۳7A'�����k̀���-o1��21hǔ��x2/�t:C	�iR�G� 4����hL��p�M%���Ӏ��� �2.fq��ݶf��E�Dq]V�Q���q���dhE��Wl�hW��u9T�"#f�/�$ͨC�I�˴�(�n\�ع�Np:�2��fͱ��k��b��6��D����gb�h4���L�{om����2���|~}�q�yn%��rJ���

�_q�U<�s�rh��ܙ�������]�����w�"2�2O�"�o$��(J���"w�8rQ�����^��<=� ��o��r�P�҉FF���\1T"�-/���Y\r$[�v�U��+�-��oi���͗��+�,n�}Ob����h��k�Rpe�8-=݀Z�q�"ДJpX��zKҖ�Lk�

	aK�
�]�����M��E���?�+!|��Q�������z:�>\C	a��|����F�1\�[� �ߌ��\q�F�f���`�����M�	B���ke�n���j�����QJ�ѩ������Q'��zd���C`��c_+M��k�O�]����9��l�'�h�����|�s�q�k,�RO}I5gW1�QP���ƥ��Ƥ�T,(�0K�"!ʗY���uu"{���dn�d.�/|@t,\��.���
��w�gv���"�:"am˯��Q�u얯��Ă��7-y�Ѯ��4�|:��k׊�^9T��M[��9�9�h��]���<����k�VE�.��V_k�w=���s��"m��C�i�i_�o��2S�IS����י���Ɵԡ�_��V�H��5��ٰ%��n�ꥯ�Z3Y��ьށ����\��(Ϸ����f*��[���n�3'hY�����QVsD�);�M��f�<����t�2i}�4�Gr��#+f*�gT�Qc&��*?

��Xrl�%Mg����ʽ�c�,�t.4����5���� k���M�]����ў-��+;�k���g����:�}���4$7�[)��P���:��{�T�`2T{a��O�1T�x�4N��fY̩��֦��ϼ��^%�E���������<k�cF0_��A2�C89�ɉ�y���-l�ظN��1.�olnv���k��U�&�Fh�Z��`R!g���Y���`��l뼷�Γ�Ƭ6<:u��b���sJ;��=6�p%�_L۴��=�Wzyv���0:���H#bܑ���&Vֹ��4d�>E�?c�/(��DB�x/��ʽ%7|1M��&O-�U8�ƲV�A��'���&��7���ivx�Ѕ�{ 3��[�Oen���1I��'K����HK+��QUn]�]�,$���?��7E�y`���7�,����J��~�t����������͍��ŗ2��1���y����u�FC1�:�{����'��c���~5�?l*�9��!�DpL�W/)�|�N����`��Gw-Q�f�T�o$�w��ѐ
�ӧ+-���Hs�!����0���E���󎮏#�feeᇉ�`����NN�-g�]�VW?����u	�������j��0s�Cn���V�	zY�,�ޒ������3t�#�_������,݄f}������~�s������c��/:Z���y�r(��������:{����T��|��k�!&f�Ċ������m��V�~�-���.��)�U�=>u�DՋ;w� �T�F�� ��
�sL��$�흛����������oު�;�󥵛��ieF)D�8ў�'B�`��T�8/����XzP	��8����6��h�2�58u��2�
=������ݼ�u��^N���i=��w���� !�#TN�k��:ȆD��,�����MT�"T�k݄p�Uf;�X��Py�YȐE�)���(���<M��R����'-�`2 0���`��J^2Z�N֒����鹭`��W���o���X-��
!%�!**b}j�f�J36O�ut���Y��T���7p���Z��\�7���;uu�<�ǘ�>�}�"��d4$�y����[H�Q���P��ezkh��h�1��u�\��M�e��2+�Q'`�rL%7��[l��'Y�=���wp� �n̞h^����G�u�Eut��F1*c�H1�(E�� �(J�"�� RX�^ņR54�Ra�.E�^E`i"�KY`)��ܻ��|���{����w�̝)�cd��W3=�f \����JR@��F��Vr{ �ˏޞȃ�F|�_m���qZ�V�SQ�:�`L6�37ڂ���w�%u��뭇���Y��.'�bHv�-at����U��nw�W|���nrQ6)!b����ݽ�y�J"�5��&;8}����Q��P��4��Z��1Gu��9< �9� �W�c���!�D�b,A�} �b����4���].-e��-LO��0�vZ#� �o#))��2�z>�]�\K
���r� /��Wc��m7�+q�"�wpvfL�y�U؏"x�zl3ei�ee���;F[�U�U�����|��i���R{�������NAy�#OMo�����5�R,N�xX��$�^�֫>kщ���Q�Ϋ4����@T>� �Vr	�{2匈j|I R��4�r@�EH�5p;�_��
($17�nw���9�-�Dj{�~c�_��ɖM0P�ج�f��)���nt�R��y:��]s@(dW�>ή��w�}i���.*��'�F\T�j/�z�Nl�,���ܐ�+� ��	I�{�\2
��&g���0u}lsn��T�e���js���>׶?�M��[�D��8p�;�����z͸o������&��� �* [�u��7�5���9-퍁�%�SQ�DH��'��)==�x&N���:18�ޓ���ڶ�ኇ�G(����ӊ�w���������U�M~<6�ڍcQo:' �n���a�0F�6�\�;^N)7i���a�M��!�:�5����/	L:4���~���X�<�_{�-h�;�h�z�`�l��ԥ�ը�����%,�W�?��Q�cSdH�}z ��=@A�[��ňX[����S�p&"Q7+�
p�����I��Q�Z�D���xZi_�z~��%��� w<(^^�i��Fx��J  8"�f $��,��'S�ǪD���j��d`���֯�	��b�Q���0�P��?� �J�H&�E�쎂��j�_&�Ey�F���"m�ѡ=/���2�y��\.�I�#60��̏c�G2���.yt����E,�� ��(d�j
8��#�p�D16���G����`����ޱ��GL�v�W���DTk�9����?Ⱥ����1P�S/����Ťo��2�5�Y?t��x��~�mX:/�U�=x�69Jb�\�$N%�
Ċ�(B�c�4S���C���G�����l���v*Tq��T	x�*V��{�J�	�0���L�f �=T��,__|� ����,���q#v��ΐ˟^¾�on�; =
��<^Ŷ��Ch�@M:<+��*䊠��[Qa�����%�*�'�;`܌�B�ؐ��6���]t��ki�;H�9�9���z,��a�@����^���z��~z�	_P^�t^d�F t!߸����3~t ��rS���['g�V>��hv*D��BPO})t�J�m��s�P%r�(�x� -�� ��N(ŏ��q��}2+�v��%B�BK�����@X��|��?��_�K��p�%(��=�
�D/3U�h(؀�Pmv�3 :��F.@��G�s�-t�ŵ��ʵ�/0�����y� .xTe'�},e"aw�	�������������6������.��vV���!�4�L[�L�a�!��&O�nG/6�<0:���g���f�}�<��z9yoZ�2nk��F�+a|w8~G6�c6)�G�u�<�"˲�0�QQP3W\�k\N��+l��9�r�؛JK�GOgI6�F$�!�E�(���w�ϖ�2��>�� ¾�R�7��!Z���xb���*��J���HN�C�m��=4�����E>���NA>�y�MXo������ �BP7^�>~����'pѝ�6�����]]	�:k�kH�P�J�zO`�=��q�zry�����6��!��S��Z��GN�����m���D�ku�L{S�$��S�v�`8g;�1��A�7�zR�Q퓟;�����O���Kn8!�d3��E��^���s*o��������`Q�`@��G���C������#W|
85��OZ��P|4�
�c���rP��S[ےl��h=M����z.�q[� RֺT��m�o;o��F�ah0_���A��oT�:w�X[F��3o��AD��7Xz%�7
��6$�=5�R�^d ׎E���9���+q~tC��$Du�E0��
��Զ�����Ц8ަ��oTP��|�M@�D�^��CN�����5��M�w]� 2�`�g��x��ax����(�)�$�����_� �م������{�aVݾ���&�9x�"P�	��S:��VOp8�̃����WIT��C�˲yqd�Q����\^7e�H�E��[ͬ@���ӥ���wN�3�;A�c6���mb*�۔TO�@ �������}^�fSU�LDe�cy����={G,�� ��c����I� �[r�1�n��9Iϰx����*�8�]��.�q]�	�|xR�c\��A�3��׬���2���V�N>�F?#���c�06��!��j�����c�ZA��{�G��!ѐ/Ҡc$���U��m,4
�����=�¿�h��34!�"��'��P�P���e���#������������q�$�W�2�.^�:��	ňXR������f���^�[*#�����	S�� &)2���/ρxF1��F�� ~�M7�Gg��n��x�mj���&"�sbGs�}����*���߶M�%,z7��5�)�W1�X�>]d�3�.���Q=%?�J�; ��p�"�[�\|Z�p��#�F�l'�+����xӥD�r�@��S!��A���]��czR��DJoQ���َGٸ=[����|ja�-�C��D��� ���W"�3�2:�5��c��3$ :=á�j�� �3��Մ�g��@���b(�LԶ�<=����ٸ�%�Bȓ��[�tZ��&�*���DoonN�}��b��!)���c�� �6���0|�����V,�O[G���X�}�Y�S�b��	���{7�6�Ю�8�cF����»�l,ԍ���t?`v�����G�'�A���Ui���e,��`*\E��<�@��/�;>j�PN,�4~H�SV����dC>}�]B �M��R�Wru�	x\�Z�Z�F�@��c%�E�UP~��F�a��:�����Uos� �P-? C��S~�C��l\�(�h�y�ײC |Oڱ���mA�n���x�>&����%�y@�Y��}	��A=݌����a��9n�����'�'�6�i�&2�����V����47�l���a5�̈́��D�;��#�����y�I]6Ρ��$�����F����x!��w���S���0�4������)�/�qd�N�FJ_� ހ���s�m���XL{� cZ�qy�+�/�"�VJ��}s����MT/���	��v�4
1�q5��t�8��vOJ��~��Y$*&5��A8��I����P�������)}��j|�[��ST�ȿ� ��D�@[hQ�� �c
(~Xh��&? �M�?�$C�!����&ئ-�혗(���V�r�j]��\๼��Z����Y�,�B�6�!T�Wb�~�8Gao�n2Aױ�ǧ$��ۭ����Ș�/���n�-cv8�s�h��J�����������Rj�l��C��/*���>�;ji�j�>����I��M (*n�+/��GV�����^���.��5v������^f_��A`x�G�%[��v��=�Ї�1|[bX10�.�ur�Z
rJ` �ʫX��K��������i�8�rA�: C'��D���*RT2�#��kk;�\��ޜ\-������U1�'8m�����ѨY3���}rH&�N@&Ƹd����`NW*>P�'��$
e�urU��mRz�t��:u��C*F��a<���s��m�:��#z	�^b :#���dol��h	����:8����~�J����a0��V9]�+��2y�4#�Ţ,��Y�$��[A���	�Z�����4a���kA�������B���33ڮ��/��"�h+Ȭ4��w��W��x�mwP�v�|�'��a��f����BxU��p+��NN	�d����Fp{X��)�����q4�bbx��~(�����P~,74�Ȓ�"�q-�r(�z�r�OS9��h]J����g�iOY}�O��Xբ��U'��ɳ����2�0����F�<%��1�����Y۬y	�#&s-�ຓ0Ћ��}6��t��9�1�������C�W�6n�"y냱Z�qۤg#H�  Ɯ����Yn���`�2+��� S��3�bj.��d�B���f�z��7al��>=���b��(��Pu��"M�o�	�μa��RTq��*o�vOG��妍���"��NM,�?��ۯ�EׯJ�6@����
`3a�`{#���ް�l�| ��ڳޛ�u!*�ʣ'�h�p��1ٲ��A8��]X9v�4.놧�j@�Y�΅�Fο���Wu����]	�6���X���VS�T(��ܧ�����Y�N���m�C�~L�߂�%�%Zo��H����H��L�dX�ķ8K���}7�n�C���\�k^�]�y�mр�>|�X��(&+�H�� �P~���|k6�׋����
�>�ᬄ�م.����>[�:]0�4n.d��k���F=���%�����	�X0�!N��8|-*��nY"�Lfe�/T��٦�!թ	�'�&g~!���}�J��8ݎg!�o� =���`J6涖�.�1�C��eC/�(gi�|�Ri����z�ꉻ��o����d�+|���o�	"6�L��(�̻����J[���^\��"��wo"�
O�R���˧x���``�i�bY�Џ��r�^x{��
H��[ȃH����	xC�k�e��v-�r@2��t�|�M�~�����i���q��on��t�oY�,��~�睅�8���H���L ��?Ru�@Ner����6��2V��#�&t�� ��j�B�O�С��"�)2�˧�5�e�B�ʳ(l��ͯdc���,�����;v���o�,��k/��6y��B��0}���~`9%��In?h"fU�@f&:�2���L�4�z�������h��&�%<�����\����*�!`T�Ȩ��	YD��#xL�B��yc��gv焴"��+h��zr�V���`����
�[u.���l��+�
?w�̷�̫Vb�
Jq
��MK����ծI������F�O�iH (�MH`���r3L�:wS:S~f �jC7^����A� {��q��PJ�f�����|ł���;�a��w�c��a�� ��J��R��[	��W�(�F���6��.{.��F����n>Xh�M˥�)�C�1�f�� rVrr �[B�AM[\XN���R� 1	��i�oy}7���Y��Nt;Gx�I�õ��m�����g�>�lh���� 6TI���ۍ�Ehu�7D0�����;��"v*����B"��)�5������	&��+,���{9q/I3�����އ�/��V`��6a��@r5_O˭��I}�{�n�^�@�_�<�Zxj�R��N�������(���}�]�<6Qu}�~�����c�D=�Ѐ�8{]�l،�/"���X��z�P2����h	Ovv0	�q;L�ݥ;W�F)9s������]?�{���&��^+�2.'+����¢ʁ��-oz�})Q�WJ����׬��/�F��2e�4&V�FO�f��'M7%\0�d��ؔ�ed�6�誂�cOS�a<���]9�XJ�T�x^*/ ��d/�
����t�b��ls���6�g6i�;��"�y'��Յ�=^�$�fp����v����ۧ�`�L)��hbd@���ꮔ�E�5�e�j/q.�V��Pd@���a��8�mr%UTWl��$�D��������F�]X�x
�R&$��z�X�����$Dૼ@ �~6x(߹���c�(���f5ɻQVm��!�(T���"zc]o,��������&R��b�zϲ�U��D��Y��Z��К~�ng�FS�S�����+���(���&��F��8�%:��q�K�.ho�V�������\	�O:�����6�x��Z"�+((�KӀ�J��h��Ou��>�<r�"j��=khcʣK��S.(�FG��������+��n�۰�8��zԵ	�]�y�����Znn��j��-�[.�jw�F�eN}(������WυwD;,��g͉�+s��5�H[�#���WB����!1�{��/#:�L�9��c���i���fz���n%s��o$�������m��=��.%腣n�S���-�ߕ���>���@/l��]�j�<l����;x?%V���$m�z��]m�)խ6yPtD�S{���{��&�9�1M����t�G`�,Y�1%��؋/S�Y(jJx��[|.I��_c*��w#C�� ��b\jʶm�[��`I�N�������N3�����h��Ѱ>�);9}�2xכ�[�n��L���T��������m�pJ�Q��4>t�����iW�u���Zp����e�O�>o	��;����>�*�I�'c��tf�{�>��H�����n�|��w��������/^����^Y�.�	[+q���41uV���(c6ЯVJ>�u�\��8\6m�Y}#���۲�F��%�֭�����"��5�[5� 81.~0��t*]}��낞K�J�dk���$*�8�;<{8H��KDҗ&�i�N�n�q��Q;n����q���gQ�aF>����i��$�<��ކ��l�./��N�;]��~e�:��Ʊy�����𳌇	^�y�_��4�I5V���u����8�=�T�mQ�U=gN=CY�\F��&H+&Z�%[��YSq�zd���/t�����ꗹ�0�O�����k�~�.�;oE�٣,`�p�C����}ʞ�!��4/Mt�4!�[j�&j����CC�?G�
~���Qd�e�z�))�<",.���C�1�-@=���#�����Y��*�"�H�c ��ܶm(ى��0@��"�T؅6�0¬����:$�y��q��>��,ا-q��ˮH��f����z8qdC;]ch����!i�Q��@�qg�YCBB���f�̧�A��#�s��u{��@8m��z�#�&(p7�|�t�]����� K���=��H+hÌ�!M��2,�x����g����I���2ܶw�OP??���>��U'�c��f��Ð ~b^��Ky6
?�P�y���)�{�,�UkƤ� e� ��5��.�|��+zj�MY�hw��|������,�z��Q�!����s4������W��.(�]���KS�˟�7�v_�f��o2�f�T����%ϻ�Axo-�$��.Ι�n�-s�"�/M�e;L��ͦ���+A��L�ժBDAT{U���`
RK�:�����P{^E���7ڥ��(}Y>`դ��^�'W����Z�e�`��r�������ǵ��A��6�&��`������H��!J檞S�z�&vL��^9�&w��J��؛���)�FOO�,����ƥ%+�eJ�����g��Oc�q��;|C���|�2N��o,e-��3<�܆�����#���:�����r��J����B����T0���O�u|�
a�\�|vM]����x��˶�]1�'V�%(��Y*A��ʕ���n�%b���v�^}�9�ZY�Z�����?�#;�W2�G�@#5`�`�4'�/[a�O�Թs�w�Ǐq��W�h��#���$7��7�j��	�} 5���VO6��N9�`�m���N���32����vl���˗|Td.;w�����^��<읱�r��:���OXT-V���--߾]u�}�8�}?E���
�y痧��~��-�?,�D��C�`�=x35R-� ɇ�ŚJ�Bl1/%녇��x��ִ�����U�/����o�y���"'��^8���?�����f4��<7�~8v�3L8��r��.S�~[QJi�{��K�ю~θ���s��0��~�0h��B*J�*2�p������.Qڇ�o�a��z�:!**2�o�����Ń�ū�2/���.�߂?�=�2U�2qc����n����DU��-��ƤܥpR��*�n^1A����Oo�j9���W�^{m�n`iްM������s
K����G7��*�4ͽ9���K" Tg�|	ʑ�6YY�˱�[�;���h���Q�9�k<@����d�u��҄5n%���ƻ(��mch���h�p`�9�����Q9�LA[q�e(���O�epO2A��0!n�f��8~p����[��P� � �A��)(�>��o������=N2��"�/���Ԥ�ƅu��M�́O%Gy�ρ�5__��<Vd�溷��>\ER׷)�J3ٝ�Ln�m� /+�/N��#��A�qV�R�%$߇]$GJ�7Cl���<���h��<��B��
��{��u½|�g�j������u�w��X�1��_�F!x}��[�z�����K̞�: �y�" �A��ƚ��@v�JV�w��+',� Y �yfD�!@@����-/���l�
v�F��<���VnJ�r�({��B���C3���Q��o#A���J���������X��엡ܦ̓�䚹9�Pu��i��˗A�tt�ݗ��C��1�:J=[���ш��Q"���:���N��E�$��6�j�xe�����2��Q��>J��	��/���7͇�q����@i����O"+����oHQA�#�����7��/��U.1(YJp(V�l��]��G��!b���3Z��W�a�:��	�C��.
����_��������guu5$�P�֥����qL0f7��8ߵZ)(���O�̳���P+���vx��ƕm�x�L%M����fR��&��D�xȡ\y>���KzO). �Y�z���N�z��ϟ@Q+3�A�B��\t4�V��n�r��'f#���]~B�~DP�A�8����!�K;E. �h�u��&�Ck�����[%7�j�ع?c�Ƙ���zf�3�x>A�g�V-Ŕ s �o���\/�)�p����?��Ck�z���=��̒���ȓ=��OIC���f\�7?ko׋-�U̏e�|o��U�tm欤, dv��;�D��c:hL����	L�;�B֓�C��1�L���%m~�ing'ũv�!�˿���@v|�e���Ok�u!��9z��xez��h�JxD0�Mz�.�u�wƱ�ޡ¼۴V�,���p{N3�􃠒ݻ\{{8{�r�Նz��eo��8�;��e�Z����[�2o_���Lq�\m���"��U-4�I�ݞ`j�S�8����m�����is�֜��g=n����S���7y����m�G�2��&���ՙ"�K��)���?�n@�W���ya�7��B+ֻ�KWG'{��� .���DA_���[����O4�< $���2O��#���-Ŵ���J�k#zR\S�r������O�78�Q�)��	� i6�(�2�`J<���Vn\���=2�8��7Q�#cc�a��"1����{Z��,�Î%�H-��T�j�#������|VN�s�����=�w��ۅ��֌�LԽB_8��NvL��<��+��;�!�;'��]Lj��}�,� ���a��R�R0Hy�}��maX+7�r�[h+�,rw���Q��{��nY�.0ԁ��|LNQ+�N�c�׬�.��i{{;�EPq�A���W��CqO��������{t�8��˱��kv!��P�hZ{�g0�kB�*�&oNu�y��� _�.�Ր7���SX�����Լd���_��r�HuR+돷d��	>�2�ڡ����57Q��$�<F�@&7o!4C&SM�Ug�����f�.�Ⳍ�P�ڊF����7��CFq���9���e���9qD}Kx{i���[�{�\�C��"����~W$�Kʷ򅷓!���\���*6['#��}���;lZ�ӨSJP��N����X�y^�&+�QɈ�f��@�^\�"*�7�q<����wl�B^����Ug\�: {�ŀ�{(8�L-bv�:�"*'�����LE=����2'Yށ<U*�:8سs&�	���/��S�0u��鑎�N�4��;��+˯�q<8���R�T�mڀ����R��e�J�C�>5�D/��;���:e����hy��0{�:գ��Pٻ���]� ���p��5wsC���]cR`'��`_�l�����;����;�ĝ������L:Ȇ��G{e��j�_���9�d�^TP4�<��r�I��aC.:���u�6�l�g�W�K*t�RT���v#M��1c�h)�<�p�d��k����0��R����'�,&�!Vc��F��a�\��&�Sa4Lk�]6⎅]��|�47I��:��i��UPל�y�w����];d���4��L�8���Cc����D�Au�ڧv��/R�&�X�J붞�l�L�t�P����%XB�l���(������+)�uJ��D5�bf���SB��K7�ߺ�n�7������ݿ;�Y裭�JroW�Ā�Aŉ�&������KWg�ȆU7��'�*n!��:<ِ��yG�㬴��N����7���S8r"g��*��M-LtB����WPJb���OZ[�����Fљ �ߵ ���|���w�R�}<�~t�
�8C���4�=q�h�pP-5u6 ���[��ؼ�E�[�PPV'�bH0�Q��R�=mȱ���3P��D1-p��� �ݟ�r�WW�����%K�v+�X�z�:10�6<� ����$J�*��8�ʆc&�ݔ�#��1hX
���"�Tr0�y�a�6��f��r&a��� f|��`c��VE�X!�۴n9�95eo��_����$� HCb�?�sB��Q�.N<��;%�dw���d9���o�1�nNY-�i�w轢�o�A�OE��=����F��k]�r��<����� ��N��q�.=�u��l��YB�ؗuho;�~eks�*�F�J��2q4 U�5'G�&���N���b%�3{Z�~�r������4~DE�-yX��������- {dd��hz{�D!0�w�l��L�q���~'_�_YA�Ǿy����'�U��Ӛ�/:&6�vȏX礆�'�.�'KWMPL�g� ��'�J�F���e}����㊡�څ~������3 ���x�n��Zr��Lo��OY�@��Xz̷6��4�$�] �&��
@��+��&��Ç��e�l����7��gfϞp+��Rl�dl.��R�I�wZ|��������31(�ʋ�;���5�"_�D.i��w���#
� ����f�����]�I��_P��:��xnC�o��?�Ր��rAy�"�W���ݧw���W��|��!" ��%"֕*�m��L���W�7b� �)��ĺ����.���- a�蜑j��n�zDn&_,E�3_��l�v�tu�Z�,*|��s���@�5k�C5�]/A��(�U:~QT5��9�)����㰌|Z�60Z�%JȠqWN|��T@�? Z�;�8{��K�577����UjQK��U���/J����t@I�UN��V�%qz���)�� ��(8Y���F��..y���<� �ğWe�׃<.�(�M�%' Dv+$�p&j�����r�5�MZ|"�(:dȝ~�e�/rl#��H	�����0�+�f���&���.��CՊ�5�Vko�Cc�+3�Hy)�{��P}]��h�R�b�j��.���/\#��I�>��j�bd������#��@^',K������㦓qg�l���_�Fڃ�O�F� �����luT��O4X(�es���b�Rz�K꺛;lӨ�E�"���|ʸ��(�#V|����[=v���Z�-��۴Jx����E~K���e8�\�{;�g]��c���Xeݠ:i��_�	7Y���D��:�H"�d5${v����[=��xų�m�kЛ��s�m�1_dL�*����f9 ���\�(ˍ<J~f��띜W�ٿ�*�oF���oP����4ǧbګ�����鍊WL�ԸB%��p3�_x8�����q����x�fF��{�8���ݘL�=�Zy6�VRd\��!2�i߫�\7V�ekM�|ƣ!�2�b�^��T��[�tUu�� �TF3��<��{۽�r�]W�?)=Ǿ�wdⳡC��W�k�p��ʃY��e:$�6���[]1��?P�������i��.��X:�} �
�^}tN�O�7��O>fg�'���؂52���4+�b�!S�x��z�/� m�=Կ�d�)�;�' ������$��^�q=�^?�!A֞ȒL�l�ך�ܷv�%ߜ�;�x�/UM��e���̃x(��(w�)�' �6��� M��&��Qm��Ǘ�[��U��Y��Lʞ����'**���v��k`n Z$����T�ou�G������>��g���#ܭ:)r�V)�vS�G���Hާ��)���+�,S3ԫ9�m���^�쾱� �<��wCnl�͏�K:�����BO��y�#r���@ x�G4cҿ��KoU�M�(���@�x����`rt}�ۭٹ��L���c�0��N��R��k�P2�\@$>�hv�4w]�B$�������!��ׄ���&��m &�6Qsj�0N8���<�89M�'L�i�g��1/<x8L��B�/�� �QP�:T��@֫!�q����W�Ѧ��n���5nP��շ�T�e�K���� P��-��3|d�/n�1C�<b���p5B�ox�?��.#�:�7'�O[P�{�K�!�F�s����d�0X�4�4n�F�����S�Es��d�Yy� m A�����m #��x2죈:��YkE�l��Y򶟣r�c4�N�j�ơ�0܍(U�b�@�:be=�8 km7~��a����z?ȧp���	L�qBF����k�(� G�fK-��Afhj_�'Yq�LoP �=c� 2����&KS��2�*�{��������M�	0��T��0��Ғ�� �\�46�פ�a�8���|R�a��mb��2Rjr6S
��o�)�_��Ю�TtH�������-�mp=�ybH�\ ��7�+UAa�`@���n���	�i�w�F�Ͱ�O8�����[��h葻���E�^_$�����ט��^: �rJ�Y�SG����rN|��R�C����w� �j3[4i�IU��ܞB�GDh��E["��V�|�_Je�A�Xt�%�͚u���9
�|_��`�Q��&j���-�NfI����'����^��$��@��w=�K֍��S��_�,��3�6���u|��a{�'�}�u��ѻ�e�̉<b�1C(b��s�m6>2[�Vil�_M��9��	<\*Cy��gUP�d��@�Z��^|yni:��j7'�i`��|R̷ɋ�\�@	$��Ʀ���X�o�K
�Lej����OS��1��y�X�E#,>��y���Zh��O[[[�|t�ʖ�zĩ�o�;��7���ʔ��zES�?j���#���z��}��\F�]��L��FY*/�G����� ڂj�$==���SP:G�G�������ny��7R�K����M��W��V� ����N����C:yS�<wG$_�Z)Tn������"������Mn5Q̗F���wl�"5�����(�^kd�����70B��qZ�ܲ�a�T4�)���2:��rj$�KB��>��/
ܡ��4u��F՛����/o���go�O�9 �T>��A����i��U�8Sp��0��iW�;��_��y��~8|�A5�l��8	��'�)���s��Nj�ڍ���|�SF�s�Mޥ��'���<n0[��N­����!�uZ����1���(�e��c��+�(|R����J[�������yൈ�J/�8;��ZZ���m��p�68hG��3u��@��0�	�E2$[�I&�׉�g�q�4(3j;���Y@ПVW��=�
�h`&�B��
����D��l?�]X���G��{��
��T�*Z�=�d����WN����e�t������rQ�|~r"1�Loy4��Dz�4�Ɵ�{��_I~T9�/:�疝0+Ss��`g�Ǐ�q�݂�a�@�U�@��?�JCí�x���1��r\Z�za�Z(��E�����L����%�̠�Fض-9Cv��փ�_)�oLZY6t�2\yd��1T��F���XH$�.��k}�c����[ԮK}<���ԤYuS�;��-�9�
�#��m��j�;p�۴�R�&q!m�Q���<
S[��*N�ӊAx�Li~�-�*�{��O^��~�\�Fa��O�&��� �a� ;t�CU7��5w��91{t�fB\B�K۔5/��1)p�����w{�6�����Jg`��^iud���Fݶ��R��3}hJ�%AOl@�介�S�ܜ�����Ef��7�L����J�B�P.e��Õ^ �;P���B�CIm���se��Z72��!������"�'Y�6�[`��rs}m��V�n`/���"v���]�U��Y��xm��(�h\4}::S�>j����9�Id��(���i(Ń`:00 ��
�W�/�_����'��{S���y�Ά��{̔�����qބ�����`�r��>D�q���e%29h��^�a�:�q3j����ԯ�V�xv����+�����P��e~(���:�b��˦ nɆn���������b��뺷�ˤ�$�j}}s��DS�
�+�f�}��q��p���c#��\r^��viD����S�����&��A��T4;�Cm���A}�x�����߰딨�F6Lb1_���y�}DͶ-�GK�¶I K���v�"0�@�G�PBSE���T.�	n��.mRt-$G �j䩟U�ޑs��������7�9ܭx�<Z��m��A�^Sw�_,s��'�-��F�i��@e�m[�Fx䱟�L�g�s��s�<���r� ���B�q?���w���M�6��#��/h����� �`G�N��=54y��������M��Aզ���g|�z�c����%Wd�I��3�h` P=ؔ!n����_��)TZ���P@���v���,Lt\�<.��w�����f�
+׹aq�|���z����[:b�3��R����F�9��)���Q��őZ�A�;� �(,8g�~Ě�CKV�I�yN�p�����^Ya�Ǩ}Fjx{{��f%j�����H��z���A2��&pK��D�+í̋��]���¦&r�k�P9hR" �j�T"W�����֞%鑐�?Ev�.e��s�5�ޅ�ل��-7
c5U0�6�m�ݺvݚU���{u���������9SC�g�	��r�(X������Xxb�t�;A��+�b%�f.���N��q�g��T��<�*��&**)e�<��+P<'��x4�f�N)�������3���@�I=}���m�f�۟_�ȟ��CG�����7�d�uW���-����",�S��G���9��/i l<�GTDD��62���y}�wѶl�!�.kKC��7����
��_���N�Ww[��+z��q��#���'�J���� �Qj)���C�޲RW,B�׎G������^\~�*>Y�*�zo>��u
��-������K�0dＯ��+��W��M7��.�_D?+��z#^FG@�r��r�����9z��nSS�v�S�bRW����g!Pb��L+�).u�6��K�=x�D�7��4n��P�k��=E�����jF�#�ժ��$�=��ސ��#�d��oViT%�]`�xC�RzkU�Ű�l�M�tN)QF"��٢�?�b��e��놮����?�rA�/0���hd�?}d�A ����s�U�$h߆$s�im���sB�c�⩆�S��J<����AHs��kR�㭳���֖'��Go�u�ͻ�C7�|7�<��u��FQQ1AG���	���KU�(8fl������B��*U�![���)[D�����~�f���E�MU�����l/��L�^�G��y��%t�]<����)_���,��0�޵�F�;�Qq�En��::YP\�mc�<y033�lRg�I��Of�`�pO��³_�X��@�����M)�8PI��U��NB��9��Ř8%C��v�yaX�6�f`@���Sn�/��NjpO8�X���X����}a]�=/ܐ����m�����ݫF�ۼR".y|�����o�2(
�Ğ������@�ߛ�1;��^#�D)���%[�EV�漩�K@?�G�vk�dK����{�5�;?��j#�a}�Ő������C1�t)#rssӥd~HI����.��y�:�>�_g���%f���.�v������~#��A�~�-#��pC���x�\�2��� ��yK,�<��*0�W��B�D�w��K*�;�ϻG�>�r-���<	�AQ˙[֯:o��;Ք��W�1��5wAc�5 ���k��kwq��rny&)�4�#�xS�0�)��k"�;�nu�$�
���e�����ζ����g�l�4
\ťL{�M��9������E�/�*���b�cR����[1v�Z����*�|�w�ؘ���>K�����u}_&�*��w�jxxx�ٮ;�/?ž?(ix�n�`w~H��_�����Jd��C7>h|�Q�jr�4G�Aː������Ðf< �|��x�����q�#$�<���b-�@��U{���&�g��'�Q����X������D��;'���4��K
F���R[M��hgx�s��u1�F��,��7�X/z�]�
d˧jP4
Xg�.��𐮨�D��"oι��V/={�Iq lޏ��:���&���/�0}�_ж��� �e�+��-��6\����X$:�s�-z��#����&��L���hV��fo���>R�h�%��Ee[�0�����D��*L�۹�q��:gay\Ո��n&3��S1d��b|彾6~�J`,x�ȅ}]6_v����ʴ������5u_�
.6@ GWI�A*Z���9@Y`�Df���s��1��ͯ���v*l�#�໘H��]jU�;B�V�Ɓ��UMyo�,r��Ï����@6nb��㮱k�Nj
�S�S!>&nY�����{_Pt)�mS�3��o-.��7-�E��k��q�Prr2������u@��$�Ҍ+_��M/���@6��\鳐̇���z�އ�W>�`�Z��7�?�4���YΦ�Z÷�.]�"]3�5�����]�6�6x ��PUx U�W֝�O�<�X��2��f���2.oXS��Q)O~ ���FKk�gec�D���v��9����C�1�c�`�{�ۦ/�D|��+��*kf�B�(� ؒx�<��̘�:��*�W�#?R2	�tx��zɯ�˄�=oo��Ĩ�����4tIv���1ј�C,��X��~{�\�s����1�@���v�����ݟ`^t4Ee��G~�n���ZU��۪f����rt�3)�q�e3@w0@ � �ן����FE]�T6��͜��� �]aQY�Rr��I��7RŻ]x�k�eA�q�<F�zP���!A҇��t�;�t��r�����:�i���l�u?�!��b����ɋ��� r��ҏ�=�0ԗ�O�WuR�^&zE/87��>,�&+��c>~W>"�5@X����=,��~�ر��W�~	620!�.@�M7�O�X�胸ۊ���E�^�WOpe��<	>'>u�<T5�5me�'%�K:<��2�����H�&dÕ�<�/Ͻwp:ɧ���~�B� t�BQ�U)��~�RO������1!##�����x�m���&�$�yP�ytE��W�#�}$��~�Э}O` b�B��h�5�ҩ�`����*����G����O���o�T�AH�DM��¯�� GӅ�;��i�����_��4�L�@��?����{���0�����H陪LJ������m^$m����(�(�������Ϡ�_	
v��ߏ�||4�2�i7�#�*�T���#eZ�ݗBg[4+��~E�u���?�;M��`��m5v�Qɟc�6`u��m�ԉNt���:į��t��]e+z�)t�i� *�1�3 �s1s�j��09�&�B����0XP@Q)��=��N��%u���w�g� 	j���w�n'�;�X%�ߎU#��������K���f��mn��t��ټs��v��J%�I� �y�$\���[�uc�b,��5[��4�2���t�/���~�Qq�f�y��ɖsF20BFa�'j�
J���iMew�%��6�w�զ�\K�1=��/[�Z�K9d=$�Sq�k� �bc��. �D��.�l�މ콹���˻ޭ	R�5�������{�3�:LR8yO%R�Vz��r����g	�	�#Wa�rk�^�ZH�W;Rs�`�~b�`n��	�[۵�
2��uF;�X��V��;���E�Ʊ�nǑ��|7����Kn4�0qx�2�
3�һl*H��8p"��#T�L��\[G�Є2��^�3Sz�hhz4}�s��8�!��!��=ExNЪi�dG�K�r=����1 7Nv����H@��uu��� ڍT�!&���ݏ/�za�T�q����u�&���9���x��CR���r ��ҥn��][С�|0��b�&�n�Owv��Kъ<i�
��C�lV4�_��nY��u�p~�10��v�L�P�Щ���q��n!�?D�@8��1�R�N���Ӱ�����P�@޷�����M9��]T2t���]Q�o��'z��,e��$x�6"���ͼ����K�{R���^��c 5�6��W����A�������M]�j�[�-7�W7N��F�j�Dj�{^�J��s��f�䬭KV��6��\v�ҥ.2D�	�Ni;>m#�L?I�9��nyOCHtPKu7)_��J_��9qFS�fF� DPċo[���v�)��9�N*�ZTWQQ����c��t�%�,��?�K*��v�%>�]-�E��{�s�L�l���w�0{۞���k��u�w)�˜�Ka�/37�8n�����_Ż  �{������^ߊG��եP��Y��Y�}nV�	��˽{�{���5��3��/�S\y1�����b�N�0E�2%���ۏ` y#��PT곑���HIA�4ȗu_�${�yy/� t�m�ked��I������jr�o:�JYY�'N�9Ȇ`�/B�>#��ư��p%|�x��Q��qYf[��p�����R*�*H�c�"!! ���� ݠ�`Q�H����t)!"% �t>R�����~���}��Z׺�����w{��ğb�/!3(�4L�J�rq@��Ò�,��YN�/��8��~P��+*��R�S���>������#���C;��ɂ+Fp��YN�b�@�U����.�]��0���f�$d��C��i||y��Z��`+ *�W �og`\u���}=_F������y3u����^����f�v��ϼ�V��Q�ٹ_=d#r��|d�BO/	��Z����$�' ��}�\���mJ\�A���&5U���9A��D���)*)]?�3ښ����tt�Ed	g �	�<
�B�ɦ釩�zƿ��6e`�Zp�á4���.�i|o���r�#]tf���uDx�F��8�\d���,L�P�Y�eA�ys�~��Ă�!^<�����է��n2n%���g��y��(��q�������k#���F!�i���a
����I~���*�U�.R>^��D?)� d��o�GK��aѹ�?+��dd���}���١i־Z�il�X��q�Nq\��'�"�j�����d�Za����I!�N���!���|����cB4VWm����Y;ͅh#�Ј+!��y��`~�Ҝ;u��C�օ�n2v��`�c �I	G��*[���c�?>]������~w�r쏍�8?�9P|��l_7�caL���.e��o1��hEj'0�$%���?N�/Q�W�A���2�
�
�:ζ��^�&(s�MʾfǬ�Q��]k�lԳ$vxK��9=SZ���Ņvj�q�#A �����db?����l�%��^U���&f%��+��x�a)��+n�cw����jq��f�9���ȱ8aINi� �:���=�������Ǐ�4�2vX��>���m�(���R����F�T��|pآ�c��<�\�3�5�<�M<��yR�M��|n���~_�����ʺ��%y@�ǫt�`e�T��k-���( GL
JB�&�ivL~�	:�k�vK�k.�^^�13�t�-e����Vd�^�.B�����4`"<�]��)���!(x��) ,5y*NB�9R���!��e͉�[L]��|��y�ӑ���滪$Wڠ�x�%��{��Hy��?-��V����u�Gz���_L����WڟO,NV�ʘ�౐J�sC�>x�ZPJ�hct9��fmm��f�� =�Ԡi�]�o-"�r��R����ț�'=�����VS��(i�H�E��[:L�����_��@�;L�c"�t2@��Б�����_�_`U�wv����ؔ��J�����<W%(h�U��]�����H̛_Y���$ux�ή�������/mY�ب��p�f������>=>HpJ�q(6��H�(�Xk7�V5f��l�P�Ԋ9`!�CBC�(i���̆��+O��f�h-��v1���]�9`ЛfW��L�#�\S�Y��]r��!��fO��d�;��|b�u�l�UEGGwg��WTq�A���hg9福���6��=_r��5<
�&>�9l����S.��g��D$�T�E.t�t����p\!���hcŢ,xO�R�b����܉@���Ts3��7Р
��V�M�#���Ę٘f��&K��^�4�k��۷��3Z�;"��즳�gk����m���ϕ��8�ɢ�4�b�����0��?��qX���uKk�9��!�Q1C\&J�`� �ņ9�ք����ރ���{� @��p�Q>�F��GHw�Y+
,������/4QSX�k?arD҈[��qa�='��G/��5����HT�O���y�\�\��p�` RJSEq"��Ȥ<j$5�|��"�{��o���wwR4�N�P(/���prFdoYr��$g�y����α��a1�`�G����j-D�)r�[���sK�T�����LWs����z��4@+��mK/���Z��k[���F��@S���H[��dd��������s�/��ݝ����,>ZX|=���̯�2O%H�CNW��*(�AHb���0�����F�Q:��2B
0%e%O��q����I�݊aFFF���+�ǣh� ��ўc�封E�����i+ݨ�ݱx¶��yp0���篸�j#�Q�Q{s�rᜆ	M/�'�.:^}�l���ʶ,�cslsBn�(�:�-�2U�L��K�ؒ2?��������8�m p�������.�꩝�����M����\�4�;6	kn99�!y�M"��S�\W��*�@@�9�o�///���{��D�`��DV��� �
��~�r,j�Z>>��m#ZePvD���,)��/����3t���0�E]$��;A)f;��K���fJRCva*�I�����|@̑����w9@l�v�{�,�^�=�88�K�en�ΰ|F���'�@�"ɲ��%�Q��7?�����Nေ�ѻ`��og|�N^bۯ~5���He��>lt��oNnk��V�m�=�\����R��@�'W�����UHт�r�|����}��]��옃K?�޿	���H���L��?�;EH5ygD�j���f`^��r�����I� ��uʯ��؏瑴r��,*e��I�l�a�6�nл�+v��46+&]��1@>q��Jڍ��v ;H.����Oԓ�6��I���~u�F��h���4o��+��il5M�f�u�"K
@4�xWS�a?&G!�X����m5�ZZ�������U���)���[x��m?׀ڍr��Ò���7У��|eh��TD��u�۩�g���L ���)�ݛ��o�iʥ,Q/'Qk�ٽ�E�CfN�N��-!YV�J��9F �t��/�$��ʲ��eJ�~xz�S5,��y��C��yh��ڰ$�dG�������0���j�\�IB�ל��tD{�k��H��UR2�Wh���-B���ùB�9��"6�;�d-s�,Yrs>�"-О��!}?��3�+�/�!H8�f>r.���w�̷��p|� ��v�X�������L�"_���B��;�v$������{�<�2ov�O[�"�����f&��{?�Dه����q��2�ha�4�ITc��N�k�]EoL�/P�A�bd�n�r�q�F��	��#�����l���/\����Of��l�)�� d��ȯ��A%�-y55��u��u�u�;��S�1V:�yO�9)��EeFd>\��Fz�,�b�x%_��<���wfH����|�h��3��0&ܑ7��H��l��`_?/ʷy�Y��Jx���2/cs����,I��9�E*�J�I�E_����� 
ncc���KI���������y`L��^��IW�L���}/by*F��4�l��g��S%����<�g���CJ3O�[Z��5��$h��:LV�Ի�W���|�tX2Һe�늡Cs����c��-yw%��,26E�:�0Ҝ�
��7��;*�	�wOyG=�!� k��OxY�-N�^ݦfP:?|���c[�QՔ�w�i������1B߂`ZmWD�C
#-=���ѯ�֓f�#�4j�Ә�~��&0�2$jd���"<�ԑ�d��I�^t�Z?�\G����q'3�e�*�uk��u��*E;=�N�6��t�����d�JnC
^��Lz�+7ė�����I��<=-e[��CǸ� �R���^ W!�V	feOpc����v̚ۂh\,��%�ڄPOz[��d�yaF�X�����	�zVSy&���ҝ#��gee6o+�-i����`_��ƽ�b���wwfC��������������o$m���X�Հ��ҥ,�Tn��')��I���Tr���&���ÝƲ��cR����hhtk�{���(����~ץ����C�ny{R=[=^=�\8�T	�����n�L]Ĳ0V��ba�Q���2�_ř˟���Ӛ�F�c$�Z�mLm??���DL����of=]E�a�U��09]��0F�Exz��n��ݘ��]�Fܳ�X��[9]�Wְ�����4��pC �YDh>�]_�XN��q3']7�`�옷�d�U���za�����con��Gޡ,p+�b%)���{�|����(5��ח�4S��G���c:?�p3��=���@��I1�y��f�j�?�8�$w7l���}+��}��G"�`M{]�E�cܛ4�
:�L3��L�P�A�q`b)�>.޷�a��Vk:S��\B�(Uܡ�E�DT���م�A����xn���Y�iۮY!���T~�>������	X�x��\͞�*��b{�!�z��!D��u�<} P����Z�;�-�*o#��#\���/k����ܘ�Z�!�X�*�GqY/aʑ'X-�x�.)'���?����Zy��,Xj-�f�L&u�ؑ	,J�F���	ׅ��c���
@4="u����p��x�ߎh���Ǉe��r7�s���ܫ��&��$a���1f����.Ї�UZ����{�ßo!��q[�u�Ѯ<���s���u��=s��
���NW-Q�݃F6�A��r�FF�6<ɪ.���߷۳�����i��VZޝ�p���M�Mm �/��Z%���?AA��}#�Wԛ���H�Y)`d�v�+��ӽ�N`/�p6h���ٔY.����u�b�r����KY�A���Ʋ�P�����.�m!�+}�$�h7��ܨ���9XៀqX}��kcN +�'���z�d��1X!��k���m�<��:PWoc��4�g���N�y����̡��9�k�$]�7���#Uv����m�j\W�^��,�JE`��Q�T�oW��A,���'�|=��'��ChRK�denњ���8� �]`a=�1��:������̗����������k߃�ۏe��a*�'���U�^��9�g?��Q�>aR�b�XYYy�[e;]f�M�w�ߑ~B��r�@��h�����Dc�������0��ɫG�_^&��Pv��ݻ"B��R|�B�F:�o�+q��e��O�\j:g�^��<[^�����/����'C�O���l�/v��Xs���%/�'%v�©� �啾�n��@y⑕ҷ;Nod$�ؒ[��{��Z"�
�X���3M��2>YG1�����#,+aR�ķ��]�P]�˅�����b�]E<Kwv��`�U}�폖�����]�ew�2s��̕i��+}�����A��E$=�P����������M)�Γ���xu�y�D�N�#8��͹�0�@�O;�ߣ_��V���$�A��+����*3혧�쵦�}8�'�W���_��9l���U]N����a�)*(�`����@+�����׍�} �@��M}�ͱ%
��S�����W��.N��4�1YB/��vP�N��[������ޠ+TqG��
f���谰fP�ll�n=^���4n�,/��	X`V
�e�{du�+��NsZ#F�>"gr0 %�&T��T`Ӥ5�|� �/���ϡ��/Q�r��Ή ��7=�Z)�}��.�C$�	��z ����-A����\mz|/z��{�9SZh*����Lڞ�q�iA��S���YH�H�b�!�a�IH#������Tp�09=�	�h@r0�=L]%nNbZL�#w���l�)�S����H޿ؒ��d���m@r�"hw�i�)�̋�2Yo��jk@�{`�������1<�L��l��$H�nT�vM\���y�My�Ie�@H0��Vҭ\�k'H�yOTF�#A�W22�խO���w�e��(9�Rn�@ꌧi���!=$��f"�7�@�!�5�4�8\��ԭ�a��f�f��ee1W�߭��>�܄Fo�q����|�TY�+�*"}d>��Fms��f�Oa��B�����%M�t~�ޭ���8Hkl:EM+
�+JÝq_M���d�-0"�M/�ؔj�[���VCb�h꥿�z)���l.�}��<�G�H޲}?�f;}�+�⥥s�W�y�h--�����ZF�(�~���?�n������Џ,"o?�Jk��,UZ�x��v��茍�U�N�k����s� -�Wօ��.;��Ӓ�J(TO�����n׈j7+Ò��o�;�`��h�5ګ|F��@ui�f"��lي��*����]��>��-��y�Wfq�㛆/�#*E���xN$f��d�����ׅ��
Jj���_gV�5ԕ���
��֕�땪�x��������b��i�)dyG����u���v>�Z��<!�)��_���Kߴ�����^��n;$%*^c�2B/���,=�����8Xq:][1����/��H=���:�|_M�����	r�b�4��"�����	(T�&N8p6&&�gE)\>��6���L�D����]���blC�y����g�A5�4�d���%0�2Z�Ӿ�ʪ(ڀ܁Iե���=�A$�u�5��	�M�}Q�d����NY������B�-���׻����X�j��a���)P��뿇�&)Eˑ�i��an���+�Mx9��tN�M�H'�0���WJ�9���vBt��!����u���6#,��G
�j�\�vm��@LU����r�sq��ߵ�;*�cb~K2�������9mgg7�������ű«�yLxKFW���ƞ�K~G\�dl�g���]\Ssa�3ɿ�ߨ��+p�LX��|�~���(���j�k��-�Y:i/Nz\O2��Х��}�7��V�.�����zX�3�LF-�^9�ir_������2�4�,�f�U�4�ǩ����ScI�i��y@����Q��NHvNN$�Ʀ�Q;��F
��6�b2/�,]}��O)|6�C��>���$"o;[.*�I���Q��4�t�b�q:d�&�PE
�Ν��(�<���2�nrfܾzu_�������	�J&�+G(7B���I l^>�{xG�r���"v�]��&?���v��U��S�J�+�X�^��d�Y��X���ȌQ��7�������[��Yvw�`}}:��,�v|�8R��ق�%[�h��:ٝF�_]�~6;y�١l���i{�N���A��޽
-َQ1�%7�8V80`r�R �nC�ve)_\��K>>��F�:��S�M��
y2���koW}J7$�<m����A^�ʥ��.����=�w��.+�bUC��}�I��f��� �`�8X,��hF&��h�#�������2U9G��YlK)���^�#RR��K�E���	/������1��/����r�7�>�EP��&�R7x@�p���ano/�s�xj�#CYF�t�f�zc�жc�*"�[�B�x	��1E�¶dIH2��Jn;_1]O�<�5W�C�=��G_�
d,{���Sڬ���-��mX�K޴iSI��0�n��{����
�TE�b|���"?��0�����|�	w�g�.�F#V��&�>��l'{�7[�]9m�Y ��%����[�6��Qr����,��2�DZ���\�����_<F=����y��۴�=(b��Vbx�F��[u�����H��\�c�=1�@{>�@_��aJ�'��!U��q8�al�ȑqz��W
s�v) J��9�=��~@Ѩ�~��N�p�v�)6�}T��f|'����`�*:��R25c��>2�&C��*za�`'$�̟�v�Ŭ�����A���.��,,�䣞�3�M|ؠ����	w[�W�}����
�B���a�"���`#�S��Ĭ�ج�;��£���0X�^�HiYq�ۄ�g�e�c�TI��
�4�M�+s�M���8IZϨ�PDr��ў�����K�w��d���Ҽ P�)%�\)���!��/**�^��}$�>/���G��;�l�v�˶SW�6�������D�w?�Ea�r"��u�K���v,e�HD�:E�tݤ���]Y�M��.�R�,�t��'�����n�|����^$e)N�E,�{��8���-_����;?-�4��߮�q�f��%��ڳa�%$Z�Flww���5H.1m��{�r��I�!l��;w���7�;���0L���O��k����9Ӟ��053#���<�)xLBb����:�) �)^��7���{��г���Ff��8&d�%�3݋Ǹ�n���$��I,���k�a�E��(��-X0��=�g�s@��8u.�����n-����z�Ny����� ��޹��G�AR�)e���r`�ᙃ��r�>J$������CO��B���~��Y�|3B�7'��t��1U�����54�pqq��� ���OOPaxA�t�ڳd^ }}�x�6�5�L��� �'&n�F�hfE
�� ����<��H���>5>&��hE���4���Uss����j�'�c̋�.0�ќ����L��B��;��<q�̈́q�d}0&B)��<h�ƍ���@�Ѫ���e��6�! #�w+&|�1J�9ި��/���Y!xF�X&(qp+P�,l������"bV�
I|h�)��ՍQ&A�e�V5�T�X�c-��f�g.�O�����F|�!!��@�xf��4�����Q��7�2��s,{��f�>�pbeeg�:������a������
��NzT���Z���x���@���-��2��}^���]�h󪲅��\�֡�1o�V@�7qq���uј$B1���d~��
~�F��y��#;[��x_|��j�hw��v�+Gl�Ϟ��k'@�� L_�a���.�I��)�l�w#Âa�c�O���8��-7X-�g.�BCp���nX8#{�9� ���HE�ջ�28!zޖF�{::\��+c�������h��ڪgnn�]E=ѹ<��S{�S!~�VLW�7��$�,��s�wtt�����\�c��{h4MVz�\�=s����6p�݇��===_à�����Փ��)���M4'��i%d�t�D�tyQ��d ���Ъ�<7�!�H��*�1D�6!M�d�ک����=@Y�e"|�#{����۱?�5��-���T�R���|��cf~aA�g�祀��y�> K�I��¾>&���#���jl�UE�h17O���vWtt�	3y���C����;x� V�H�G�Gr�����[G��J�op�m;�a�g��ҬR��=;����8��B#�@�c��1�o�n+�+҈u��7�b��8�SH�*k�WN�G�����d�q�����14Wֱ��lM�Vɢ��˄�S�a?�]����>�촶�����*)I�F�6��fؼ�4�hn��N���}�\+QT5��?�:�6��t�Tm�D�F>�v�3$d�m�V�fb��<1-M�gv����]��������JryW�:hh��x�UtG�?A�"���3����p�6��\h >ؒ��y7�j� %�)ioz���6�i��K���+�c��Qe|B!�bء����*����Փ��B�Wh�N����K�������'0ݍ�6��L��?N7m$P@�1&��%�'�FT�(��	:M�?��2���U���}�����k��� ?%����U�ꂉ�����������*TcҰ�R�/J�\��#pB�1U"*v'��T��H;~������-����0����=@}	��
ВA���>����=�F`rF���1�E�|(�SE��m�@����6�C�rtrR3vV
��|��sW�;lX�|�	_Aֈ]�3��i��?b���q!t/��[�����m�xs<�B@o������zu剷�� ��u?�Z�L��[����?E�����"f9f	�����A�8W5���>�jH�޼���y��h��OW����P{^��$�"�:����X�p�`Oqo\����`dQ�Ճ����C��6I-'�bd�-?T�e$���##����Kg�b�iy��چ���|.�!�m �ސ�wF���{DpP��q�%)��V^�́ժo��XҚ���:��.���w,�#A�<� ��9 G҈U
�G���8�0F�{d�i�6��J�0@^<�>�O�LA�# 6�����=�U��r�?��Z�?�`c*\�fFR��v�A%����� ���zК�;6��?.���ۢMS�(3c��%� �*��-F[�)���g�hy�f3��Խ�6}`x��/��:lO����Q/���n�w��bn2|��2�W�1��*�V&�Tَ4�Z&�SB�!x�{��E���b.\�t��r�;�%�N���m�����A�'T,��$hhG�=�y�hܔ�]��������rG�ٌh�_J���^����.���ܙ3�Z|�Fb՟ _>-`<�٘YY+:y�鍓�'_^0�j<h�H�[0{���~?m��7�g��I,ި���������I���n<5��1�����2�.ށ]��_�����
b�,^D�>tE��X�,�8����3�����Zئ�_jeq��4]ᤠ/��C0����2釉�;���V҆�R)�]� ���0)�d`�i?dsO2_������)E)�NI0w�%Q#]'�|�`�	��Yc�j���eה;�3I#���e$��r<���x�&KW)��Y�Wa�+��B	�;<+vF&B9�n��'ɽ���&���{ϕD/�����L()�hG�3;SE�RXx�WY�P��k�g �M���\(/	N�W@�`k�2xz�{�&���=	z{>{�Ī���x3]�DnS�5��4�VQ��R�m@ං،T�����4�`L�&���{���i{��S_��a�W/1�O�]�`o�w��Gц�ڒnj�+�D8HX��'f|�v�'jj��>p�5X�M��� ��|U]�B��K�6rG��b���F�0�#""\Y@�HU�����9�W2�\[��)���1�W�����梩f�ٙ��D��¨����m�)�����
�Qs��+n�זC2���������.?�aw�B�:����L��6,��w������x�VS�O�C���YԺ�=f���[00(�~Orr�2K����L��X��{�K�
���cOR�-����� * �֭�4�t\&�]�� ⛅O�
�ذx�4��f�(�߹uk-D��)���� 8x���͛K�*C$]�ª�u��}qNN�L*ku�\6�fJ�#��=(5����Z~���WBq�����/_qv���d�y4i�RD�Wp�c^�R[�T��U�q���ۏ�F��	Fb��ѣ�\gÊ ~������7.'�~~��3�1Ug� BQ�n�/�i�_`�9�O�I�[q�yR�~���H2tv��/��	�e(.��E�6�!���Pr�L���,���v��s�;]�b��z��0[�G՚��U��z�?=d��-#����\�2)2?�N���ÍIxM��s��son�[��a`�c�ð֧�2/�L�����7zA�Z?l�+H[�vv1U��۳m��W`�'o9v�ϝi1%0�k��F�b��zϟd�qzg�N҅�{aU���LR�`�`���7@��T���M����.��'D<yUR��o>�=�Em��?rL(�L4x~bo���(w�����6r�N���I�NEr�B��8m���<%��[��'��p�Iw�/Y'7P�%�������x�e����f��Sw�и������;��Mu����X����Ζ^�l���t�ȕ�����3ݎ����,��R��^GȪ��n݊�/`104�_��k2�Kx���8�n$%)|�Þ*���m-�"�zX�R����.�	�Ô�2��u]����v=!�`0������ß�c�l��,K��i����"�+��vc�I��\�4P�:3SϨ�ÞH�L,������"r:J�8_�Wd"tfEF>�L����� ����p�����$Yq����$V
�C���2 XՄ�)�t?)1���B�B�b��l?qq�7��V�>w1���n3O7�W��@x� 嶤-Ex�*��\������[&��7� xE�8D��G,�h~ZNP��M�SB����Y������� jO�QbN�e-���H������ `%��`��8��d�3$!����}*A��;@�G�l%\�.؄k�􉲜�<^?W(~�
�m.��<[�	��i|a�.S6nKӤ^�T!KכvڢQ��YM��a�y��/���$���������6r�b6�7f�Bv�'��í|����v��A�h�e��š��4֍nÌQ���K��G��,�Pc� ���ާ�Aߪ�����`>��q��"�Y�� $�ԩSy��||"�rHp��vb�@`�1-�����|����ĭݟ �xR;��c����^����;X]�����%��D��
�MF$mdl��~B�L>��&����&��0H�a�)<
���O�W��׫�5��*t�=? @��yk�E_���욨�+�q�uu~i/!��&�}K�`��m��ok���iʴ0*�΅����{�f��07��J��w7[�t�C?����,lYdAp�s��I�ֹM�F	�
,|����=������6���.�2���5y]�֮X��Tj&�d���*��:,�ȏ�9<����%u�.j�]�v�e����a�g��5m�N������jٖb��_�� ���:�2�=��@\"���g���KՔ��%��|}�fh�?FÂH��'\#'P��4IF��?Q��ٵK���<��)t��SXTTt��<��6[������2��a������ק�] SB����a��A.)z�9�p���Czk��X5���R�:����Ae�]���7p���
g��a^���C�����7�?�J���_��K]�W��G$��t�6ƪ��C���槭xpU�4�ʻ_g��ϱ./u�Hs�w�{M�����ux Q+��Ex
�2)�u	H8� S�
�t�/�7(_�����SkQ&8�Ç�Y�\+K�Sj��d9~u��\�q��VG�8ѕ��sr��ج����֔��\kJ B��
%�ӌħ��u��[�-MF>%v�y��^�ڗ�<?�4Bb�c�����aEz�Ios�t<:4-7�_lҮ����!��Mf�?��_;<Jp��R����x�w5��/��{� h0 �AJܙ�C�H�%����"�y��$� "�òt��FO�q����� �:��(�����<����]�W��>��.�LSK�,�|�o�����9�M� ��<��*g�N6Z��.���	����ծ�|�f�/�{�t�X��?��6»���Z�.�w���tϮ�.��Uu�����66�%� �Dn5�3��tU{�g�T�{2�D�E�2y��؅m��MN?u�����Q�U��<���c1{-�]]�!��t�zuz�U�<�5V�������R3NLL$M�"i˙!�ś��2K�� 9 v̆�u�r/�zI=H��u1��͕�0�т,���i�������b,�$*W��=�@� �O ���q�ͷ_�
�I�8o�z�VK�!�/М�S33���0�od&ӜMZ�AfھZ�G�lW�5��ķɥ;��V_"�v�͆��z�~ٹf�,�}#����ov�WZ�nd����a�������Ӊ/����������arP���,Tc l�tf����`�r�4ʋ��QO�ż��b���>H�6>->���C@j���,��e�}))�������o�myt��~�$dvq��^KP�L�'�ج�m�W��b�p�O���Y6��NҪ�-5���G��NM'����j�J��J{z���%6��r|�r[����f�����Aڡ�,���f�C|�y�w���/o����޼sl+�L�� *^�n���2��%K��)R#�4���2X6��֏�}9ߤ����+x�2.�abZ�,`@��4T/V���%]c(a��7<a�f�邚ȶ�S�XRK�QG��a(�3�MX�)S�č�:qi�
�����R�v�ik��rt5�*��'��v��aǘ�.�]�/ΑNL�C���:����[ Ɂ�sa������>а�5��0׈�/�*֫��M^|(\?QH�P�`����Ç���R&OA�cͰe�5G܁}�eD�C)�#6�o��`T����l�����y����@�!����x�ei�5��v�lW.����
���	WApG!�i֦v��������L�"���6��Q��ӳ?�-�Gn,22RE P͸�PӲ�eݲdH�K*"���c�����C�E�v ݸ; ��]�[��?�~�R���nA��OҴ� �q?"�thy�s�dn���E	iF�hrrz�2KM0:�@KeW�3���3LȚƋ����?.V�Bp�x�315WE���3r�\��c�/z�~>`F��ggٽ0��[��N`���S��P��ʂh��>��?ءw�(Z��h0���)Y�399�{^hrE�������%��"�������ץ����٬gGy����j���]Җ%&�	K��MCq�ef?F�c��_�빟<�4�����o�0!k��վ�2�7��2�s��`��?^�J5Vx��J�c��Y��lI ����	=�@��e��!���o>*C�<r��?�h�-Ja>r7ֱr��������S��vE�m�h��9w�)�{��]��_ʿ��߶la.׬��#�UbXG<_���d7�h[��y��7����$�rcQ�3���J�q�d��:8k��n�Fe�� o>Q1�HTR����z��ʪTzeeէ�Ƙ�߀_����b3H"�yg<	�N�%i�Ƶ����A
��lŚ�z�"ۑn��{����~��Ƃ�*1L�򆽎�h��YDx`��Y�^ܴy��#X����w�B����ğ��mt�R~�r�����+��y\����j-�#��oE�q�yze<�q�&��DJu�Ԙ��� &y�R�,f1x�4"��s���29vb-2u�ϗ�kע�'9�v�vt�]���G#v����4����	�;+�Ԟ"�_x��={��H�c�^��Xﾚ�D�ۀsC����>BySS�=5|7��Q7�R�����i@�'+ӳ.�g�-�BWE�ZѲ~�,�9�ng���=:\�2�;!3$k'ç��ꂠ9�Ֆ�硝�툛~~H��kݧr3f�u�8���^���jO�{-��o��v���@V���C�&d7���m�]����ɑ��Wó/����qi����W��d�nza>B+�e9��lm�bz@�;��o/*\����RO{� �*���"�y;�HY��t�I�mq��T"�K��t�,�:Zl�dd\�ZZ�@�:���콵��$t$X�_Cҫv[�$͝��@@��"���U��`������odM^(n�V|hx�j3�@E
���Z�IiF��U?l�{m�j<����+�~0s>&���q�R�yk����P'D����Wc��7~��⪅`I��ɧ�6��'NDG`��>���%NNe�8$`�x�$˗��� �Ng�ö���px�4GG�վh󪘪{�a�xyy9:���t�����^��O��_B] ��7��#|��B��˿�W���2-�����i�31�0s����T��(��u/p�`	3�G�[�Ҙ]����`/��o	:���	��Ǉ����rz=�N��N`n�P����j��x��\��ҵ{u�W\��މ/����v��� ITh���C��� �1[Y��)|xϞ����p?�J��d�G�n��&��mYV���7�8�B��l��4���T;0�����~�ؚ�Tx3lV(u�?4!����f����V����
?�=@���;u��e��ؑR���yٌ�kƶʍ9m8_a1�A�ѳ����s�� �Y���9ݤ��6�f�T�d������a1����Ax_�����^�i/ͻ��s��3���@`
f]�Y^���q3������s�~f�����8���ǹ^:��_k֮7is��sj�)�|�mq���Mw������ռ�}Z�@<1.��fz����i���^D�����R���rN�Ä<�[�M8��f@��_���d�� ��t��ޮ(�����_���_#R�O[?mgcS200�_p4�ʺ���m-)`���D����0̰3���i�F$�uUXn4pk�$3'}�	w�}���bڬ��rcmO�'{ܖ\��Fg� 5�X�P��?�l9�FUj�Ȟ1;=M*�Q��$:j�QUA����x,�mH�~�+ى���сr{'@%	*���	�zp X-@�8����C�nq���#Z�����C�R~�L:
��:W�ֱ5�����c�3�?��^A�1�v�x:��x�E�r���	F5��X�.�����8��'ؓ#F�qc+�'�" *� ��T��~�V�<f-'�:�7(]Y6qsv�Gs�N.ߠFq�`ǆ�y�6_	��c��9]�D�ښ��{�Z4��Ar\1����M��ã�6~��l]���uia��l4т����9�]v��=�ѕ�7�k�A��JQtJ���|ie�����l��ů�ܾP���D=^�D���,]o�dQ����)+��řV�?��[p�hZ���o���Kc�Q�@�}��Y��P�����FU
��h�2���xg.ʄ�p�R�� ���gNoA���+�����g[J��4rB?���X�Nf����Q��7vyɱ���,-����-�q���e��:������xX%q�;:XCfaayT��+x[zYĲ_��J���,c�t���1��]�(W��} ꖜ�Y60`�V�ø�:"�T��Q_H�o�N@�����iǡP�hX���X�Uk�AG�<���V\iC��+�kp���)+�z@ب���e�X�^yNN�!����[�WZ� �)s�ssW�e<W��&���,l �ucc�t��-ȭt�����U �.�g]w��e�Z%�G�l�IN"W{w���jQ�xL6*���P�|w��y,�~�L��Az���zÇ�lj'\��;v��m0&�%&&1
.�t0v�ZRE�]�䴶��6Ņ]llؒ��׀W��p�[a�=�l�y�Ȯ��X�|8}��@^�*�z��ږ��
sW�9a��̉I�����1!��%i���� �ϰ��1�4ܯ�V�h�����8��ݕ��Z�\$i�����a���缼pزߠ�<p�N��g��<pK��{��s���x����E[g3o�Azz�pS�
ox��\��[��Z���}5�w)�&���=���9������ޫ	x_�^�>Ӹ\��$��߻A؝�j�����k�I�Z�mڷp������]㛛{�������ݗ����;�R��~^���/����&�e��z��Go����(�Cڕ���4�d���+�m"�����B�Q��c^|���J��׻���BB�`�����ɰ񁮢�\��A�/�;v�<�å�������sp'{��%i�����tZt4������?8�Pe���>lQ��l�樯�M����&�?��'L�g��Nxz$��fUد��z�Å�A�q��ә]
 _i;��ׂb��r�&/O����g���K����9U[�j,8���Y?6�ћ���H�E�]s��=x��eJ�ȧjr�-AF��i��˯�s3Z��߹�ٿU��9��)w	a�-Z��ˉS֔�i��y��x���V�wG��G���b&=n���j*o�tPTT�Z���J�w<G�w�aL��s=�A����}�Z�2d����ǞkE�d�W}���_�ҡX�	E����t~�K����#���*akN^ay ��i��O՟����q���w�|�n�ڷ�3&?�p��3L�M?O_pD��ʥ�nJ&H�b�9J�ܥ;��'$�Zw<�}������c�~��s����Lѝ~o�����=���c;85X��Ln��d�o�a5�G̛�q`��`\�������ԥ84sڿ]>���汗Ns�]ͻL�U�/)Ӑ��1&_Y���}�(���#nǦ�=;�+�X�_�pџ�?��K����O��8���w�w>xI�v����I 5Xܟ�.N덜�b:{U/�o��9ⰵ?���>�{�A���9N=���B
L)�Ռ^3���wa��gnf�5(N��v���-O�s�x�=hI7�rf纏����W?j�0>������/e��-za:�b����{�k��������5ΘG��5ȍ��l�vy�V�7��1&�_���j\'P�����
;S?�m�k�gbb��4pu�{�����8u�FF\#bMk�Ӵ����7H�H���J��@���٤������`���|Ϟr?��̣�����-u���g8�K�D�]A��#v��_Ue���+��y8y�,�k��f��l������o9[2��%EWռ�7d�j���d�CSk��w�9̤�OoR�]���\dpD�C�tD�p	����_�s��I��kM�7lؐ�8�6��z��܇I)�G�v[F�O�2;�����*a����g��fh�!����p�'�r�˧W}�UH��>�rwE��cU���6?����0��qk݃+�Zo5�ut6HV��L�n�������Mo9�x���1��^��?dF��ҽ$ey�I�i~������G�!p����zS��)KO?��*��/c6��� {�y2F)LU$�Ar<7���� ������٤;����8��<=�����w��eFe���[�Ԩ���M߶�%K��(o����7}�?Wi����Y�����3�b��W�W�d��9mC_�UT+1�}*9�奤l���'1���Й���aw��g��x�x+h�5��uKD�nc��$��W+�z���K;N����r��
�g��A���D��-��k�v&q�m�-Uˈ-=�Ƨ泵�,cy����>x�-���~:���yzp:%{����gk	韖N�j+
��=��b#O��*��𒳡N\��w�4j+9"vҸ�=����uG��;"��/�V[['���	�&I����s��ǫ��6���`lM���zIQY�g�3�iv(�?��u��˻�i��.�R@���oUcM\\��9�������C�*:�����a�+��z�Z��G]���(�LO�tsVAd�id��L������)σΪ>���O�ˣ/��>����
�L�����=��e����ۼ�,3;�j� �?{Eo3S�p�F����7v����o�Iφ�-=����/������4ڜj��0�.�6�����R���p��}	z�jit��_��$ ����!Y�������`~P�m<�2c���8�$�k����x�n	Q��޼3YKA�Z� �����\�յ�~����t���<mӮ�<�9���7�x�ݹ�7^j�F����|Pz�9��{�ii�+��T���:��>���r����t�qю��M���A��בg|�s/p��!I�Y�G=~>>��'���&��g���Zh#��\�`LؽyE�VU	��SJ/�r�@k۬7���v���&''S�L�cZ¢������;�ͫ<�*˃�lb/�b"�1
�4�����=�I��= 䊨����,��ߨn�D_������p,����T�$IFG�
��le�gvvFh����l/�+�!!��MIVFF����}_�����s=׹N�����s>�w<F8DM�b���~<s�%��������Č쨳�S_S����"֓ٓD/����<7	��<����Q
m����hC�=�K�~\K� Q��7=e��{:����*-#�iA~���}F���hD~6Z����>��IG�:�������/�����b�2�ѽmQPD$�������@g�@�ӹI� [+Oi��L�� <��L�zg��S)ޫ�G��=��o�����ks��T����Mon�0{s���-���Or��h�X����:������r��N�_�
F�sTA�9^%���f�	�슌���zeBu����������{�K���oԉ�B��=��H�.O1F��`��Vj��~G��T_OQ����/�[(�NVp�b���+�MO�w�/<�Yj��C��Z�����b��ϓ��n�.r�"��"�_�$�IJb[����߅�����Ӑ(\��9�vs��P=����oԅ��F�B�kK�n��L�P]Q����>�}��R7�
JK �x��?=%/��V9p�'�q7z�ɉ D��Wo�{���B�}�6!1�B����)��|���)������mm7��4�Oy���5�T7��`?��8z�<T.^�(�}`>�m�sm�.^�"���_�!��gzĚo`b��־_��Z�������c����Vy�-)kG0�x��,��fa�#��	�iߕwB5~���^�Q��-�8����s��P���S�"��c���5���Nc˗��6���q�}�����pl����9�i�����n�����h�b�2~��'u�Lt���@�h��q��06��Y�H��R�zg&�*����)��1��)���	��o�OIVqfLN�%���v͛�{�g�����i>~���"�{��彩A�נB3��5���k?��sO����f �L�����I�����kP��U���������U� �Ag F��C�k�]���M��������s?�kfr@�:3_L��W�'�q�B���`T�@gg�6ɕ�J���G�D��3I�-^I}}�?�����
��jL�Ŀ|��#ÒjR�i��؜a����z����/7�gU�6��s�,�s*Y��Y�<��:E��W��P���{�����賓�����߬�!p�C$Q�nN�W�j��Y����aGʫ�ˣw����{��FMvq����Xx�E;!G�^A9�p�<�_�mp0�������''�B��|��!R�eN���}u��_	2�Z�p7Qx:1^t������f�&A���,q�ש4ҹta�%����p:����߮��<�
qz����bu퍊�D������Qξ���݇�޼��*��K����#��:$�O~{�ܽ�@��!�ԏ8hC�������{F��L���Ui��k6�rZ�7BЉOc˶|=e]��Cc�6/�D�H��{��s��S�vΏ��~*ė�*�����.����aA ��C|\��Q1|��9K�e
ܙ[�2<-[O������=�BK�����^*,g�;��;�`�����T��cK�<�Q���D1��t'vxH�߯��j6Zhw�`�6�-��P(���K��\?�.�����{�K��4<�Ć�,36�}6�����2'���y����������|q�}�&�ϼ�ӦW��Ry��lB���)�	��p�4I��/�c��g�M.���&k�(�?(N����isy���Ə"Zn!��{���:��Ӹ�����yj�P]`]r��O����$^B��+�A�C�,�iѨ�o�y9�$5L��#�	���zc���_��`�����_�ec��W/��1�`�>����$�`������:�
O^�SG���������f��L_�����f�4��H%v����/����D�|�F��k�89S��N�1��]5��:m��!w~6�_ ���q���2�MW]M9LxAQK���l�0G�J7Y�I�~]=��CJ���p�������Rm�D'YG��q�YT������6'7�!��f�Kh_T��]M��|{�o8����EMI
=�����_����_�4~?�@y�%lowp�c޸��S�F;���=�g���z����m�����w_k�jre �rӆ�̷KX�.�Mod�s�r'�� %ѻNb^���0\Z�.p������en�=AnR�lC<	߶���x��LJKο*!� 1#�U��M�cHW�9q~��qΔ����Զ͡��L�󝕄7U�'2N������Iݺ�"B��(�Hcؐ�cI�}�R\�C���f�{��t���
\�?��ü��;��P_��QL��X�{�ɵ��j�i D��,�[�/d��hO��9(���؟}(Â�?���uʸh����N�r��a�����'�����sE�ox�:�[��5��Kr���i;��;��;�)��w��G��	�~U{��9?�Sx��v-Ƿ*�p�+ �0!�1��묐?������]��ݿ�xl���G�|��bhl���Im��� :,�q���$���_�o�
��4ϝ;�,�9�O�0�JjN</|�^ۄ�\.��:�ȥY�B��h�L{�����1xE\.ؠ��k,c^�������V�7�^o�/���$�{��}�sR?�h��*�����Y�<��\��d�5֗����7S�>�ct������m#��W'P�p�����z���TI�"~$�C��~�3>|t"�6Y=U�nʈ�c�`�h����@j_��,���`\���X� ����c��qζ���'Z���6�A����d�6�o�=˶����&Pz�,Y�⟠�����P���Sh%*ɥ�Kr��[�xب,�J*̚�����������9h������v#�<�%B@�{��鹶	%�?yT4!%E���T�h�V� M�J8�>һs;3��I	י��鱵�t�]���ӿ�%��cup}}��Νݩ��_|�!w�����"sߌ�{����'t�8=�;�a����h@�)bzi��u5���J/yT��C��A��8�!G�Z&�*��<���7�Hdй���i������O�l�����'�ۯ���}�;y�Vi�M�b��fT@Eo�Mz�+�d]�v��d'��<��|�&�����W�v��W�Q�TU�{=W��<��ɦ͚9A"�X >����neg}_�{Z�]�'��e�0�#�^�r�#:>TS�co<(Uy�QP5�c;eX��,�B����=Ē��0	��P���9��Sd��_Zڨ(\�W~HR������K=�CRW'9g�(;ز�5���^*�[X�*h��Ə���lm$܍��ƅ����w��8��q*?I�bf#��
R6����ŕVT�XW>Oq5^I~=FA�v���CGnj�,��[���-���8
W�a^�F}/��z�MT�d��㕸�Z����OD�3����K�LF,N�9�
(t�o�'���Maˇ��-n�D�	�k�.�G�Ug_m`/>��v�)I:�$E�Qfއ;͆3�10ɝv���NZ&ݬb�QQ�i��i�d�S�{�	��&
'���ړX���@�J��U6��u:!�VYy1�����
���֥�q��|���o7�.�R���㶍�����p�T�St��Cn.����ȇ6���Ʉ����\��WJ� ��^�*)��e�����jGЕ�@��G�3N��{"��ݸ��ݟko>��|%�jw\��a26���l�7�s�J�6�]U(6Yi�:zݐ��/[ƺ�V��m��$�_P�NR�+���1$����~��8K}@��(���L�=�:Ÿ�FE��o��:��u��WD�B\�I�/1p�P��ipSnu��u#����Z�d�Fvj���ŵY�:�N�y�uG��|�j��=B>����$�mk��D��V�� ��[���4�;��'�h����#�� x����.̼��K�]U@#����vR*��.""R�RT�H]69%�5���$y`ʯ�����G%���^�/�7��rȰ��q҇�;99�:�^�e
�<{�ӱ5=��|T�%�p�`F*�ϩ��5�_�ܴu���!K�x��N�����L�Az�f	�n������_��o<d�&��[�y-�455˥qцN��>=��J&?�=���*>���+/+����-�3c��&�֪����s��E�v��l?3�k�PH׸o������(��c������z�C�$1ϩ�|�����2һ׼��{�4X�cu�A�ʜ�[v�:黎�mVn(��u40������H�uu�)㹄�� ��}.s�j�L���J-v{���ч����:y��os��-R��>ny�v͟>�*�U�ua�6G'7lYg���N��hP�]H�uU�v3�_	?���~L�k-zeU�A��ӽD�;3��"���	�*�	P\���x�pQ��f=��I=�mY����$qo��Ռ�̀��Y�n<���z�sdt"��dUԦbo��N�v�	^���&^o*6�ލ1�^�-����m_�����q�%-vzj?���j��ێ��IM13�_�u���s�-|uyhS������������F{8���Ƥ<�������=�?cވ>��yû�;m`m�u�qi�/���#Aq��kV����j��g\��7�ϱ��'2,GQ[gm����u�֓��2��x3�x2�ʆ���-�7n��AJ�%n�Qr&�ۑ������}/��Ctr<���K���/=E�V���?o�<�u���V���O�I����w�����E��ͼ���̕��=�� rvlل���蜦{6
�*_���]��ݳ�ؠ����I̸�����m$\8�~���&��e�Q�r�N�DҞp�-.u(�M�n��I�	��ڢ��`�ݜ�y�l$m��-�3�!�7ؿM�B�|vݎ��faeL����w/6���pr2.e7�۵������h쉼&sV5YH�b���X���K��#A������+b���;�(��!����n��Ι��:�7��&(�վ����%��îD����t��b�0)�t!�&mllB�k�g-����	�h;ym"=Τc}���{���bC��کjj�F:Ž�A�/��]b��Z�_պ족��D!'�s�U�L6�D��Pu���C��T
��d�K�/���:��������DH� ���5i't�f�4�
j�_�8_�L�9��Dr����L�b�~�'�z�)
���X�ʪ|���^�K����ָ52*��)	���0RڄN�ٻ
b�϶-��y����:���+N09m׌29�Pc����D���H�Wzhg�Wz�_�3�d%w���Ҫ!5��W���o����T�.�g�jRn[�PE�.t����iY���K^j�Ƅ7����s��� |岃��MTM��N�r\RU,�Bq
��IZ\����1ڪZ9.7J�R�J=�O>����這�C�4 �1���	�	�������:�Ie� �#�%�s�b�??�D(��h݌u�5(p��}���OYaQ��)
\5�'�0=�kd�1a:ame%.7��1�V(��Ԅ��P��j/���0eL��s$�Q�'x�@�|&-N������E�?ST� K�BKo��_��Q��ڐ����P����٭&A����{|(����5�m|�j6�'`X#�����>%V�CR��'�;��fAg@�p��t��ri�
�ͮ�^~���������IҒ���ȕzK�L@g�u��&;}���).|�ϑ�	%eeΨ�O��:;n���?%�2���,��&�m�)�7��R���D��"�}�4�QH/�"�p��+�x��6���}.��
&ٳ�������7L��Պq��i���˜@��$�g_�����L�M[GOq�	m�{����,4s���*Kb�o��/�(%�/-o����C/6�����ͪl��*�@7��dt���(���V��S�a�G^�Hlm.�Snm_������O 8f���[�����:ۿ��S��|��궷�b?D5��:�[�+�(���-��P�C���U��i��恱��E�~���Kl�)h���Ռ	��q��s�%?��R�2F�("�X�$����+�m�	 �+���L<:��uks}�xK���8�3���e/��ۅ|@WkS�i��Xp2$5[O+�����g�U{e�2��?���&3��)�I�h�du��]E^��'yau#��ln��he\S�#��<Ċf���7����'gʇuꆩ�;�57X�c��zM�,����:���V�S/ֆ��u�+Æ:���`�s̑=w�f¹�b 
���{�k�AH���	�4Y	
	�f_����<�vUa��'�����`
ϟ�O"�����Q0�v�6�� �8 �����u��*�!��ԝGQ�D�������.��Vsf���x�+,c����L�m�`��]Xm�]~���<��ْlP�S���T����EM(�j%r��9]Brr����/�#~9�{D8��U��0�*��l ���������I�JA�A.�YNql-�ې�������??\��i%pRr�W����"��PS�10�,9U�2�3�Z8���F���#,\�||ƼǾD.��N�ۃ��
>�ɹJ�J�pZ<\���(:�x�ȍ4�6�W���u4#^N�+2��.0�����\�-��+�l<E���$���c�ȇO|M��;�[RTD��\�ͽ��)�$
���t���O�K�c�Vs(���!���7π��7x���{��onڔ��46<��T]w¹��eEd�x���9Ӆ ��� ��yⓟ�����X����K^�ڼ�_���`q~x�r H���0�[���2�n*�|Մ�e�8c� Gm�Q��|ǃ&��Vd��w싱r��3>Q���}����͉<��9J��d?J�̛�A�,�ϔ/�����1�Ӛ.$#3s�'Y!�)�ZFb��2g���u�pa��ӛ������EW9��.�����.��v�e��K`�y2��}}}5�����T��7�W�HQ��j��@�3‧����i��� ����
~�����:��8���x�����9.VS<�~&|j����f��.�ȭ�L#޳�����$�ʮ�K�H� R��p ��we����Z����Rkgj6��O��~;��s$��,J�h����8J&���5滨��Y�§����]��Y�1�1�3����p鯿�Zq���KIu��^q��S��&�%�nLHH��>�?�ArQ�!R57�Q2���M��Pu��w='��x겇 ��a�������`��6� ��7d�ڄ���!��aZ�)u��jA�=��$$�'&�����@�&2mK��h�0��P��Hm��[�H9쵃��N�;e�ϡ����7k��`��!�r�w�D`�S�S��Ԟ�������a�d]����eLXYp��D��P����4L_�
 <÷:MJ��\v�nqE��1�Ǎ�ޒ�hfWb�	K䧝���t9�ʏnen�)��L�R' ��;����;�]Cè9���H��SKk9B�k��ݺ��|c쉰O�b,�ߝ��8�z�2����+�I�U{��M��\���)/S�ou6mU��:���¼�a��n-pR?�Sy�
GJ�Ebd��ZA��&R,�������Q��ĵ�/�
R�s����+ks)��/���:�?�Ҭ:^x3�S�<o�A�C��2��������{V�{�M-��4[����u_L9�qq7Ƒ3|�'m�`�2�}]賓%~�Xru	��>�9%�y* )A���������ǐ�1���]#)tk���>CU}���~�Q�x����b�5����2����3��o��5���J���g���ůt1Rt�,�l�1gᙳp��:u��?�)�[w e7�W����hjjB:(/�Q\���� 57�KjP�?�yb$��ai\q�r���̝(�<���� ������#Z�e���Mf�Oc�@���<��� ��ϕف�ԏ�l�R�(;?��k�۶�Q��!�b,'N��^�|m�?��S6���T�������b���0U'#�� �#�no����_�G��iUM�Zm��ˋ�9���VC��4u���i����lQב�����L^�Sg�k�V����լ,��m����E<p�E��e_ӺT:?=P��~m_B�L��W9�<is�+U�Z�<v�L��dʰӞ�q�c"���Zw��5P�w=�z����:�����w7	hF���~<D`�dChh�yc�S�4�N�(�u����,&��{�v��Ё��'�n�esi�8���� ��Q�|ß3q��$���a��B4�	 HG��O���ku��:^j��K�,��i���m�����AZ�����W�1�4�/e���6��S�|��}A*�6��ތMq�B�K�ē����z:>�l�d�"�zV幚T
�e1R��������l��S.���\ް(Q��k��X^^~=J����`�M���e�L�9���7�4�<�#G^[�Tm���y�w�K�0Ĭ!�Mԏ�C��t�:��~&����F���kN�W��,�{j�X�Bvz�=nO�^l�2O/���.��t9
�۲D>�9>�]�����hsH���%v��V�݌��-c�?h�}��h�
�B[��<�������c�AcA÷-jek��"�p=�A������64����V��|2s�A�s.�旑E��js붖nK��f��?�=Vȉ�C���)ᴸb:��J(�W�9��|Hh���4�!%�p��ʰ�B#-B*5����=�_�{qq��.{�H�����X�������/���5��%�������K�5֗��~H�խ�yl�-�3��>�a�H抃�C_O�~��ˠ��arP2A
3�V���@���&���:�K�x�����E_�_L�a�zU`�_F��+���8����k��5^�:���($�N]&����SI��� U�j�±�k��h��J!�66�Ї��M�	�8�} �O��ϟ���kg�i  0�_��n���l�˰�����k)۫̄�m��?���.�ޅ>s�a�E�M�co���**^3}B;�\�G
|~uZZZ���˛ߨ��͞�=�[��h�K*�N�qb~�����@Tᦣ���
�W�e#i�ND=��\c��GK��7�<ǚcΙzx3��'�hqY�A������Z\铓v'C\��3���9՝��%E�3��i��Z3[�#��-�;��D�&�|___,a1b�DB��\��u�~��T��d23E����9	Kn��c��%�N�n/��VU��k�Y�k��(Ґ`�%U,��)�鵅c���=��R�P �G4�;�۽�+�Y��[��~u���Ի�\;]��]��v��U%14����Ǩ�y��	b�뭭�ϖ2V�vd(�>2���.¸ۿ�J��UZ�ײ�@����C��)~��{.��g׽���sT�����UU0o�?��8�_�Z����UnQ�LNN�MǧO;&K&��/h�YWV6������E��Y��G�e�B$���zn���K���l�<o�CF�P;1�U����yK"���<�,�<Fd-E4�i� ��Y�j�� \ԏ>���ٱ��x��u{{��~��B&�{hԙJ��ȕ�ohU}� D��?t9o�Q6�rii>��r���/�qg��v�Ѝ5�������U$�b�Kf�|�(�x%���w�>66
�?��/�"�v�yϯ��de��2�е%��@���qr���$F5�1	z1[����e�]]���ʪ�����֜ԏ8�(��~� ���sysK����&SJ[�SYvv���]�x���s(�U�����?����n�Q��by�>5'�+��?aaa��9P���Z[[�R�8���V�6��CR$�_��tEKQ�S���`��e��A���s� 3���c��|@�/�QD7{�ױ�7�eL�ϯ�����E�{���`����ٙ�4��,�m�k+�}ܧƤ������dFƟ�����uy�min�SYd���4�͝��;�\�#�@9��W{�:`�zx�Wo1��վ{��Nx�M`K��0��z�uȚb��~;U�:��G����y�>�y�A�8P���ۋ�l��6Ŝ��G�� EEEe(̡��Qu��畼?ޕFu5�.Cm$f@KEb]��I��nC��/I�]���ᜉ�	��^��111`��ri �H7~�d���KY�:%������7IY��ĵ�$���9�Ž]Q
�Lz@��y��R���
��w�WDcZ�K�~kk��sR���T��(��2��WVZ�U�p�ޗ�0O�R����YJ�h@���oj���WR���YY�����)0���ͥw���S��a�sW��(�=Ĝĺ�+��:;9b���MV���瀨�)��������u�I8�I�s�֠4�ځ]����xJ��skj����0���Z�^@�o��;�"pl02x�-�gve-88gZ�f�~����/2�ɉ�\NLLLPH�Z���.6��i�M zK<-�:����s������Z����=�7R<F��A,���IO��a"CjL"��E�R)p�����#p�YB�j�}��{�h���!�G /X؈KU��vB���Av�9W�g��uujri4�����^GaH}x�&�����Ǐ�}�� ��G�C�A�xΪ���ru[U�l��'[3.�>]7\�Ǔ����u�>��������`��T������|�9	�{z��M'�N��\N�|E����%�1�'�)��f��/�Qx�tϔ`R���MĊ��w�~Lm�f�+5��CĊ�l��*�mi�S�e�I*X���r�8k}Y����p�p5��sݦ�O���M�%���|��+�}}�<���X��g�uPH�6�'�أ����g�w���y���o�Wh� �����|^�6�¡�������k�4'�$"�b�X���<������9�g�����]Z�=0�lR�^+A(%�,�]��_j�_�{�Ճ�j��~>>�h������*����AyF�ܺ�Z��u&���SQq�|�r���3$5���Y���3��n��� �������6b# ��1�G|w���� U��= دP�;��s�.�L��.��M���ʻo�(�Cg�� �T��L�yS��@�|�'�~7��`��Aon`��wȐ	@wM���ߒ0(s<Iذc$���.*ػ��Ƥ ������%�2�F��`�-	�A�~��j��3�������%u��[	H'��s�a�ڵ�f�9�,G��i����i����>�ַwpЄ2����X�a

B�댸Ujik�Ր�7p!� ���m�:?]�]
<\[k�ض[�����O���v�f�jVu�a��G��� �p[@Ʀ��aH�'�#�}H	*l��?�*�+RZ��9���-������ʱ��?o����YS�u @��z��j������A�h	:��*�[3�o7�(c\L�59��>|XV�A;���2p��2a���U�M���A�o&o<�.�pd?\��n��ek52��1B0��)��p������q�B�;�Vj�ف,��fe(P'Ooog��#��?W��ϟW�8�v�ߴ4⍃���(�|E��[���ְ N2���(>�?&a�f��Dt����Ç��zMJ��	#��oIpqsG��W���&cX�~��գĞ%�E�{
�A"zx|&��������cccP�_���]@k�1som���Vr��x㦋���kk�Nõƀ��H�f���#�`᪕!?P���%p�����8+�:�ekvv�h�Le��^�g�k��P.2�ձM���90�wΰ�"�Y"t\�Fy�w�����@�w��̴�p���h�^	�(�� :���f�&&�&������naq�X��N��/n:
.:
�5Ӟ-EZ��و���4_"�8Z��#�)����+��g��@�C�l]Z*<( �2F��e�/�{�N���q�*����7p��<m�t�D!�o54���k�wq!��YU=謭��Z $±c� �3�n���~p �M�:?�z�bY*�Mcf����rn�h	{���%j���89wv��5xh��W����y���������q��Ou�5g��!ii(��S���3��/�9�5�J#�/⣍��!�31u���>r�C��ݣ?yR�=�<��P�R���\�w) ��^(p�����2���9~���t�.Dc	^�щ!�=zgz0�8\3�v�Y��u*�����9A�}39�8�ר�Em�j�nnnNMOR��Y���mh�[U%���M[����kG��n�9hkU��`q^YI�#�%>�S�ҫ��Zr���
����g�D	�|���g�޷o�ǟ_��KKY����_�4�sRG��ۻ�����ghz9'?_�['����ܝ==Y�-��[8d���Y�?�X��Ç=㗑?����S�;~0���7��,�>����أ�:�L�2B=I*����ZO��������U��oy�2�Uɮ.�)�$��Ii��CKa��� �Ǿ����
rgsw)�"{:Y^]�s*ZL\\�9Ǐ+�І��6� ��0���G�}a�c+��˶���SSS�SCP��"`
v���ay<��!K$����fp��&JVb:ğ�B�B���Ag>)L�w���� �������'/�xH�4��Y(��便Bl�TK`�h��:��*��X�i�|FF3p�������q�|����*-��b�J��|} 'Q��號bd<�o��ȷ����]����;Q������i�!&h/:��Ǭ�J��ݞ&���:�Os��f�?!!��DDr�I0X7�$B<c���n鹼��%E��Q�AL�2��*�S��zϗ#�����:B�7��>Wɤ?u�s�U�e�7�����F��o�^^^^��yS�=}��ȋ��xZ������� ق��*I��yH`.=B���'�,�r���D{����ث��Ej|KK6}����Ȏ"몠X����0U�$ǌ��޶7��+�"&ְ<'#����K�������Ի�C����)�*t�D �h���9PM�ܪ3�va(���f*݃��7E���t�Vx6<��������;���j'�;�p8�m����ϐ�JSGL�򅱒t��U��NN1���4Kl�q����$I?HUnG$�Jؚ�x@�e��^�`��u��=`,�7�\��6?[��!�E������{���t��4`X ���!�<�NS�~uV��+��W��d��Q�̭�P��/����� kD�%?��ohٶ%k��F�$��kf������ཽ�s�TWn�E�A!!��o7��yf	��Ş�k���v��҄��3~>�Ga�,�DaD�U2q�j�b>���Ô�\��<�Natx�J�k�"�]]]�..��o�����":���~t��ڒHJ\!?91��*9tgUV�ࡀ�FE9��(����(���5��������H4`G�`�����C�[�h���X���a:EV��ϭ�-0��{����'��v�:�H��hiI�pcHJ��Ȗ�N.��Y�����Mԏ�O�q�n)*�_u���9��� ��0:�IM̌�#��F�����L�jռ�G�s��aSH����4�ݍi���@���o�.L=�����^ r4�����έ8,Ouӎj h�g��߿�]�a���rre)G{;;u&y�g�7�=��|
�n�ۛ�h��''�����V+I����?[�����$����Yp���Х&}q��;F�y* I0ߏ���d���Ǵw�.��c=�A����E��[�q=]CM�1K�A�߰����ʃ���Н׾�<]�:*�����a���J �	��'����y������9<(��FJ�6wK�����F?��]�S�-� �7X� 3F!�i��L�ݹt	#��w�''=PU����B��EK++�puH6PC�xL�km{\z�c��]/�#�]DY<3\g��gF���#���u����3?>�sEuZ����s��[[�E���Ԋ��0z�m�P��P��}��J������eX�������bԷY����,c���"Q}a	z�҈�1kB� r��M������A��� �6D Z��\�H�Uշ�04��?�ԦV�81�ʖ1of*�7S�M
t�fw.��_��)�el�mM������,�($j�	��Qƞ��ݭ��a��K��1A����kʘ�Z#�v�cd�WQ��O�"D���,
ʰ�BK(��&^m�f(�����v�c�/0v�����ۺ���g�ߑ̺�����|�7�09��]!��LPkOd�#j��D��	��A�*�/�9L�ǙX���A��/�3��)':�"g53�KKˏ-��F*�d����Ff��ؚkT�&��ֻh�D>��7����>��8���ȣ5[k�hyճ���6E� ��>�6(��ԑ犿�e��=5�3�9�����f���X�]IA���C0����_�@�A\����e-z	����/Q��� �|$����:��+W�i\ �uMok��k&E�=�7Q��ϋ5���`��i����~.��&��f�w����>�\E�Oz�z;�.�e&��V�j����oq��G5ѰWkz�cx��|v.�>��H��[�2O�ݽXk`-�*�� �֝�Nr1��!�'��?7(s�Gqk\��Is��CL{�1�x�a�Z���ZP�a�w�/���h�q��m��}qt���e�������j�`�p���+J�fDVm����p�n�	(�0�����ç��.b,ht.����7UPb��[�{Ṣ��䄺@�N}�-EJ������`�h�6�K�v�DV~~7��[�	@�ܤ !�+x���]�w���u�&K��@����ۅ��ۻ��8�r�@_��b�ȇ�	�i��nG(_mV�p@�߃��8���C��]Bc֔��%p��E�H��t%�_�e�AO��o�{N��P1�E/6iq�ߒȇ"�*��g��7&slQ}��R�#�� �E<�GHJ*�-�G�W�R��^G(?�C5~]CC_��1������+o.��u��6��ǀ�K{�����41�����:K$�X��M�� ����t������5&��d D�)��CA�P�����Ѧ1��8W����i�hU���ap�-�������|��]�or삂���W���v@��ywJ2�|�W�, �6����l������C�@h����c�n�����}���@��j�,����N'�)���{����Ԗ�Vj��
��<t$�Y��_��x������B���H@h���MQ����~���!�;��O�m���%��<_X�9�"�!F�zD?6��u4��S`�$F��F���(�fc����4�d�����h+�P�'EQ >���#�� ��A�P?�I��eU c�{.�.����#������B�^kq鴙��V�JKK[[.�B����S�l_3w{�1�ԉ�J!�P�t{�v_���0`ǨW=x{ep�1z�y�T������n?�����&h[�pXt] �h�I�$S�pKKK)<(['�{kO���/�)굹�-���";���d���2�~��~(#�3 �zP'�	h7�\\ 9�����ugT� >��Y̨�3��`҆lz��*2{
F�dU�ߛ��	�.���l�u��r��b��
@#��
����D�)����\k�H
��MF����u}hEjf�&�v�[�A�� ����E���0�=/'G�y��|��P�秈F���+M��s����ǏOe>��g�F{�� �e�F��(1��B-�|�\��!������!MU9��{{����������l�\7�|�+gaD�2ꐉT
�¥li'�<�2�6*�e	�-1��F�7N�ҁ ��qvg.B��J�aI�a%ǼX�1x;�m�7MF	�X$&ϝ;0-��6}p���!��X�q�-c�]/�؛���53��w�Y�T�h��s�\����U]@�:+���j�T�<�QM���9�����
��)m�j� ?�z�w	qR/�&��^���,��_�T��S�4�
�F!( ��6�9� �ޠ�@?��|2���P}��J$, �;/,�uV5��\�0�?qҭr�7�l�Rs�Jhf���n.U,���)����Iw������*M��������+uۛUc��
�����#�����_��Ä��Q����~���7*��p��%��7M��b���^�rJ..����H�������(�"�����ꘑ,-� p�U�f+�i2(WUs�����1f_��yxyM��&��Nr`:A$-��4j��a�Kp#�Z� n|e%p� x��8�{�s9jm*�s�!���7���y�H�q��HzUj��`�az�+�C���ZÄT6f�Ez�,��|�ׯfb1��.
C##/���@<�x�`Y�#µ$�$�_adc����ը�ӧ����j��lS�t�V��#�}46��ꦁ���3����(��E4���glчQ��%��IU!4mE�cS�[b�B;������%)�$wb���m.dT練IU�F��4�C�;Qxٞ��lm�(d���+��W,٣8�3�V-c�d@NqVT�^I��=��+F�x�|XlH�|�T�m���Kx���1��?�.xr��]@�*�$ IV{�r�3:�k�ϸ�~7�\5`!�_ -�z`����������S�&���O�F���+���c?wa\�m3!R�/����
jH6�ps�oxbD̀|��UUU��fz(F"#n��r/�N��!Cfac��>+����L�aG���/��U�a���Ч17r���(� �s�ږ?6h%���1)�?�1�U�WG)	+��+�����G�2��2q�[����m��
�1�q췿KQ�Ԍ#�s��~�� :� I�=�7���Y��2�7�.�9����d��p�7R��М�F��y��@�o\"�r7&�쓤��e9
���}������P�Wi��%����4�f�b;Hߵ	y�3� �Fh��GtF,����W�(v0��޹|:�z�}������188853��C�	!3��I��9@�y��;��IG�ST���[�����`%y�/Z,hZ��NM� ��~ q�s�u=�+�l��5 ?�9iiW���#hB���?tvuM���VQ��,<,<|jidBW�^�+�k���x%�*���Eg�3yB��9�]V��:+���䐆P�(L�ʻ�����ZTPD�i�fl����O��h\�pL ����{��ҁ�{�o�����e�Y;�3��L!�G���&_2�燆T�ˬ�`oN^jΡ�T��x��"�E��Ў�D@;��^���^�RK�TMD��àD��1o\		�b��ξ���h;���r^�Z	�D�A���I�L|}�
!nA���\��!ڛ�����[4��W� �K����A�L�n����m��<,]]]�#w�;;:,�1�@k�x��F��~�nD�Х�߷$�T�B��<ף��0@��k�g�*��+���M83��XF� �e#޸�w����JlZ靆�Zs�h<۹�Ś�R��HIؚ�(�5aɼ���%cE���!�U�%Y��h�{�p)[��B@ݰ�7�����jHH�S�B�c�%�4Hj��LN��Tf�7Œ���(=>�]b�c���zF�ӈ�E�3�Ä{*ʈ2t�-������H�4�z���Z�.W���ʰ�-Jo����&3�U�}�����%(�ă-�"��i�*́�\0�T����=EO_����8mF+&&��Ƽy-�|��.דQ�>tB�s"p����@4� �� ��c}�|zk}.��7~�r��VRQ��X]�����<h��Rmcn	���KK�K�*�1-c?7{0�*D�x�ҥ����]K�H��@7�@H$�/\G�	�ߛ������堼�?[@
?;$�Kz'�I�bCĪ���_�ҹ		����?@�9��q�D�B��Zً^bI��C��Z�����D�:NNX����y���0/fg���Q�����<��$2K6�y�Ə���N�����<~�?ʼ]���:A��mCx�|C(�S�/˙2�V	E��:�ќ�Z�L'@P:�u���)(�k���x� ��cn��!��&�UU����׫�S�R�/�{����'�k�Y� I�֙)ņ(0a8A�JH���a**#�ZY����$J���IEa�"Zx��XE[;���k� � �*���}3GV]����<�1��04[1J)�Oef��,*���EzffD�~jCb
�kN��/����u��� 4A&=|M"�!reW��59�a�:��hE[�3q�f�Yp��Q����������^SU�i���
m��b�DY	�2��8裷1h�֮�������H}���gO0�*�ٳ�PSR�;:���̱}��}��� ��`�;�\ �����wq��/ ,��^WW6PA-�,��O׉�R	;%�iv�
�4ik2a�<��k_x�I���EX�z���:z���+�ߒ��Ё��F�C�m�3jM7>uz�|������������|*�!�=0Ѩ�b�NOF�Fx�)�ٖs��[?T�U� x��Mc�/g\�'!�WOq鶕Z<�ScBL��
��vu4i��u��1�:Z��#�n]�e.��QҠs\��Sªe�0����G9`�3^đ�:���e;����%�To��c%�2�QR(�Ch�"�<��)�H�2��IHu��d�L�#!eH�B2d.Q���C��߿ǽO�:gkx׻�^{o��n~>��d ʮ��u�� �&�����`0����u6__�=B1�>��2\k����v�����p�@D:Gj�oŮ�گ��|(2�2��7߾=����'�"�e�A�I�K��@�Y�����`�qf�YY�Cʱ��i\~��&�_1o��Q�t������\��_����{䨪�<�QDx���ȿNnT ±L����6��?ξ��k�(:��^�j�Z�Z��H�~�9	�����9�~O $���}���š|7X��Fz����>'�yc�b>�)[�����]w����pt~�/��?�E��|��n]�n~QӏO&
�(w�C0<,Xq������\�"tk^9Gc��e]��{��B�/1�va���x�oh;�7L���ϯ�a�{qm=�3�Pm��`g�|� �2�8:�y��O��1��E�8�2���_s.����1�\ �~{�{������WRi-��;�O�� �*=,C/Ni;��j�y'��߽Gߜ�T�4X�� ����\��~����?ο�~~T�oq�o Xஞ?Z������l�-�]��Mk���6\�Yl���-�/`��¡��v"��z/�+���1^�u�!�r��	��3��(Zs��,�0�rL�=��-�j{��u6��y6Pd���f����$�g�C��J��>�+~�C~zE�i�w?�~��º�#G9o
(m	:�2=��ȥ��3����Ą��rS8��Eb�R�6��M/�_�_��і�Q���x�Q@�qq*+W��vÎ�1n�;#w�Uε���������r�^j��a�!�5��=З�dR�ҥQ��ĝ`��A
(���� ��I֊�.n�ԋt+r����[�XPH��+w� @��#~oU9�	���4���r=<,,�I�p����M��׿[_w��n�=�z��b��#u��#�m�_��f+/�	{.���ayG`mO�����&�e���U�M]����GTT0(m2���jd�H�,m=�R8��0�� ��|�9/�r�i��v��{��&#���a�^����c��=Ƶ�cƖ�%Me�l ��!�3e��5��SЊ���T�Q�\ �����Q��!��bCu��̻��¹�/l�����:���he2�2�x�7+�GQ,�����\��|ZȔ���_`���7���9�+�:r����ߖ�"�]����Q�yY����q##�OȽI+u�v~�6����G [�^x���X��p��-��m��{���z{<8�p��sO� ����������p����B1d, ��0�*@��ó_��f�@��4?�V�qz%IU͍���j�`oi94 &���D����RG��|1�X��.*�@/a1�m�D���eהk�$覴)����b^)[/�:���n��(�������#���
�Pz�Gutt4��6t��?���yS��&��2F���� ���ϟ?ҹI2��U���C*1�&?�/?��B_-n}t�-y9�,N+m���:Y��Zt�`��&x_Z�������P�U><\)���*������9B6<i���^XT��It�M�����`��G�_��{������s�]ʡ`��X�ƃ�ې��~6�6U���������v�����|b�tXm���h�6Mk뎴7i�e�1�_'s���������
�>^v!ݼ�av�!D�
H&�:?S��Ӄ4�OB�K��z�'H��]{����fF��+�Ph�z_�C�d]n2A�__��W�j{�h��8�"��r�o�����}A��3��Q��m�6l��7 �p�/��'�]�g�a�em���n���Y��{l��yI�0o�}��̸��&���o�kd�U�`����E�wYVF��b�g���싘��j�*߾�1�KdR�D0���e�_����:t��r*_��Ҽt���ކ,��o743���Դ�W����P��@���W��� L<��G�.�&'���	"�p(�?J0���@t�	d,�?��+Cr"|�a$�BƤ�8��ɚ�ˆ���p�ݗw��Y4jjk?{�����i�v��ޟ�x7y<�,�E�m�Y�O�6,�/y#˕=�Z���n�|�BB����.����ĉ�0Pp�-`6�:KB��7:�~<��ڟjQ������"}!�ئ�7T�5Y"���
	�M9�M扺 ^լaa�T��o8��M/،T��w���놆2�y'䖵��c&�,N&^��-W��M��*�q�+m|l`�u�ǏG�u��J066�����%d<��2;����nA�ϐ��ٔ�LF��#�ƪ�� ;��@,ܻ3�
��5x��K�`*�m�����4���32R�&|� W�t���܄D�6�g		���Y��#�4#�:]����lxvGv�����*��Pů�eN]j��/�~B�u(�����9�D�l6�khkG��jI[��x�L��f`]7�I.�����p~o�������6-��X>k�Һz/�8�YE�ӧ��c��4�͔2�<��]���ǚ�����~L4J��
�r�Hw�H���X[��q���T<�ܐ�Pfr|���(���{#cno�s��;&�n�wr�������*�z����N�AѵL;_�8�������Fr&o��Vsf�ǥ��_��ʲ��Ns���*�Bׅ�~]�/�tL�������d։���B�v�7AWrr�w�z�GeUՓ���@�jsv��p������l�H.�9j�j��t�=`����A�w �p�T�u��H6����p|����^z?���O�t�k_�Z*�:9��ɉ��5ww��9�ZL1�J;�
2�����艺o��z(��'_^� �p�4x�*������s~w��F�P��!�d:��G�M�����¯�]w�J��B01�����"1��&$�z�����6(�Ι~�S˛x4�(�������79�̴o��Pr�
��g�{�%�M��rĐ k/E�{�#\ggh�j�g�iQ7.��5��kn缩'@�|llL��`����"�@G�ɜW�Ź2���E&�MK�M��?��:�����A}�'~�;�I`��R������h;��{R���888t�?����^���ɱ�ɾ`�9jjiu���E,�������x|����rSM��Ǜ��k���e'K�P�L��y.�0^�U,P���j�U�����ɜ�Ef�N�v8+���n�[L��)+���p}�js�l�R�����C7zHQUՏS��)�����+B2�i��T$�� �=��UP���*��+
j-�Jz�v)�wl�������b��>�X��׮��ݵt�>�w}�a�9�5�)�1�eÆ}��K+ǆn�q���2��[2�&�#VC|۳�=t�Л���A����2j�j���6ۏ���]#�c�0)V�2|���Fp֔����,?'��ԏ����1ժ�~E5��Ɇ	��?�	4�2����}�`��T�|}}G��'�����(�'{!y���F��Z�j�,X O�O _��Eb���	Vk�D��8َ����1R���bd��e��w�T�ģ`XR������g�T�P�}$fQ��nk�@���j������h�		5�j��#���/�p���M<����Yk�yv��%R�n%�g���U���ޑ�����)��(���2|��]�T���T��ѭ��Ј��\B6䓊t�#1����[9!�c�&Mf���ڴ�IN��-<���t��󜤶J�l�xSW��u��k:t���V��F�K�n#1��߾}���s��#p��t��X�_��ű�~��:K��&.�S[�G�jq	���� p��T�v<������G]��k�l1�63��U�d��6^J�)&��b�הzQ?x�#���ֵ	Z {������3�f���D	II�H.J�K�5�?��*a^L=��!oN#7k	���M �p��,xeޒ�/N_�$�G3���iڴ����WQcc.n����������}�f���@��ޗ�'���{�]@��A��=���˛uɚ8�N�������K��`��|�B?�X,a�׸qe�-}��*��j�����)�	snY ����=�s���W�+�5c�P>4��[ׯ�r�W[]�{�#ŚF�����V,�8�[D*X��9H���ɡ�U�l�:�>���������������g��}ddd������
P���-x'�=	�`�CG���cV#������ݧA�:^ �e��`��K��5d�		)ӯ3<p�S�����g��;LZ��� Y]m6g�w�y��%���nZ�p�YCPx��� �����"��=�@&TƦ��G�eFD�{�y���Zy#���1��n4���=��Ku��F~�OƝ�9W�w��~qJ3-Z�î����/پ|�Y��	�Dq�����[�frVX��5��C�y��O���]����n_��v��]]]5<
&J��B^:���u��Z��$�L���|���{2N	�rh��ƲiP�R|a�"�����@ ��V�]��ȹ��R7:�?�a���ۛd}g|tT	�5��ԏՃ��ѵ�U����V$�g��`���4�
* V�y��3o������q�_B��whA�'<n��Ө��v��K&��#�*H,\M^��F���;{�g�$k��>\
�s㤢5�ߊ�5�{m����>��>�N�Ie9'��&��U)��E���#����3T��o��]Z��o�G��nDMH$.�9�?��i��2��\�p�H� ��y�y�*ס��5<�0�������1.��ц�@D�]�+�����6�����h��x>�F����O@Nl�Ui�4-X��3�^^�]�^GXL:�u���X)�4ɕ4��/|O)�O*H!���k�b��[#=��[H�}����emR~s���N�R���#���='w�.�'��4�w��D�����]"�����"y4>r(�k�����$��E\�		g�j���Y
������B����_��𥿽ie�WXX��yi=jB���Q�@����V	��9�� �l���0������'%���x��#��> ٳ�b�aӏ������u����8�<S-+��j������ey,�y|�k�f�!���\BB���`m���u��c�]- �C�ŧ(/]�x�cﬅ������-JR����a�=֗��j �;���Ѫ��n8�.u��ߥ�8TF�K]]B[��'���V��.���W��z+�}b�����B[���K��ן���KKK#.iij��^Y���P�5��OS�ֳ70��c	����ۮ`ۊ���Aaa��˱����{�V�M�5<s�A�z���_����t�O�������p)��;!<� V�P�<�'^?���%k��ȑ��uN��l	��V3����g�"�H��2Ӧ�6�U��C�?�v)�;�):R{6������X`\�4#���U&���&�8��s7Y��ϒ����Սq Nv�r	UF(�"6���h��>.[|�#��R7�b 0�K�ܼ���|1Xb��$99�y'/9��/xxP�~v���7��ߗ��_�!ر��� �^GȦ�/	�8'F@�7iD��h7����c����F�%V16��D?Ö:�ɇv��}��gz h!YYY�8�xr	��'Q��A0�81
���3�q��ڼ5ܷ^@��%��[�"�(^h �8W߹zI'=��d̩�$H�0����_p�ׯ_0l�7���m"��R��X�7xpX[Z"+��l��p���q����l��H��ƾ�Cy�쀛������27��wCI6��[��b$G;t�uyrŴ���&D��`��CDt��2���DF�_���`t� ��������IwVZ�QQ��u�^��AgXH�蛬�G�D�!w�n��������	��3����}��$���M��}����%��?K�0����w�Un��ԑ�.w�0�~<��̏�4��]	ET��cX���X`cҰ��(qXY9�v��#���g�%?#��� �a �n�÷����XƷ��� ��IE�MHa7����n<$-l�dݯ���/�:���DA���=����g;���Z�u��E&[���V'�8Sm�D˭�؁�`�NuC�������)���y;i��KǛmR(�6.�Z0Ȑ!���Ԕ�\Ν1�inum1b�Н� +w@S���~�`���С�����*f�o�_ ������ݳ�Ȃ9���<u�N�"�X�����'j�l�v� � D�3+��	��+H�(���kK�k'�Q<,�OS�&67FI3FJ��9�b	�|#~�Q���AT��e�B`�׀w��g���!�PH|������L]��뎬>˳v0w���.	���C��� |��0pi�b4\5߹���(hC;�RL�$'��9i���L���L�p�DP� 2�s'HK�gnB��Í㞆,���s�G����YDs�D�v<%Vq��+@;e��G�M鄼��""�\��g�X��=WX���i/^�H	ω�Cx��c�u=�:ܲ��q���h~O��m��XOJ_) r
[8�	ȰZ���_*lNe�jR`u����v���`���k���2Q.Cd01][[��U4S�p���X�h���i�w�$��t��UR�2�yP�#�l�F�r�yv g0��Y�mZ~b��j�����>��lf����F���j�C��2`N�[BU���G��.~�������5�D�E�ߗ�{�Ҭ�GJ���?���2�P��2	��{عO�29��J��K�.���r�+>y�R�&pA��Õ�h���o޼�O��
���ڪ�7m�'�����b5<��Q�}Q##��
��M��
�� E�X	�Nr���̑���&�y $S�����3�}<��˗�%GBw���ɂ!�K�����@���������'���7
�c[ed�pKi�ȏ}�;j���aR~���HC����i�Q4b~b�G�}+q�O��_]�S)�~�Y������֡7ϴb�jj�g���Ǔ��	�V������0� +�.H��s��0��l�J��<�;6Q����%n}L���~Uy��]�Њ�֛b�)>���.�7����V��j��$�22�$&��n��H��8@Ӵ�L]�hUjr��
6ρ/?�t������&�n�5!����m�c��_�׳��v=��߿���"�)���J�5iZlx%=}W�^J!)�
2M$}�M���E�+�����&dd� �0N��|��B��ӳ��,��/��iffV�C�Mț�:��:_�ĉG�E�%͢�C�g��ӗ%fER���p�3��G��Y��%���,�?Sx�"��`�f�փ?����ſM�CDV���`���0'Q�E�cz���㫿��T�hhh��i�.�K*���}M[������o;%����m��pVٸ���Q:70�¼Yl1����� ���g��c V�x��<o̴���i[��2B��C���Ϗz�V�$��OF��e�3�9w<	YS�=�2U����|�lJ=�y*�71�1~��72:��sr������ѩ�1t;��#s>���]�87���oV  w�!�+���(�f���Z�RF9xuﺶ�l^ o<p�ӑ�I`EK�qi��.7�,>E
��I�F!VB��{[��֋vE��d����5��x؁7:�.�x�0P7�Q��˗x�8�Ltٴ]���F�Oj�)E^�/�9׬Y�I���	�_���G���2���`R>~��~���y9��MC�3g���l6/�_�b��mp�	-#��}����OX�RQq�zb���?@��C�-P��4��:������iȬ ����M�r�[��b�-�F>4�%�@��&�v1�犾����Z>*������~�� X��=���)7�v���������n��o+�ș�^�Z_oM=qW���ǉ5�H�Uyt�-�IA�>�>B__�G}LK:5�̹M�! tOO_��ˌ=��eۻ����Eݥ
@��<��5�u��ub-�T	�B����x�=55<&
#�Rd1���
�i��JBN��0`[�͢^J.$]������(xCn��9�:̇�+D>i�ֵ�T)��y�Y{i:�y����ԅA/�V���I�K���d3�]}xs���C)�ׯ�|�soI�o }���� sC�+;�N�B�OO�� #������[@�h4��:����dރ�: }w�|�se �e��zhL���!���X�t�ҥm�� ��Ӭ���jj�D�����\^��Y~���L���Ԁ�H�8��ׄ�6 o�$i��Ջ��q�s����$9N6O���Ҷ�������������<����wG��ځ�� X޽6Z���Gÿ�|!�f�q���]Gbb�y��GU�4���Ŧȏ��wT|���~��� d��D�5A\�g��V�gu�����6��>%%%�E;33�Eܐ��?c��H{j�,�"c��ͧ��{鿅?�,>^KO/��4 ���S�!��].$��}&�KAwvԙF)ρ�K���Z<i��;�k��"4�����Aj9��X���k��sg��[�f�e=�O�EI�x��9#�x��F��۹��S���OLO�nkk��g�/���<�o`�D����Yk`�*⫴pה��~�Xё���ӬC�/�,;u/�� �gΗ������ƅ���%�&��a܄��@��w΁ �޽;\]S3&��x��A������MP+�o���:}�	 ��74�Lc��Ç�{a�sO�����i�����=��-W��t�}�(��!�ce%�37���\�WcX)�/��;26%-�4 >>P �T�rz�������x�!l�����Ss�˚��M_� �Ά0���Ξ?}� ��,6��i���U���NH���(�Wd�n��� �&iZh[��*�V�Ķ��ŋL��hoN�)	&#�2�k'Տ�7-���3K=>&���Ke��v��%�	�K:�[�bKEm�R���M���n�o�=����?>9�J��$�my�������iI�A������}e��
S��R�E�w�� �u����G}F9i�����"F6T��rhh(���wIH�� ����R��b�r�.�>S|��`�%�R(����݃37 �m[P	�ھ}W�'�z����P|{���F�OD�G ِ��HL�E�����p��8�$����Iv�)�3��H�,OǤ2����pIl����"a����C��N`\Dث�}}*`�M����;��׀�������������Íۍ����(I�!.G��hL	�`�QDI�m{G�Z$ԗ����9�ӴӦ>�����a�_k��R�@h`鎌��T�@�"0�������+^�)�潸Q�ބ!<OK_��d�]�O�N/y�h��O�t�O���ˊ}�K���q�΂��,"���=5#��k��U-���N���*GV~/���?s'sM�`ֱ��^���\�깐�׹�x50.�0Q~�3#�&���v�`:h7D@��Ǐ�.Z�$ X�0?�Y6���54.�i���V�^=gI�� �?}��|�x��*�w$&)y����=���###�E���v��<�v��6_E[����P�?AF�ٲ�a ���S��=HMo��E����]�B`A��f��u��=z��s�mii۟�F��T	<��1|���8;�XT�����HC���f�wgg�z�H��7,S�O?�^&�4�ge{�����/y�s��u��i�sg��^�L�#0�C#}�K �c�R~��e�"#�*����[��k�瀯!�R�A��Α�D`¨`C�7/�SE�|��W��(�����{&��<r���R9'}�����2-6�u�2�>\l�K���b#sY�� f�VF#^=o'�'H'�*�9��n�Ց���a�Ϸ?c�O�q��*�#S�������^F}���#h׺����K�g�P&CO�0�:r>�ii1qq%�Zb�����kJ3;uʲЇ|y% pPv<j:��
�f��m�ٗW�#X�a������ů��1m�SX��9̲9�Ep��*�]�:��<�Q'W��=7�pd$���;�DcHKK�	 VU|��sC�,�4T��Ĕy���P�X���f�Lu!���)y!��S��l���O��� �F� �� 	�Ωz8�����Ga��(
H��)��ɉ��4����E��T�Y�p���M�=�஌S�@k�v�'��̮�*�z����\�I�V��{a^��*�j�@qկ�<��U��<7��R��:	��%ȹf�Y����O�JH;p,���[G��r/t�?�Ek�|I	��S��ZSw4��'�{ׁg=��?��J����C��ҀSXO+�k��w��ie������0�u�%����OwW��$�2n�U与�Y�cl��KVU�­�}�����ѪT|�������E�����P�*X�dA�^�禔377ϖ�fX�>�~�L< T	*�!s��VP>.���jJ(��D�h*$ `ٍIj_���3�]��^YWW7w|'��v�B�)͗OF;������t kb�wn 1(-о��j|�����7�ֺ<��F�<�*�dFe2�GC蔊n���o\�(|z���0��L����I��wt�Da(���K���zD�~gC<�e���t�eй��C)%ϔkr;�e��`ֆ�'��O�fFm&E}��/�hg�p���[�<��,�����/$��0�xb����}9g𔨇�b��&�X�kC�r���n}S�ԿDLtai������kj����������RƘ��3�����9���P�}~���uS9Ӝ����h-c�(ط������
d>~���`�u^�6m:}�L�*�Ģ�;��3�����x�᠟��T�=>D_&�����jp�,0b�����ɏW��H$�&�<�/�j�6H?Hes|
qP�eͬsQ<4��9�R��K��;�j�#�����',��ڦO���(�ǎ��6]�k}
����]YYM�U���?6A��р�I��<
�]Fb�,���y�hO�q'����'/n���75����.�b��J�HB�a��8�}ۄFA����w�ϟ���N���9� v�]�1\�X��q�d���o{���|OO�±��S6? XM{��(U�3Ȁzěn÷�|Z� \Tf_��Aa��~��Ã`��Cŧ~���ߓv�2/��K��)�L�{��,!s��Y$�S�	j�1Ϟ�c��5��ꘄ�Ւ�Uߊ% �D�b�H�"}��#��A������� _�w���`ݾ�+�WlV9
#g[�0����O����ir��������s��s�!��0���yE����-C�8 Rn:,:S�
:���ӧO��|�x�1�}Hc�1�.վ �A!!�SChӁ�1��l�`o`0���RWD�ْ�>_,|a�q�=6�,&������D}N�(-qѵtk�|wA�����b��H\���Ш�u�m6��pnb��}�Ԥife�ڽ��G�z��-��t��b���ׯ��Ret$�#0�\�8�1I��z��PaZ�=̡Fό����x�YP@�	*�Z�{���P��|���|�w�ڋ����;�^rs�1/{*fq��u5V�
/b&#�c�=D�>&��2 4��(]p~�+Ȋ���K*k!X�,���A_a#B���޽{��ٽi�o,�Z!�y P�.lV�����d��ƅ����ץK/!��kP�4��-������E{v��$ǭ���t���h��\|��5~v�E�Ԟwj�K��K�����Y�VKHa�
kc�����C��P�/�����s��B�I��M��ÿt�ط*	��s�(���2NY���|r.wg��&Ar���s�IJ:�{���l�z���F�/4��<�y7s���ظ�S�>���TFc���? կ�B+Q
PzCZ$XN+p���_MuZ��`^FNN��Q��b�'��Y�yY��C��\��N�)���>�ym������;�T"ы�K�s��5�5��tp�D�/�X���N�\U���� ��a��@�ކ��[�</�\Tpr�Ԣ٫�F�%)�r" @�&ا@��s��=MMՄ�A�=v�׊���������}�����k�)�i�O�7|rjgq�k��@��R��&oo�̆:�˄�T�7����ƀ��c����]6w��-y���D��=x1|um��P��ġ��xf���	y���3u!���߂�0�z��ΰ��|J�w��4�'�ݕ� ��	��Ί��~2s��lć��
`��ҀI���<�|�_����&���\�|�1�K���)_�hx[��Y�V�*J���>��@��z�Cw[=�F����L��xtߑQ�����߿K s+��c߾��T�(���	n�~d�6��qL̡��x� �p��'�)���+_ZZ�UP��`_�(�$�Ű4��;\��2fyio�}�I	�������c��s�%�>�i޳kh�df�dfEu.8f���57�]G΁���U�1w����y�y�l<S76N,+S�a7ܜ�|h+�9=��x�O�8 FX �
�L��V�b<r�'q��)���>��^�"���� ��8���C'���O�뾸L+���QMh�����'��Sċ9�c1�l /�~����LPLLO@�W�]f�I���t��˗+���r�M3��=Q1l��:l;���` �X�2�A���3�#6��a��T�Wޫए�K�����;��-�o��� Г���p	<s(	UG�=�Ԣ�lܴ|A��u`����Kxf�ˬn)m��'�}��O/ߺm����k\�(�8��14�0`oh^����'��i
�>���z��B���w�p�pN�v�� �m<�>}���ns���#)�X�︊���=W�E�B�qW�Cc���L���N��;��|����lD�ٖ7X{g�	�IO�!1V56&�?��O�1�}������N�$]��r����:2~�������3�z%D?�B^'7:Y�k���� ��'b<��l��S�U#��q����@������EC��!#��C��'ΑU�*��ij�k�4�i=�8���bA��tڿJ�KZ��� ���MSȾ��9�H�RL�b	|����/���ȿf�^zo��]j[_�H�j����½]�q���N�'�2}�i6��c �rǁo�+)IU�׺Qp��3M_�k�y���̰�:v,���M-]ݧ�M�:�[�7:Q��!1�ͽ3� �½vVç�I����G%�����p���_�P>22R&��?��P|�)B82!���df�g�ͧ�Ok�%�~S�����)�|�����f�����>&�|Y[r�������C^������43sjǘm#���ϙƾ��OS��%9
 �⫪c4�����dUWV�_9�'���H�#�e���0':����y=��@IԦ+w���#�Ꜹ�FΛ;�����.~����� �VS]I���W�;S���591zo��7��J,���qjl��*E��9Q3ā�z�P�W��c��pU�L�x�=	嬬��!.$���X`V�����O�� u��)�z�\�#��E�@�1�GkZ�[tlG�, �<Р�M������]��ծ��Ճ�^���4��u�j%��
�z*sC�'����)=|c�!�]�~��%B��|�Y�zW��ĝq��p��[b}���EZ��˵����Wd���*c=cUF��w]�Lg��>~���<���MWel:	�`��S�l���`Π;w,���=q�)a� ������@X(7��#`�a��z����{��5�������t�]߯���+�q�c9�oii���,!1��7�
ֆϝ � ��RO Bifn�=l��x�ڢ�Qh'����6l��̭Ӛ=��G?�
�C
�s�����	Z�l|�������l�j�'0��K�cuM����;�Ұ��_iS4�cJ[��ǋhZ  j�U��d������M�0[q��TEO/75����XS�4��.R�gJ(DOo��������5��I��TjF4 l�ܹ�[��}�����k&-~��$�����I �)0�[�Np�Fn~^��G��_�~[X��\Fo�'y���{ϥ�T���թ���=�\֝��X�u���L��c��/k8Ԙo�$�tܽƉ��7k���ڞѬ�o�! ^�u������V�Q=��*�$����<<^999o��9��HAf);�����ʰ�&�3;pz���6ױ�"��x�.[f�ݯ��?0|l#�y��Ή1
!	��5]qn�iI�5�	��wc:��܆r�������D
��4,hd�5��%s�����l�5k�=z���Pw�	�ԛ�<Pq�5PM��Qs~8��H���&G��k=�V~��%k���Z�*jk�"""pN[8�b*��	��,/��t�p��Ȟ����p�5�uRΑ�$��� �1+L���(��}���W��i���;w.�40&%�R������V���/�x��T-��z4��}��W�h�`l�SO�Q�[j��}r���(GE�%K����⒒ѪBBk݆N�ʹH���AdR� �M�T�x2lm"�C�3�}b�yb�#�ի݊b��10"ҏl>y7ٜ��E��H,O�����~u�Z�5�<��,i)����5x�'�%������/��F«tAL�I��
.y`���-xuC�9����c���'��I�^�Y������z����w��?�c��,`�.�'�3t2{����Qk���p]� <5*㷆�?sVC$�w�^�����8��|����97{vvw{WTT覝�*�'!�XWKT4�L��eR7,=��/�X�f�*�	g��o�Y�8��r���-^-_'~|��tU�����h``��qWM���Fe*!�[*���}$�}j������|���S�gL���;�:B�DqH�_������Bϟ;�������Ñ�ݩ�X�/��_;q4%
S��̛���*���e�r�6���S*��Wnذ;|�������mt�Q%�$�f������[K�^������jM�8؍eY����	���sr�'��=�ÿ$;@%�!���]�}���t��v�n�H	�ft�-��ڧre�{d�Ђ7d(O�(V��Ek��c��ݴ·0�����7���@��������,��P���ɹ= �P�m��[���ÿڎih��.�;;6�!��8oi��tDޕ���]�%G��@؍��<�����*��o�!F�kǚ�����8l�OD���7tfzWӓ��&1w⢸�D��G}||�<�v���&��?9�CNN.�x^���������ud/x��r��&���N��:��t��.j;/��!s��IU8+feY)�-1�a�xkME}�j��Qѥ�{O�˭�wk���+g�\��O�t['�]����F���J���h�0���?_�U�] _
a�lr������v���G]Z���/�ǃt����m��&ɐ�����͠Q�
rs��<�P<]L���U��}h�|F��P
�+Dn�/�j�-�"?��(�����vq"w�;Rޱ�"����'Ё�}�~�Fy�OmY(��j��lrc����������I�u;��
�	G�
��FIػ�߾��V+Ry�!�j@=5=�]���]�V��<�!��D��HEc-K�m,s�0��fů�i��8�
&��߉��:���������ٺ�Ŵ��-�E���ƙ������W��d�+���8�_4m���<Ϙ�N�M�s����':��V�7��xr����C?�����y/8�o������Ԣ����@�bd'0�M���w�ΰ/^\���[�F�1tL{`�<	�C�-�`�R�'s~�#�������g��Ƿ�>79�[�;�>�Ym�R��%rw�[�~�N2R_�T�E���g�5���|IFfr L����^J�p�tG<����|�3�9:�}���u��Z���u�GF�ۀ�D/��| ��z�*��8�������|��h�&�D#�I��6���f�)��I���</�.�lE(-Zsi�v�!���iEc���{���@���� ���_o��^�y���+�d����r�W'ˆ�Z�[�b4b�� e�ޏWz9���HL���9�}Yפ{Wk�ހ"�Ы_oI�#����d�N��)��#$_[�Z�U?��i��1��,������ϯR��?���C-̟.m���%����x��s�T#fy4����kݸ���ϡ��bA����ɿ��&���֎T�C�n`�x�LQ�|= iM�?����/}n� �* �,������osfR�qп�5��Sq�I�GFG[�B�U�,K��q��	��L���L�Rt�<��0��.���J�po�QX�R}m��,D��L97��Q���|v�?6d2J� ��X=�r���d��5�t4��3�V�!h��X�SP�a!6���6�"Lf\B�.���n� ]|cq���o5���0
�iu����?�����A��<ΒK�½��	���\��+3!u�7����^0�-����s��A���߸��K��<�MYD=��@9�ļ>dz�3J�G�풓#1l.X~�p�p�~+�O�nW7�V���iI�2�	����$1+�WO���:3���-ɉ��ʐ�Ŭ (;[f$ɰ�gӯ¯�gct��5�t�̙�`Bc%�S��%��IXkc�>R��wf ��i�Mˣ���	��3-������6�d#��m�xӔ8�e���;,8�fz�.
�м2��9Mgr�^��n{�Gm�����?#k>�O�:X�ŻThsٌ�44-&TN5���?��孃@~pG��.���NL�����1�Y�qM~�m!��٘�ɷ�'��j���8�r:�X��N��-�m�8�6$te��*8�c��FAo�m����� ��0�6�XAw �?�?��؉���&�R�=�>h�cin�8	���>TU������9��C�2JvLq�t�m�BB��?���.���.�E�S������G�SI�0�L��o�1�?ZH엚^~P
�<���@�UZj*�@h�~��S�J.f"�^��Mw��N��5�����޸v�Z�?��@�o�8�5�8]�
@�N��2m.�Q�G��ZM�*�9%A��\ܐ�}d�1k���3�Xڡ�>(�R8[���%�	�u����V���:{�0�>�i~��a�;͙���������刍߶MM��@>�5H݂ �.t�"�����GsY �p�C.Ғ��t�^�M<�-�^�5.)����JD�"���|��
�[��L�3�m۫�*#�N6�	{'2==��^��2ߓIwILe7������y���`Fƴ�H��2*8:p�cF���Q�u�uLBB�Lt{o��8��F�X,�<s�L���bH�+*������~�.,X���}���OH��RQ ��U�s��)%��|�4E\�oC#Qm�k�;%�!օ����7�2�K�Ȉ.��6oR�M��8���Be J��dN}�FH<U������v[<}���^VB+��K��n��=߿�`�M�
�<��8�룋�ݳ�KXe���������*�Q��8u���kl����_/!V�yoA80*z�5�ʖKz��Y�g� q�hR=�����=�{cc��NvO�.�P��D�mZ�~�z��23�a�_�P�}�_2;����|�j7�#{&?d�>aaa�1�n���i�ijr-�8���!��;χ�ڐ��`�z��0Z�2A4���wV"Ȯ&N/����jz�$�
�L��&�M���眜������{bFL+�w�}���I��ro1(x���>�`��Q}��tEC���]�`dF�$(I�7�fJ�*Fjjj0�mF�R��*���zW�&4w%N7Tlkj
Q��Y�^���u}Dq�[���g9tDMk�-udd���ɽ��Aڂ'@+�b�t�F����ψ�l������қ\"�Tl�tT,�6�|�hu6Ǐ���; �@e�_��L���0X��zw�h��<�����+���M���c���] "�q�_H�de]ݪ���(�uK�O���.H9x�!��+�ٶz�� �F�������߿�  *FFn������ G��r����͞�?���l0+k٠B��X:-S�T��"|����D�=|�s�/v.;m.4���i8Ԉ�ݦhllL�hV�0���U����*�]ӟ*Z�Hջw�>�p9�������'����ʜ���b���9=0� @xA�ϟ� 5앥��sgZ�O����Q��d�{�R�VΛa$V��W���[b%�hق��B�W��9���iS�t�t�fP0õ'�"�;��A��z("��P�THj����7-`�T�ȝ�����-�M����߮�6w����/�K��8)1?&�˯US�<���\L��.�8�笀�r��g���}o�Vx�����!u�~�����L&�s!������h[�\�rl�Գ)0T	1{| ��>�aqέ��K����D���c���V}����!�!e���`�LN�.����w�]eZM��[j_�|���� ��@��ݻ�-]j�ċ��%o􊔼�n෯W==-{n{�L������*������/o����h C�TZ	tٴHX��J!��Ȣ�(d	�BNjZ�'''�6�웓�cim����677�ئ|�ĵ��7�OFc�>�Y�����8�t�>��D��<�Yjz�N���ģ�`�[!�E�K���>x��V����������@20��@�f��6��py^n��	���^��0�ǃ+0:\��o,\��ld�������t��.2�,-J"�#1�_��Ѳ���B�Y�ظ!zC�Y�B&���i��u�G%�\bH ?I.ÿp�̫%m��O}rA�qn�q��dkkH���00�6K:��_XЊ\~��[����n�;@Б`������o@+��s��n�A���&e�/����V��#���zմ���@}l'��K2ՀM��T�]h���O�N���d�v�a�" 
>�� <�M��]]^���0��ջl>5q.�r��-��-"B�q7����P#`����]�adOOߗ�S�&4�X�D?�����|M����>}�E�_FP��B�l8<�s���u ;��e�>q[�&����x�A=��"��í��o��ˡ�r�\Ļ|�s�mK���F0P�B��������bw�������mWˮ��7f?D�gF`X��*`��l�Rg���:x�D!�� nr��6�7�[�~���g����-y<�a3[0��n��>���Ba'k��e 	�.��\	����I c8���L��<g�i�b���zj2��́���2A�b�o��6NhR�޵?FDX̝��4-��)�MgO�?o�Ic���7���_��Jy����jժ�66��R�2N���v9�PyT"a.��k����\�����&�
�B�T2;�S���I�<ώS�Dʔ��$���n��3�e��3�w���������/g��s�^�Z�u?���¸�vsV��0]�jK�=�qp�p!�9�����\��$r����� ( a�{Q^��"�9J`Zg�WM1�UeeM
v��ia�Imu�A�� `�/
�X̢-�*�C9R2�>�2ӚW�-��r`3sss8��o�'���]B4Cv�^^�d
8~��OY�cT�)���y/� ����h��oݷ�>y�d/Á����J��-��X���MB�~�ԃ!����u�Rʏ�J[�d��OP����)���6�*�i:���|^�Ao�|�c�Y���ӎW�<�ry�-e�Hi	�ŔNH*6t��;���A I��>\�'��Lu�&�@^���-�����wu�u�I�a#W@-��34�wY�ms-.�6�nhbT�jaT!w�3�1�,IZJǡG��:�Z�v�a�Q��k;�I*�O#S�Xhw% ���4�CSwc�Xx�i��x(\���Ҳ�j��ȹ^1���
�5,,����w@�9���1�8�%!!KΥ��j�Fr
-q�%�����!�:�_�F�W��)Sdɢo�9�������e�e�s	|��W��k����,�� ��̀	d�$t}��5��]Gk�����D�x���|Ȉ#w+�'�!++�OmP��ò�%����16�\�Wu����R���S9����0��Z;(����y|ͪfa�Yp#���\˹~�$ƗqdM:zzy�ڄ��WS����7cjkϓ��Xr��� 3u����G}�Ʈ�Q��x��ִ�tͅ��=����l���~�@�Lk1U|����GC� <��.-=�e˂���?e``��(ר���]�lvB6ݼߕ�M����rճD�q��jvߑ��!�7��(��T������ݳ8+I����	qꍖ={�����ft���*�qqq�x1$���8��r��EY��+��`{��:�:�q��&^Im������7���-.,���@+z��������t�+[�J�$��a���'wRT�BU�x�:.·w�&�S>�Ҥ�˷��kt�Y��N1㗅�/*�����K���9�g�����\c��Q�eEL�����M�g/0L�#I @�B��!j�OIr�Ww�������M���N��^
�#����h������I7�/��|r��w�L�<A�*~~
�YB^�͐��/G]�6�^�b�l7��ހ��&k/��Vn���b�uh\m0��4D)eO����[��&o�hyww���Rn4e�UW��xU���x�w��ˑ�%!E�G�� 0�`h��Z��XA�A�".�N�Yʓ��k8�tB���餴�a�s/眡9 ^0~��w�_�6��3F7+S���zr?�)���⓾�l�<A\��ek��g��Ţ�����Fm�]��0V���+����ԥ�5������gl3����HW��;7��9�). ���/�E|�);�f��#WUU�_Us�^���H�E�i=�n޺�T�IyM�r�����[�eg3::�����I�㫸!��%ෟ�(���"\���P�,���bZcT'�Ny� 0�8����7����O����Ʌ�,5�(���!`��ٳȶ����&*	R���ױu66�=��q���%�]�aE��a ��7�Nn�~��l��^p�]滇�b\��R��Fݥa���m��\w'���$/�} /�H�1ta���ج�f��O^l�5�|�^l�YS�\ t����@�cR;�Aoˠ��T�:ʚ�1O����--O,�����q�C����ݔ�S����SP����"q����a����~�F����TUV�ƒ��o� [��i�[@Bnpὥ�]��2�����X&Ld)S����,��/�5jи�+���Sa��--���\��qǉh!?���C�D��C�Qv�r��7��{M�[����7����.��s�n�̱jԨh��?���Aު�7t��3&���w�#� P蔶G"��@� �a�v\����_�(��"ۦ��>7g��аPW`�U-�`�]ܖ�R��"OKؽ�yX�.���L�w��z�|���o)F������5��-5�EFզ?qq�f���<1������ |b&����GiC���W q���
q������Y:�~?nk���hB�235���4�EȺ����0.��o���`@�}��$��quu��y� u�d�P0lѩ���'�1;�*r{�ې��w{z»x6��J8�����B����(TmC�	+$���I�ס����� 5�a^o@4z������5333����yy�p�3�zAƅ����d͏?��&���O��3�Z�G�[�Y��k\�-��Zs�Z�N���,)'k�b�Rz�毄�dPu��ٓ�
�8�"bA��$��	�>�%��i'CC��C��ۉ��� �DA�^�elll�+4΢}���' xV]A��j$���b��)u��-4#
�%���^s���U���*�5�E�j�7��fh;#�Τ۵ ю�)��m�=K^���-�h،����(�j�}����-�B���k�T�\�y���^�~�ݘ�m�O��!���2V��G�#�����W�I�M�B�d�+��E�p�M�.���^W�3~��n��D��dj���?:
M�Țȼ��Pʰ4j���_^.C�ۈpxP5�(� ��f�f;��.�d��SVV-=�	>� �H�@��W�7��D��:�4;9�6�󤘘�<"֢�Z�#�"{�����	���f�\�HY!I����������y� �,dl��
�@7i/-�,W���?&��pp�Ɓ([ �-;�w���d烇X�`�e}����P.�6�$�����.BJ�CI��@࿦"�-$GV���5*K���͚l��ic��_8;5��D�~��D!�=kћr���O�Nۑ"\�����7�����GmB�w�G���P�^��*�(��,۷C��GE[$	,��i���Ve� 	0j;�r������5���``N�0� ႁ�<�Z����D�N�iB�p�%�R�^;;�Hy�[��'7�SfV�҇�yڨ�*!UNQ�y�Ĭ�3hܳ�ewvv�@�nyz�y��/�y, Yʏ�t��n��
�����@\^C�Ӌu?pB���ID!;����܍������b�h�3;�l},�����F��Ƃ�'����(����BhZD��A���D��ᖁ����^��A�w7��mも8GCk�Z�g�q�^PXD����Ӣ��,v�����G�!Qÿ�t+�zv �sݸ^BRtS��.B�H\��+�L8s��a%W)��I!O�0����$ ����=Z�E�u>���9ȢI�aq_lEhl,�e���l02)�}.쯿�"�\yBE���3�H��ʲ>n�0�a^(�ښ�h�̶�R<�1�v*�.�#E`�
�9'׋1Q�p� Ty+����Y���Ť?�Mc|��ڊs�Д�ɔ�ag!�S Ehs��� �	�����ؼ9"*�S������CD����m&�g��Ͱnjg�^����6���yӄ���ڹ�&]%}��O�HJP��W�������:��[��]�*��p�^��a��B��U��'=�k�^^KVڹz�L��>N�s�R�:$3-qf�a����ؚ����
l8��t��$�~�4n&x�̸����������;�HJn�d�����_�˫��O���653�DK��B�	y��͛n�PfoμW�1�d]�L�{������U�zzhi�b���|cpA��7�O-1 ���/υ�7~eQ�KJ�L��A.x/p*ـ��o�k:fAL�'�����d>az���_��
p�4&�L����׍�࠱��.��S]�A��J^6��P�]��4����~���YBY���˗!{B������A0�|k�<��Md��틻�!�i��	a2�[�����K��K��j�s�!�F�3yS�@�[:��y��9{ԯ��Bl��7멐�l3�B��_�>ыI��W[�j҅�F������,6���4i֕�oa�e�s��Z�����օ����ߵ^|RS��E��8�o=�ɵ�&�lVW_�%�SJ�����%�CVRJ�3�.a�j ����)�������	�� eO	����.[L�S,B�Z�9��>݃,�5����ӳ�F�lS�9�/����ޛ
�k`p����t��i�	~|�ۓ���(�J
/[Ԛ����P �<� �ŁB�DO9�U��׃«�Yy�{v�G�r?�K�ý!>��� [t�|���( �-"##�{�F�a�h/*a��Gi77�pj�o�/����Cv���>����������;����S�����k��D�����`��e�4x�y!��3�����Pг�v�_��D|$rr����4�ir�HS������;uOI$��'��č{N��g��v-ҷ�
���fgvJ�l��f;�t�G{�ns[y�:l��+�&�~Z���~�:�����ނ:��إ��D��"�wڜ\AcM�VT���o�� {tK�?ioH5$�p�����{K#�&�X�������fo 6�Á!�9�����t7���W=��+"�^�����p�1�����	e�[`�~!�5�߸'�vm�a��;Ӈ��Nn��#e͐�\ٺt�֨����_B�ۏ�>ccc���{���W���b�#AP9|����4�?����٥Pg��)�d s�g�"���v�>��M�o|�����/>>�v�"�8B|�Kym��*K
�j�)~�;L$�<:0e�󬰰���x{U1.,`^)&�����1�>Pboo�-y$������Ե� ��<���(���s~� tZ]�ABF�C_����O}d��,{!�\6�����!�]�^f5j�,:�������H0��"�wKE�,��wo=G0�����F�[��+/>F~9?B�PPP`�i��0�֭�?at6&&��޽{��D�� ���؃��F����|��w�D�����S�4���4s;��g�����_dU�:�1Vp����D�3r�/E>U6�<6ߪ>�!��a'�+�U���T�&� ����Y@@Ey9��0�|����� ?Sè�)�b�}2�6�"�o�q�b�~� ^Qm\q^0\������n�=��p����T�5MM����A����<<&�l�^[[�Lh	�o{wP9�`WIH	�`n��f��x?ga�`l7��c�!��+(��R�A<���Fq�Q�`pk���OL�n��r�x���uȫxf�جg�O֪�qH���l"IP!�ߐ��,�~�T'vAgvrH)^Kz��ا��HY\��Kb~
R�����O5��^B`����=�|)b��è�T������&�4?
���%,H����/E�����)y2+����x����D,u�3@^M�L^�0�=R�
�;
L���'���oH��Q�o�q�@�sI0�����n��r��&�	��@�0Q���4Y������xw��9�/R>b���3��_<�=��HoTl'�N[x9u�<#p������>Aj�N��_�S@��W���v���<�����D�^��
�1�_b�?���$텪�Rg��b�� ����!��=>�UңL�LO�Q���_6XEk3�J�V�����&&&�����oU��cV-N��cU�?�a0\�Gyno&�!o���czv˝�A4Z`s�Y��旇�ώE}ݯ�F'N?��K,�%I����Z�C?�qx��R6npݕO�F�W����?jѼ�
��8��e` ʄ�;�~$�dAU`���l��>�,P%м������׽W�S#�$���H[����羢@���|N`���`CJ��y������U��V��U�t[��y�c�pT�Ƥ��D,��غ�С$��Eqd �Ԗ�D\��޺�)��v�lllf��D��6��a�����VC�嫄K���v��X���3�Px�Y,H� �U��⩥3�@�i��"Yd i@D1���G��w =s��
ѣ{�]�jR?�J@r�]�Kl�U}��m(b�s|��XlG_p���駿Y��5�l��]�3���oZ��'�4:�@y�Pk�<��i=֓��xwŧq�����%�JĎ�Y��X��G���3�r��J��.��/ y��B2>Q���v���p
���:��S�_lH�οU�&��N��fVo`���n�ϫW�p},$|�tSiIUMM�Z�ɿ�����.]4
�.�;���+P�!L�A���B�C>"���R��h��q�P'�}[�	MR����Y�� ���>x)�Č��At��Kn!�q������5�G@����p|ρ\C�1����,���;�531�0C����p�0��fL)�8'%%e>Ф
=Z��#�^� �	�g-��T.�{�����d-�D�"�2 �lOY��"�0v�������d��h�]�iRn�9��k��\�&L�y�?���f
�\����ʪ���Uʹm�v����vN�<yY1oJ�v����-T�h�VJ��%h��ޞ�޴A�c"2��%7�+���ӊ����ۯ�=	�6)d��c��&��"�B�����#�T��ROT40�222����/{;˒��gjKn4�A���|�͠�M�Z�jk�qE�G���� 0��=y��jbLMM��^/���1�|6����!~RA��xG��Dnh
��(�@x�TZVSS2���[}rW����aFډ� �%�l^{�6EPI�F�'�H~؉�PJL���o�h���|�8	����sD�,� i�6gcc�)���P$�P��I�yMڹj�̧����|�f^J?9�sE9A���`�@O����o�>��yyx�b��b�7���m۶�o���f&��&p�U����O�O�4�)�@�����d3!�@@����4�t!��jT}���p6�
�Q���$
��OdC�F�`�e� �>?9"��)���
�7�yTP+ ��V����n} �G��Bŭ�1=Y֙`]����.,l�Y#h��s�QMooo�Tcmԥ�Lđ�6�al�Yq)�� �`^�P�?FR����^?�PZQ�Ѷ���}�.�rU�!S�o�,��|
dW}�em�����q��H����ʤ��V���
��y�" c�p������3\[b<d�2�A�ݾ�8M)����>���K25���-�+��,�;��؅����T�8cc�;?����~q8��\�x���Sȴ[�LZr=JB��.tv��ܔ�}���E|�S��H����f�ׅTVW����Z��[�6i!���ë��p�B��.���鯯/���j=z�����R6�w��Hun���\�=��X�
V�폌�.p�6�b��R���c��7LSi��	�dJ�Y�|�/>]��p���SD$ip�W��I=ڑ7Ԗ�vao9��q��dd8�1<<<�QRb��c�Dtt43y�Sٜ�;/d��9�@E"6f <���s��m�st��O�w�����	2��V.���� K�mO�7�56k��<����W��!Q\�E������L�w��	�����#�.�h�b��8�!>�'ۉ�Ɨ��n�����3 Ԏ� �@� g1s��\�>�>?�=/�n��-�z��'s�w��&]����R�I� Q{w:��@@b�X����i�jbe�tK𚇡֜�o��><��K�C�-89q>�x�c)v�������<�O��o(�H2�*B�:��hW�JG"z
�rqad˯���
��8��g����$�FGl8�h��R�$�F����y��ā<r�!�0 ?x�j�z a�o����@��c��F�<��OVS�#�%Z#�EPK�\L�t/V�����#���ő}�3�qf����C"O �	����5 �WJ�u�J���D@I���t�D��a��y�S�Ne{Ǿ��!нʴ���)�K�I��G9zo��W�-<�]�/yK7��{֋�)	>~vWȤ����Uk/q{77u�JjL�r w�L�06<i�@�Q.��K�Uf�_�t���+'��Sa8�e�\⃮z�]D��g5^�3�y�l��8�S]DǑN�6�t�@����^�k0c�3�i��#^������O��N4�X�R�f7��@��Px���VEA\#"�{lԧ -hP�UsM��l��mhr,p}���,��=�>�N���'9��(��$dV�ӫn�aV?��_װ��v�7�.4/$�����	�~R3~mV��UĎ��ԨUG���d�2ż��>,=]D���en���92�4�GP�����mO�۷?�E?ĂlSN�/zvLo�O}^S�zH-��8G�����Y4����q��.+6�0�_�h���
@���c���H�A�Y��!6���"��HM��&�~"�s
�� -j3�LԬ{�q˻����Ǯ�@�0\�Ϡ�����!ߛ'h�QAA���*�d� �F�#8+�y)���NN�o���� �I7h���Xz��V�Aќ���fͅ'}\�zյX��& �Z^�/vٺ
R�e��\����`�NT��zl;|�o�	��t����K'�7�S7
��ޜq��0�/���i2@لX�*� `c~S�M0(�K���x9`i��
`,��X�\]�>��Ԯ�����m@"}��F�JJ@
8�gq�1h%��?�(�ع"��i'�ֳ]�!�?�W;��%h���^t`� ��1�],�����qJ	r�����H�>_� ��<t���_��͋( '���y��=W�����!�m)�y!�y!Z@K���9���g�l�
�C�I�5j#F�9��q!pK����f�t�sF,PK<����]f��yr2s�Jf�U~����m�S�L��o�+j�=���d��ma�	��ܞB��B����z��^�%]PP��usyMӎ�%����vf��APǖ��s�|߂�C��x��=��t@O��:�kY��)L�0�x	���o�fpQ�����}.k�U���D(pg�THB�'4�T��-����� �q��6�w����)-V^�W"��|�1������x/C��	r4`�����^�\�wI̺���von�<���6"�	��ː^@f�N��`p�bQQ�UbM�f�#<W��,oNw����s�AF(~��p	��ϑ����;u�N��^�u% U#�|:]�A��m��!0'=~�U\\�5g�^�10��� O�k����P�^���1ș~�H���X4���Z��5۹n�*Uh��Y�e�c^�QJ���{��RǪ�M��F���WG+WTW_1e��I�������q+R5%�I�s�Y%V#ͅ��K���Grc���ZGr(@'2/�Б:�X\�[�����M���8�%DN� ������9��O�AD�W�*�j��vs�XWI���=ni2�,���������|��a�@䍍�����L\���<��J8�= �:r��@��?������3����1����z�������,[^GF�M��.��5�G��������v�k1�C/]���ZgkApiiF�����W�g$�<�K��8�E��X��\�t�~�Q��):0�8��'��H�~��#�]vX�S6�����\����/���逵��b�&^�sL���2��!4�cѢ'�h;0�^]����x�I2�cйZ�o��O�S�Ĭv��!V���m	�}0�g�����^�*�@f�A)"�~����X�6]]]��w��M:ρ6Y3)bi~��.�[�wcmt����E4@���qڝ[x��:!�NaA���_�*���3j�g]���r�*�a{���I%1s� �\~GL��c2�)� @��-5ʻH`P�qd�� 낂���E�L��}��W		𿙳�c9�UA/B����3຀`������A�+Wn��DFF�^VUm�?��	��U%%�����i���^ 
1Ԧ[܍�ٞ��@� �Ԭ������g���:ǂw�Y1����6y� ��5����]#x�~��A	��K-���P��t]}��t_�Ns��ρ�|�JV�0�D�����@�O������6��M�J�DP7��'�B�k�Q����Q��H �_�Q1�@GVU�;�ׁD���:	'�\�G�(�^�O9�~��D<	j^�|đ[�����j#0���U����ٌ�P�!0������eho�eHp���y�j����~C�Z�q�� @s /�7�.s�'k�kHOK����~{5��X�g?	�`�4~�� ,�']�l��q!(m��~꺪��g���<�����ׯϜ?_t7Z���
z7�Cڸ���d4멯/s���d��4k��	�֣˷;8������<�Ĳ��g>vg�;�:��a���2�.�=����#�˗3;��E�/\�|���
'� ��w&�QVq۔�j����Z����S�tQ�N���׎��y�3h�@\���d���v4�˃�n�]�߆�?s��Z��g�(��*��?��ϐ���7�oKA� ��Ѿ���#8�0~|Sf7[���,�~o���w,m�QCY��(E��g�����FG`J[c��4v�1m�5+U)tN(��|��֋�ڛ��P�����ձ���*'��h�<�Y�G��/�ߔ)�(�G��Wb�{����3�j�Ӵ�YRt$�aЗ���T5�h�$[�^�}���7�f�TY�eo#8�h��%.�K�t�9ٴR�1��x����z���9�a/��GM��3�9�؊���+�8�V/?#)Q�9"�S���D"��X~�t}���q<�C%*������(�f:������MOOo����6��/�T��JKKn";�m�Z�����3�t���~�J4n\�X>�	�!7���p�r��$.�L��u�k ]�VwP=p�'
!�������H�:9>�w=U���G�l|�I;�oY�&�^;�����ˍ���� ^��i�v���7��`0�l�XT��!@XD�f�8�m�0�Mu�x�ML�@uZ���Z��C8�Șiܯ���3jB��TM���b�V��I;�,�ö����L��c��uc3Z��%@�C�TL�
�P�Ĥ��<ΐU6��ĹҰ�H��{͗�!���\��љ���S8��r怣�Y�P=$
��7{V;�9B������ t����C��s=��~��&z*�l�p	�#��'Xv����^���'6cS�9@�Lk3���9V����<$&�n7Z&>�}��.B�0��W":r.�1���F��"՘;�FˤLȳS���h'�NՖ����>ק~��:#7��8�Y�|�#��؏'��S�C��n�3u�AYV�C�&��v/�N L���뛙ͺ��PjÅ���W�&�@"�O~��j<�~��s�)#����!/<7�6�@}��-����� �M� ��Y]W�,d���nc�:C��@s #s5�����M�M0�	ҳg�Q�PW����ꍌXs�[�v��L����e�3�������"�`����ٿ�ĥ���|�^KSU�7N�Z���5((�)����?�0��moWF��'?b������%��$n�q+�z����C<P���e�õ�����}��F�~)��
$<5�ŋ�O�91�+�jA ��~�Ձ��"�l���\���:d���Zl`/�����/������޳����@�+����\��`1�_�̄�pc}5�AC��爙�m���6���i��/cx��is�j}��ky���)	!�a-x�$ԋ��k>�z��%j��ުS:4�pB%k�� "!!aiuei:~�&LEeOG�ZX0��� ���_��@�<yb���G����!��&b��awf���X���܊S��S�b��KR��)� T�x"���dTF� �>b{�M����֡ͽ$R�E�H�k�q];<
$�	��e�/i��X�=�kq�^Zs�����_�3�-f3���m^뺝l ;@�/���~���w��xrvD�sy�ZG�;�&&& ![�{]ʇ�К1�	+�~�fD̘���藪�$����\�)��?��Q��5(j�K�!�n�i�p-���ˁ��ƥ�S#]n�S�<~��͎�v��
��¸����s�b����9}r����_#o��YV��/�=� @��b�K1��4Ϩ����aI2�.�ʄL���~�.p��9nj`~.���_`Y�`���^�a.v��YX޺0td�)�1\7N�	�~�5����0eO+Ld7{i�z�+�;�4.��"�e\T�ub�o��������)�=�ů��E���`�����9����p�}��@�sy�'�=���;]$f���f�(��|��)��T�
�_��m�#�v<�ي���aX���O�P&T�,?M�g��.8�n`�?{D���cf?��.��y��Pw���_�S�-���U�C�<��M3��؁��o&�S��l�\�������|��� 
P&�R�@���`xv��9�L�^�j��4��kl���X��'��tEFs��]W�dv#�ƒ�E����C�q
�>$��������y��.�[���s/�zJ����w?|	i�ܶ�G=T�/�~/hQG@��ʂG�ϞH�l����?
� uCX�C@>�����H8����mm�w~X���Q�	��o���f,G�փ�����8ÁgS��뮀�Re��!wʤ*U���U�d�'�~����q���(�<���7����g�j�[�N����NX��
�}�����t���z�M�6nz�f�|��2�x<�!�EKϨ���]\�ݵ����j�5\d`/@���Æ���A7Qkk3fPq6�f�C}�ϡ��B�/C�G��:����H�����yj>�\�������
�f��C�,qf���P=N�^)?��@1SPy,k����i��CJ)��:]�	�}��%I�aLS�nZyU2�^c��k�/���}��������J�P���t�_�{���\mv�]���K�rgY����(��R��H{X|g��2�N�K@jXW���XI�	n,�n��������zf_>u^�}bN3�G����J�����20���O��l!����ƃt7ˊntww���xƐ3���{..2���V������^��W~i��1*�����?~\.c�ӌ����}<�8H�Edd����w:�1�}��ܾ��#�bﱟ��EB� n��%�bTC|��Ѣ�}nf"��]��+��8'������fև�K���U�pch$d^�UD�>q%i"���P�����}��pHto��C��\�/�鯫n�w�Z11��JTN�|�uc�#u��/.E>��ˢ�����a�!p4��#�4p8�e��l3�Ɍ',LOO{�S��ٗ�\�y�\f���]��x�Uz��+t�z����)1j��Цd2�\���i��v cπ�w�Y��"�J����
7�М.hλ����|���DϖP�����������#��� 0`�'+I�?����1?���nsQ�l�[�W3��y� ��߸q�l��#}�$(ˎqMʶm���R�������Y�mR�vp�ioN���}9����ǫW�~����p�8��ˡ�=\#�3����Ƈ����Kԓ����2ǉ��:ũ�N��}�xN�ߜ�V�l�q6��5��Ά�U���]$>8�����s��mLa6e������ 
�����)�۳g����c�aX�9٬pvv�3�)�mk㵩����{�Q&-���LK�g�ka�3 δ��R#��BT��T�o�b���4���@��-�_�1E�g����w-��;��9jZ�N�F��e>l�b�?�Vw���f}�9 ��=�Q��3ý���Y��+&^��F'7���|K��\	���Z>ˠ�*άn{�����CY�ǻk�|�o��2���R�_B����E`t���w������]�O� ���]�d��+�W�pZ�3�I���#d�������W�0� �^��ō
�z£3���b�������K��0�[��w���}�����W��:��7���8�5#�3�n���GO8e�X�ۍiǶ�P���#'N�H�ԖPn� =����0$����o���Ϝ��>�#���\%�"�<���T��׊	%�7�������T�UWo-**
_��� �1333�a����Qn2��GC����X)�;w�|��EԶ�<�^����ge�����b��<����<��ێ�'QWF�5뭌�̓�߄GEFU���V7t���1����a�UR�Qז��͎'���b?,$�d�8�hǈ' =~���[��5�J1�)?R��,@�+�"�UMS�ה:�Gj�O�x��|�n��x�i"�O��b����n2?�=,*�b�f�}�]0�3���f�r*�Ң�30��LO.�����������:�t��OF�=����8���s[�v�/8?_] ��ҙ�hl�<#Z]YɄŵ�
iii�x��� ����?�)f}Wz�D�^a�*2uNtn�b蛦�w�20E�DU�N����-x�Nî�����N�lV�b����啨S��qP$�r�gZ�������� ��/��il��n2:1��׊�>��[{"BA8���l<l�aVVV����[���Ш�����y����	�A�@1��Q�M�RF� ��J�6<_�zv5����	��E���~� ��@��P[�,(8	�U��	���Err��N��i��R0w������ˊmQ���|�ÿ��u���se��©ٍUY��MȔ\�j�,2q��z������O�C=��m'g;��K����]Ij��S<9]��Σs�*:�h��/��H]��N��v�P���ÍKH����R'����9�Jo�8a֫Py+����J�(^R?��g��Km���=D]��i�wK�����=��BMx�iݺuq��'�}�w,$��2>*{|�o�n*+��y!𾿿?��^3�>�t�F��N����t�q���K��oH��ܸ\�0@�Qg�?��E�盪[=҅{VX\�'��)[�I�[c����r����]�^?4T�l���-����>��L�Х��c��:��J�ˤ[Uo�z���w&�rܘ۾�i��ֲB��"JlL�������t��GT�z�.`!���x��I�m�9�wRn�ō��QWN�����L�޽y��A*����q�n��VT��C�\h��f�!b��'��!r�"mGݨ��7;��3�:ϯF��
��d�a,�$PĂ�{�F�7�O�RMt���渭�[F��y��VP~xf�	 ��{St�u.�ݼy���z��v<)p��QZnE�7� ����A;�����eJ�=z0%���8�����������cc=���9�Y~��]��@�����{w��IWq�ؖ���y����H>�	��	���ު(̊W����Xu�u��?oK�@�Jʚ�9 �w0���W��ek(�}㼼�Zx�3�s�n���_ܷ��w����ϟ�X�K�������U�`a�S{H&�''|�_I<|H=K��իxH�E	���Snge�%��g�]���R�;���K�Q˴N=z&*l��w����׵��B����f;5�O�x^0��]ӫ����oRX~lY
���p��Q��'Oᰜ�@~c���G�wv ��9k�D��@�>	�K#<4�A�C@���-<��q(R֎�#NM����2J�����fx�4�-�Hr�����S.��T3Ѯ�y���K�>�zeB�&�g"��0�	lO�=z��)MM̓J��$������^�O��o����2aݺ�1��?[��Uu����C�%P���p�����G�3�B1e�?0�a^^� 0����o=�J�Zu��ƻ��H=Dp[խ1�6���\\����}i��J�g~܃?�p���s�#�2g=Z���� ,�q��@����BɒkVPٽ�!�J%z�K����ȴ�
{/wR飝���?����w����]��*W����U���w����]��V�8_�V�����A����׎$�OLW����ΩǤ��4�+�61P��������$�_j��K_��@�ܕ��-ZMG������w��+�]���
y���!\����+�]��
W�������w��?Vh���@zL_����=a��pqպ�߈"��M�-��IwB~�����G�p�o]߉�)}���1i��� PK   vOXS��lG  bG  /   images/52445b69-20cf-48af-a05a-7b7247ebe25e.png @ΈPNG

   IHDR   d   k   ��'�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  F�IDATx��}t\յ�7}F�wɲ�&�r��b:L~J��	�nBI!�jNB�7c�iƸ�ؖ��bY��:��{�{GI#K2������Z���{�ٽ�}��#HӜ������ZH׉tM�+�.F�|> �b�C�&N���wC��1i�{nn�Yiq���%����0�u��}؞wT>��~/PT���C(�3!��o<�˃�N���y�t{��4�ލ����m��j5򽖾o�q��G��V^�q�Ke%�O��o.��:D�f������.�P?�!D:]7��S��}^B�\�Cǐȥ�Խ�<#�o?uj�b�X��݅�[��\�Y��EQ�DbZ^<���Ӌ�=.�.���C���U����wF��d����Gtz�P��q���l��	S��#0^d��i����6]��J���;�0�	$�f��~}����qc<&ڄ��P$ǘ`�k�au��ъ�+\�:B�^;r �����f�����}�O�����2tڑ���?���``1��` ��LŘ�a'}_��@i}Z�<X��>f�|:��p���O����M�x��?���Bc�b�����1��E�E��M��G�F�0���'����������*Wn���L�Ӈ�r��nL8I�̘V�O�%R��u$�._��D[~&���/��Ĳ9I�5���%��PDX�4/�J���xG=�ф�ǉ'S7W��&�D��w��q�������t��X<��iH�ŚM�x�hk����Ex���1Ak�Ƹ1�Xq�X�~*/}Q��_-���RZ4̈7���*|���j�@]�tx��M�!�E��``�xl��T����'��gb{Q'z�%��:&��e]8�cq�	c���3q�O{�����``ҝC��@ݝMW�t|���kl&�8<���N~�<O]��6T��O��8s!%�"n��$�+���wiQ����=��x����1=�ݿ�5="a��Ӈ�=v�q�r`c5mQ�I]�~`w>�	��:�I��Xkd����������l��)s�j0;݊���0�ˣE�Հ������&��e��Ÿ���'�4�n�F�+g2$L����t-eɸ��qx����{�Z�-~1��&I��"���z�KN�$t#7�M�X��*�}ͩ����Xt�T��')>RQ�(8�"^�;}���سs��3jd��w��N�����Y���x��_��1��3��T&��C��U�:z<)܅s#k��h�G�*�5�d�z�l��Z<�^	K�R(�_���	2��[}$��K£�Lťe��V/�pxtL�Nb����A�4�d�����ɤ�����C/�`��<|��9Xx�fR^q7���Z�:+y�����h�ݍ�$�_jډ��� �V�'"��l&ô���`\�_�@1�ӣS�A��vꦎ 
�+��^���"B>�e)���G<xg�\Tu��]��u��}d;��O�;�H��x�7�q��%p�m�ES�܈^p{���*q�`���6E{Bb��:��1"��0���z�W>~�|��x<���9A�4q���K�GpkͰ�� >��e���|�m�ํh"���Z�ѦH
9�.���p3���z\G02���8��in�k��bNr����Y̤��i��z��o`�-_���7�c��V����֓t�sd]��c�兙��4X��6��^MsP�H���:_M���"
�i�M��7y�0�{܆m�z���ɝmq����X�R^��L�^_��6����jH�5��}"kz%�{T��!�iy6~��>��at�� �eu�/
ѻ;�ĵ 5���cnp��pjpU��_9��}:��E������7�q�ɗ������L�e4�$&�r�K��\�kɵ}fm	$�IO����B�u���aQݡ���O�N��GoN���a�e�{M4kFR��ߏ��)XqR*�z���M5�)�
`b���W6;QQ�˦w��"�(e�v��Nߝ}�+�����{0F�F'1/1�j��Lz�.�킄b<K���c�4x
#�3AN#k�i�ш!qܛ_�+�:�C�˻�Ƈ��)Q����A���'���DRH��B�_����S��U�`[-Ο���>(	xʧ�� ��$Y ?="U�m>�ˋ��'Oh(�%��-��w�)�_�,�0L�n�渟��Uw}O(���#��y����y�w ����?at� �fNM�������Anf��j�kOc�䰌���&;��:�٣�1F��],~��j��@�w�#x��@�c��I�����j�����H�� �����/܆h�SN�a��Z��~$��qcv����X��_\�V_"*=Y�tG"�#���N3�8!���.�bZ�ZR)��FG��<�R��|�on,��c�~"����{7�	&���n $B�C�=����[���/\ǒ�Ev�C��͌c�5���qQ�W��.V��A0�~�!���0Mfu��Έap睏Q��5�Vu�҄#L$�M���A�r�����pE�S�^�k�lb;.�Ҋ�P�z,��w�8R�šq�N;�&���������"���k�7��na0��.���l&�߆�#^9��ኴ��H2feA���V��sg::���"�U81��5�9N`��uDR����vrd�8f\3��j�c�H�4Ԥ���&5��턀n��7%a$��t%�K�������K�f5@�M���	���0�Mj#�cC�⤇jZHh��|L�2��Y�����[�I��'4��$e<��	v)�FeU5Z[��II�;w.�Ƀ�'�^\������!�~��Sb%�Kސ`�i��!�إ�;�VhM�|S%�)���1����p�����~H!�8<}�"Q3���_7�A#���6�)2E��B�NoS`w��I��sN����Ln���S��j����S���ظq��uẙz<�+Q��C�����6`J���Mͨ����8���N���O��_�q��V�u���<L��F���y�:�A`�N�EA�HZNH��'����͸fb�4�{����Ѻ�6+�����I���ݎ�w݅�zh���2��8�G��$V)v#�"#)0���ө�@�1�n��چ��v�.�2
!!!�����u�Ȍ����I���݁��"P�d�6"��.,H�&	�� RQVV&�0����+�y���Lr�a�n9Ig�%�r3�Z�!2"��̀b<�zRAkL�E�nf�ٹ����]�ӈ��m����͸����k����Kڑo�˘�.�aX�>�b����;h�or����I�}��i�	�"���c���]�N%�؈��v#1̃o�QYY���pA�ͦd<��EQ�P~@�z/~�ى�F� �:���WLH3�&.����:Vav�����3;��*T���1Q�a�5�`����&R_���s>yX�����C�㞻����]a�*G�\0�v�C��f�3���Py��m��;����V8}������{[�ˀ瞼	���=x�=F�a����1���E���g�>Ԗ�[�`��G�hk��!'�!�jkk��Œb�jE*�(��Ո��Fhh�,������.	�BȐgǐ�k���"���6����'���A��:ȳ�A& hƀ���:\V6��:'f4�h��K̺���4ć��H����w�z$B�<�{���ꝍтk�����^fU�Cح&�z}9*�q�=�U�A"�Id�JQfU���4E������߮G�-{(�����K�u���jWM4�M���(=��\#k$�Z�������#ˏD&�Ν;a4���saN%�ȫ��=��ZZ�PSTG*��8�.��_�����c�X���vW��X sg�[1Q`�SW���m���^@��b"���U`f|�-V�M��^"�A�M����asi��y"��]6�[{�pO��Z�ʋ(�9'�� �[�+��KDJ=E�"O��Оb
�w��jN�ɸ-#�x�@Ϫ��ǈM�3���\<�a	�ɵ��eJ�N��0,]����hnnFMMM���ں��n�zE�4d���O]����>�}����2?q�3KZJJ��FV���Tv�<�R&���EV[���5�XvW��� ��9
���I]�IxY�8��ɹ���a�h��'�3�{��U<U�6x�p&.!sp�8dV}࠶n�{6��˖⣢�X>����<p�A组l
g3q��N����i�|q��V=^:<�\���<��Q�EP�`�p�݄Ө�Ʉ��d�����`����33��j���@Lt$�*��a�W�_�'��3����PM��ʌ|�*�KL`��6�ӦM���.�(i5;�C00,��K�C�\�U�w��)yB�Gˌ�ᢐ�ӟ�%\M%55�?��0�~T���1KqǅY8�m�sM@J����iO#n|� ^�u6�}F���N,C�E��B<����&�gx ��1<P��53�N��43߱r�\g��wք��:��Y�t��~Ւ����ӧ�=hjj�����]eX���L�Ĉf�G'">>111��v��!v�����y�+{�����k��r񃻱����9�g�g��aZb���ۧ��S�Sa%#΄h���AQ6�L:��q���q�WUA	"�nX�I)�.���_ߔ�>܅t}!f&6#!�!�cB���v�P��ݍ�M���2�=��j+�YU�Q�@�j3a��H\��Jq�^$�;#�/F*����L$�۫,BH� �T@�'�͊@N����;��OV{===�*9��Aa4:H��EA01�İ}t�\��|���lߟ�9	U��zj��ٮr���c¾�8T�'�K�⊓�q�syx����%�cD���+�������������]�h,��ʚ�Wc����Yix��1�6&�Z�?�)���961����8dF:� Î��&���ꊉ��ew�������5�Lbw�������I5�%�vx=���Ӱ
�]��}��$EK��1��F+߾Y��k��Ł�)X�m>:Z����R�ԡGBB�Z6/JBaU'������!	�;0=p�H;�ܾ��J���d�fSl��J�:1�^5H�����:\�x*��!�=�6�ãPX?t
� �K��7���Z`!ubиeI4&:�f�G�L�Q�g���~I�~�b��̸{c*~;�#v^�� :2��#���PX]:�v J�Y>��l��q
�j��A.��4�=���|��c���">*�`�Id�U'!&vD<�]܊+ۍ��؅��$� g��$���A��M��H�6#9�$���iu�ᶡ������+)��p�L��(��݁��-h �R����a$2��ܞ������#�W���tiAY��+ñ�6T��0��~?�j��_�cQz�D�i�.�³Pa��p�	ߔ����|�4��o�c�XLHEG�[ZPΌGYQoŽ/��7
�oAz�t?/[׷9P�hCW�C�83��ة�cDM�~��.O��������ש���R*٭%θ�$��_L��TM�	�FD���;����%C.������t�2�޻���SE񦤱��j��\�ÿ-��KGꎧ�d�Q����5'�N��+�#��\DD��0�s)ح��W+�7ե�$�T����Fŏƨ�H[?��z�Q;#��U�%J yZnvv�<��f��g���/+`#	�����f�d��w��9!�M�i�Q��t## �D�(�z�*#"�4�MO�g��'>:�g�ѹpa2��I�۫N@t��=�>)-S\�ÖA{	�KT�^��7oY���p�T�-�D^�E'e�b�k�QQf���V�o�,���\b�޺2u�����]G�A�?� CÃ���[J�Q���s�ղ�S�>^�3�̕j�{��CfN^ I���Gq��K;����xsS6�m21�&aq����k����C6a��N�K4g)�Q!�K-��Z^�җ'�Ɗ��xG�:%]lL`�����.�G��7�iyA���:�,���KJ��h���_�g�#��(knb8^V� ��Y�$3��E�	)a8��L�/���]���Tl��?VS$� ���Չ3g�I59���r�_�Ҋ9Y���ؖ�*[�����U�,���K��ޥglO���~���vm�W��C�S%)�7.�3�������mw̵_����{�i��eɟ\{�cFS�3�"���'�޺lN�\�����6,���֕)�E(b���둓j��q���k���LI���щYdK���`N�l8��w�?��	}�V<
&
s�4v��j���2�������`�Œf`���!��y�}�o#&܈坸�ɽ�I�]���w�Z���o9?[��Ug����e�<��j<��4LN�1
j�bGXJ��9p�EI7����m�<O�v�Ɛ�{¸H���P�1�������mX�a+�1Y����#B`�2��M���`cB�w�p9$�� ���
AXU�@�U��(1�L�]Bz��נ�ڎ;߬���� ;Ʉ��]�Y҃�x#�:1N���n���Mp9�-MV��_�y�����:e���������5��z�`z��8�ⶹq�����]sd���M�ߺ��ʍ����&\K���2������R�s�ɘ�b�ׇ:1%݌�X#^���O���������h��o�Q������F�Wo����YN�@ijF8VQ�gז�b䵓 �A�@�u�9r��Bm��o=������Jcq�f��<k�������������h�2�&Fa�}&Oy�ǣǀ���Ա!�?>ݤ�On�-hw��$~<���|��J����?�v1��Z'�olb������z�+,z"B-�?R(���O�(��F�������zL�p$-eܔg��:�!�(��5_U���M8gnr��p��w�V�]�[��O��+n�	B�{��p���X����I��	ab�{�
���գ�g���$�s��߶�$�X���pG$a劙��3���*��;<�� �W�3D�=�դ� �Di$��O���#i���?AH��#��6�}���@'�T����n��0�����k�$6�s=������P�Bj�� j(�i$-P"�w��^-$~2��(R`�+}���Q���|�F�����%���O�.ý$��Q����Y��]x��P�����#G^۪e��;d��mPr��x�V��(�~�WO��^��+��Q��ꭱ�1[��[�� �vW�Wr�˅YO�,���ipN�s	k�Q��i�j�����<>����W�x5�?�w��%��1��������_d��!l��j�Kr�l�����)�����!v�$����D�h����`Nj=���t�F�S��ӿ{���R˕��j�U74{��w>��e®�$I>r�,-��bZek����HՈVv�VtF��-zP��FsϊnU��*p�}�'X����HSCcz07�a�K=`@f���u�0:�x^��+�\���.�Y�7i혛� [�V.��h�.?�ې8B�̡ɝ7��&�AxT"��,AS]���Y�H����0=)J��kBzB�}z�Zp�`�l����6r��W.4�rr>I��ȡ�>C�c��k������e�'�ޅxGV�����D������@ȣ��dJ[c	�ǎd���&5�c��Q^^�5o�[W$"]�Q�H�5b��d���+����y^�QdG��/R2r�Jס][Q��{$`2)�{�ݍșu��]���C���O>�G;"����(�z�����?���X�������Ά�a�:�ځ�D��f:���CH+�;I�]�R��WĬlra�o��� U.��5 ��k�p.��si�Ɉ�����hn�v�ⴋ~p�$H_�d��Q��Fc�`%��	��6,!q*-��P�q����G�El2�뾃h��F�����䨱΍	�����β|	Z\����a�X]y<ny���=�*^4�Y2�$�n��q	'?�}j�kx�1��^�U�+c���1v�}q�z�V���P��:��E�cdyoo�>q�<j�����od}�b����A��ڰ��P���]:�^�݈������w��ۑ�3�^�����/�4�Zes�F�#��ȾG���rv�O�2�|��O}v`쓟�g�#|����΅�,�:]/�z�gG�X��#}��*A/��l|��x.<'�1�Pj:�����������/�Swn�N�G�x�?w �����.(هm��G�7��Ӄ�Ic��6�]�H�ԣ�ņec�B�ŷ�}
��6.r�I`����3��z5 ܶ�k�eB1n\Q��YY6RbC���BVx#�Ԣ�� ZZ����;B�m���������2r��|��A�v����l�cL�~X8�)�>9\�x?J�k�jmF\�x�+͆֠,�z��X�sM��W_����&�\�J#&����/+�`Su$�$�3(R��C�φ�:sR
lJ���i�Vz���Eqq�!�$�I`����=�6�߾@u�5�'��U~B ��i2���[#�jwd���\�2�Z
�(�%��X�n���Ip���`� p8(�k�1M����m��u�M�đ�4V���V�#xq�t�"}�����,	n�ꠘ�G%�6%%Y�y�q� >��4Ԛfp	!��r"�j��}�m�C?T7�v�2�u� ����ק�>:���m1�Xm�p�f��7����PY �ޟy��8�2Խ^:�C����	lCڐaS�t�C�n|�|�Y,����#{�5J�hp�$4JZ�$�d��DR~��6��B{0.�=�JI��q���{���rQ[+�Z&�J`�U�4�.�d�]j;�b29BϿ�Hj�H�ezb������\�#*��G�aS<�-6$�X峓w��6m�#���+ANL�$6����1B�4֯g���ؤ�$�ޭ�`�ybL{\���L�*n��r��+������ɡX���6U/X�*����6̘-�ws������Q�:&RR��|_P���7U�L�iv��;K�iVn�t��aiz%n��d,�MCJ�I��C��c�*��x��L+��=`��O��̱�����d	A�ZQA��ح���,Y���<$$���k�`����}�������U�����b"��fn�hV�\0rߕ����lttt���	0;at5���{wt�Է8൵���������7��4�ɉ�8uF6�yt�{�	�V��k^)�럮�zm�[��ywVLa��U��ݝ�ǵ�6j	a_~Y'"C0G�`RIG�T#�LR���;Gp��<�V1��X���aX{�<��QU�=��c�⺾��'hٷ�WcH~��'K �Y�^K���f������!51ƛ�}�z���V���ꪫ�f�bǜ%�HzC�!��#��	ߔn��X�ǃq�ODb�L%��x����*�׋��>����sU�ɹqG*jga����������,����?-��Ӊ�N�X͝}[#m�&b�Y����e'�T�[=�{r�{���l�P>sy����>��ᓔ��.�G�����z�E���݁��6IH6&��,�>|;.b!.�2�	�\6_�m�c9L-Θ/�1�g�h���L@}���E������k&�gO����w@ؐ� �Ӛ�lH�ie���& 1��}��I_�Z�`�R`�jÚ���5���n��c�+5?\�m�a������{:v�	Y�N!���8t�d��s5A�sظ�y���N2�mrtQ�E�.��ו�qx\by�i����=���l��NL��?� �ٸ�+r˲K1>�U�
�6k�=�:6��*�����FRD������h���Mr{��H*۽&��V*k��P�0@ko���q�WA�ؾ�E�����T ��e~��6���o#"�O��%禓�z����^��~�ٰMѨ�K��B>8}��W
��)� ޞ��ǥ0���ά�����jm�##���x�*:�g#���j
��w���1�d �?9���`g}��P��rK&�(��2~ߘJA��_�{�|��^%����׌g�C�S0�D~����`����P��R���5Y���"�r�uo[#����5�Dg��$�)˚.�o&F�I/D�~�ф��w�&���:�!E{X�w�Ӹ�bCy&�h]H�x�М����!�׎~��12T�8���>���<5v���b*4H�3�z�����O1�C9P��%�L�m�������I�<}�NP*����a��WS��E��iDe�M�`.L�Kj�M5x�\���5-69^{�9c%��8'V&���f��7$e�jc�Ks
0;�󫰷E��k��32ˑ;Ń=u�x=�`���ks�j�H����Oh�q���N�A�Z��r�'iW��K\�l���I=&���'>�/��eH��F1��}B佘���:9M���Ͳ��	xmc���at/������Ζ٠�I��!�$��A@�?ҎD��x�����0���i�,�D������mv���}��}85��F���(��LfN��������[0A�'K� ���%)����D�� �Uu����l�ݳԶ�\�ۢ�=?��h�6IB��ϛ�(�o٥�*��w�k!�Q�QD`<���|26�B�0|�Ȭ�(��������"U|�Pv_1����!��|]S4�ґuꖚT�h�"��q�a=>����ltN����3���ݰ�I���6V��D�1a]j���X��C�/������ѱN��\�b�9Y���4\:�i�(x�xZ�!��uX�ćGq�x���r��[�u	sU8�P����G�Ǜ��Ɨ��p�ꃰ�[1��s0>%L���J�=�D�3g'���)6f�p9&���pl�����X�ֈ����]���\pf�yn�Q̛n����}��~H/��%"+.�TD�x��x��j��V^
���4yP`�Ryy�>P�O�Ցg�����$��0T������I(&�2=3ߒL�U���1b�l�b���K�5������:Qc��]���t9�����H���}����.��G���!5�U;�Q���&ҿ����]i,!�h,-���.�*K#mf��*L��������ڪ�㊖ Q�_2m.ÐՋ�&�⿿�Ĳ�I�B�a#�4�\���|��#趺%0L�4���ZIZȑ�M���Q'�+&$�����h��Dq������p��:Z�0gtm^�$�&�[��Ǝ(tهX� �tػ�k�d��a�+(<��O���ƒ��()�d<������>�cd���ru_�R|�[�������$|N��x\�O��=��=D=i�p�D2V���\d��j�kH��!5�:��E�`IF=��k�7�Z�O@$0<���3��\��gHm:�R�ID	�~g�p�F�Kq::ݫ�����"b\A����?!T�37v8���
Dǘ�r�X�8Ϫ�u"��0����s�PA1���7^��)�@?���VA>9��/+3`l�#b�+���"!S���=3z�E�ƈ�b�`k�J!C��Iѷ�7xN�j���ZBh��f��6�+���)��/Z��K�`���)r�z��g98H��ȝ�"#�dw�%u�5x�e��1���ۦ{�~��Wv#��Mj��V�HQ��0��8c�T�U�?�z��u�␑5�W�Yàk٘��7plL�v��w��pK,�57��8�p�0��)n�TY��=����'��p2΅�)�#}���_��pJ�
pz$����9�yָ(4�s/�4C��?]>I�M/����*��WOƆ���!G�կ���pˠ��\�0kJuh+s��GR�*�KjX����^B��^�LWrG�Y|�sr�N�ڰ��opI+o��]��Z�d����d�ڭ!���Z��ְ���\V'�[	��~J�!B,��ɹ�%W���w[�سpѢd�V$�Z�"<G�����R�8+;��.�Q����%{���%XBn����$�?pF\��1š'|�����[�b[�j3���m坑r����fc�#�bGaK��n!�'�����1B ��o{��>��<I�����R�/�^��#�ҷ�\`��7�����܆���&�E�(���r$w��Gd���?������j��("�%��iDnN������z���	�p��.��}N�$�B'66)T�L��SS{~s�y负#'E<��A�|�&l�NGiu.8�;<Cq�f�ŝߝ��i��IZ��tn�h�d�!ܬŁ��cc��5�qBR�,φ�F!.a,�k�Q��ug��#o���g$�blz<r�MGWG�Z���pV���{���8!��#���&>ŀ�U^�}��<���^�-��c[�"���m�N�k�T�`�r����ad#�8T�%�n?�&ےFꏝ��VL�=ƛD�Q��_�.��&9ڌ77Vȁ`MV�:"�=f������"��o|s��ɞA�n�aO�c5����y��1m�Yh^����B�E�U;�������S����P[U�﷾-���GI�a	�"���GE��(\*6��|4��΃��^�]ݯN�?ڮ�����k_U)�9���y�$��}��Q{|�*6�U50@D�&]~F ǁK�U��!�'l3�޲H"qn���������3E�^�րmfí��s�'�V�p��[&������Z��X����gގ}��A�4�S�%���Jav�������"���iz��!%E�!�_��o�|7�[�t�~n�[U.>�Y]c\9�om?d�&�����{ć���V\�!�!�������^�HҤ�w�<�������U���u�p�Y�q�p��/���m��v$n��ٴ?xl^c5��.jԻ�J����wlg�moB�1̀�g|���["ʥ���-��_���z:�w�Ą�_���!��[)=�rT�TTN����/U#��*'iUXd?��g�K�u�������3=��I�#���vY)��AR��e���T)�^�H�@�1����/��}g.҄�S�$-�n��F�Sg'J������|�k���#�s�����+{��r�[/��p�Fm��t�%K�%?ƹ3>�4������͵?�(L�1�^sj,���7���4v�{l�&{��$�j�{�����$	��!bJ�1�p��7KDzٌ�Z�}�J�G�U^�.oF�{2.҈�)�}�=N��܅���,lE�`� ����I1G����W��F`kA+>���Z1��I���ϭ-��r>����kT�q2�p��
(���Xj�V]2z��'E�M���dF��	�xS�;񓓞�eH�틼&\qr��X�p<�^	�:!w\����Ӊ�vmp������}���I����l���l�ۄN���N���8@�����1#�����N��C�B%�9onfeE"�(��.aw���O�S��܏Q��w�3��V������9C�/��s�&����#wF�|���_�8R}��~���
nYBϘS�v���0��4��l���1B>��Kk9��:h�+B~C���د��orD�F���(����C&ne��Gq�\Rg\ƓO>^u�Gv3��
�qX��N|,	ɉ�����e�cl9�|��$	*�8��M2
J���t���#��\���ʰ|~���ņ��n��$��%�X�~���ii+/�(Ǉ�n�%�ݴ�����S���wʛf8㻈D�W	� &<z7/�B�����Ie)9x���9IѦ�;s����O �d�[T�-pq- �P��&`Zf�cU����%#l�2�f�hr�Hpc�9�#�~no/x}!�q��}�ɹ�]dȿ9�&�˓[!�+�<���s-VZ�l�C;�,R=���r8(S�&����{^+P$���Ѫ���+5UX��'�����f�#�6�[Y`R/+c�WVNv+Q���_׊ڽ��b1�lk@cKϰ���q�4;��će���w��]�dӡV�/c۝���5|`
(znƌ�FL��1Vy����D�w����*��Q���릓�^���z�+��X��s�9ż��ב >Ⱦ�Ɔ��	��k�8u8����x�D���4=0�ň���0��̈PTiUg�����,����/eč�I͘�\�Vow'<Q��G�	��OM ���������%V��y}��>�T�`Ѵ�\��Y�Y��Ͻ����HR��������f)��w'"�q�X{4���JX��M�s1!V\=%�_�*�y��謱e�Y���r$�8a!�އK&aiz��}�V�h{^Ο�*��@���Sk��)�|	�+��p	���Ԡϥ�t�\�`-��=e��2�O�]��ʥ;W�`^r�r���WD2Ax�k�bhpfV)Ρ�_{H2.z�ps�����G�hVtV�܇�[9��Μ4�XNG_6�P��"��X&J����' 9���=�>b�/���%iՒ��[ތ��ѳ?%�2��9�I�5�sat���[�ϣ��
��s��\�ksJ_j��`���M����xo����^�\�q�O���h�1�5<W�!��_sxro.����~1��rm.�����듹F����Bƣ��N�1�d��2�z��p�'���sO�s|�U������G�1�(q�c6����bp�M���y$S�Ŭ�9��A�fTb<!�J�������WQ_�������3x���]�)BLF긘V���׫��`�W=.�v��C���DB�9��/�1R�4����o�4�U6��u�ߢw_��z�q�N8���8)HӨ������1=>�k�����4����Icg�v�'��T���K����%��ɣqW�\��+�~Ng0.�/;���3&��A����2|F���u�iʷ�
<G�(>��99�K8ܥL��0����L�'���QGf��j>������LR�2���I/���'Wt8�?ջ�Y"Hum��^F������	�J���Y�aB:��_�8_���n���+_|���	��<^�k��Nύ#IN&@H��qz�	�}~�Oܷ*Yݶ|�I���>X����v����&��N����`���$Daͭ��/�㹫���0�Fb��N�9���#�a\�Z���ϝq�@�qiP�d�C8������
WT�A���ʹ������K�tB���:㣹BX��He��JQ�5�bk�5n���-L�-"[p�~_�/���w�3������V�y+;V��fV?��~����{-xL~����
���)�'�q��sU�1��V�p�<�ң�J0o%驤�	4T[�s���ArZ��c�J<'��1�4������ٻ�WJ�#���n�85�S�8f\�4�KWL?A�����I�mu�^v��~��o��J���3wm�J����D�N��M���CV���T'}F�'αE���Hϳ]�j|I�6��"����}��|"�Hܦ�G�D�a����zS�_�J�$v>֓�4�́��s
����7
rt����'s�$O�J�jB���_fb��*����kΓz�P������},��+G[I6�=�
.���<���w���I���."u�e�l�Hd��_@\�!��VR?��R�|�9%Ld�쿈t3�Cv�Nz��&�Mg��B��%�p?�@n7W����ɵe]Έ���l��������CD��~��>�����2#;�ؗ�/�=�l���v�����0���@/ќy�,�1�J��g�n���f�γ��ø`�ȹ(4f	��Q���=�<�{�w���e��ǐZ�S���bZ�iG��X.����u0�n�B�fC�q���i"�Y�
I�r�X`Y�]s�B�Ș�!J�A�'���$/��x?]�s�?��	�I�V��[�S�S�$R�1�$~�d��q��	)�:/j�=�`��N*���$�-a_��2z&���fr��^���}p_ג����D��&��4�������<����ܗ���LFN�x	���`�B���ag�`\�6z�q�q�$�]HZ.Z5g�6��GD�H����4ϕp���ߴ�VY��2s?%��J��J���iV�jA���}���>�@��
��<�K&3QL$)?�G��í�9���}�Mx��Tq�XD���Ҙ�����:���D[	���(�`�<�����r���`!���ר��:_z&���ϵC�S���޹��9�����	Es��`��aԫ��]�_�ϩL�8�i�^��!�#���Ջ]�8lsU7{�#�L����r�)s��z�<������~��,��T��B�Q@}1��[b=�����#G��J���\`Ԑ�2���~�z��9u�����7��ڐ6B$s7hUUG�sPb�7A���N!�]`vZ�B��5�[��� .��7vcǒ�c)d�TFse�jo�T<��|�`d�{:y]�ꙿ|NKƗ䱺{��>��?��o�/N�>/'�xE<٥���R<�}4���p���4x�V�<A��;�Q� �X6n<Y� 	<Qz�s�����I�|fn�0&ĐsU�y3������O�7Wf�'�p�u�qf;�1�7�ƛ��Z	�W(�
�y�Ag�"U�<׾��Vv�^-s已�(?��QJ�C�=p`��7���%�4��B��&���������S�>&����*f��(�ԟU�n�|3Z����������gn�\���w��e���!]v0T����ҙ�`t��c"�ҿ��S���=#�ɳʚG�Î���TOc��1��D�r|Sߚ�:75��S+ނ� �����
��.��e簺��ۃ��>e�.�h��Z��C~C�s4��	�~�D�$��{C�v��3��z<#��O�d���#�(��٬�Ug��ŵeX���c"�z}�Ȏ׀B�0�^��yq��i^��5�=�?5�̈�o!<܈�%cGQ.Y��?�V����45k���5�C�K�]qJ:����S�xŴ��&ﾽ���G��iq���gK�e%���m]��4B�*����}@�
/�_B�z�b�NJ
{lB�y�P�8�{Ax���W��0M�Ŝ�Q�I��q� ^lb",̍�e�y�w43.V^<V�ay��h��XS�-Ei���h#����݂ 9ӫ�K��G�Z�~YB����^)�2V^��ux������[0%#\��w��un^��+~���>+I�o�f�������-�朏����������{�o�p����Z� �:�IJi����������τ7�<y����XOލ���1�>O�Y�0�מK��Ŕ�0ٟ��:ٯ�ˣ�2����������6�Q�jR?s�Gc��F�'A�t��
>@��)1h�rJ߬)6
x�.����8=#h,��}/n?]���?�G�a]��u��^d���%+y����'a�&���67H2�J�Պ�D���&"���=r�Y^Y���w��𤻹 !+9D�����C�+�C��*��F΍_|ɛL?[_��~>�i~�^��յ�I�������΋���o���������\9I���BG�f'�~�i�CQSu�/���_�od�-��6�C�'�_���s~�z!Mtͦj<pU��8����͵�9<���L�ͳc{A�T�%U���rǭ��?����CO6��s�1i�Ao��C�:H���t��2��#�d���m46�6�f�I%
3���⹲*llw�+���7h��cޅ|Ѣ��I��O?
�C���P<�u�?���M?�Ͳ���N���u>]'я��}�0*&̠���5�~���ۉ�բ�����p�;7\�õG�w[~J�3Qݞ�q-KRAY'�1������k�1Fy�9B����E�yFyOJ��["*6ؚ�1Ǥy3S�zY��1��S6.�]���~s4����;)4/;���c�X|�:�Ds������.�����9 �K�    IEND�B`�PK   vOXإl˨6 �= /   images/734bc482-36f4-48b6-9076-7f88fee16b3e.png�z�W[M�u�B�"Ŋ�ŭX��Sܭ+��x�R��k�"!@p�w$wwr�{�����dB�ZÜ����w���I��ٳgx�
2�Ϟ��"_�Xϑ�|�yk��m$U%�=�M��3�@���E����3���J�s�%�KzY}i7+s[g':m[G�g���	q��������ҸT}���QQFR�'k��e"�+� �����ӳ��,F꬚�,��Ʌ�#�hIି}��b�z�EK
�DP������b�A�P��n�����m���:eW�ν �>j�Y�>����F����"���0�Bh��'��KL��w����ۅ�7@" �]�����d�dr�!Q�/�Zp�;+��6�͐���ú�t#�ENR��90f'Xo�H:N(d"?�φXs�u���y� RB��.��i^�&�/*:�g` ��@�7����q��X>��i$��4�~��VH1���J6L[<�w��bH|l�����W>��#������:;>"g��_�%��wq�s�7�"6��&<�����w.I���"}���M�׶vΨ ��Mx1�F���lEf�h�59\Α-c�_x}�����A��$5�5��w?�oj��"6N��_�@�o��5�o��/(���`�Qo\m�:]��{�|I�(��M�r�s{��;O������
�	��&�'6�-�}�.(t(7R'-��F\T!�8�62<	���}]I	KW=�c�WM��pE�7��߽:��H.�k�;�u ������6Pn�3
�~x��� �S�Ťvl�)睝A,�ԟs�$l�ӔJ���#�����^�߸����Ň_&n�ܰ�g���e.S�3����)��w� �އ���Z�˃E�y�r��C��c��a�C��Hޡ�,#��m����DY��bdbSN�h�����`��{G�@v J}���5������^Y�f!͔�����M;T�,C��itu�<~�҃���8��;sp�y6jӖ=�'�͋������E�"�ע��/�~�t԰����K�}U�a�x��'ǲ�.��+v�=
K�{�wTA���y	���"ȧ�'�(�}F2��i(Ac�V7��Ѩ��ӗQg�*���+ZlF�'�m6�g5�����±#J9L�����,�!���#���ߎ�V�߯�u���#E�O8n� N�	4�_"��z0w��,�E���^{�C���K�SJ�þ�[�hTN֮�O	�������D�1�i8� _�j��}�ˑ�]�٪�8�۶�LR�{�<��x�����Q6;=�G�/��t�u)O��|�]�uK��9~�ps6��]*�" %���������`IYF�Ed��:"2���e�ܳ�}��x�{bJ�3��~�|.
V��6E	��A��F��x#�^" Λ�0�򸨃��5�&�z�LGz�:�הi}��P���Kj��*ٴ0Ǳ߲Jd���{w�K'J�/��0�
�8��d�F<�xX�%�&�:��i��_09�C�����H����
x���>|�sj��(�pN��V��T��BQ5�}��{{���_w��'Q9��:iu8�m����H�
�_�泐!��wj� ��?>"����&�k?�^�{�q�ήQ�k��ؗ��q��>5A0�p=����d��`ݔ�Maۚ��c��)���xҫ��T�6��V�]v����v9*�¢�B�h�S�U�I(7E��a��	�i�v�$�hp�Ĳx����z�|\��q�D`��p��:����c\�Ө7�%ٹ�b(����|8gFh-��W�����dA�^�D�O�ФS3#5l�p�y% ��>Y�N�\n'v]L:�zo0F��F��a�MFƑ3��<�_X|Ll~e+�:}m���t��Rc�����DP�� ���0?���'���'�����J]�셿iU��1�j���^�w�I�?�ޞ��k�̥�\>�N&�ʚY�Zqsz��
^�a۸uM��	^y�}�����K�:�4�Z�J����x#�a�{@�wV����U�1��P����T{����n:�2�׺oU�]G�pf�]be��6��Fʾœ�;�����L�����	�������Z]���J?iڻVˁ,+
�)�"\��/���xŨ�l�aע>	fZsr�
r��B/z ����k����MQ�s&%,6 �;�
*�F�lǷŞ����C*�pr�2�z��i���z�����ƈ0��|�7��Z�6���j"��:�v�1!���멚��	
`�_��i���y�@
m8>�M��d��`M��uL��̨+���$(dq�Q�|���J^���(7x�����3OϮ�{khK6D5d��̱�zU�Q<�<h���)����k�"���V¼d���jh��I�k��o�65�Ww��tť�Y�^�9K,���Χ=��J���AL������50m�~�����l����� Hm1j�S/�[(��S�?1��#��5��gr��ۋZ�}kA���՞ 3ׯ�����@f�I��E�����&����[�VB�(��A��qR�[��L<�Å��	�NNy�|�p�GJ.����D]��Z��U����#�ǪfᎺ���9�yV�cg�'�@�M���֖՗�Pc��.���Neޔ��sl_���$(���݅��bs���W�M_�S� w��:3�\�f̽���0�Sj���ME�J��|
��a�r�㱹�UNbgO}�()9���翠��d�QJW�"�5�2��,Xl2P�'1-��d5�&T$OXQtT�w[�d�T3�{���� uTֆ-_�	ؠ�'��4/ֆ���u�o��h8ؖ��yQ�x���L��!բ��j�4�9�V���m����c�6����7�ዔ��zGyɯ����He�"��v�f�y���r/��V�}��l�r�n��ͭ=��H�0@�j��*E�A�Z�k���-�s�6��"̓d�8<f"�����W� 2�T5�Es!e\PW�+8�"�w�;U�Q��oqyC�#����Z��D��Ѱ*ܫ~gmə���!V�g),��DN�F�/m98aǅ�np~s;��h���/B�.��'&��cT�C@�=~gR�D���1�90��^�T��gɚ*˼<��=�ё���B3h|�$�7�0Ba?�h�� p>(w�;�嘃�uRS�}[
o'ܼɐE�MF2�1�'�����2�Bo��/�?ֈ8����e� ��Z�}��B;U����\�4����R�JV��:�3���4������+�| ;�)�Lƕ���٭����`�n�DTj��i���]퀅��*�P�$"b�W�[k�2>��6�b���u���f�I%�.�Ȫ�5�p����=dQ+���7��Ww#�ijdd4�2�𻁰& x)6b�bG;d�-[L��MI�X�������o/�Enk�:�����Y���?���$�	��X<^��'TX��]��.T�[΁���zA�C%#�*ĺd=�{x$~D ���ҟ��Dܮ��c������;�"#������{hm�4���]��1�)8@�x���V���6e�V�KmDӌ`|<���>��2��Xzw� �K-��5���#-s��\�(����F������F�Ƭ������.G�֋��?QF1�Zi0i;v��|�|�
���tN2=P[L�ݿ�#/�3��5�/�iJt����G3�Ԉ/h�ݯ�W3j�����=k�v!gq��!R����V�#���	c����E��J��Z��l7�f7H�I��� ���� �x��\���~�>#Nv�pi���aS��/hA{�l\aW�#������������� p�\�V]J�Q���� ��F;G|��H$Ha�e�t�#H�Jj���6��җ9j�}�8aʭx����cp����lT#�Y�_R�_
���8~Q͒�6�/�H������h8~�*�k��WH)&��\�[-Q��5��=29��l�%����m҉�6w�-p|��]R98�nR�x��6Us��й$�Z��Z�(:m�ʙ�����Tg&����G�ru�%�L�;;�5#�ݎǉ�Д����ۥ�&���6�d��>x�����I���y�3o<��4{_p�]���<
V��u�B����L#�\ĕԐ�g��\C-_��P���u\�S�)�JR��D�Oλ�`C;�}w���D/���&
-�@d<$� Z�;4bY�®��y������.Z����$]Ԩ���{>>K��Y�Mƹ}�?ޝ�"�u�81�_j�*^�}k�O����\ؼ1��tŝ�|s���G7�K�w�|�=�4i��+���ʾ�ޖ<R��E�gG�x{}���\����X�N��W��A�U�!T��gu䲢l��`Z�"I�q�|l��iU��b){�QxH�s��Ԋݦ���U��_���Ey��Eo�~��b�Y�y;2d��G�,FFtb��Ӟm�/��yImEh�Kp8IXa�*��Jz�W��e�{�޶'����8b�4����J2��O"�GX)�B>"��J����8��_�(�S��ң��y�\�Oq�˥)�3��P��3fd�X�
�MιTl�K��T�;s7���I*��g���[!OV>	�����X2��x�o��>�K+M޲��R�C�����W��]�I�XA��J�;BCH���-_��dѓЫ0��x�Q�F��O�F&G��	��k���8�Ϲ�|E�\�[������`��9��f����a�Ͽ �1R�; ,:���B��Ff����rOՅ��"Y�rv�F�3`�g��ӎ�o�{��� �T��*���H;P�~��w�Y@.eKj����IͲ4X5��$X��ݴ*90��x�,�,�]��]9ѹaj��1I�<� ~��z8��:���q��f*�j�$Xy�uV���m!�iH|)�#��hIY�Q��'��ɘ�N��XL��X�c��8���o{��Z���}���;�}�Dn6~u
�W3Gq+�I��|8����$�l�����-�tx}+�t:m�R����)	�����)�>��/2�<�����b�OKw@�#rH�r �� ~�erA:����vڷ���b���b�k��W��o�������\q�*o�����'?�3��*&�0�����wq\�\񇌐h����yzb�m�gn�Xn�/,�xt��sdyM�6����ʃk/�;\a�$M�#�ϫ{?#S�?�ܪV�JX�6��{c�_��1�3U�m��/3����"��F3��t����P�i�c��錫�ϱm�Y奍��#�
��&�(L�eS8��ؘ������4,�Q$�w��O|%�t���a�Zz�B���)�_�3�M�K>_Ҷ�����[ÿ̣O�����:�e��HK�N���H��Y�[ɸ���.)\X���RX���|�0̠dZy�N��]nlq�(�hD��o/��j�e���~%�g΃�����]����=���FĶ���p����r����|�gL '5v/�gc�����b��|܅ qȬO�;�Jؒ�L:�8ҹ͌��y�ث�����e��+�"bmO��^E��}t�Zp��4O�3��SR<�^��lo-���/�7K�,�Qd;2r�a0�Z��x?�.h��3༮����o�p�27k����:���q��F4N��������2����d@���I�d����@��VU�)ϬF�������"Ȩp�9.��t3DI��)��We���l�r���U����P�w�/�廚�ØgH�DN-n�W�:e2�w^+4Ȓ����l4�&��A0ͣ��#TE�j���y��?8ep�w�|��@pu\^����s�z8#�շ��{wc��TzO����ޜ9�����r¯	�S�b�j=]�ֆ��l�q��Q	�������̬B^�������C�)��Pe�Q�&�©�*Iw�нS��y,���<���k�0D*�YvK�+і�H�$�1��
,T�\L��p'A~��`���q{�ned���5. ��A��0kZ.S���0k$�w[��n�k����H�phuc\��N�U޼�Mb�%d�w&�x�I4k�t�ԙ���kK8m�7�F`��uJ)B�N.��"��7���`ӄ��-5�jy��h��ч�S ��������,�Zg_'S����^?�z]Ž�D��j�>�fx<��lS8���k����O�g��� *��kq=h��.��|�#"�S|(�~������!��Z���U�m}�B�&|ܭG��;�g��F>8�;x@�tb��'{�'���Hz��ݟ72��\b�čE@����Rj���R�1�`qαm#^�QG�N�����32�b�"C�(�`S8$ ;��W�v%�F�u'�jj�����L�Z��\FKf��n3�6��ɴ+r�X��z�g�!bٖĥ*�#�{��8=i�W�}W5���>�Q`:�Û�U!�}�$G�޸r���R���w��f�V��A>1��!�v����b�Ы_z~eP}���d����㻯�WO�Ln �(Ҿ�p����(D�v\BE������}n������q��Z�0,_jc�l/�e�w�
���ڟw�}�*S����b�u���|���./FE���� �!����{B��5��C�;�R~X�]��ɖ'6��#)m��5��FfSǾ�-qI�����X(޲���6:�7pmCA�W�+A�WV�������.������1Caȧ�?�lX?�i�<7%�Da|�+�`�⾲R$�lʝ�._���o$�4jl��	d�6d�+�$Le��4N9F�D�: ��,65f�'�h����4���l�[>��3!�>�y$8=��Ǆ �C�k+p[���Uk�Hb�U/W�G�5�������1bBY���/���T��p#��x~n����h��ݚ���K�e=����צ���N�@B.G��m <�?�3ÌY.[���أ���".f�vrp���nr���5

[0=N�D�,I�}��F��12�0ӻ��6'�,�����?3���=�#˴�\���c`Z��_���L���Ɩq�m�"�JRD��h��ˢ�*�Ǧ���3��m!ԗ���˓]C_�����#�~(7v"���+۶U2��qMK&����k����@������c�p0N�;V u*����8ק�������]��49g5�#h��K	3��$�R�� VpfQߩ�ӟ�p�+�5������^�3o��|��;ݖ�ݧG�\�F�C�܅;��ʄb}f�����f-eǂ�Ҩ�@�Gͦ�V+�K~3��XQ��L�͕pk�(CN'��k�<���SJC<6��g�ϣ�Hlo�l��A��)��]�P'�	��~]L��޽$m�ۃ��[�4�# ����o.�)<OG��Sv�et\-�㶩c���Ϻb:��!����)� �Ś�Xj�+c�ыL�1��������܀��9h��*-�N��&sj��Q���O{jG���1~fv7tR1Ur�5����O~;\�ADC��=��At���n�2�H�K�-H�c�~�E�k�+��	�_ �Ok(t{��M�U+�9��� k��'�[>U�>l=RG"ϪM�W!�G�[�{���u9��b��5���iQ ���?�c==PmJz��1:++���1~�ŘA͑r2�	}<�D�>-�n�<A\��&�*�wՔ$ �B��ӡP+ab��`.�g#S3����7��9��F�k�7���il)�`���9�s�8�qr2�NuM�5��0Ŏ�O���Z6J[o���r���DB�X��E����9������zh��jG���ZGQ���'s�>��&�r{
b�w��;���R��$3l��;U����a�I-Q���#��.��C�q���Zk?/�)�%5�9A���ڟ������a�T|-�l���}�
$W�Z��s�w#L { ��)ᚇ#�����
@�LW0�$����	���-L��N����m����t�J(�gm��_�bT�eH�U51�\!���)2���c��M�B�q���ۡ�,�.hݷ�C�[���0�e�l�/���(X!5������2��ᐄS=.7��d��>�9�#J��f���z��#�K1ȅ��ǣW�������MZ	F� G���-�We��f��D�9>�����O����z)�����}+}��~��`v�*��})�ϿJ+K�L�*�\�n��^S��M�+��\�1g���}�!.x��"�Ь��u�u���5����wud|�ah��;�?�gЫ���5��F�βF�rK+K���t2&����z��lԻ�����G����Js�'o����f��������8Ώ��iA\�H�]Z���1��Ȝ�m���>Ϻ��F=���[ק�BV�q�h���*#De\W���]��C�Y�����py���6#����R�@��\�P�2�)<�Mg����G%���Ge������CEyK�|�����GN�8��+Sk�?u,��԰���@]�<l�hM���g�F�,��1S�ld�&_����'��oh-�1��`ib�F
��p��\�p�ߔi��oj��SZՆ�a00Kg���+�?R<e~�(#����Cd`�m�"5�e��)� ���az%S�հF�%~؄�����!~�

���5YV�̺�Iv�׍�5t���]��"-��O��6��^�T�#J���L�V偲!MlQK�p���H��uc#|�A�d@���?��l�q�o>VR�N�D+��Ʒ6��fY�ɲ惘��nś/�5�������Ċ����8�Z�߸�l{Z��Z��O0�FOcw�U)�1+��B?U˲}�>˼�+���g��VBI��8��ӗ.p�?�:�5[]БilQP�q>�����t���^S�����aD���wn��裇��9�@X���f��p��2 �<�ͳ�Q*��?�����7�5_��GUH��;[IQS���T��U#ʴ����~�2��L��!���&���܉�D�%܇�)T��!R�����<):eT}��N��o����A7�io�][.�����lׅ�޴��R���Ph2jM���˱@'���yk5�9�bƄmG�����Loxc�K��N��A�%�&��F���f�!���$Z���� �z�KM�y^�����a��/[�;��������Ƹ	S3쒒7c��>9���v�M]wۋ�����w����m�,H���]O~�՚��JTcu[�Tm�y���2�?��|�������"���b���O���=�畬ũ%߉�C^�������:Z�@'����!�ow:$$�`y��v���t:���ր���y�g�b�F��{=6�J�뜍%0��c?�ܝLSTV���
�ɽ�Ǚ5s_�dG ��A5��9uT#���H�CZ�K��gK�Ɇ��65"�ubݚh�YڹK��:���D�k3�Ҧp�(d�s�hM�2(��� �4(^�7w�2���_�H���4��{����H�|��~��I��b��և�+��X�]�0�qV�l��(ټ�?�?u+-1Ͽ��&��]�� ��1��n��	l�F�a�\��kYZz���������{w<��R1�cΜ�8�'�WV�8�j�T��oԘ�)k���фK��L���̎k~V�#xjT�Js��0da6߉�u�T��bPcɚbb*b�̐���**�俸���{&��� �{�=䯓���(�|r�����];R�F�h��.�^h1��c]��U1_��tn��[��H�TjD���+�w��
�����$7g�l�5G�����%&�RI�w�Cc0񕎰�!O[@K�`��Z/F�+��	�R�r+=ѵ�OA%�tKb�/���0Hm{l��9�zh��(dB ��(�hZ:q�|D�B��=��)�u=k@:�c�J1{:�Ԯ��f�N�a]�#�ߨ��hd.JYP�������_�8n��ǂ�T�Nfҟf��5-6���[�?����������«ȓw�wC��/�;�J�y���|̓���I��)�/Ze@�K�fv\��ghs&�t��$��I_��(�F'�	�CO�����q`��C13���
��-����C1p�m1m�TKM���c�~�U@$�'5��b�;�'��K��aC5�P����L*2bB���׳��?<��|��Ķ���-).y��Ȕ�;�S��e���KC��iё3�}�1?n���﻿��+�Q������8�J����8V��C����JbJX:�(l��$���7	L�C���A�i�	��)����j���02GS�p]�ÀU�{�K��Oυ���L*��bާ��ݘM�5B[��剈��9UE
15T����ew�Zl��@	��:9Γ��O���R�#��e�Ҫ�x�B�+`�s��2����*�Ȯ,,�
�o-���-�������1@U㳯nhh,�,�;�5�f}��{?�v����X6F�!7m캗:�d{��%�U> �AẦ{P��p[3����V��_)�tP��G������щ�R�k��,�n�Dֆ�k`�5EBꃞk�pM��Gy+]T5��I@ֹ��G_X<�d>�t���q��v~�bw�"d�o��݋<�!�߾[{j¶��{ʲÜ��.w�����>$������h�I;D\t�
	=�4S���!��j�7��O�5y�5�TX�ӥ�Hd�w`�f�TbnS\ ��\ƾo1N3�YԾ�x�#m$��x�3sv���]�����S�^�^F�A�2K�����S$U����͉��8|z1~QI��k�b�,Yl-f�w[~�e�aŘ��l$���^Ĵ�r��n��[�\����}��}��O[ݚR����}Ն -��w��t�m,z�����`�a����o��~%��_���譙ϛ���A=k�{�^��m}���1�\�pj��C3)&Y��5�����s�Fl��[�>�#$�Ӎ0bk{P���W;$n�\(���=�-�nz���$ݺx+7��;�=��g�5?�Qy��-�_x�#ٰD�2g���a����^.;V>A�ק�IF�	�������m��z[P
�c�<�Q��+�f��AY}�.��D��Z�x>ԎՆU�'���mv'!�G�C�#&�w���;.�(�
���ântQ�G������U�ϟ���v!ta�4����8A�O���Ҥ�ZPW7���Q91�(�[�o_�l��j/ΜȪ��LN���.�][�A��A>/JH6P��8����Ǡ���2���{�B=�遦.��)�e�( �X��~��&���Eg3i�zj�_�>�5k>]��?@6���H�G�����̓S�U>{�s�����~�n�j�/5���X�R@�!�.��1ү���,��G�+/]�ۯ���(��Ú�{p,S?mc�" K^�������3sv�^~��˻��qH�Q���uql�N�C{cu��^WO��c���2Ũt#�m8�*K����%h�RƟΨ���@×4P���}@NCv*e�~.������������p���5�ͩ���#�]�T4��8�i����e&��1c���S��{3ã�GG�I�"�hvE���SxAX��&Q��.������!F�G*^��q�L�-���:U!����]b��c{Y�)~���9#����
@i�e�^��`ixp���"��>|Aj��F?�Gţ��aЫ�.��ƁM����ʆ��j��.5_��ޗ�W��dy-��R;�Z\�-���L�h%_�l���h��]KU-��R����gz�M�G���D��M^a(�_��?�!��
O�~_l�e��K�畞|_pıN�Qq�3���1���Ѓ	�W+������'��N��ߴ�K��-)��@I��)���b��l�k��|�����wv����m�r -��S8||
Vk����Q^�����tȤ��T�ۼ���(\�s����.�%��~�"���3U����u<�{����rv�;��Xh`�=�K�� a�r���2��Ti��j�K޸��jkٴ3�11\B[��"��`��iL�D�{<��*��*���t��.%��<9!��VJ���Or���2"�o����$к%d���Ӹt�Uݴ��:&��9��<Β������ �)�3���k��/3?)��L�~!���Ϝ�ޟ=�m����\���]�?;w�y�a4���x���D]�/�����jBؑo�䟱D���&�^�n�����D�[����&�E��j[3n��lh��׫zmV3�F��O�����T;�`$�=����c���^H�!4t2�ϔf��#b�F<����`a��[�Ջp¹bC�`�3'{�� ��E�����,`�#���=��6|X���8_��w�3Ɨ`O��9x+��1��J��$�ch��u�#b�Lؾv�K3~Μ�����:�\�0q��?pŬ���=�9c<kA��R��P���v`0��l�{s���n}(�7�Ǳm���rJ^SRBXC��6������Ȍ��d�-G��y_�zN-��?2���"�/h�m���r�դ��~��M�@�G�*P�"ʠJ�����pz�}���-`}CR��>�6��O��:Ψ�"$��G�Q����.HI	E6������O�N�}�YOBM;�c�E���l�/o�������H\����:ǿ6x�򩽔����1=*���=�w�ƞ�Gt�,s�y`��vqv��~���>�gKXy^U���\���P��/���Y+���rǌ�<��<>����%���$���00;9�<�{�.�Ԛq�k$~F����KM�dv��-{bA��RuK��� aouF�Zr޹��MT�A��B��(��H��%66�����n�D��GKd�W�?]V���o��>�Q����M�6���՚*⠌�S�>S!�ur��1�~��\9نxN��v�Ȧ5'�'b�����@%�qs~���3����T�g�)�g��j�~c�]��G&�Z��:͖r���$_Ѭ^��Hl��Gg���&d�/�SF<^���j��l�T��k=�c���������x^��`[���N��T);}lf�w�����֨"��qV�8�q�ڧG�wP!'�m�����^�f4=� &Սª��}8�J,��+̈ѳ���C	���WoZc>�@6 ��<���k	P���(P\%lܕ%�1�Bo�_0�����oܾd������ˎג�/���z.��=:љj]M���A��F�h�����^�^����h1>���S��3����q���<�0�+{�'�z�~a� Ud��`�d%g���w�#���C]����ѕ
��sj�"o$����i-"�����H�殪�2�L���-vѳ���V�G���	P�2�;U��PJS�
�4?�������r�u{є�1��ΞoX���������v�-=�&�=�6OY���P-(b*��V���Y�䅁okDf�L}�,��������R�B�3*�����5���1F�S���X�M'��M����Zh�q�[.�A��h���ٺ�k_�J�q�0�;;�~fܯ��3'Z�z�#�q�H���5�f��.�Xl|`�F@.�Q?�i�y�8����N��t������+�v�ӣ���|�Gqr.�'F;��.d$<`��8$�s`/2�����"X�a�N�R4���a��q��i�
�@�W�\�6:�w~g�kֱ�����v��h�gZ��y�昫�����e>M�S E��c�ִ!\k���s]+
���i�6������[�������O(:]�g�l��u/5_t�d��	���y��"g�hӂ�#�����|��/�u$[.�0��=��ܛ�i�v�_�L�ї���z�� ��?�h��b;�>����>E����N����������]�gi����?z5�7��,����c�����ܱFh2���O�V*���L�� h)C��B�k�y�G����/ܧ^*�,�szSdZ^�{=�_��/�]�l�?��o��+�������֨�b�;R9-��8��0/q��};3k���Z�fC�ޢ��}��;�_�~+�[���ȎJ��6�����R�|0Ɔ���+�2m���{2�ټ?���X���! ��v���Gf�F<���o�=#�6[xjbBۺ> rZ���(\�9�~���D��f��j�[�� Ŀ�j���&mb܅$����H�oJ�U�0:�F 8���3.�,Ch1��E
�o��e��c&�t�t�pT��b��B�HL��^yl?�h���;��t�-�$�~���o��U;�� <Ӄ�I�����	��f��m~>	ٹa�+�#�+xp�11� w�������7��$�.&��>v�5��$6��~�V|�Hƪ'��f��{��bS�����n���`��S;O[P��2��G����jN�Ŋk0�X��۽�7�(��y��`�r���%�m��2"����`S�V'�%
�3��Z��:2kx�#e����eV�/�@�3E{^�R�;�Fz���`)��� �^3D��8|��!~VX�=.ߒ��w���,�q"p��f���S�K�c/�O�tM�ô��ǜ�����s��`���J��}�n$��>)8�bl9��5��~�͈��p���-E�}�;�`1��q��^�o�%�WP��.F �۲��>�j}�	��<B�$�RdD��@l̗�����n�pʿ[;����A�"&���XN]oKzӅ�*SG�G��UN����H�hTM ��еWY���T�w�V!��7UJ����+������ZN��[/ ����;�K�*r9�]и�v8o0�uNS�Ź��������g�l�q~Yz253�$$�l���[O��������tO؏�ʿo�Sc�_S���K����
���i\B�z���A$��Ҧbi?ay�9^;;�Xs����>öU��<� [%�}t��gTW0�i�A���'�}��w^�v��/�"��pc^�X=�f�z\݅׿��<oʠiǉ��z������$S:�I`�c�7_��P����cbK��A�u�B=���^z�|6���iO�����Z��Z���T��e���Gzf@"�+�B�KC+��=a�܇�����\8����8|.ZK���u>�0�=��ڠYr@��G��^����%�v�а<_��P���*�_�^�R��@!�gp�#��}qS��hǽ�s[,�����/��<.N�K�1f�;е�q!>kN��P��a1�,�Jm�V��
۳�'���@�.�n�?.A�>+=�����W�z�X���z��f'�z{�G���?.���4�l�ثz�Ks� ��cp��TB�aȀ}0��nwd=/ZaM���������龜�lsX��?�.�V_��<F#w~, o`���X
���9�³X��n[㝷>dT�P���'���m��b�M�Mq�uo��7�ʠ흇*,�t1o�Tik���틦��k�[���=�W��5�ŪaRA�lz<"��.���q��3x>��f_�*sR�k?�yՔ��lC��=}1��at+�w
`>yK����%��(�9ϛ�,to������?����R�3"��&�ɠX�9J�,2���򻅈���G)��]b��b�M�SU�pe�j��q�6�r�Ç�|��r�T�j@�oK��i9}����T�8N�/��`��~��iG/�K~ț��	����iS��S���|��"�`�x*��.��U&$��&Ĵrٴ2|�	8
"2�^���|ب�
���E����8+��[��<&,7�$��A�e�����QE�=ZCCKŌ#5S��
,����d�V��aDi}9���6�B^D�E_�E-����/�N̂V3So���rH�V-��{�g��~�^ʹE�i����կ{�p4GG��jYhf�cdwk�0��pJ�O�z)��4�S�6�'}��Jx��0Z�c�j��݊$�j��z�X|�v+��lm3�q�����)�E����2!^LV\�{�.Fi�kt&:(JJ��%�+���K��p6�S%ߋ1�M��XQ*�	�cJ9�kVJ�Q<nv�L��vկg�qw���6/�3r�vA&à-�GO-�G����֍������s �Y߇g;!��Z�����,�h�S��=�EyI������gWTPg/|ڞG]����$�tR��[���<��rJ���a'dє���z�fx׹}I�{�FDj�WU�U�z6*���e�i�wf�{ �����B�$"jR�U0rlg
Ď��hf�<5���f�U�x�jp���aH�
�(�H/O�
���qa��]�����^�Q�����V_N�O�"��@SK.�o����|�6]��4��g�<akH��=���ۛ�=Bl��-��9�{�Ϣ���6�F{���l7wr1��\�R$�ɼǄUs�U�>������.�l���L�^3W��,�������X�j��M�0&[9�Z·��6��Of���,Æt^4��q;.S�RBbh�iV�!�@�0�W%U�������6�K��Ҳ�2V�\6Nnu�:Y˶m-��m�ԉ������~~�u_����d%�R<c\�`1�9D�j5a�����YH��#:�,��G�}��,n��!y��y�9�WF²�H�j���r�]Ɍ7Ha�[�T2~�5�VU¹F�h��7ֿ\�6�/ضed9�5 �x������C5ڵl�]�T�;�U�-m�bAO�i� Z�E���e/�9Rnu��{*�ۦ'8*�"�k�I�E�(S���ش�!��;������u�����+�g���"�{[䄃��9��Iy2?��x)���1��t!U��0(IsCiEC4!0Ecm�q3X�B��.�v8����[B�ie`������n|���Yg�K9�@nC�ZP�z�+YXc�_�����䕠��e�~f���:����JuA���Y{	�V�j��ǘ_�C	gbӠ���U-��.{�4��=�`\>.r�w�Ȕ�ru�� �,k�Qc���޶�t����V�1�fp�Z=��e[�����:�?��.Wd]{f{'L�G�|S}�DnA>w��i�m��ro����p�,��p�f�9�ţ�!AG��m#���(_�((��I�C]�p텬{�jt"�`��n��'��^s]/�sW���	1��|��.d&�侑�|����5eA��]A{I���3D�L���k�x.�Fz�b
¡�	G�x���!�c��(�[L��g�g��J�&��2��,ג����2e��8�3×��΋ͨ��+�\�������L�8
-���/!Vu��23~��X�#�x���@0v��wt�E���WsȤ���1B��j_M�MՑ ��[����!�NW8�ˈű�7�$[6='`�w�Ξ)�8�M�͈e�
RR��J��p2?�~�DU�@�HִNI�|��Y������5����v]O!���<`�|�C.����e��p�_��r��H����H��lW֬,�_&���766ĚO����u�.��n�VæQH�����#ҥ3̐�D���USms��k��pި�e�8P�w�``1)���!L���	Q�teU��E
9��yI�s\+�J�ԉ��J伎-'ck��=#�{�BRJnxЄ�?J�^Vz�� C�괉R]h8����M�T��]p�\��V�+��u���Ԝ��s���å	��W({��tl[^~��U�J�miN��ϲX+V�+�C\E�8��U�;�Y�3�ߟ3Vɀl;��T$�CI!;��:���<;�Os�Y���f�:��<���J3��Y,��oOD����7�|��Y۰Xbd�,>�Zښ�G�U�����܈z���(�hp�ew��bWG�%W`U���|X��u+�lk��S�k)ˈ��:�x�>�^���mϺ�����d��˄�ocFլ���B�l�+��J�tY׊��쇇�׳�����¼v�5��f|�(�`�zξ�i���i;ޙ�m��ɿ��bk'��Q+������P*S���߼�P
7�D��pZ��a�uVN�L�b�)�z�(n����V#��F�����O8����YO�}�#������G�[�i �C��.��}o*�HeN����4/���'�� k���NDUM��&�ќ�X����).d�4�Ĭk�YJ9
��ݼ�&�YR�X�A���_��L����_Wj�˛�L�W�d+�z��	 ����0���-��(�	�
�<�%Xw��ʰ1f��ܔ� ⅾQt�AB�U�	mgNN*��������+h��n��k����|ު�w�oMDY����ܥ�T�jE+z58d��@�L��Ӏ��P�͓�\DՅ��J�.?.;^���5M������ʍ׽|��B��Ar�ќ�@^��Ɋ?�B�
MZv�Dj�&�T
�l,���GErr���W�4�)�p�3`E�,]��["{\��ّ����X^�8�>��ý�3�T�7r���q��â�I��`��r,f��b2H$�!�� �o�HQ>�{��<CCV����7ʇ�8�hV+G�Hw�������r����a%�u�Ll���{�X!�e��L����Y��O�H���KI<:k��E4�T�F� ����?yC	F'�˻��1;����`
�<�����p��=��]�	���A�<��+;�n�����̊i%qw5�w[�6OE�b%-H�2C�z"�{\�:p�Ҟ�fL���_aב�*�T�ّ�DN=\���S�U�l�xۣ߿��s��-4�;��!�S֗��c���d������df]�*�ٔ+�Ԧ��C�-?W#��:ᒖ6��_�\濃d��[���{S�	p��\N���0|�E���6����"f(����|��eы�k�0o�@���D姹<|�e-t��)P]>������\�B'���4�"ޢ���$���&���OI���Jk�!�����N�ǌ3��	c��_�:��T��mRY�8�F5M��m�p��k���VcX|x ^`�]��z[���P
�y��сz����F��B?qq��pC������cf����`�ݒ�h1�C\,�}uO�&��'�P��^1	E��/���hY���j�)p1����yO�$X�}�T��3����I�Z�.���Q�s2@���Ġ��e�&Ơo��$�c�|������v�@�,$����#�;�s�������q���q���[rb��a@�<���O8�C�$c�Dc̱�Z2��tZO3=S��f�7|y <m=~ڊT�fC���^��0xf�򺦑�r�j\3V(o�&������+�l��f�Dޫ\@�@�Iib��X~�w`���@e$UE>�'R��I\�<��dyXVu�z]]�nR؎~�}��օeֺ���Z�������fj-�8�;�Z�=��}d*�
|����O��s��b>��1��������#��}+>'�}l(�>���d�w	����@��g����^Ӹy�v���en�t"E��}��k�cI����
�3�?~jao���F�H6�j����!�Ю���8��^w0��;8�¡��J }�(C�
l�m�;Q#��k�� �Y���&Z�ѻ9nS��l��^�S�V���٠��b��Lt�Ht;? A����A���C���#kV�,p���q��_v�\JwZ�Yt!J� �/����{3�,��Jo�[���Y�:h�(��u�a�&(����3���R-���n�'�^�N�y�rr�6cNz�kxT���6g���wG���=�1���e�1��&���5_w���P��A�� �{)����t��D7���:���fA�CJu$��L)�$&���
�~9��Ex�5�O7�85�;X������f#׭R�����9��v�772�]�O,��HH�3:��l4Ř�c%�>qՐ[���������XAp ��r�]^�fz�;C�ρ ����b��s����C��-��T�u�w�Dew���O:!�^�$T6�}�*M�����S�P���>��Ui�$�?��m�n ��KG�
=W�ko~���@��xğA/�[�P?�ѭ*�@�L�Q���# �US�Ui#Qj�Bcy��fDx�i}�]<�x��7c�逎� ����c�-��u�)2@��h��ɉ\qhu�i	e���|{ig^+B���O1��9ԃ��_{(	8	�~��1�8��|>4�F���װF�ݍ�Ǥ�\ױ<Z���7��@��@�3rs���5��)��/C�K��B>�n��yv���P}�a�b������q�𛖺'����zn-^&+�w	���p��z��Gw�b�vԕ� ���i���t�pӈ Hĺ�0IϩC�2�{uZ���61�S�^{��t�h��@��ų���Yg��;
�/#�qS�e�ş�{E�\&C22��a�\a��1�w�0D#@)��8�DJԙ(&��^w,��:V�Q�ج������ނHOj�S������O�ܹTyO�	^���{�IĘ".�$ԃ�04�� b��P��T�B�H��+�
?�*;+y�Z�>rK�k�~��88&3���'u=3������||O_����뉷��'k.k��
Y��3eSW�[�t����J㻙�`R�%I:-��Ֆ9�l8���&�����LDU��[wmæ5��$��|������G�֒��l雷��虮��H�P^FR��{>��Oc�'�q�N�=+7��=�4eSG�$Q�V�*���Fq��$�R{Ԗ݊�̾tx��7E+��o�Ӗ?h�v��l���1�Ԓ����Ӿa� �����츙z���!.T�%��gƫ�˴n�D:C�{`g��d�Z�����|q��-kI�y]�
�_l�J-�w4���Y�gu��X�w�7�q&�l�)��q�����R�8���dS#��/�P�>[կ��To�����9��҅�鄴bk�v�OEA��d�3�~���U��W)����?M<,]�l��5�^<W�.m���hr}t����v-rܝ〄���m���PQ���;ރE}6�teYUZ�s��u��b���ā� �����&l+?�~��1+I�R+����f��e��5ʹ��@��D����b����9M��3\��Bce�z�T͗*1_÷�?� :"G��Yx}d��H�[���$�Z�B>k��0|D`�|;iKf$Ap�򼎙1K�Ig�8kIa�v�uЩ�oW'2�瑂f'ރ<Ls^�E�ҍ5�K��0G�"�\�R��x�!����(��m��s,�~��gN��1��8�5Ս5������-�XEY����vW�pӎv����Uw`d^߾�#�^w��i��Y6����S�O�~���ԾT�vƂ�n�s�^�@�<2gLli�g����ƺA��*�oC��V����B��s���D��E�=b�g�ԟ"}�q�G4�LDJ�-MI�T�M���d8�����X[�l�?F?YV ��~`��uZ����|}d�O�����|]�x_�;u �c�ж���ee=����E��!d/���m��Нl^J d|(����4�ܾ3����t �*i��8�P�MI�+0��e�/�Y����v�K9s� P�lG�I
á�G�LT[��k691A�/��-:d_�Ę��`ךbͨ�h��l�C�)PFr��AB��]���y_�m�>����b�>�.�g�j͹=Y��g�d�*fH&����ro,�,�p��XE�T�jj���#��y?$`Te��(�9tcqy,2�O�C/!�v �6��$#��bQv��ȫ�\���-N���DEVux�Q�sSN썫t�~�3ފY�T�0TT�Nq�*��FD�F���̟�.���%�1p'���'|�D���Gċ��\ج;�I\n�D݉�\>��m�^��roQ�W��O
�yҊg�����	�M5X�9�CxZ_��*�u:Er��
$Yd0�sx��DQ�
��)�cN�l����+��U��Kl!\(���$v�1�3�D�p-l�N:]�xl���p�w��:�`pD.]��a/"�'	|7t���
t���{
��,��Ql'�.�������j�$���chb�Yv��}Ў�Ģ�`�I�W��Z�X\yr'�<˹���J�T_��ر��Ȓ"���f6&k���tKj���I�uՍ�,��}!��;�$���H�{o9�7i���,[�Z��fU)+��� |�M�JT�=�1,"�͆�=���H�� Ǜ��|�4E$�h����������Ħ-���X!y�����G1���DË~6�P_>�aV���?����h�5��֏0-7��X��������xzldZ�\���%PB�3�Q��m�f�����ٛiQ���@�B��Oq�U���+��!uO����xT����z;������?�ʖ�~��P	�G:�P�S�������ٵ�D��	QI�t?��F>��V��vM��,�mdܫ.��{pE��]�3�G���ѐ�.hxH�Y0s�}?c+L����2$2LsIp�6��H��fR�<~A�cZ`*_*ɯ��!�0Z�U-a��t|a�8Zs�j���1���`�ȷ�[sՋ���]�SFRk��/�4���EX�����E3�//7۫<WRl=��F�� �?��v&�k�(���x.9��T�-��y�G$=���05�<i���L�X�?*iĜ3�z��; ��X�W�bt�2q�� K��/bao�	�fHn�0�1�[?��i���9���[��������>��DM����w�[����(���5}�;�F�8�ӧ$��OO��g��/:�����o�.��p�N�olٽÊg�ܘ��d�s��,ϙ �Q��If�t	�ؕ�u\��8�ޑUds?9���l>�w�k'��Ӱ�I��+�&j�y���.Td+"ߥw:�.��l�T���2V5�x�\�n��A�����x������s�c����N�C�'�}�X^/?���Q�����T"lN��Ig�]U�(�sOR(�G`��o���������T>ɤʈ��"���<��\m�� ��WG�ǿ�=�|�\��c?xE�.o�R䳔s̽W�K�o�����P=׃*q!J����;b�H�'�Y�v�+6�I�Ӊ�[�u��f����->ȫP$m*��{{>�iά���ðb����<Yڍf�۵���A֮\���mI���+IEl��G+�V;���4=^ɀ��hI;��!51�a���E
E}��~H�������I8�.;�uF�UFy���a���&>����LRJI���[:��Æ�(n�%/؟��g��J�<��V'�'��{���.Iօ�KB�my�IQǙ�gu��NDu5g���͇�M8��t��/��B�3]5�9ښ��ѿ7�������,�wTMx��9���?��bg�銐�Ct�7�q���v���,h��H���p�4�3YW5�|�1�K�#��,r=l����-.U���@�<=Rsi��d�IНV;�u�%�(��-��C���iH;6�Ti*9�!���mc+t��M��G�bST�Mb�3"�H�	i@��L�fY��,�8�O�<�]��6��	2�/�l��sh-��� �����J��}���Ѯ�LWk�$�YI-z#g#6����"S%�����P���v���^X��%x�ъ��|��2��wG��#$zf�4���d7�� 
��V�W&C5
!�3>V������ ���	��/"��)��v�Kj¬��N]�~5�a�G�zt��;}o�����N����v��2�fN�wdb��鯼�<��IN� me;�yH~c���H����h|�V+���_�G�E�º�v2� ��إ�@�fӾ�V)_�zB����`��2�����WL19Jj_�����D�{瑳d��o�)쐁�����uo���Z}P�:~�q
c�����PIkX�0�$ �1�]��s���)�j�_������[.W��T�7�D�^�xɩ@O��������юQ� 7���,4�+��a!>�n�)7~j���y���g�K˜��� ���N+��W胕z>�1��XpC�C����[:XF��U��D#F������Yg���8���U|ޣ;]5N�kd�Ue%���K�^��ԍ�)�S0	�C"�qpd�߰��#aN)�8l,�S�ϥ�9Q���2{&�i����E��C��\�ͥS ���xH�����?	�M��������a�a�9����91��L�(�����-S�8�#[ߡ�k^Sբ���B/��{���n���z?�r��ũ�n������*w�g}��`pڌ���e��D�D\K��
��jB%)�)鿂ǯ���E�����^T���ꕐV���t��������v_×}��U-������xBoH�_�=����^�z��f|j�+�L��i�/rv�V�&`5S7�7�hă���+�?�h�&l�c��`��:g�;X�3��ν?F�i0����b�Ym��F��-s��*�`Ї�_�ټ#c�	3���Py��3�8ۄ@T֫����è`����	:���n�-��qӅ����߸≺���e瞇Ԇ��L��s�\fv&.�/�[����,%���^r��J���uIu��Wh�G����@^N�I�����K���SU��ߣ�X[�L#B�_Z�ҽ��f\��_�c��%3b�h��Q{yM��V�ߙ0��ug���ӗ=��!��]D���ܾBd6�k|@QV�뮌A�����nP&�f���nǍ�"w�>W�{���_�Mx|����K÷p�{��cI�1�<�;���,N"�)I��i?4�j%�-��_�\"՗ud��b{gQ��C ��I;�wy�S�z�!�{Q��[�2�U���Vp�}��)q���������a4%S�V�W��gͅ��4�N� �)�e9`���6�8ɽ�G���{dW��{V#�q�Ļz斾"F��F�b\���!�!��sS��2v���y�mj'93 ���):}>�
d� ɔO�C�Q�Ğ��)ɣ�~Td�ޠ7�=ddb�Dr�����w��QŇ�[��m�8z�9 ]�Ule��Y�sk:-�78Zs��l*����,qݵ]��X�;ۀ퉉��%z��:��I����#Ⱥ�76	aBe^�{m×X�g�M��z��С����fG�z��ls�Wg���[����.�gN��#�l��f�=,��@ܽ�� �J���-�6ꇃM�Z;���9Ӫۯp�����d'��x#�R=g"��[�1�}�:=�@6I�n���j	����D�NW)�k�՛�&��(G%	VS�[p�q�	m�V�}t��J�gy����滂��r9�tYF��g1M"���	�9�I��r-�%��O�Np��e��w���ܙ��z���mc^ڽ5�{�)��/�ӱ�v�y��bwMNf���H+��Ӧ\`��H�����5��h�y����Q��Dj�s���������k�n��a9v�x�_����dB�N���[��C�<-���#��d��G�� k���G�Fq��f���ب�Hubr��˴r�q�6H]WL�"��c=5pz
�Y9`��o�K�^r�ݧ��{��[:Բԇy�1��cwQakP��B,ke���i| ����\��/[%o��&i��5b��}(sV�i�;��;� �o��zڪ<ԣ� k�A��?�.uz$N�0	~u�`�)ϻ�<�V_�b|�y͉�"J�8�ԟ-����1�t� *���?��X��4�(�M�~�ǒ���z@3�&�a��p)�`2�~��?�p��pJ@`/��-���!|�K�M��GSM���7ߤ<�=�b�6����D��吵���8[#N�0�{��\6�bo-�X�G&���<���=��bV4��(��Ҿ���縥}����J`O�V��ב�y���_Р�DUM�C�|R�������4D!���Ë�����3�4Ԡ��i������!^��D��hI��@F.�4{'β��5;mE����AY�泿L�Ф�Kx�ǯIxE�����V��4�@!��曈:�'�7��"R2=��<
C��u�TBBRh�H��+4b�	e�A��Y�U�7Խ7ߣ��m��M��	I��e莉=�ܯ�;�Q����`��a��yO�k(�%�oyE�@Q����*��e�Rݶ��͂�ݬ��~��_�4^�@�.������|V�>�D�}�[8z�ҭ�o9*_����1�23��(�������O2C` V��������jġ;��A���I�3�}w�,	2/J�O�6������ߝ6�X�DC2NWB�D1>�	xɱ��`hHóa�J�������܉����^��r���}Ӹ�L7�Po,Yݲ�ŋ<�%:xrU;�?E��Q�Co����<�%
��[�;x��P��n~)F���x6S���{��j���z�'�bA����0��B�P~J7�/��7 ����{�hW��8�fr �i'�H��6޻ўg�������[��
��ϧ���a�|���I�H���v�g�"����&`-j�҈�+������4��Kq��e�����dԧ�k֮�"[Irhb��CB%�@j3�<5��Sq�^c�N%eӴZ.�HO:�Sv+����qq��(���4Q���v��C��%��\ʽ�7/$E�F��#%�?��ck�V��i�e��D�u!��ܟ5'&��R	ȣ�8��8̽n�����)�������y�w��6�Qp�c���^hC���K�2}t	�_9p�32��-�5��Q�e�f�t�H��6t�^���sT�]���2�7�'κ�b!�b�Zq�,�����2�j�'�C}�Hb�[��E�����2�]�TT��Q�y�
Fm'o}��S	����������D��w��3]�u����C$`�B����:;�A�C�yr%}9[ ���G%7� �k�kL{�T�D�ݾ\=}Sɢh�0
P�K?�Lcm-Ӓr��y@��2����9�Ŋ'N�8g����qƪ�E�(]���Td��:��_v���"d���SL�Ś� T`~w#	����o�r��P�����75��1�p|C�b���z�� -�qN��c¾���^���jb���t�j���dU��b��SG%��E[H�36�������X3w]�C���K�������Է2g;�̱�ZhjƲ�_����'�Ý�c`�2g�y�=���?�t��hWu^�	_|�s��R�G���?
*/�-�:(�NS������\�Y@+��ȯ�}�R?G�xz�"Ug.��*��~E��歲�*�f�N�_�8�uڨإ��j<�O�@k��X�����-{����.0'��k މ\�>L�|�;,�[S��;��߭�U�p1$�^}*Ӱ�BS�f��/�PK6o�����|�jh]�ƻ�6	3|�lw�ﾯ4J��՟{ NSn�����a�M>($iU�~,股��ݘ�"L>���}�c�~%����W���/g3��{�U�e�̋��|��&��|�/��gSc�}�3������^�	�ݣ���s�{&��3���r X�����
.y�'��͕P�єp�+:6�]{D�;��a�����1��%f�A�wP�����H����|~!����"����+a���m �+:.����
q66�W�htО��F\�>#���z�ݿb���ԣ��)�Gi�����PuŴ]2�Ϙ<����XF�^A>�E���t%��n*�*�_��ӱ�l��`�}4��X�������^l�)�?�D��a�nb���7�۸��K��C�00�"�a�{�Z�|��Э3`�����޲%�� ��ix�H�,*��qJ�D �7.�%W�9��Ѽa�`{F��+�ú�I����i�(1��
�뫈z��{�1��iy�6���wj�ZD�X/Y�Ɵ�\�_TyX%a�H�J�1�#-m��Ch�o�l����ݻQ�����WI�5|-�L��Y�@�z�h�B��1��e-ś�]d��J��w��<p����T�2<2�\Xp���0N2�'�SK��+45?�����[���R��XL"��?�@�<j�X FC�A�G���NZ��D��Nh߇ZJ��$�L�?p�L5�5tZȹ�I�����ʢ�u�]�&��^�Mg�̖ӌ�p��	�j��O.v�7Ɠ/��0��
��
m���퓵�I�i��s� �L~��MB+��_R����� /E�J���k2���� A�Ew�F���)5�E�жK�<�1"�:>X�2�c�*�:d�@��tԬ�v�1�5�ҕ�'g�����F�:��Iҁ-[c��[��L|a�fC��/�y�0Y�S�v	S�OP5K�a���ak�Q*�f�N�S���z��ˬ�t�����|��1��
t1�R�j�jk�S��� �2H@���|���8i�,�*�4̱� @�;���^��Yo�Q�B�����> �E�Ϙm�h���bL��$ЅAg���x��0=d]��^�=X���>���K��o�Y� h��7Q8��X��n-3>�����/R���Q��/�����^�`�!p���{�ѯ?C,\O2���X{�?r6O��@r&� ���(������%�Q���m��q��x{��Gןa�^����xne��s��v�<������;}��	����tA���x��,a8#��Y5�?��0H�-I����6ݦ�_��O�Q�蘅;�%�cD.�5%���O�,�I��%�hިF�ՈJ[��d�� ���5�Y���SP	�q�q��nm�5�^х�Xp��s���
S�pZ�:ڼ�'b��A!Gw#G�nOY��H�9��I��z�H�/y$���0��J&����/雦��FgFz�W=~�����G�����qdEdd�������njJ�[u��&����Pw^1�7���rd���$��P������y3`��y1������؂|��3�knQ^�W-.Yd�ص�'c"�9��Ut6θ�˭&�h�{\���P4���$�zZ�L��O���-���?���7S��u�Q �������iĭ�����8EZ6xؿ����א~������e~�\���|��@k[�� �K��Ƭ�u{�r6g.n�� !��e�Td;�b�#��'t�	�͸Q-�)�?h����T�����c����آ�΅tb7��rU���Ͽ
(j6s���=Y-�5��^�;�AN����Ntu&t�"�<�i	ہ�'��]��,��אV`j���o���?J�v�_�5$�s�W��f�9���^-��a>��Ά���z �d U �ܮ`�1^����"c��]�yh�\��<բR�,�y�k��#��_���I*k���>�ן@n��%�k��>��ai<��Ժ�7Ψ|�Ez�R�QOqd���0:��$��Ik�u��y�ty��e0NimKS�[~R]�Z��^fj��Ɵ_�)
D�t��s���D�H�|�ξ�
�$s5�^���b�X+�r��ҔƬ��U5q�6���pgd�$�q����t+��%��{��we]od������h��e�@4�X��R��OfԆVp��k����o�=�Y�L0V���H�hM�('�"h@�6Z�V�NC�=����W�C��D�7%|�.>R�ךϻ��/ɷ���m_�Uڕ�r?�=`l�l�˻���%�9�7�<������32���J��'�	�y�=��p��2���ec��(�C�;)U���Y>��[p"�7Mh�pl@���TշG\��T�v��9y;����ˏ�q*����<�QC�f@c�y�~��$�>P�$���i=�������?+w�=Iiiѳl�_2�a~՞���U:���RF̩�����2�p��A��;�nλ�l_�QYU=]�M��@P�)6�=��a�ʑbbCX�a֘e��B˅V���@���%Y�qzwSLRǝnG+s�ªi���NN�As�&\̃N�-�e�oJ�a����ÊW�V�D�n���������O3l�����g� ۄ={KwC�]�8��X�0� U��Oؚ�?����n<;#�=P?�������$}��<�3a�5f� ���4zqY���a��HMp����w�ΛW���ie#P��������+��2��P:�>����Y鍭��Zֹ���,k�ER���wX؛D5�(��U�V��N���0�Oq�	�&��OFC���_�G�cT8��+���9Յ�F���ȳ՛�(�f��l��'B��
�~���D��w�z�7�^x`I7~�'��ڹ珇2�1Y�1
�8�Yveu!���}��נ>�],��'#=������m��p�)��hY���)�tcExw!���v��sp�6������%߃�Y,���jPaC������fo ���q����{ni���m�B:ꥍ�Y66�x�C��-�&�6t��5χ���dxN: �0H�~Tڮ�-�U=��$�˥7'h]�s����	� �KԅE;�c=��SS῝��AG��v÷��n.%l�B7i��D�Q�|T��A�qL�PY��s�%���hZ��B�䂗���`�.�c��35�E$�����N8:Z���DPe�v���hC��L9au��#ߵ �Z�ߡ�}MQˌ������������'�-���U�{�����I(lY��J5(RB9�Ϙۢ�g�K�d�b�/*�Uø�j0\�uwm���AE=[���x<�ض�{��5��uvw�O�\��^���_-[W1ӏE���E��/�ѧC��]|�΅�\UYO���2BW�Hf���W�v����^-�ԁ��&/N&Ѡr1�$���R]b��B}�1E�����7mx_���U4�˯����71$PR�^�����0��5�J��F�n10�q���Ϣ�e@�����Wj�����4΅�p|��ʑ4�L�)E�|����ˉK%�����9����$^>���Vc(�A��J|�����G���
��0�,'֑=p�����0tR���Ol��d��7F
�Ln��dX�z���]�QD�Fn���ijJ�o!�m���**0U���	��7�T��,��l-�]�&�V2���/�f�$���z�cc�K��L	d!�V<h̓Ȱ��vw��v)��z�
Ӛ�i�n�A�M��V��<�ϝH)��v����^��U���xfoM{(�<���[�Q�ί�����F��Y���k@eģ@F��ܡ�h��"��F�:@{5Ze5C�]���N@�f�����?*u��/�Tf-U�ıHͻа���_�T�M�Q��;F\�<9�ָ�#	\��Y�O.�v1� 1ݩA�v�oY���&�J�)�c-�a����M�_545-�-pg�����LRլ�Ą��`�]��rvH���W�32�LQ�F��M�P�}K{ {p�;���&Ԙ�o���>�!RN��7�C'���tl�@�bk}h��飈�9.iv�}X�ڲ��M���j,�(��dK�_y�Jv��0:��@Ŕ��Ѻ�-Yb�tJ)Y1�I�G�n	����4z��'�l<�y�؜�&^G$�!v�!��[��@��pC���#��g 7�{@d2Y�\��R��+����HU��@Z��|���`�f�"�Laϼ B�W(cō�m�S�s���݌��Ǧ/Dj���S�%�m�WH&C6EGuR�Ή�������sR:�1���cJ�%���f��O%�P��䈮	��Y��x�Q� ��M��'�����ϕ��b���	;��� �2#��z�@���)\zlul�_�T�-2n�c�zm�b����������^���I�+�Ljk��4	5Zb�~kJ��h�܎�Lo�z�����h�����ȩ9��(>8aP��8P�y%p8f��j'���$l�x���*��q����
��V/l��j�E�,�M/�0n���$�	���o%��d	��(�1=�65+�H�u�����d�w�)-;���@Z�ݿ�[�&�RB(`��h��#<]a�,;���o�7p%�E� ���1���@Сl�7@={xU@����i��Mzx�J��o�_��s�a�i�c:�.���%�����ja��V�*��Ѿ`0%���[ٵt��?�w^�r8�a��?�2-�6U>$�X3�Ӫ0�uB�efʣ���9h+B�Q]"�����9�z�d�=����x��+AyȭO���yj�kٯ����/�U�XS�Ƚ�<�[��I1e�-7�f��;J"\[��y�^(gA��rXSH���?��.����E"�5�֦��j�Z����8��~*��3�b&���%iv�YLt+o��^�V� ���z|	��Ep���k��se](8ŉ�4�3���WF�b�M׶�C!�5���?�N������
�0�9������p�9/���.�:lɢ�5�+�N�ڜKX������o*���5�8.�,-S@ãG�P�Ԥ�����@�{�N4�]����}V|�R\W��;�<M ��_�&�jr`m��#3�dX���(�jh:u{*\9�&���Vb�7��4���ҤK�
�2N�P��Z��t����-�h�x���S���}ә.��(M^�\�} �.@��3��4^`�,��b���I	���VHy��2���[yF�%G�����g�/��W�7G����Q�����K��Cl�"�$����T!*�vّ��S�/�N�cn�2n2�����e�����-z��;�l�ֻ�{;<}\�&J��#-�F���]pm:�|:��{]��aq��yp�{4M��2[��o���&����=�yU��	9���2<>��]��xR[n\E��@G�g8���)�-�Q@��@��y�ؒ��µlؾKb�i�Qm��.����֯av=�����>�>�J�5U��A�u��=�Я�cڱ�&�b�qcQ�$����Z�F/����$N���9.]r����\���zL{A��2�x���}q��7�{�]������9j'x!�i���[�2�17D�vd��s�^{��|ڥs$�3�a!>8N��g�4c�2�t9GT�\XBY%z�٦��,��rs��V��C{�\���#��Z���;�r4#nb�#F�p�!;c�Qm�-b��]]�}�mU��	ݵ�X�Tf�ϛ��9��GY�0E�X�P��6���BF�������w<�"��/�S�����N�bQ#�M�R��\udI�|a��O4�&d�s[��V5�U��'w=�'_��D��㵣�}J�4+���=�����&�F�;Xs�%���[����tj�}j����3]�]�st1+�G#%���~�:�f6F��o<3��
���'A��H��HH�A�a��\�hӈ�-�U_#���h|w�p�������懘ݫL��]�j�"�^��^����o��.O��`���Ɣ-և�z(��Y �u��KB��e�8�[	���+t-��A������=��t-�;���c�}�������Y��0L�ᐭSO4�4&�d�w�p�I�o�ב��&��v�̀�����'�j�s��mOt��aal�UME�~94;)��"vS0�%R��[�	c+I�)YWB.��NE�����I�
��?�0�+Y$�O��cw����G1|O����W ˀ�x��t�vL�긹�J�[���Ｕz_��xKS�*�}�����e�m6X�7YQ������m�s{N�A{�n��@tر��h4��d���(H!MpI�������T1�9޶W��_6p��?��Ŝ���	�������y�/���U������wXt�Y&�7�z�nMX�o����힭=�u$��?'��K,H�|�����?'+2�	:��'���Hil� )�BjѪM�dpm����&L�k	UZ��]:%)���g~�����wf�?W�w��H�/�����?��&��0�y��$r�tm�iI���r�ZR�*��r��z�h.�C�F�*��HM�����N����GI��G\���&F��KA��j�����z)*He[�D0�ȍ���]��B)����笓.�u�KO�n1�����ז>d�M�_~��ɢ�uz�3�P����L^r�ֆ������>�p�Y�o�_¯����8F�t��h����K���UC{a�ӫU�j&\V����Q4����/��������mn{(S�ڳ[�mT���vL�j#L�fM�����/�Ä������蔈W���t^뵡B4`�h]�I�pI���8i"pK"��[2�3�.]|;^~���>:���~�Q'_�Ֆ����\߮�!ᓔ4ox9�\�k	����=�#��|���<G��a�̿���܃i�,[��VqB]x��A�3�����uH��ky�(ZFc�ǟ6q�����u�����/��#L���Xs��q�a{�L!WM8���|Dq7�M(�C\���8���#Qi�S��3o����Q��e����X��Qs&|��Ħc&�]���t `�����Hu]�@�"������!{n�}孿��v�8_|��B|�-��֛���&k-6Y��ŕ�H��G�`i~�#<#2�%:�ҷ<�뷠q1%�A��*}_vg8�[[��Ca����. Lk%�����gz"4�iA����pYm����>��qk�螗/n�ύGQ�j1��9	y�W��#:V�G�C���֫�[��S�{7�3�Z�������C�\��e�QH�Y����И��ugYe�����=�������������`����S�D�ۋ�Jq/Y����oas{6�,5���#]\|��$.~�b����>�+��#�������i� @EF��1��xZ"Osxv�v��hW��s�����zy����ۡa�ɫc�m6�gf!�E����U�o(�2�] ¡y��f���x��Xt!��ξ�.�~>�����O�	W��ڭ�Igi����ra䢓���&��H�,�j�B)iN�w�%7Yo��������'�>���x��<tX�f�w]�P���me��xs��2�	�Lu�$UF8�0�zo�Y�$��B��W��oA��!��j%�8c,4"�熭
��t���Ѓ-u݂V^�e��42FQ�mn�+��^���b^躜�x���m�Mv����`NA��DS�WI���	o�b�q�%����wpRU�����)[ �WAAA��`��-�7T����j��ލ�b�FM�1jb�b����]�m������sg����,�3��7�4d�}����<��G���#W�����dd%΀I��Z����<��rҥc�g�a6bQ���y>�|�w�/�����ś�~��3�G�=-�h=:��u�u�L�GǹE��ap?�k\vӣU�i�� ���vĎ�T B�YP�l��`��3dH%VI��X�"�kp�YW����������o��?�1�LRn?��Ygp�TB��M0A��>� =��j1m�X��ז�,�͂����7��gTK��2D�~�t�j�w'2��ܺ�K�xm� ��	z%=����ۖ[<����'K���.�B��"�&�k_w��{�+�ݢ�ȅ7�ddV���p?H�\$1J^+
92Hu��_����r��������.[O��[O�A��Ϊ��6��%La�Bn�%_~;�w��d��Z\�Acÿ3*�i�t��I�;ߓ��V�{�bb�[]�������[��r6����в � ¤Y�t��Xc�0:s�Cq��2���7ZR���"<�����Ҋ�ё�5��TP)�a�L���_�g��ˍ˿�_�0��+1��i�D�_��m��Iv2���8�!^O��L�@�*���(\v�#PP�oXuD�Տj�(5dm�iV;���}��Y���<af7�?��\y���j������Ǘ���썡�5�z�4��9,(/�[��J2Ê���Z��@+v��T��W�{��>v{t�,����1��7�H�\�L"����Np�VI����|�Ɏ�}8����_u�~�<�zn{
���8("����k��<t�m�mL5Ds.�"!쪈�#B��j@ѝ�_
�rj���b?�������#qsG�1�W�|VX�?j��8�D!�"�Y~1G��[U����_:��(�&���_OO�~wF¿N����Sԙx���#�YW��i/�`+@��D�4,*gp
D0��q���O���5�<�b�
�n�0낃��D,��@�����σ���>��ւ��lL��އ�ï�~���������~;��m6�(ų����f���z���lH�4�sv��.<�}��W�߁)�)G�(S������Y�ѹ?s$���0��u���}��ã�-���c�{�fX�(p�{�Z	/�pFz� "����-@��f�)��eg���FَpyF��)�G�܊�����''q�e���,�,�3h��;7w��뉬�,߫Q�r����_��B{�s��JP�1PD��c�^�M�d����'qج	CF/4:�T��$P� ��dun!��d`:�R=�/�*��o�R>�1���k�]x0��V 	�ZM�Y���u����.J՚@VH��$3�a!�""��L��`ctF��_�r,&�Ub^�-ׅ%���IU���;Md����--Bҡ���-�%.��B��Fl9e5Ќ����"�
��)�G�5�A��R�Y�} �N��DyMmX��2��}p���M��}��x�_w��i-n��D��KUEhZ���Z��c�s7׈�R�����g_yT������y'�=&���C3{�d�)ٲ/�(yR���x���m������__���n\��}���[v.�#/@Ns9�O$<�cp�?�=!�i;t���B��.[��[���r�^���G���;sWP���U�B�!��9����3�X�-"{��Y�5RM҆uW_y�ݷ�4�����G'����)PD�gâ]p�l:f�,JF��0���sd_2��i��c��HMN���g�^�d��8���P�`��Z+���4�a� �� N���hi�B�f ��72��8�$ئ��S�#p�P���Me���A�6Q�ñd�lg�,�=�^��o�/"K���D<�xMp� �h���-J�*�0��1�hV]�~��q�O�Q��B4֚0�߂\!D��S���Y;mhy����w�S۲pσ_�Ix'�w���ϡ�N1e�5���ʂLq��h=�Z׍m��\B���7j�Pg�0�_3ܬ���fx�=!����Y���p"�Q){���G���o�'�O�KoxN���q����EL$n�����-�5aA�} L=��7
DԷ�6���t�Y.�{w��h�t��?�SԅB�!�3��)�)�Ӭ�?�E3�����ր�}��m��5��^x�f��W=(�("�3�f�E��v�]���Bs����Q��X��%-VN�U$������e4W<'�N�҉��	�"&v*���
N8��#x|��v��D:@��L�a�ёw�D�C�?��d��D̊����o�k����a�(�Ȱ^�p"|�/�j��)�j��p�ע�j�s�e������hh�a�!ێ����m!��(�鳘�2�:"��`�H>�or�BoȠ
1�w�.>��ȸ��Ug�+[ �HD.��1E�n�E%ɠe�_$:͹>}�«��;�D�B���x��`���	�ZECjaX�I�E�"y�Y�0���+����p�OnS�DA�w����9=��֕�c&U#�XB�	�G���ef��{���-�$�|?��q��{`Ġ��a�H4v�6gc�x�B�A7�睴3�=�N��֙G�uΜ9��ОPD,8ˍ�̈́u_l�p�~o���&m���nO��8]]��^�s_z8dWL
Z&�:gF��	ׇ)�;���Kt��"�=&���c�۾17`u���?�&+,mQ�bqXU�>�2K�d+2[�	������9N<�~I�~�n��6� k����5��N�GFMYBX4�)4z-S��68�C�X�h`�^��,�{�⪛�0�O�=Q��;������Ͽ+?�oL3Ӧ��1#��Ѧ��C���3�TA�G�?C��D��Efd L��j�g;3q��Gc��/Ti�u�j�b�+!���
LC��&K6�'N��
�^�Z�s/�=Y������|:��k&�i\�n��5c[�P:�
�nB456ɌUU+��7�z�jB���#��F.(�3��)�h/֚��[a8E��Q���g
��ys�������ј�J��v���p85�;'�r����6@���'��Γ��5�>~'T �
���e���W`�E���Ѝ�2�A�<wB_�Mű�8f��|���Ч�CEƗ{("���|�y����e�}׍��cBU�t#8zZ��˖$�
�7[и��㥚I�O����wޟ������]oNH���ۭ�i���$n���q5�ĆFG�6��Z�	]O��:�$DȘO��x��ω|?��*Dw������������3��DL��2�Z	�O"Ka��(<h)q���
���V A��`f6�ȧ�G+n��0�v�e���%�<s_h�{�3��7��e�-SlA���W)���Ǒ�]��o	<Ϗ8�&�p�Ah�^�Չv�&	�9��p"Z\�<�:�p�P�o��p��#I}�4F>���p,�d-��z6��t^'�sk�>A�>�م��S��VPtق����Dd������E�sN�ǝ�Y$=�T��������쀕��kxD*�����h;����f��0�����"Nz��j�ڻl���w��2��s;���j���<p��u��r�6vb���R+�{�!�d p�pVxՈ�~���'��p5��N;N>��Q�ݑ�'�®D��R�a dd�Bz�M���ψp��9𸹽��>[;o⍷��܉�[��L�����cچ��ݖk�o�E�U�wB�8g6ʊ�T09�8h�y[�5��7��p�?��^UM{W�TES45�̄TgA6�&�O ���i�rhظ��'d�8�>Q��{���ġAkF�S���n���umjE��X�����z����9ؖFgCr�&א�ZHy��J!�Zt]�[DY����j�_^/)���/�'�Ĵ�GU���:Y[�ιR�D�0�B�52�'6��e�w�̣���a��}��1��N�mH�u(td�?�O�U��IS������m��]���W�O���@a��"�=��1q�Ň�"�E�.�f�
�w'��X�Z��n�[I�d/Є�n��ᝏ�"~'ꑏ����*�pȾ�G��S�*�&b"dۖ�|Q�Hw�q����hk_�|A�jZz݀J���]t7����e�����'#���o���S1y������C7�E)*�~sb�*Q+��Fli�л`���w�qgކD��:��sN�I��s��2��x��rs1�(�5��Ͽ�����4�{:R����&��
F*��3��!]�.	gТ���$��c������g��zE�����hjnD��M*�sKI���yJsE+�YjO��~�]�x�_}�_��j��Pt�g�5¤�EC�%!���AQH���6�E�?ң��>�N��w8�������Ŀ��t���K�qHi��LW��'hG��Q�B��0t�y���q�U�kOУ�����,�w�q{�g�m��I�^�r�V��݊V2,+'�_m���Xt��D��/[p�Yw�mޏ��:hk٪�����-0�<m,.|�ȶ@�9)̦�t`�	R#���O>�6.�����r�W��(���Q\u��p�5VHDW��&dA���\ht�eYz��z9������{m�Knx����p�8���t�L����o��%^F+ �,\��?��Z[�����W�v R���S���J��ri��l����zä��t��P��p,�梍(���!�ץRE�*��T��^th��3/�5�~�8t����He{Nv�Y���
: e�NS�0i�����k������'�A+4�`�U������5��xd_������ǉ�X�F��s멗�6#�΢*Ai9�"�=���;v㕇�kiI�hV$�ĀC�0�(tLN�K�W�/SPS6�us�p���-c�ᜓ��wނGVV�;i�|��
)G����A���b��1Q���W�����r1v����xN<d+�7q4�V�+��6l�{�gt=�V!��B�(�l>y5��އ��o�@�����!�lV\J�E�õ�n�4u��o���r�������Qk��2�z�C���`�����$��6fq�H�6v�-�﹮��묄Ǟ~
�N��i����}�����3��E�xou��ډ���2L̞�F͵�cg�CO���m�9Vһ*`ƚ$2M�Z�1/�v%�cڿ��hEO�Qg܊KO���4@�=)P��}й�+=*��|����˹����?��ZM����}�!}�6�Mj���4陲ߞS�7�h@���O��aY�Jp��t"j�h�٠`1��J8���:ҳ���c��d%��N�P�CG��kĈ2�x���p
&*!�Y3��T��X��-��g]�'�2�K��T$�B�]�ȥ8��0n�n7	���u����ǁ{m��^��ڔBl�Bþ{LE��(�F�qV|�Y�̬:��$�E���t\}���Ep����?���8����"{>��@���Y��4��b�.[b��Jذ���k�i��|���z*����FTJeX��x���IöqٍAVC$�|I�>�w�|���Gd��2�~ �4����֊%{F���8�;�S=�[����S��`�= ���?�� f��8�1��2t���p�@X�w�>;���s3��=��S�PD|���t͹m
-�陛E:,�n�3�02�Ļ�8�`iLz��mȸ���5:4m_nee�ڈ����a?��Cu�N�4F[n��P���08*FЌ��u������e�(9���!�<��ou��/`A��C�oA�瑱#�+H4�c!�h�	2.�hz��k_���3/��9#jK��whNQ�in���y�4��(��8"�ل��o��˅>j_�+�7��꣊H�Hּ
���39�6���D,�*&��)V
{b­�_�+m���mhB�	���i������;�=�NM��N�~af����e"u5�l����@B����AP�i6b��Fp���{��V��q�Y�cP�QVDfq7��R�|�Tq�n�E�%���Ҩ�kil�
)ʙZHz/b�_��uс�p�5�t������_�Al}�u��ŵ�`~��[��&�)�{���Q˩KFJc*ǑME]�h/WU�5a b"��1��|��>^П��}���W(��iȨ ������66A[�j�M���Kz̈=�� ]ǡ3�#�H�j���~P�V-��g6=O�暱��&l��h<8�M(�F[Q�k�Y�MV��d�p6x�d�\����ǳ/��Z�K����c6��_-;d����R�z/?�!c�> /��	�ƍ�{d�%d���������,g�V�����S/�������Ŗ�W�k��<4�V�lt�Иز�8='�ާ���{v�gI�g^���ٟ���L���5�~ko��9hn"#�
��D�
�J�?h���W�4���?��J�[N���������l2y�Ɔ�Ju���C�U[�dI*��*��5H/-�R!��r��H���fp{���6��422|���CN�Uz�MZ�VmB�H��Y(�����Y�1��V�l"�Z/�z�y=���w���Gs�߰��'�t5D�b�Z�x�Pp9�ށHJ�;��f���BD�']��7���[�f��A2�}zn�`��j�!\;�J�*4����Zǽ�����]���b: ���!�t��V����x�a�֔u�fe��>�2R,vԴ��y�3�:���Il���5�Yb23 �Ϥ�<�>&I$?�x�5p��BO����pf]�/���~6�R��ȯ�d�D�}N�ÅB�!�#�QA+Zဩ�����_��G_���>�����/�h����O��PK�F^d�3K��R]�J���*��.���e�|�V����܆2��|>�RXF{{�C�W$���;o��m�ܶ��##�-�pm8�R[lۅa�(!v=��D���g0n� �^�/t+FK�B46�F�V�!�X�c9�z;D�Kp����d\���A�v��a���`dD�S�(�MXг�WAs�	�s��ĳoԅ#�{����\��R�Z:��Lb��I��K����4vJ=�~��!��@m`e�N���#���壺8U9`���0�� ��H��T���A��h9�<o0���j�+�~G��M� &��@Xsi�h�
�v/taӢ��pm��Y?�~��^ނjK�6(|�PD|��E���9i��\��$pu��?گb:�8]}[�8ew3�~���[�O���mD4>232,yxF������I8c��q:(�B�iT�Ô�b�~+����.�Pz���ٯ�'��|�~�ݸ�W���egX:ʥ6RaLċ^�}��Gr��m7[��W���ј3e��7Y��[Ű�G��,X���F�8�'�/����>�#W�H9N��wB:�����!o���������H���z���4�׆�/���!���p.��8������R==3R��-�1��3#Ljc'᫘~ĵ��� �"\��8P�3�u�.tT���,N,ǈW�p�;}�-LƟTR�wEė?p�e�:��h�����+�B���$�F�������:�$S&W�Q>(�P���&2=��J�G_E�!�r�m��m
�M��PN�\.� �!X9���t�T\g�O���QϘ�sN�"dd;�TdӲi��D�]Q�M�i�ဝ����>��M��ws��_��R���'����+��RMܴL<��[��H̦k�k�u��,GI��>ڑ~̯�LC4�.��k���ۧ(U�-���1Ms�Æ	9O��5����b������~��7�{:9-�M�����`�6 �8�t�4L|�ʰ5��3����h�lkj�9�vT��T�6x�v��^�i��~���9�iʤ�+��ܛ_���{P�N����^}
ڔ����YX,ܮ��1R�D�PD5�+H8�("��H$�(C�M�s�p^d`��Y�~�ѿ��VZ�V�C2�z۪*&��A�!D�2Jc���S;�����񿽃�	� r!�J�!m���4Y_	����눈+Wsm��
M2��ԫ���̠y���'�k�
�4>��~��>�k|��K���O?fr��~���}�������FY���DG�ɖ��S��G�-Z��n̗O>?��F
a��x�y�Y�tN�r�p��-\���^MD�k��7�?{57^z "�\�Rgd7�-�Z��r��)AR|�a;mz��W~���.��-��wEė/p������4�,OJ��p��E�;L��	Ҙ��$F���O�q�V�=]B��\����pdC{��/Z�[m-Kpm���ց�!���[C8U�׌�)O�$BDs���ܨ]�_��z��ZT�H��nҐh���$�h,Z�:�4ۘ��0<��GP���F2��P��hqah6��v�/�4�=��97�?zu:���j>��4��Fgē�x�CF@io�1T�������*+��� �R7�4P)�����'�IP��Q B�V��R)�q,y�dNmaeD�i�|T[D��%~{~n��GD
/@����h�堼�w]B�xC[�nM�����8�ZVP��]�;�"���N��v��[r�$��B�d;��2\�lA�����7+�����\��`��b�0�4ړD� �'9�����c"C�!']�j|����J�W��
��	1�MH��)��k��,�k.N��z��$��=�#�O���F`�N��$��5�R����6�;qU<��E�k ���(�E�v��x��J	znVh曲n$<|�i�n9��A����[����H�
{5a�h_�h�D�#�?Zj`̐q���C%^@+�恥��,J�]��}V�O��z!��a;��"r�2�C<�t=�G��c��#�4�ɗQ�`�갟�g�)͉���uS�!�E�jFV�Ⱦ%��Q࠰d���A7�t/���4��R������iӱ_���k��Gܺ@��� ��/`N�4�~��;o���E���ʬ�
]��Q(�7>c�L�3!��r�}������$ .��>�_�z[.M��$S�g��kD�4�b�B�4�(�e4�G/�:�����:�s*]?�fU��%��1QT*%��1nU��2����B�c�$�L���8���P�jm8W�v�at����&�@njl�B}�X�WKv:�;5�����c��zC{�R]/��C�8�U�Bv��ID���1�Z�<��.��n�����Fd��V��� 
K<��Ǌ;��������?m��^s���X�1_>Pԁ5N=q�]o���np+�����وS�ޡ+�`7r�1�� 4e�Ό�dGh,6�Ti�O���?=�'_��oږ�_wY�'&L�a��,�-��8D��Ѻ(�a�8�?�V�c��#�b�MVE�O�T�dg�fiRl'�y�sl��*x�o�lVg[OF�^L"������k}�:���g��^����Br�K'E�����D�{5+"^/�m�� P"e��Z�W�4��^.ן����j��a~gb��|uI�5��z���sp���n�oTu��.�r�$�a�y:GU ��a[f4��#w���c�
ͼg�V(,S("�݃�n���z[�Y0�����A�YyN?gϩ��ᥰD�Tt��s*�.���L֪���J{�%0���q��/B��A�~+:U/~� M����5����)'/��j=���;gc�MW2&�ȏit�`�hǲ�
�.��k��A�z2ry��fB�Π��`!�fQ���R�F�)����d�O&㝮
&`)�Z���B}��X2�Xv:���7~xa�E;������l�NȵC{I>�p��cP�~Xo��%�aE��7�$@�W�%�=o�AhqX.4�����2e��w<>��|�Ga�A�����8����MYc�ޮ��|��YH$�S����uR<(3dk�8"n�a@c�G��f�����
�zH�����!}ah1a��lX�lP��0������]����:ZJ�64!����0�1`��ӆM�Ё�P��v�	N��~3d$�kߑ�ຼ�|�ٿ���S\�. �B��ϿI8��[0�e-�Y4_����tZ�:�j/��0��Ä�V�W^��-3�2���6�Zfjy�v7�p̴^��^�|!��	��eEĿ[غ�u�8`�M�.l�5S��l���j��j��e0y����4�\ђu㩦ñ��ǟ��N�:��o6AFuCpc`�6���LY'��&�(�D��7>F��[��r�8r�vRxH��f)38m��)�,M�]�æЃ�{!��}5�s�X^ܶK�?��9�l�U�A�e������6��{��Vv�?�L��,=�����4ё1��LU�5y�0t:7��~�������{p�)�`ؠ<����G����X�`qMߏ5�
W=l��p���̥�����_��wEĿC��O�o��l���A�YF�a��Ry!rM���dT\a���]��qd�(�`�����8�;	�/1�"vhfV�p��6n�ʖo�Fx��uU�^\�{�=��O�I16[�d��;ddx�;,l���뭊��x
=m�e"⮼�R��-���3�4����둼��j�rkHmm-P�p���;��;��4:�X7 M�s��mU�C���2�F�����У���z�Ǟ~�8k?�m2e�fAf�*t���O��R{��I?�g��/��!&ⳡ�L���w�V8q܀���|�I���I�-f�\�6�eAX��@W�e�4��̽�ٯaY9,�_��� ���栞�D�ۈh�dV�R5\�m2�b$�.��ޜ�z׼&Iǵ�g&�-$	�LO7i~�e��\cU<LD�>���ֶ2��-�X2��U�m����b�%ۮ?"��&�~��B��T���}�[�v�ֶ��r�HG3�"�S��8ix^��z��rr�d�?;��?5I�Xk���>;�:�z�:� �ir��Ь��#��6��ŕ���6�p�����އϼ4�]�x.�L��"����Z��}���:wXd�/,����ɏ��!�*����H����l̈́��(�!ι�v"��Z����hj�M��@�
�ˤ��kF5ݐ���L�M_}瓨d�[0J��s$��Q"�
uX2�ѡ��kh�u��p|��<�6.�h<6^8�W�l] N2��eHB���ￂ�8�a�D��!�U4.����|�
�����`t��L7�āE"&��DA�bxj�W��`���,X����]	��.�·��11h�p/m� �Y�Cg�i�މӎ��\
�K��B�)9�;f�Ï9�4���KHRڳ�U����+C��{�g�t��D?@�\�,�� ��/{��Đ#�|����f��D���D�:0� y2�c�Ob+�e�=��?i�)a
��T/&&Z*׏�g��/���W�����ZtO�Gχ1EC�;�b�k�L�(�h�.SmG�4�����u��B��l���"_B$����P�|�ѧ�r/�aTU��8g�y�v�Z������l�>�{W[���LE�d��X���4�T�����,�`�l�g����q�߇i����@K�t��BKe�u����P�]�R�����q�ܘCgl�ť��3��q?_%�эPD|٣y�5o��zc7K��K�&C�B7"�`�y��Bh�<���q�~A�
�&XeĊ��{���F!ÓϾ�&���eH65�г����]����f��p֝0�(,�n]�Ùs768���kq�X�i��=�y�/�W�x��/鶯[���,ݐU�I�����E=a��p�Bߧ��:��T��	��4Sֈ�zY��������/~��ǌ=օ�^�p�� t�D�y��»
�+K�R� J�X&����t��S_|��7�x���/ �.("�l�)���s���~��n�IPb�	�(��9<��k��/�B�a��oFģ:tK�7g�L�C���BAE�{<�zH�C#�MƟ����v�i���鬐q8e�<�܇5O�9Yf�5G�,���鬓Щ /�ƹ�g��ԗ�T=c��Vp�lGʇT«�i�72{؎�Q����9��-���Qhk-�W��Em�0s�^�1�h�����G�t,��ַh5�x�%���֛����MFoLuӑmC�+��q
������uZ��_�M�>}��x��^���UEŻ	j/;�)4��6ޣ_�=:"+�la
�
�n��с��x��\y�P�f���}�����bC��� �1 ��2U�K���� �0�<�t?�V1�J��a1HݲF>�r�F%"���ǌX�dΈ;�r�)ɒ�	�[U7�z���0Mq�&����̚b'g�葎uƏ�{ͯ��*>OG��ɡ���"Jq�0d��F\6�e�0�A����W��$���#z��Z`�M�\K��@�n��PXr��.�&�Y�|�8�H��տ�3�=6���[�×�T����/;Xux��6�`�z\���%�/g�ǹIP�>�������
����?�#�T���8�a��:z�76����悅��DXH�Zf'K&��%LC�j����)��5F[L�������`�ň��n`�vD�`�,j��UgLUgDHgm�B8�]������ Z,Ϡ��W>q�p��1XB��y�d6�2��4DF����'P��?p�yw������~͈C�3aY����M�l�-4â�9���#��L�L�4S����v��S���_�`!��|��Eė8Ck���l5�k]0B#r#�h�}�-�;��8脫����-߾	��CQ�����3��{:�>����e�	��-��F2���nˊ��L�W\��JW����G-����d�!�M�T�p1:����'㎉�C��������y��2��DcG�N�)c��L	��α+�mj=3pʤ�pAH$<����UC�b:Jh-	B����/B�� �ŏz3���Pm��P*�'�.U���)ȶLg�As4��ې$�k�t�A{l��ѧ��!��y�:
K��/<`�7ѿaR�n!�<$���6ɔS������ھT���Q�ͣ:%��7Z��96����m7��D�h$�9A�fR��4Y���>X�,�֛����G�2��l����i��br%S�|ei&�Փ$�ߞ}
���}F�O�g�&:2%L�d�'	qQ�&��v��T\���r��k�k���F8�:�@�Li�P�*g�z��O���`�Kn�y3���ڐɬ���5Dq
K�f6V��Lˑ�p�\�~~��~���y�������6�*�~�уI��hҤְ���2,� M���jΒ��ktC��A2 S#B��p�w��9_Aa�P��+�mC��yp�#��j��a����/o_�.b"�����k�Jt���L�i����Dl 5c�'��0B�M�K��lAO���=Hd�1[r)���jT��,������
���?k'��@O*�XJ�1G��08��k�V�cݵ�׿5�N�	κk#�ӆ�[�0�Й�mUS�LL��'�G����v
��~�g_y7�9t��G��N�`E����W���f�N���4�j��o0E*�6Cՙ*R�eJ�-���+��������/Ѭd5�K��w/��v��춽��cu�t2�L�^�,k�:T���tt���a¤��Jz#~ߓx��Y^R�I���2����X�5�lOԙ�Z_4�x��N�	�L�R���^Ͻ�1�?\f1ED"�aI�����FQ"ۘ٦��w��ڃ���O�E[7CI��Ɛ�w&8�iH�V�gV��+�I*���h}J���^��Q&�l5ϵ�|v0	7���� }W�M'��_�x��������L#ؖ#5%p>Mj!�K��&rd<zeT��t���/��βHpw[��]w	����N����n_�{�}���>�=U]uf֯���4����gق��^�`O�����4seE��"��,�0�Ǝ���tr�x�3�ѧ�d���9�r[gY���o}3��p�J�e�t�<��M?����/{����vQ���C&�ǚq���!�)��������m$��&��O;���'��\�DՒ�yR���Yx�M�`}�A�3*�$�M*�r���g<��Ʉ���f�����3�st���ӫ��ѳ
e76�V[H�l�p'qN���0d<���W��m�ՠ-z�֮Tu+�A/D[��x�~�-
6~�gs�+Q4�{�}r�Kw��U�hb[���O�w��l_�a���E�2�
AE����Ca 3�#	Á����
,��s��'`�� ����;���^4�YRG�R]��P�ހMMO�װG$�-��
�m�͵EX%�����d3܁���e���˳������$)��y��.�v��xߏq=��h6j�:�T>g~�wc\�%�� +Uu1��|��Ͳ�Ԕa3L�`LC�r`�(|��_2r1aFb���K�K��zPSP���C���T�B^�I4�f%���%aIr�3χ�a�� j�G�G�n�s�sP�;@XO�_GPT�\���3��?�hb��:��9�n/!��f+�Y�f\�y��T��M�D��9��
-��ʨ�.�F'.k7:"G،�l����ó3gau7�ℤ��&�Һ\2�L��� �"��"�:��6�sxO�<ޕ�K*S']�$�������T.Gz��0��s*s��gm��]���t�sߜ��R9����d�J���Y_�F���9	����^���J\�,��=o�D�$�������Uf�!O� �b�Sղ� 0Ǘ]�h+!������B?�4� w�;�S�g�V�5玎$�nBcw�$y/��l��M�>��N��ȍ����5����l}=��'0�'��f~<3�>�K��V����{��c�c|����1���#���`j���MLy������i�}p��7�&\~;�T�_�~Z|&�M�������#�.�E��r�%���	9�[4l��&������%���,�����`]���KP,k���-p�%��q������ �����:�����0�I��kj��1�h�))�g�K����#�'�c�2�`�ࡉ!���	��@O;T9Y���se��W������;Mk*��c�)���8R����c����3��o�ȠH+	|s��UF�ϻ]K��Ȭˬ�+�R��� ��4�{��v>��i�_�[��;!���9q�&�"%:��mJBۤ�:;�l�<���)	��c���ڔ��CY��b�i��i4E�[N�O�i�]$�Dy�T���n2r�\��S2� C?�Ʌ�/0��o7sX�
P}���:�������-�
�#���<F%��鳴�yy��4G�ݑ�5&n�6��cG�yz��mwz?>jG�X���EBq�U����~KJ��cM6��65��mF�N��#��--�r\�N�d ���ߊ�c�|d����]V��� D6�8a�����5Z
�l���"�IP�<���\��y��%/����'t�ʃ�%V`��7�-��*v�K���3�|��Dp24��a>�ε>�ُp�o��-�P���GN�_�i���&���-�cw)g/{��[���B�u���f�b��A��֔����Ũ[��O��?~�Ù9o`�}+]��k4J��jݜ��9Ӷ����#,E�5D:K���A�⿯���ݩ�����u`��<7��P�D�$j�(;HR��Uś�]��#�QЅ.p�'����.\E��_��O���p7Z��̎�L�m1��"���4�����%��I8wSAR�P��}��t~��(��?1��o��e��EVT����O�}����=n��<���%G�=\���/c��;�[��)h9��:��W�Ъ2톄����qt��6T9��|�J~���L���Yr�##��-0+b�ܑ���y��7���|V���z`��Fk�Jo/Ȧ����%q������<�k�'koBء�+,�OR�ٗ�7K�h����]�[��I��_$�e�z�$ӈt0e�\�od�@�p'�| ��^w˖���86�d�ȋ3��,&����fk|�+,�6q��M�p�(�Vtb�^�c����mF��8�(��4�C��4τ��0#�)�d�D�͆�/�6����?O���:���_ �Idp�D�%�h�x� ��U��i���2���;��;�4)�de|<l'Nj�JeHg���0�A̢���塺SQz��|���PFX����px20�#�Q�܌�.�>5���.g�ۛG9TW��զ��_`�=��oP�A�?�F�Eѵ�(��=us�s=��^��L�*?1L�D�S+����-d��b,�A�t��5�gY 9�Q�U�@P���!*!�C��Z�+J_���^)f���iN�� �@�~\ֹ_��a�@�^&�ؕ�e��a�r�T4j%*i��[:A��Z�'����6��kI~�	�Y�����dY�P%�w�:�T�t��?�bs8㽇���P,n������[k�?o���iZ�m�'��U��t��&��e��>���ӡ�Q��윁��9��1A��k�ȅ�"���{N�F2�xr޹$I���E-��e��9zg&
r���,��wr�Q�=�˅m�P�f�2��r���~.9��Պ�����ު'����`Ǣ�pMR#�B�!�DTa��H�'qa<Ì�	Q!!�����̫;�8����^�}�\R�[z��-�K飇bV��U�O���Y��.��|�����IV���}(1��̭�����m}=����^�X�m^������V|��
b��l�v�(_�'�� �����D�Qiv>�TRh�A_�_����E'�/#ߝ��~X2��/V�d��~yBS<��$< z���/uS(L!C�������IԎ��8���(,%߈�2���~�n�����)׫�(G�ʉ���!^Pb�IÏ����P�x�ιA6�6û
C8�V���>�w ��^0;�&�](��8�|�:\����C�����}�"���8Y�����y.�,JL��4i�49�:����Ռ�I&ti���}�s�i��b��9S3��qlsD�U7!N��!x�:�:�����1v�KĊM���DH��dn��ú�:M� �77#���ŋK�Q"�G��\������3Ug��t��.��\�%�՝�.athx�?7��?�\&�n��Xz����]8O �i����vCq��F�M������":㚿cj@��8���#��Ox�Q���E�~�5�� 7T	f���j��o��5K=ځ���cn*�1�?������z��G��]��j�e�R��bw��kEHY.��J(P�Q s��q��x���5;�������ߐ�ϸh}�qfK�H�DӯJ h0���i����Z(i��.6�_]7���r����9��J�"DNJR*J�X�	�_;S]��˰�$��������?'J�T>�:f�o<D5��A�G���~U���Q�J6�xާ8 �=�@��Dyȿh;��m�qJ����������v�I$`��*�d��5�/�/S�~��G���л�&5h$�e�nJ���	[K�Q�5�.�����3&�9 ���vD�*�`6;����r����D:ۢ0)E�B����N���j��x	�槐Ϊ_.�]]�:��K�G��R��ј�r=�.��K�6U����b�������޼?�T��|]�b��r��,sr}��nh@���ȗ����s�G�1!P%*		N��l%sm�6�؎�!�o�{K�ty�GȂ��KN�e�`T3{�����~Z� �v�ys6�l�E}M�pζ��L���#�3����UqlnG�o��s�Q����͉zź�r��!�e^� Y�{�;p��a�#*���D:�W�������-����5`�Q}Jl<�r"����xLVX;�nD�D��q�3ޟyVpߙ,�ݘ[/�w'Rt��(�u2�ue�3e5��5���� Fc�G<�[C�R��u�o3���>rb����E�%.i椊z]\�k�b��S��&M&x���x�|�}|����vr�c\����H�hRm7��S�H�(��K���w�"�1�%���E�y�x�*��GU��ő<|�_y>A�"��FJ�u$�%�'��F�]1<`��1���mBÿ���iK����y��&�j"w�Q}�]\�X�/iH�+��|Or��bpٸ�rk���7�'�����R��4:m����䤌݋�����]�ǖ|���p��b�GR\����ye��o7�V�1�9餔�z�s k�)�i�L�����M��_�!��&6a�8B��%S����}"m0U��o�M���[�@W��f�wD�ǂM���T˭囇���&<�le�?Q���}n��I�Րq0��ž˟����m+�՛<���v��3��f�n� G����c �Q�݀���BP�}��)�21��O?�R�D"Ol~��ͬ����d��:*�P�$P.b�p�q&(Imv�N����>[��۩���|x���K�yB�5n�Ǥ�{Ӵ0
�%�̗�J��i�A°K�)�(*�c�j��W������;]��EiQ��SH\���Ij�#����~�!��>����"�}/E�G4��<�F�J�I~���ڊ�T�1������)��,>�٣�"h�*�L֎R���X����ӗ#7�KI?�Y��5`��(e�g�f�������7\��@��,���"�eNB�R�Q �PUY}�O�γ��4�&Q%3ǭp�#2�2�R��!�u��?+:��:�-E$��wAC����p���jx0(���?vy0i�8 (��gg֬���h�j�a�:�X����on,ڵO7mD͆?��]ݶ�liX�ZHW4������2c�R#�hy,�3kHE~�n?�PH�u���me�fI֊JDD�����ǒ [C�J���m��?%l��F(�%�� �sAZ&υ��#�;K����t��Ʌx=D��ʪ �~/]�BQ� <�i�q��ӅR�5�9��g�7��ڙ���.�Z��2D  |��P�INL��zq�d��u��� �kA��[�G�i��2W\�oT��ьJ�F�n�qįty���D�=��ṔOt��K,°��&�`A�7�.�f�}�'t����͒�����7�%���[�.�?���l?���S	̰�uXc��ff�2����`$a�J*QEi}*��yv��3�̷��l�2�1�.��ey��7)2u!<���O+��,)�l�wM����*�o���z��7���8�C�G,�/K���J�^%�����/,�CO��je�Nf��׬K��>�������j9F��W�C��XO�at������>��O�2���9���w)�o�5��%9�Z��k�D�
��Ѭ>�qH��Erb����͉�����#R~=w&^7�$DY�=ĸ#9N痼�'�MPZd]BPo�r�6�PY2�R7���z�i-�(��4�$M�E�0�yn��4o,{��ʿ���x�`��B��?<�gt��VT��&.� /��N���hւuƦ���6�h����ȟ�8�n�$��s�[?c}��ߋ]��<�G�4x��c���%��j�R��Y<W�"�U�?�}��V���c�xbV$M�п���-�Ԥ��=.>t�h=��..w��8���(Sb�$��QUn�DN@R)(R�c��ؐr��#��>'3��O*�l�e��(��CB��u��~���5IdqjF�A��0��W���QMwq2<;�@\�d�1x%���T�?)!��vW��1&hd���v}E��w�F,�B<�i9���alɔT�!��h����i �PYi�FV1_���>�W��1��Z�ȇ�v�m/GvƮo.F�B,句���#��n�|SQ-C�Io(I��H��l��&��k���< M�#���8�@�>����!y�F�0�q���tz@0W�0	���<�F��ҫ�R�(�D�Fn!c5������O>�/}�Q����w*�c8	�-���&hB��f !�DpF*4˼�R���>�"G��(,������ϛB������ϳ3uj�ي���3q\���z�Hc<�&k*����$�,>��XlA�f�Z��e��i��1��|��`ہl�[P��d�+������d�Q8���}AD(J�c9��kVMO���p�P��~N @'�Dne�^�҇M�w"�1�*�>Z�Qwr���z�GX5M?N���.]h�!���F�$X�T�12v���cD��`!ƫ)i�C�������55���|>׻�w��f (c��cxԃ�G"��G�[#(�h�'A�~��h� l� �].iU����5]��l�O�����GH�n�βդ͜1���ꙺ�rdr��<�W�8m$�uZ��b��J�/��o���b� ����(P��\ �\�
���(�moR�#h��~��D��t�����^6d�-�OW�a����j�8"Y��+�6e��u��z�ƽ�}Ή}j�ԉ�Cs}Vya���=��>�������J�8����6�X�d�1�n�"���c��mt!Xxֳ�	C�`4�,)K��Zq��|�*�^�]��Z�WcA�0���}�<��XA�%hb4k��}�xֿF���*&q:��h<��Bd`�?ɀ���lc�#��H�I�e�
Y��L}1�f�Z�9\J�-U�/�������P=�Yn\�:����������*���M1c�y����Dޘ�������.!3��sz�<�?�˰y��ɲ�#��Hc�xU_! ��x�O�aX��M0�5�g4��3%���y'���EIa_ew����n2~T�d��,s��3Ж<���9u��3�K�Ғ��S,�F���
Yf�,��U]jwl=T�'�c2�IF �Ϯ$�>t`\-�A�IX��̢�aE*�X������ ww���g�:Y�N�� oH�*��$�Xm
��o(�k\M�H�i$\�"}Y�<�v�y���Zh���`:��X���sJ]�`�v�����B���������_[hB����^@."C��@�^�~S����upIT��)2�{2NNƯ���P��)D�5�PE��La7-�=`���+�7>�T�r�郱���'��al㑤#��!�[N�zނ2^>l���"�����n+��`�R.[5Q�)��#����H�Vs�BE�/�&e-��y�})jTq#�e@11{���g��R;bb{��^�sm~��*Y�|0�
L�0o�̉E��@hA��Ry�ڜQތW�`G�y�a�V��^����G�Nυ9OO{�
1.��L���[�(@��;C�Զ 2��nKKl2���5��T��1�ڒ����l�ǧ��WUH�h�u��{7�e��4;ޔ��j�z�=I�8;~�}���Rʯ�I7�$�3�{�0f]N{o��^&���r�0OlI�8�#v^�A��[y�����8O"���[T��o<u�P?�*	G-�g5-��՝�1�֦B����U�BE�n��91�� ��:�FFM�p���:W��<$M'��]"�F:�ЌJ���JFǕk�&��?��|��R��+Hy�~oGUOSQ�����o�H̃-i�Y�/�k�gx�?��M�k�"9���#�'{e�^��kvvR���gc
ݮ"��&n�)��
GU$�=h��]�9�EZ��ۓLA�fJ]HM�Er����B�/"pO
��B]�ֱMd�H�m�I&�^\l�-=ao��(���!��q���e���(<��l�B���
'�ٯ�[��H�E騷� �Mr�"�G9�!�s;lP�Ր9��,<E��_u�5��w����n�A�a�E��5�n�I�%pW�YA��KQ�۷�Ob��g|ʽ��:܈�)�\O��� ����P� �Q�R���s�x�+�*����
R�&���S������QH�XD(���]Mc��]����Ms)��_�f�������DH� �J�w{�x�7���fq�}vm�咱5n]�e�2�_���U�%�N�B",�7��|F;5��<��l^�M@.��n��ߜӃ,�ůFU���9ܞ�罯"C�7C5D�x[x�I���>tdd8H�_�m*M0�5F�k	�����!�Pt���m�A�4���IV[�O�W5�h��|{^���W,�#�l�'0>�A+��Q�)\���X��k/}+6[�w� ���xYMw��v��#*|��t��?���8SH�߽��L2ՠ����"O�L��G2&����c�Y�ܒ�dU`�؝�9ǵR�>y���a�ſ���␤��\�~� D8w�!��+�p��E9ߏ�FdGH �$�� ^s�'Q�yi{E�]6XT�EKD����b>�q%!-�8��=���Q6=���������S�xu8�x��c8>��r}��4s)������@*��͹��A����c�����ES5��16�5�pY.y?����V�\��4T�ӻ���`e\��o�� >�T#���O^��^�0�W�w߻���~��yq��9�����\8}|9�蛁���P�D2i�dMs_"e�b��S��g�ɞ�#;���~���n��|u�m��pt���۪*D���[mD�2˂(�R.�)��I�����n�{/�k�Eei����}<��p|�[�X���(-Q��j�;a�T�窉v����`�8��%v��U3�����F�*��V�QLP$+<H�%Ӎ5���+*�*J�tڝ�*�H�/D��\|���+�&`��� ��~!T�)���s�ܑ<矌�(r���*�mӧ�R/ƞ)��y*���|����k�|�p���|���>���I����E��*�����5cN��<i7p��g�F���QE�����'�Ӿ���Ţ����4��?T�2)��I��"�����~�YW�Z����u)��h�k�f�;0P�g$��-a�0r�$�E���a�$�D����By����3�'^�/�#�>$�>�uE�d��`Qc0l�׃o����:�q+�
�-�4�s�?��e�/0+ˉ�|V/�u�]6E�tRcy�Wv��1��<�d�m�Z�C��%]�Ɲ�����*4 �%��Z'yC�B�eW%j:Ɔ,����]mX�~�ʴ-�ց���a9l�dX͆�\�q���� ��g L�!W~�E�\�y��ѻ
��J�b�@�?���R|`a���o��Q2�9��,����>i�Lڬ���7^qPf1p&�K����.O�IC��J�9 ϑ@;�o*J��i���h���H��@!2ݢ�@�Y�Y��@����4�����ì���Xi���c��FNji���!�E��f��P�E��6C���!`�A�A�1� �n��\��%��#o���������a(��[�u\��+�t9��pv4��s?/�cI�?�'m��:��4�D-8�<C)+�<X�8���*t��U@�������[�,
VBJ�m�j�Ie���֟��O��E�����3���p�M�Х"U�h��t�mr��&׬Whd��}�>��*��㛆Y}�=�Љr
;P"��`�@�����S��fܗ��h��UwN#��k���M�2�a����i��i���yK�.Z)9�&.ж�$E {9'�`O �E0���B������Z����z�>�}=�������8�+���Б���:�8Y�3T�jЏ_L�%Ky�Խigʅ�P�Nԟ�����}�cJ��yO��������S�⼴
�^�� /$���4��k[Eq�㟹�k��Q�ȡSɔ�RF�����)�ۧ)��/Y�sU�(�$E�V��03]mX0�4D'���{��N�?�D��ul�U�R�4jV�yo{����u���j��kg���;��U{�B
Hy�3���_�ƤBBt֬%/C�f����/�ʢH���x��
Up��
���
�J��B:y@�څ�m��u�]5x7��CI�֋��	�Vb c�5��	P�=/��XJl�gI)�����j
|5R��0�ݖ��j�lfAA�r���%x� �%4��b��b��� 8M6��&�#.�1��S���*_A�.�y*���|=��G9���n��RB�q��Ui׿	�xṠ�L;���X��X�bvl�A�lwu�=�Q1?���r!��!���8M w��w4D7�N::�CVM�E	/`�0(f��@���$&�a�2��q��A�q3�O��([��A�B�C��S>�>�QKs=�0nO�'9�c;�8^��T�d��J;d���#�U�*"Dx#��4D&�l��i;�d�|�3��J�D�;��];)����5@�엪�t1�N�Ы\�ϐ+�GYO-���*�͓5���Z�~��C���w3%�b���68/�-����&��	'�����V�
T��9�cX�b9��7d����=��L�[
`N%B�A���J����-Ϩ�7t�L��e7�_l����p<"�J���������D�B�܏��F�$z��,/x"`��Άo慩�����2������&��׆�Jְ%M���{2��H�����7�=6��k9����o��(p'��	���)Ep�(�Z�:!>E�Ҩ��2���"20�Fᆳ:c��!�L3����ߚǩ�eL����2G�oT��ߏd�++���bw��'�����L�R�P�Hަ`���S���x��x��0��g@�y��h�ֈdK;�+\��E�_�[{P]���72c�գ,~v�cR�0KwcL��*U���~�r��̒@�֕m���",����Xsv�eW�boe�����g�C�/��W��ϣׯ�]��e�#0��l�+&w��;ĵ�����Ћ��4�%,=0�L����2�z��':����2��v�e�cd�z,����|᪬�~�~�ꅜ"i��c� �LtG��aco������3X6mX�d�_�F.��e����}�7�����1lػ�ǎ[�䤴�4��b����?��j�6Re*;.�,MG��O	D+2��k"�/��d��}�&�Y���4��+�ԀIL���*�4v��#>W!�lԶ_��b�����;#��\C�Mp+��+����ޑKF!ςT֜�ι
���#�F|��������J1��s9����?�ƶ*�Z/=b�$��Iq@�LF
�{��c2��Lh!)�@��iV�d�w���KC��c�j�����^u�iz�ݶ�&��ֻ/q������&(]q�Y����*`����H��es8�q��h�t��W��{���<�X��T�YY�lJ_��o;�@�����V�n{w��¬ǳ�=@m��b#���������,�oB�FZ�����C�Ԧ�i����k��@�/��xs��ez��(#�lޏ|�4cc���oq{Y�ru�~1u���yTV{�����PF-C9B*]��')��/L���k��HUe��	�G@�.)׫�ݪ�F��\$�J����$p6�ĺ��9ʆ
����Į�:r�mf�����פѱ������G��Zv��q0ӻ�����;����"M�x7ke�R[t�&k��3y�v<���(?^�`��\������iӻ�D��;��Xlj�:�����H[_Cɑ:D���?��S!�K��bx|�)_���� �}Mn�7|+��u
W'elA1�<3|���8E�8h n׭�������Q9�l[��D���ɡ!r���˘Om��y���޲S�#��Sl�� ���c�?���8��[�!�K�;��4r$ v;X���6��N�ëoZ�
g����z�4���l��4�o�t�lk����tn�)KHK�ɮ�,�j�bC<�)����p��1�֟�VDq�5aϣ$&�5�@�%��O�d�jî������$s}��{�n_��q�������@ό���TB�j��=�T,I�ߗ�W�;)�'z8�;�|����.n��φ���fJZ]d}_�./�n<? =,vS[Ӛ�Npk ~rV^3��*׮5J\��7��9������4��9����y��*ȡ�q7K�2Zr��6^75%R�Edi;D$km��FN�a�7ʪ�j������%;3o�3�X��s20=:d�`�T|L��|���j������xy�ᙶ@�*�S�����Y�`I��p�5�t�|An�qܴ�#� ���
Q��ҥ`T�(������E��~�o_xx���z[�ye0҃ESͨ�����u�P����,\�2r�AM]��\��c8K�f�����뇆��ہ����P%�R��I����">Y��44��ֵ�_觍��Ր�2����O(͓��ː �HК7�!b��:�V@�Y��Kc=��3ό�8��(��`E����[�C��b�,L���<��E�*�!"�N��H�0AY�u��y�~?�}#	�o+��z�E$!���%ÓX��ʨy4��~rc�ǔO,�d��3�h��'~�1�*_��|f�,w1�0�1�&3t��fÔN����&Uy�Zб������(��0%E����ݩ�s;}�Q�6&���g�9/�"f��u]�r9��U�_�^}��L
8(#���Z:��D���@ueT�C�+�\D�(MG�-¾��̄Z�$Y!ĉ]k�Q@����$��)/L�|w`����Nr���D�L�#�:����x=�/��ï�[Δ#���S���*�X|+t��ᅡ1S�Kq�+���ncr��y���f|�5r���/t�/�H�G?哺�\S^�%q���Z��2�K������]����5yQV{�(�߹�>�e��خy 1r�hݹB���r11s{C,h!�|��s8���J"���.:.$��K�Ʊ�����/��-w���"��4�y#^�C�5J����o�s�<��D�#�N�l��u5�qЄ���	a���lz):�(�m�ǅ�=Ea��R'#������j��V��Hı�ȓ�L/u��X�\�]��͠O���(�n�n��@��h����GV�B�)�Q�ȋf���@��*Tَ�Ekە*�����Ћ��k�>X��.mPhx����~W���3��
���Z��E ���8��y�W�A64('nJ��o��AP����)SV�؋��9���K	������O#jx�(�(�}�?>شł���v�*#�6��dK�i���F�r�e��#Y,�H�bO9�F&��Ԛ���-��.�Q>a��D���v��ʽO�\u��x����q����#<���~7��P���EZ��h�߄
կLˑnR�kFO��m�>R$�Eb����nef�jI���:�=�MUOw�v���e�KN��R��s�v��|���S��,����|�D��]}�������.�W�yX�(�EjnT\yK)q�-ʘA����*��l9�b�PƤ�"��2Fm���ژ)��b�K��SȢ=��?�A��!�i�����NJgr���Xk�h�6�� ��~�5�S�>jU����\%��8g��z'�46}U1H��-+���6Ǒ�m���D�j���JY���o! �UD��vG����(ܲ�E��&"���_��H��.{�j׭nk#V�������qx%���m�9�Ab,�@��&�`�y�=3�!H���.n�7F�u��s`T+��@#�I��]ӗ���pM�BgS
n��23�勭�J�M�G�h���\׊��}3���z��ԺB��_�N�@\ف.a��<��� /�(�>�0��[�����n�T�[�d����p����SDO�V�,���e��A~�F�^S�s�bw��,�MGF���[������ಕ<e���=jTJ����[/Z=J��*|�Ǿ�6�ř�l�~��2�i�t4���q�z�a��@ }��oBf��LWe�ҟQ4(y�O������?RG�/D�:�_듏����*Y�Y*�~�=\���� -h1rP=ĵҦR�Ԑ��sxdf���_���_/��w:Riu� �w�G/�����hP9vvΟ�6G$�,�y�Z~��0�O2i��6GU����܄	������<E��V;�{����I��~;x�'�I9<�	q@L[��lt��+U[J$�O;U��^h�NĈ%"�t�����3h�Xp�w�q�y�%�6��t���w�
�~,Z��&�a����]p �21���f�TE0����;�|�EG��ɵq�Q�BM�ᠬT��ޫFG��c.���` 3G�ʧ�� ��ܢ�,C�y�!�7En�	ؗ��P%0��Rf���Mh8��Z��cޖ&����9)�6u¯������򹲟������;Ef�VN��e�=@oKq蚎�n`I0-'Y���*�sɪ�uapyl^�3+gw���F�؏و&[�pG�g@uF�����O��*�E���F�i��wo��4�i��Z�w�&��/��`G<7�\6W�TR9��%!���>�!C�6�xF�D���o��n��rS�+�F�$��e�Y��J�Pu�yn��(`�KrbC�&P�ãD� ����G���M���_�b�ߢ�
���^"a��p�vr�m���(��*9E�?а>�L�ϡ�V�n� ۾�ah0L
��*�ɣ��Q�u$( S�%Z?BEr
e��c&�3P�-��󵏞q�W�(�c�Mɑ��屶�Q�l#���B !/#�_�pb����4h�j�� ��;9׽���Eo�hw�J�qF޶��^u�qO�]����BbrkN��پ�R�S3��2IN�dB5��~_���!���,ل���ĕF=4�P�DßZ�be�ކ�H�ee��l�7�2 �E��UL�3���n�pȁ]Q-`np⦈q���"���r�?zEiԃ��h`b�13�u;(�?���,�bNv�z>��0��IF���G�7��I<�Yd�S�w��ya��y�*_D��1���XfYf�1B䕌��́��'�)��Z\	g�iA���Q�bT걇�n��0�T������;�Q��'Ȯhn
G@�h�#�@��A��c��ovto|R�0_�m螀���5A�H��o��|�UH\` f@�_�^:�E"�ͱ�[  ��2v']��p3���]� J��G�i����۞O�>>��$4��3�xai,R:���J������\Z�;oy�\#10I5�R��Vu;ԋ��u��]��k#>�������������e*f����%���'�e�}k�n�bh�D�\�0���=QD���Y D�Ñ�w�v��W j�{;�!R��Vp��u�C�}�ҞA<@ �����I�z�V�=^&�&k�Ү(sݻ���"a��������j~���T��)�ڐ�aA�)�s͈���?�,YQ��pWd��z�S�V*���t*>�Jd�Ӳ��Y��}�k
�}K?�4���:��
���uN���a4F���m�Ttwn��������^�Q�P%���R�lEP�>�b0�c�$�������n"��W�ۥC�/h�g���Io׺/�G�6�7`N,e�M��K���`*���7�X��AHP�<�,��ہ����M���$g������6}Hː��!|C� �VɃ	�4[�t[X�����ϋ3��s,��셲1����D����%��P5f�>M�R���.��E0��ft�G����M��?V�������*GU�Yf�*����=v>��W���e7����l/�_�)'���; w���"c�t�8e^��)4��,삂�[��c��_����A{
Z�I��f�N�P��L� � 9=�KR��
+��v�l��0T7��8^踩{q�~{�<�v�c*=ݟB�RTL� �H5 ��4�v8�ɝ�j��p�f���A���z��QK��C�� �����*ve`�������ˡ�8��]�g��hV��E{����CY�p��\O��kZ����%�a$��1���������^�'?�X�B���ުhExP�aE�@�v�Z�)����7�5�!���W�"�p�V|��c�"w�����nU��ғL.�)�-�F)#�wz�Aw5 ��QA1<c
�ÈAQ��Z��g���򜦽���`I�R��YH\z�uʐp�xo�T�\NCM���U"�ʢ�%[:��oX���f'�b���go�+ڢm��n�4vc7��ƶ��I�Nc['hl��>9щ�r߻������{r���q���TB�,��W�0Cw����d{�)`�3��6�#k�F^]_3��R������T�#_��������N��[*�H�H\KDצ��/a����-qR*���9����ԉ
t�^��S <_�uF�y�=�u;p��C����c��i{x�N�2����6$��D��H�ջ��yPR�������w�WJ����ʍ-Ψ�ԻI��*>�'َ�/���](8���ߡ���[���D��P�X�ɲ�g�Y��]��t�W"G�Q�>�2a��>�k���ϭѮ�]ӿ��$���P�{�R]Q�A���n�#�}��^j1�R軯��a�Lam�bƲ�a���.�|�'X�ق(Ep"�a$��~��G[��g��w���c�NM�R�����B?X�`���: `����-��Jl+�Z'���H�97�uȥw�d�4t4E��1%:�F!�#Q�&z�����F4n�店4^���]�����i
&;��w��W##��B� Om^�M�
gM���`m,9��������� �� ��[P+�"�|�#�7�3kG�VD߄�M�޽o��vG�1�ʃ�9�{"�^�_|�)�g���Y���m���7��:� �I��?@]�
ԏ����T:|u:�TS������R��lQ�o����OH���v5
��T���kK�`��������K��j%�T���\S�r��Q��'ƫ��'H'�0q�J�_h6�Ve\qp�Ig���r=��Y�.���H������Yk�t�����F���bZ}-xf���0�U���*+�2_&R(��Zpd�pF�UKy,�����J�m��ת�i���X��b�Z�ߦ����~҈�EI�EG���יFlc��*���^4A�#z�j��tn6����ϐ�����&w�?�w�����+GR�F͟��O�76amD��U�7�S��YQ�gM����[�Q�k�Ϊ�׻�x-3,���Jg��rM<`����ᓪ��]���<Z�O���R�O/�mǋ�'�F�9�8_ٺ�n�m�t~ܼa�CM���q�ڟM���c2K�8ѳF?:?���5O�_������!�������W"�u��J�;�+��Y��v����rL�q����{oi��؂���N�s������ub!�"@:�UW���o|�G���C9���Rf��[��?�.'�eA�_���&���wEPa塋���]�PCm|�R�nOԯ,�VO S��/�.t�f`�?�1�7��P�DY�dz�$�:_�,��p���~G�o�e����:c��^	/�ö�������'���و��Ozp����Խ�!	`��l��:n�(�?�Kd�H���&�=��G���p��

�/34���_�i�h�����<�|l�^�r�+W��m3)gIH�TW��f�tD��,6�D�xۊ��gNS���bU��M�Y�������qWD�/jY��c�%(��BiH�cz\�I�;A�_6dL�o�Ƥh�4��p�|��j썀K`Ǫ�.C�	]zHiD۷l�gc	���̉�;�2i������o�ے��8��:�����"�v�8^8��v93�6�A*BuF�h�5ڒ�	0/����/,��V���g�� �U�B�+2�P�LX墥pa�2��)�̢U�7�� ���%&�_a^U��!�g�A;�Baִ�١(Ez|�5!��GN�ͬC*j��["��5:�i�c�=�J�e�]�X��"-�ϛ~#�)WVH��ڊK��H���� �݇ ��71A�}rRAgiI�[��,�.	E��w �T����*���L)����7���9��A��'v�O����ѧR��BS��>�:���@=�!ve�5^�2���SƚC���-�7�m��T�t�+h���A��U4�B"͂�r�Q����<:}=� A�H�������SR�����Wd·Z�<�K8/4F�'�>��"!�������$*ݣ��ز��������,��p��5�;���������~�,"\s�~� b�c��P0�$�+��ܬ>���؎�f��E�E=A�I�x�2r�?��.�������ZP������,�Bxi�짯M�BA�o�0��2ȁ$�k��� Vb�Fɋ-W�#�¶@��S���?�B[
u����UU+��~!�%Z(�	����
]5�zڂ�U�@;F�Q��9���&���U��b�v����&im���6]��r�a{�
��:�*R͝���9m)&m���"աo��Z���Ԭ{�:����$)�CA�	� R�J����9h��;������*`�'�4Uw�dV�b�@���C[�a�9�7`d?�1���0[��}1t��X��k"_�U�M]
�$Q�F�3���:It������d�28mK0����u��d���VcVJ�K������k��[��~�H��'l��Rl�����BF�H.b�J�V�����n��wH:s)W-��c%���V%�ma�*�;5@�$���yEI�k�|��(B��|�mUȤ:~7*���<؝��!�� ��_��::Q$�>di�;1,=}���W��	?��C׍_qN�s��P�L����	-���2��`n�W����)�\�=���!��_H�~�ȥ�<^��#S�8`����G�n?��%?c�����f�@�͘�o�'oɪ��i�v�n�[���)uw�����0�й9�z�t/3|��ى���ٽ��!M%o��r2��g�����:�53`F�o����*uiO��_9p��@�o{l6����p(OD:pJ��<�7Y[?��v�hL�v�[��l�#��gF�k��249�ƃ��z��
����@�I�@�֝�AԤ�_��~� ���?�%��H��V�p�����/8p��1lM�c�H��1�̴� ���>^v�v�lk���=o�g�[�ƙU�g@��!q;խ�qܛ���]7S!�:.�{�F	�|�UF�����S�����W}г�����*��ᑮS�R�2
a���GS^'%i�w�5w����[�tԡ�B��f�����o��
�%�@EBa�U�X�b��}��Ͻ���h[P�F˶�0�E]c��-(�vgo�B�M�㶆(�~��g��E�n�����(���4待��붽M��7J)eq)���l���z�-80��AF�^sP��;J�!�s��h���� ,��waD�������GBvJ�֨�V������ao$I��ܴ��ޞ���P']��	� ��n��Ǡp��kj��)	~����~�(@OO��!\���@�*���H�����Q�B����;+E:�l�����wo��y�ԣ19��{�FX��f�a����X�r���.WiGbAA|�8��E|{���MZ����C��!�)��Ԩ2KV��y�����Q2E�6䓜E��7���n�ݷ�;�I���;n
�Ǔ�z�qz
��z�H{e\�n��|�9���7O�+��8���/I7璌'Z7=&>ezy��1�3!��}I�����ܦ�g��7�6F3��ȱ�$s7�GS�����PB悄笠�_��F�&n��&F����1�3���r��C<��l�چ�1�7qDD��[�[`�z�t��B��WQ4�eo�G)�w(
>��ĂR;��}9mL�mʒ	3l��h9|��G�^q�(U���]!q{� y����l�Ċ?d�����Z�� S	�3�����	4�����MZ���z�� ��r
�1n�7���j��F�J�Mu�w�$���76��!칀��(��[Ȍ匶X*�Ķ��N����I{�r���*��+�L&GO懎m	m�X�	甯\f��Gqìf���	�nd�������9�F��"�q$p\��y��s-}�fm0s��Ҍ���[)���nO�l�G����j��fp/�����		��!i���`U�f1��¢�VN+�v���6��n�˞g����.;��b�^:���Y91�3�ܙ��'Q���C���a��W���D��_Բ@�� ��j$�\�lo���$9Ů���Y���I�i��PQ5	z��,�����2���e��&�ʝ1����R7(��������7i��1�B�p!o��� jE�H��3K�r�����ړw���= Ki{��7��q}�ypq�����z�)�hX�UG�ɩVt[�Yk-��ҚZe��^�7��x3�!j�� �΢���Z�Lt�����[KL�b�ƕY3P�����nyܩ�)j^v9/���Z!X���5	t����뾶�����H����$���u���BXQ�yi9���F xъ�x�|����}ݾCQlvU;'�'�R�͈/ג�_�M�5fȦ�0Z�\_K� ��^�r7�g� �ٛJ�{��J�g��V���ragl��k�&��@Q���F������Ǵ1�v�*��"��ٺɨ�VsF����ߝ�>�����h��jz/1��*z{K�TNQ4�_QLj�Mݪ��2���W�:T%\��b�|#�0�R(x[����=^~1Ձ��i���� a��sy�]����]�٥CZ�2/�Ƶ?#V���ø��5 ��;1EIbG�I�--�g䣞� �)=��d-Zi�۩�A�{s��t�l���#�=�6��\���ZE��DY�b��Ә�~���
��IY�n�Qn��L����6���]b~ٍN ��w�3����pB!�
-�����+~��F��\�Ao��%��*+��љ���(�9�*ʽ)+d��U�Y��L�l�	;ߒ#�z�x��.��g�'��6-K#�Ud?�|D�M��c��n�����KipFw���-)�a�'�+�%�f���ڍT� O+2C^r�ƽW��=���5��u�6^�hS���?�z���o��ҹ��G}�
����J�NP���NB�U�.ӯ���~?�?YL�|=P�ll�IE�i�hc��nU�+y�T>�����?7�F~Yu?[Z�� f��N�
>�j
?���)¹��ؽ6ρMe%['/��CS��J8������Y��݇�-�r��3h���pr��[s�+��}�8n���@cR*h:�:#yB`�d�}w��RI������7Qmm��#�Mh<�9��� �yF��]q�8�Io���# #���dÒ3-2��Kʺ7��Ɓ;�7���0�i�w$"
���O)��	r��O��g����F�ˍ�&��5I��q�@�]�TsU�=z"PTR���[?�ki1>�h�e�}��0���]���6B�='�2t��*���z{���@�һ]0u�?$��@���&_��ggy����X�2���wR� u��63�HA�A&�gQ����gF֨�N�o�M��'�
����$������Y��W~�Lv�IK��a��$J<�_�h;�ow?=H8�2Yu�qcVz8���dX�vcx��2o���[fE^��O���J"]����ha���k�����[܈d%�^�v�|3a�H�i��R��P�P�;�)�����<�;���r�Y������s޸o<�#��)
��EVh�x<}��^�I���.������2#������3
S�4�d���в����7ME7���i!=�F��e���V*gF�z��?ʙ�un����ڍ�uwb��=��=C��*߇>������}��u��ݿ��E�}��ۃ)����}��q��I�Y���Ƽ����yoߊre��K�Ͱ�Z��-Q�=xg[^g��?������k�Z����g��8	(�5�e[�J�����<aV���a�q��;q׺Ք��
}�����9h�-�����wGV�d� �x���h�0YN�6��:� ��>-�� �)@uh��QQIK�ݗ:ҋɷ�2�����9��R]HGu���E�ފi���3#S��{&�
����`%�1�vQ5��|���/���e��X�Ԛ� O)�bLY>�*��Z��΁������Cq�� L�?�gR��5-���p��ZC����}P���SV9��/l&���ę����� �{٤�Y[�~0 ���7n҅$��>�)X`�ě��D���y��k�ݒ��8S���w����m��e;�=�QX�0���e�GT�2<&�/����ܸ%��+X����!U��3��t��ES�a(���vK�QK�	����FO�:�!ΜΔ�`�/`�����ǫ�3 <����G �K�;����BIM_y�ؙ�5�sn����s�ēt�Cߜcls��6���H��|��z�\Kr,�Do�B6}�Dd������q��S��He9kb-�S<{�ޤ�4���z��K+��	ʼ�H��c���o��H����H!l����iYϞ��I�$+�c�3-�����l���0��1d>����C�N籀�J����%����孖@q4�r7~v��b	14���)����	�����έj�j���ꐢ>��J~ȡo^����`d����'��Q!�t-���������Kvk�<9���z|�!M:�Dt��|�S�gv��s�6�\�u�}���V��&��dq��Az4>��Ӡ���f/+��Ok���䑪l��s`q�)�z&G\ C����t`���!�P�۟��Dx���_��r��nJf,��o]H�&"s�e����`��f�kd���s���Uj�(��Z��ߕ��q�ԟC��D��#�Dъ�Q��	[����M�j{��Ћ�����=3��D�����^4uE'�G����a��As���R6#J¯M�nv�fY%���<
�CIBr����MM�%o�^�*�g�j^��@%�$���=s���(̏�����ҫ���$�ͳ�N�:F�R�@/���X*���}?`̪�d�#ޭCS�YB�+��r�Q���(jN�x��E�&?듼N��.�i���U�%~c(n�~�֓��Z��-�q�xm�VN��jb%��D]WZ�_�%��D5`J�)��l�b|"�p�a�k4uS�$c�0�BY]�/k�n
�O-n�?�kkM�HaS �9j��6Ӭ�n��hT�COb(mk�.�s
Q"!j#��D����P�k��Ma�Su��<�U\�3 I8p�3�����1������ԉ�EK�Ê�!,�.q�؊��x&�k��������O�ꨬ�.u-m���}�{a�M>>c#��+#,5XӅ_�RC��^!DB��w��H�6+QŬ��0RU�����B�b��V[��UޙOJP�t%m����+j����݋��c���~�>�D,/�2o��rfƖa���$LN���⇺���A0@H�i1�M'��d�CD���;�Y��}qa�E5 ,5�ܺF:�'���1���M@�"i���i�UN<3�ښ�`KQ�Q��ܭϧG,f��}H����ըc3��8ѐ�n ���сH?�e��I)��8�d(+�5,��ː;��K�Se�Ma�鮤���"+�F/�*�������S��KA�n}!���͆��rP�/r������0��|�g�aH��資(��;��g��}Wbp�����Q�5�>:��:64�#��Ӵg�;e��T_9_N�W}��&l��˔�����2�5�1邥���?��Rsje|��X�Yǒ���x�ʉ��>��:^ˏ$i;K��Z1�b���c���(���Ed�~,�u?$M�8J6!sgj�א�w����D0$�f:.A��g�-��_K�􏵠�R!GbH���Y��:Ӄ����
�f�a*-U���\�����P�}bd���.�K�=�.������|��PV�N'��3Uq=}hiՐ;���Nt�]ծ���|.�G����i� �i``��׶#!�N����0C���fYs�g�V�B7���Ê��"�h�����n��->.t�)Do�����o�4P�-�-��r�.����t5*P��X���c�T�,ؓ6I���X�����Y�,F�jr�Ҙ�*���yh�ʁ���^8�?N����P��յ�lKUX?=`�б�l/��`z��u0!����Y�۔�x���-6S������%&���y�P+?ڂ}���(q�+�-(�K��y�`s֙!f|1v5��/U0%�tV����J 1�W}M��.�����|@�"T�@�	�sf���e4��lc�Wɪ�Z���B4���zMa]�1�'Pd�n@�?�9�P�i�@�5�Az$^�;�/3V�-�V|H`8�RF�Gs��)3[���S!�����oľ~��0������t״IeA�s3�+{R��K���4�N��|\ϗ���6�� ��%dU<_��7� y;����0n�}��7���,I��
M/ߠ)5Ɓ=W�M�k����4�DQ������$�a-�R�����%i�7r���=���3UZ��>����-b�$��o%I��7�k�	��l��7�㋟}3a�5�h��.^�1!u$���EV�<�뙘�հ'�.��D$��㌙�]~n��M�4��=����v���[�Z���<�Nʓ��qe��ݻ�M��=��nw9X���D����<θ���au)��/&��6�$��a8gE�5��H��������ȕ�ҽ��#��EWQP�	�W�t{���)r��ex;�q�\�N��9���1�<���*a��B�w�I�����QC�,�]�>>z���$�.�a�=w��� #�����{b���S�5a\��:oqK�����'�un��;lu��s��,����%�GTԊx����]:D{;h)=�]1��8|��d׼���v�W�PȜq���͕bkO���.�9��Sk�'�����-����LK�	R՟�|�˭+")��Dj���4��06��È9m�'�I-aiv}.�����y⣞U��/�y��~��,�n��;4����bF��~��{:lPU�e+�������4��T Ё��0eUIc���J���:��:������9r���$ ������S\�[��]	�#;�)F����O�18D;<��^�#�5�]ŝBxE0�b��x��!$�5̟ ��CS����҉�d�1�/���{��Ǚ\m�K�ռ����0*ʬ������~�!'uvV:�L��(��e\�f�Ԡ޽嗚,w��ڏ���d��':qV��E���r�)!'F�eO���9�B�տ�i{�_�dH����tx��i�X�}�&h�,�9�yM����P�%+���x���Q��#����Կ�G&�ݎG�*}���]�,kώ7����w.���A�	M�7�����;��#���ԓh~̿���Gv�par�/ ���.�&�v�cv�����|uƃpL��
��r���t��H}��'q$$�..Gn�@܎�
�,�j����⚑��Rq�ա���xp���(!�ch��U>�8��!�Fu{�=��%�J�u��Q��u��~�I��L;�Ȳ�t$����b�N֐$��nW�_#J��(��t'�ġHt�_�w�Z;M󊃰���* �J�#��#z	9��39��i?Z�~�7����κ�8ϓ��E$e�g�_�-n2O��ir"�Й>�d���I�}����{e���h�ʸ#��!<�<���.���Ɛe�H"��+ۃ��QP�����I~���m&�pLm��i L�aF�
q�E��5��zx�}���E���+�_�3�?��w����(uM�$�쿯��v͹�]��({��&G��̬��U������:����.g��g%��.-u�mM��^Ъ�|?� *�:��R.w�]�cc��v�	_�C@��  ^c���A>��|ud1:d��ߎ�V��ztzt�ﵙ!h��7!�}%��'�����K�g�v�vv�:d2�`�j)����Gwt�L�Si���՝�פ��f�i�ͭ��o��q۹�a���ۿ�e��RY�f�Ñwe��G̀�����*�ֲ�u��8����g`i�`V�0}<��h���<�Dާ�"�*ن�\��oS===䎿���Ì^vq�\6�$3Y,�S������X�ޤ���$M6�~�]��0$�Bq�U���pq�%�y3_V;�쉬��8�`��i���Ym�F�r����˓X�C^�-�PW9֊,V��֭�'>gh���GRy�jaH���)ʴE w�Hl��Dx'�G�FόZ$�j���h��6�"�4"�i��?j�0&*!|�X�P�`N2�EZ?� :�[L��7'��M봪5#���6&*ϙ\�12�%'$C���12]���ek�������#��;L�h?��Ǝڧ�,�K��ܢ��Y���J�O�O>S��^�&D��=���J�D��z����x��l��usCW��`$ݕn��0̮�V�E�ו"���Pj����]�,���{&A/�[ϛ����ݾX������o���%�s�%�6���b�TL,jU�_����X{����8o��k�i�$u���X��)T}Y.�楒�&���T�F�F]l�BRFb�V��?�V�e�c�c��T0rx7��r\��}%mR����B�E0^Mͻ$���p�����䑘�U���,�k���!{^��&��`(ʮ�PѮ�m7��s��ws�9
>ҁ��B�]1�"��g���\�e.8��с��\���b4ȇ��ETζ8�xF=�ݟ��Oe�#I
����.S��=�s�џ��l���ɶ���N�X1YbN�3w"��ּ�n���������ޑ�����Y?_��l�v��������blWӈt]�z�v8L�Q<���f��pI����"'��c�y��Y�E�1f`4��O�ޭhHfJ�fjE+��{��W����B�AK^�RƷ�{_wVA�,���Qz��l�#^�G���A|G�A���o ����	ӂ���'�ܭ�i�?��H�t��^���yv��s��k <�	m(��|A�ІEj�-�6�����4�{��%-&����}��j�פ�Nܾ0A�*jq��D��P�:�L��q�(��|yK��a����uw�6��г��j���ܫ�(^�/���З��z�A�d������+İ��AD緷���wB���8���E[8j����=�7�%�9zo�����G��A\^�S����%�]_v���/5/4���4�Eϫ�"�g|�l�[ k@v�Y��(��o���M���T��D�����Qrs�+y�t��U��ہ�lHH�vo���]���~qp]s]I�.V�I59���|!A�J����pd᧨9^a�L��&��������:ǝٞ�A��JD& ��/'�H`�5�٠
=TT�u��s�xx|�wÝ#NiKc��}���'�.�ͳ0/>��{���Y���wե���0ssc�{�漙#3���V����b�9��Q���]e`d��%�2���u�gq�n��M���1�<�Tq���O�z��M�f=�z?��mE�x�g84�Hnč��$7/v|��|�6z�Kk�}Ox@�8��)�F�Mbyl���P��و� ���+��%m�J��}	s�P3�\�d?�J�Id��z��|��g=1�A-6|-׶����C{�S>˩���h�U�&���S� ����a�J��ݝ��	�d��J��x�����8)F�K�H��#�u��u����)._��r�X��ƫ�(�k�Z�9��+N��4�x��xX��O��	t;I=��X�7Ub���3�����?�ޯZ�V����a���p>g5��*ؿ:
E�1z�r���t��}��7��T=r>��o7J���/Z�P1;x~�j*�1�.�{[2T!͸� U�V��Yҗ��7X`�5�Y]�n�~�2�.0FȈ��Ld^\�:`����-e�f|���2�r�У�7�^�8zA+
��"l�)FkG[<��՝r؈� &�>w8�'���N�&I�\�'�"N����w����a�/g֤��	V����߄����:K[1�X�O䚛T���fe�5&>����@+#Bᯐ-R�<���a������l�<��¹�b��0�,�ӱ�)�!nҥB6>3�{:S@�Ka��b�R?�Vۋ�ન�P�%ъJ�N�Ba��ܑ�`0RS�d�W�^��m��/�ӕ���6�0�N ,�]��UXz1�D��6V῜d��I���Z|�l���o!���r��{�r����9��O��]Lu9�#M�Ia�|}��:��vVpI_-?���7À��dGɖ�8�%g�}O����Yn�v�PՅ�?�\Q���vr@~4�|�dD^�A�ݍ���Kbf�kצ�7���k�+�ǻ��{��a>8]�ވ ��ѯ�xf��^��%%�HΈ2�JyіNi�ރ��r�[`<C��6����չ�WAfq����`brN/c��W�Oh�;�!��Ǜٱ��.p�#�6ப��_'��f����tg���|�>e��e����l�Ua�?v�����&ݬk��j��,��Пl��!����s���k�_J|15 �X	����'�g�q��Q�ٝ�3
�cp���W�̳�M��,�;ϛ�����Ղ�i��&8�1Ǭ�w�6��r}�D~J�Y<,C^�V(�\�B(���C�����	2גkO�9�\�Z�=1�<3��S��݈�q���5�q�VK�i�66[�[�ـR_���y.�X���������$��R�?�yz�z7\6�5�eJ7x� p����>Q�:�fM�2lw��E��#h���.��������a�3;��S�R��O���I��}�Y�d��@L���F���*�+���G���?`��������pCz��zO�|&�F�x�9�����~]��nx�C6"4s�YB�v:q�������+�<CER����m����ƳV[:u��{�Uǝ�'r���'���C�:Oqn�R�Pn�hS�e*�L�(��W�c0hΔ�@��\�;4��A�m�y}�W(�I�X?��wS�
��b��:�AZQ=<g��e=�i��Z8t���f��G:����a��2#�S��`2�� Gku�n�I�9��P�>~0	����:3��Pp�D3��~�2b.n�4%������뙑T��[��B�2�/n2^��5�1��]n�O�����]�������e���=a�"��d�\d�~��^ ���+]�'��gnJ#���+�gg��	�6�&
(I�	j
��¯��]Ugk����U��hD�m*�!�D.aٙm�NG[y�z�!X�_H����������oh��7kf��־S  ��ul{��X�b��F~Š��y
(Rc�`�7c�	���LGk�����]^�&�]Ϳx6���$<F{��l�crynE�;u���G_/ӌR03��Ǭ>�ށ�|���j�;���<�y�ng�[=3������y��bz������:5�1�g����['�H�+3@q��G���u�s�4�)��(��P��}�E�m,&/��ы4�[�t�f�pa��Eh��rOǹh0�vhg�{7��"]M���@V��ϕ�ܓQ����VѦIƒHloa-Q����7L�g�rr�q_=`{�-�P��;��iǹ�z��ݖ���C]v�����`h�&���j*����]�'Y�Z��f���.�V����t����)b\�ǚ��s��ݐ�'g�W�b8� V�i,lY+�fxi���S�o��m�K�_*��fv$�Q�,�%F��Z����6��&:]K\yz����|\�Go,kޭ��~��%ˠ���ٲ��*֚[�WϖQ�Dihr��BqeLѝ�Ϳ�)�zv�yu��t�=V�#
4x)��l��(���
Z�nB�.��X0�/ :Q���[;GH|���F&�/{���p���-�M��.>f.�.�^|/���ۂq�+��xr�RQ�ߡ�Ճ�$Vb=۴�s	;����S:-$&p���|��Q�H,]W�혱�Q�l�Mq<���#~���x� ����U�ɇčpoF�0��%0`����)�ʙr�y��Mc�t���#����xe��z>ƈ׮�����{�>An{�j2�Ӿ�䝗�@�&K	g��"�'�?�E*H���l��wx��J:<-v��Taa�CgN��[�[k))Q�&1	t��|'�^^��W�&Ȥ�X�IGxh~z�\���F���F"b��aZM��o����(fOg�Gj�GH��rj�D[�A�5���V�'ɱ�Iǀƚ{Q�ؔ<�Xr���u���T���%ܪ#k����C?��Hx&��Ṩp�F=k��v�pD2��� 0�����Ϫ��!��)W���%޽5�T$�Y��#d{���^��`~��&@�LÇ��9��4�	Xy�^���u^�Ѽ��~�#��N@�s��L���O ����ӊ���j"�TO5��E�c���/\%m���,x��7%8s*J���r�z�B�y�����t��M��L�݈M�}�%nu&v�,��q\b�1�p<|��<�`��>��5�n�M}<��}d\9ر|��0ii���^ӝ��P��tn_!���KS�
���{\/�Z}��e':��4	Ȃۍ��S܋�0#�b^&������C�ݦ�����8�z%x�M[�2N�D��� ��6±���%�r����|����LPu	-�]/|������H�s�&�m��H �T���Ű��C���n^�J����T����g�J<���s�)`�jR4�fY~Ci��
$�o����\�i
 �/�--\���[��䶡�cS��ڦ)S��{|]��K��yplf�ْA���zҴ����q_�1MRI�j�|{�Ұ�����/�H�V���-?�&��h��XC��(;yڪ� � �͆W���9٬{-����C�0���؝��9���l"Mj������F(��� �1n&��^�Zn���R���~�ȬC�W\���<fG����xO�KUC�đ*Gl�b�#yu.O*��5=�����Nj�Q���i/䮭ֿ���u&#�Z��n���b�'Z��M��턦(�u.�X��e��_o�!�b�wߘ������՘D�(kT���e�
� �n4��TL�_=?Xe)"x���S�wQ�w24�ּRF�x���% ��ena0¿�V�<�;Q���'���v�!��r�?Vj4;���;�,�w>#��(С<r;�'T�KVO_rз&��A�P9W��lW7RAy@���q,�<�A��m�#C�+�Mz����qDԯ�X�̰�cB��uZ��[䣷o<�;���#N�.��凨5�}*��M����H��"%8�%4V�B��S��ϯ�n/1���qD�Q��b�T�-^~�\yD��&;lpb��@��;cQJ��aN��bU/U3gU���ry�}s�"����	m��KG������﫹k�ܛ^E8��$~h����~�!k/��������kom�9�.GɸINp�-����6�7�$>����-��"K`�#( ��<f	|D������g��\/(v�-�acZ��_1�/Y5����Ǌ 񱒣f�f\����9��i'�[��i~��xu�i��;�x��r���ն+� ��n80��':�#�6��7'�� �4W�Gfc�59sdu[$��),ԗ�4f�����"���<)����aTC~=E-�}O(����Ѝ5.
�����8�z�*�aJX<�s��2�1��$#i�D.M�~Ka��eV�t1!BO�nL�g��<�h�o\j�t`�d�' 7m�,o�V7}�����_f��/�(�й��@ aQ���S���i�3�k�D���,ʅ�������7�Em�1���z��O�𻱉����/���]7���;`%>/�ɚ#�����P�<	��^��CH�~�T"�#u��{O{�7�JQ ,��u���m?p߯�=]Y��ً���q`?/�ub�"j��<��C>C� 9�vl�`#j�r�ȍ����KR�Txk��z�E5.ƭ��)F�V���T�	X��N��/��iW��6<��Cy��p̝�8��_��v~�*��0����o���Q~���`��x��\���Ovm�}��9�.���*v�ɦ�{�%�@29m���"]�s:��R�J��j�¶���&����������5i�j�9�D��Ic�u�������a��p9ic�� ?���w��G�p炊G�L����2wD��F�AO�UQ������� 1W����!�:[�J�x8/��Y��y����	�]z�%��5&P�ƚB�n�8_�5[aK9�nSY(�&ݤ�!WI���8�����Q7����I�@��+��8�M����H�~�����ʸ���m��N�a E��C�kh�n����k�B���_�������4��{����>V�"�f������ewja-W��e=呇+թju�٥WQ���"x�*_�p�}%T.���m�xM�L`�S2�AP���T�HYF��+�r��W.�N�����VU�������I�����׫�p!��s-쇆-�D�Q�`���e�{u���a��~��5vNۃH�T�� ��+ɆeA|\���� iW-���.L���+�?0�΋����τq�!0Z���(ێ��_��}��Ą�.��>�H?�G��?��\�?�H�Tp�o.��ݨ���^�'��-�����3&E����:2���6����1��Q���?�nS�N{�C>0fX0�P��`I�P�����698]��ji�Y�G�jÐ��?���ق#I�\3��I�����م��@�� �Ǝ�w���<(�r;��MF��/2�PF W�kq����9��ɘj��s#�7��'.Y�:a��/�:������3d�r�x۰嘺���c�| :��V�h"�*�ZhQch����/�*�(��~�Y��'�~����]h�ڹ�z5n_��������k�IIރ@٣Sׄ�������=j�D�U���^��ǌ]ol���{��E�_�ܯ����������@����k=�CH��k&�%X[Ӧ~$�-��`�G�Q����n	�\�]o)��S�\d��O�4ҫf��I�0��i¬P���f?������ :�v��Y�⡷>�ڸڨ��b���$�91�c/�+lI 9������;�4�86Xs��#v&/�C�B�1��׬#	͞�i��s�rbk��W�'�5@��[֤�}k��C�����΋^M#r�c���}.��D��;U:^� ���3�]I��-��f�m��^���/��3Ó�M�d�ܟ��޲Q�f���^b�!�q����{}A��� �������Cϥ['��PV_$b�����g+�3iw?�G;&��!!"���^� �iv���r��N����gK�/��җ�˻��|���޻���(�*U6q�󉚜��3VXs��@	$Gt$�K�6�H�#��iذ�б�e�>؝\c�9��G��bh�!�1&������$�+�d��ZU_
/���@O7��d�&�n(1|�{ëRP~�>�ӳ�afJ�C�t��:<FtF}��+�7����np^�yV�o����:IF�`���gk��N��6%���a�磩8���q���`�`_;��S
qUI^oc��?��l|����	Iw���{.?���f��M��N�~�`��2<d��ɶ��0�B�se�^ɹKPW����B��z9�v�o���b�C�ow��;��Q
y5�v[�(yx~b���`p��ZQ���!��Ev)����7Ϥ�{I,��Ovd�$�z���2 2]Ƴ��l�/~Z�ȝ���?��]�c�O*�כ�&ŐG��*���Y�9)����-j���|m;�.d}��`��r��]j�i����n����atN��E��oPo�'��X��jUhf��,*x��������
xʅ�P�z���t�y�VQ[���	�|�Y�J���\�ѓ���Y����MW�t$��o�X��{]t�)!0�����}��-���48Y����۬Y2f�9 ����Zet�ǸYܶ����ɞ1���0�tX�p�uO.��^-�).
��ؘwE���I�G>�^䝩IY��.wjE�zO���i�[�)r�V[>n�s�C���p3|e$��=n�*����#E	��l���NluY�n��å����ERYʙ���������1� ��do�]8�rWH:�i{�̶���[���@7�?Cć�p?D��}U�K|wCbQC�)�2��R^��`u�d�����u�D�J6��w�	�;��=��B�tw�t@��_}�奏�%��}�����������[�)6}� "p��`���J����8ꥴ��J���.4�0j�g��mA�=�r�->�:��Ӌ�������_=Q*�w�\A������G%���$=�'�mzu�ݕ��J�g�50�+�p]\�����м㰰��N��;��Y�Ë��t�˨��\���ڎ�"�1ٯ8��x�0]���	�t���t�3������xkF�(K'��9OI����ըß����2�ۯ�qɝ�J�١yF?��	�Ȱ�l�[��<�����7k���P-�;�8ITxZCL?-�p�M�ےT���/���Y�%��>FNt�ɤA7��d>CҊ���П����Z�"��?X�ٛ�r�ȖN��/@4�q:�탦�֙CS�C>����|���%���9��G�q�{KV�f�if�f�Z���Z����ehɊH�ʸ�މ�z����}[F���_��S~�@��ļџ=���	"���Ԙ+1���;?"�����:ΰ��n��f��
	�{0�5�.P�����6ٯKx_��}���Ȱ/(�d�mNe����Q3x��n�dc d���mqlu�¨l���R5r�C�I�~p����%�-ב�U��.�{d�Q�g�ݶu/�f(���~[S��2B��Vi˥�����҉#�/\�w�X�O�:���D�ѵ�ea@Ҿ�II�1(�c:���VY�Bpkm~(v_ߗ6���%����#��u3f�+�c�>�t-dZ@>}��2��E��k�(��T5C�(��j��F�A��5 ����U���BV�.�����x���Wn;�Cϥ;��O���w�}u���_	8��`'
�ى��DX�N�$:���i��@�+%	LdOӦ'��0D�,f>����9{�~'�:�w�O��_��RBA2TYdO���L�����6i>;B~��J���	È/~�$jS�"�k�H�M�9�
.������!�
���9@�"�V�lǼ��7����>M��Mj_xb-�^����1>�׿����W����=[����4�&�UҚ�畦�F|�$�������)��c�7��C�U�E�^���I$iPn>}�{ے}��z@<�u�A���q��)
!�=��M���7$)�O�sw�Ň�ࢺS�Y�Ƚ�o�K��9�~��
�:zn�L��B��-�<�v�sf��okktcS���ĥz+���Cֶ͜[�PXu�UF�i2rOYUš����%ո?L�f���Ŧ�jx�o�[ۚ��������hv<.O5a?>�[`�Ω�!�]x���?�֍� O"ZUWGlkk۸���n��jV�԰=�n����h[2���}ߤ�m�&�>z�ζp�v��!�C*�tLy�5�ҩ��W�DTQ��ȃ�;��:��vr���c��3 ���wcO��a6���+L
��S��׸�����B5�칵��BO���3]ݫ\%0~�-��nl��{�t9�����+���z��e➥k� ����6П��qf�Sک�����mï�Iм��}';pH����&�N�S�-h��}�!�B��AȔ��R�ǂ��~����	6^섳�Fm�2M��ducU[��f�s{���-U�ir8<��^by����u�w�D��#����=�e��5?�_
S20��v�.��T���Q~���?�t�����N��4�*`qm�a����Y{���O���z̑��\渲7^��Z����U+904F쾱fœa����vn�`[)�"��I�s�{=�4���C7��PP��U���s����h�Ŵ~�p�
�+��s͎�ަ)�>�1��0�8M�{�T]ǰfT�o�o�m�.���u����Zz��֖|i�M�?�N�`�%k�']ѭ	���c���C�����9�ա�\,��vTX�G��jeA�ƙ�F !�������}^�.�~9e�:�!�q�W�)q-�*@Y���]�����<m8���U.o�#�q}
�e���!�s�����2�R�9��?��>�o�#s�}�.��2ތ�3z���{�zJ��p���H�*����3��ڱC''�׸����%��[_@b91P�kB����ȱYX�{��[J/Rj��>]�(��lA��g�&Z,�S�'j�ĺ�z�qa������/>0��.�?w ��$��_�O���\��Hŧ�ch"��8BL=��|o%p���d(�U(�u�i��uz�|�̻��څ19��qr��wB*��0��T���S���a�f���+��� ��yM����πm��Fw����<�pq��^y����ܾ�_c@P;����.��p�o��f;�T�;��*&ϟK��Q߲�FGE�������vJ|�=�-�f?�}�T��fN��0" VV�:��k|���%�3��s9�g��V1��?�i�ΗU� ge�q`�)��ԁ�=�t���9��|h����2��'Jx΅15�g"�t�:zz���uB1�q|F%Hk.�i��[QY�Vɘ��f�5�x�����9��ǧ��2�0�HN$g�Q��y�32�z�&��y"i8��Kf^��[��U��z�id��ch&v_�AƹO��:5��ַ���X��P$��#�9⨿��G�	�\qi�4��!�Y[� g"��>�c��'��u
�W|�#%��jE��e��<-���m;E?�qN��;�@3d�L�q)��'x�n���W[s�,kxp����k���9ѥ�|&�Ȏ1�V�6K:t�d;l������Ǔ�F�p���<��9:�灞��LS����r�	�@*����޴�o����L4�[�?'���e�H��,jg��f�x;���$���&��8F���2� �j+[hW=c�:��!����ӯs�v���F#�ʧ��Ĥr5�<TM&́�0������+)Xݷ�"�y-�9��8`L��=ߣ����sy���1�55�j?�6�.	�@�q��#��_�6�Xm��n�4�������P::|�(��%'��Wt���'��Z��L���G�@~W��W�
h0�.c��?�b�7��EE��~g^Rص�ɝG� TG6/�4TzB�iEГ�nb�FU�C˶pҜ�#�'W �Ⱦ����g���1 �(�t�`a�5Z`��"J�Y)�LR�����4�x�«�F���I�\m���fU��SwI����`�x:'�.�]��O�$���`���K(te�&G�LA�^�#�s)$��u^���;��b�Yl��jh�����C��8Ơ�D�.HԶ?�>�XI�T�xuY�����������d4�����Ϸ��:+��Ы+�����Yҡ�"x���g+<�u���;�A�vGC�/�[~��3M4�$�ZO]j}��x�G
xշ��M�q�Ax�����nF�kxT��s�N�%���ڶ)��1#5��Rί�wX3�C���٠���!�F8e�Ҧ����uN����|q|�fG��E2`=����X)�b��Y{^�؃���-�Νj�9c?�颪�j�jYh[�J|�����N@f���y,=!�˳�S\� ��ű�{y�sP��_�
����e."2BX��0!:����F���u�¬o,+�\�r�
�CYfHI�_�,N�Ǧ���,�5ۗ�~B]�r,Xhr^7���Ӳ౪���j=���A��p=��7�:/�t��wz.~y���A���C#�::��9z���n��z5��ٛ�w�%M��w�C��D��g|?)�y����ƴD��3$�CO���P�7�;d�mR�^��@�F����TV)���.A�}���w�1��o�S�ŽUC+�g�v��y=�>>�R�򁦭�i�0h��>�E�j�S�7�7�4����W��̒P�Z1�>�TLı?Y��MwL��˻����n�]���*��l����'�_�f@ ./���������Y��$2����'�'�������Gt��L��;�<�%�<|��KoD��:�@���J�Q|@Ra�ct�3�!4*>��~1���6�O�����V��XP:�������ǔ"�1.4 ���@1�ϗ������'��n�TV.�e;&��7/2���#t�N���!U��.vZ��0���Yo�}Y��\|)ܒwb"Y2%��%n�,�C��B�\ݾ���W�K��f��:�"���ӛm�Y�h����(�Ѱ�2��Jyc��N���k6@�N.x�}B�Ϝ���\eCd32�H	Vh�2Ӹu6P�&ۍ��Xw]�7�T��|(U���Q6Rg葤 ���̈́�VYDU����ٽ�n�� �Ҫ�'�0iB��Pt�)*��[�=Џ�lҵh��7�gJ'����U$:X;O�$Y�}�_�S�g����~���|?Ps��UP0@�I��l�?{�v�V{�ٔ�p�,�	��tj��D�T� �I��$e��a��K��,bI0A^c�:[�a��v�j������w�V:��g�p��n0n<Ǚ�t (@������hTR�H���$���)J�K6Q!bU�Ui"�����o�U�~o]�.ȰE��èZ�v<[r���vxE�Y2�a��fk�MU�j��70�:�j�F����6p��	�n~>%�骹dp�Q�`ֶ�=W�t=�>��о�	Çd�OM֝��ʎl_���9�i(5:�c�FI�`��F#���x]��(��v�<��c��OHhE�#6�G�#�yr2 و��������8�W�Џ�8���<�w�j����Jd�>���m_~DZ�����C����2D�|Q��P_�^�c1�t2��|��C���C�� I
|�Z�@ΰ�a��B�L�`�6�x��a��rV�CE�Bd�D��
���[�SpR������%��*���(�]��I��3Wf�@ue��Y:�"��
#�)|�ۂ׭�Z�ЀB#~����ʕ�`\�&��e�-�� �l%1�E�̄�y�<hhA����ҭ�/z����x��ZT؆����7ń���n��$QA���'��4Y�p��f��QV~d��z����L�B�NԏK�+j���k�<V����gwa�鳨�	f����I�����+eL)���f��C�?�YK�j������R����g�e����)����Ğ�j�bY����E>�����9��`�-Jm�,�������m�]����+᣹�����Q�����4��?W�*�Yh���+>��뎻8�"���x	 i�����c)x�5ܘ��V�&m� _<yҴ�l�գ)���0�U���A
�F�NT0���s�|�����Kx��g2����6ĸ&]�S0O����T�j롉�;��@2�P:�^[���~����d��W\�m|Ҡ!����bki�ib����C5Ӌ��
Z@�Z�NP������o�f����0��6ϘxsR&�~����0���	��r�!YhRGZ���@1=�,�v�D�'����v$�Z�^2�a�e-HE���c��(���ϝd�+}�B{?�`�]iXO�*'+�KjVW�HZ�ձ��d�Q�q;)r�mq��y]/���Cy�7a1�V�E�:1����4c�����(�z���X��L& 8̶��z挃��U@q�]ҞoH�6��r@�\��"�i��2̢A)�G����"Zrr	���$�fO`g�j'�����B���YA 5i��y$�'��/�qQ�Brj΁ƾ���(���ʲ�W9Aގ6���)�GHrM�/4�Č�����lw����KJ+�<{�u�޼���Hه��eb`D������48N
2Dr9z�bWf9f@��e���lG�uņ��pf�	(��]LyTZ	mH'��]6�I)�m^���G�۱G�gְ}=��[%(ە�¢�;��dW�9a��.�I�i^�� �?9�ۙ��ǋW�_���q�"C�XA�9 F[�P�������f�** 
�a�7o�I"rY����K��2D=�¿�߱ͮ�޷���c�տ�G�W��r2*���S(G�^��:��av�ڋp&��=�;�,Q\�!g�+oUa�b��.wT�yb|�|ݿ*yn����B�*�Y�Rـ6��5��^��O�اb���h�.�T6A)�ץ?_��
�Z����������MW��мܹ̚(*�X���r�aE��u��5�6��n8����L2�V'c��N���|�|�y�I+B�2�P�Y�A��Rf���6��[kq�x��j��1�9r��L-p�iX�/t]Ϡ5}$}���(��♯���]�7��C��w�*
u��5Ѫ��Ap��+!<���#���r�=]�L�}��a���]��9{V���q{/0��;Q��tg�%�-�J$L��$V|^�� 7�N\�F�*ʙq���p^|��� �~�s�r�YqX|���@}�M�M`�\|E��������럩�c�_� ?�,�Ӳ����[�%�Rvj���,�^�-�p��ߴAC{w�)ݯ�Q+p<�u�G,/7�jz�1+���a_�W{z �l��i?��Wy�;�;@[:*RQ��UK�|�'+_VaS�b��N=I΢4쩼�G��j�R�Z0�1D-�ϣ�K/^�q�{�L��Q��- �H.=7:�OYD�_�gJ婢YeW�t$i!-���ijk�X���V�J�V_�� �x���hk�%A�U�� ,�9������F�ˡ��6�Ԍl�������x&4<E�hG�@A\�$g�E��Զ��9Q����||$]ޏ�wѫ�/����`_���߲�,�^�O�m7�׶�}O ;�=� c��Bx��@q��v/ݢ��(�8T=ݢq]Y]�s�$����������&|Wヾ!���)�e�^���e�D�x"mb�t�d�܇����s
��͋$8���ʏ+��G.]�U񌃧7Cƌ��d�@��Aʠ�O�)E��gnu'>w�ۏyr�
�b>Wx<봺���"
o5�"�ׁ�j�:�q�>�W�&O�ۀ��$����җ�k�	����P����uq}�@��wj��i��vg}F&��<7�M���'�-W�V,ZW-��+GbԶ`R �� G���K���4���c�N��OŤ�]����B�*u�$Q�C@=��:2�<�xFhD~��J;{���[,���)�jV����Nw������3��oHj�pZ��6>��Q��j��<�S@����T\�e:LT�%H� ��șN�8��eП�i��S���f��=�cWcW�O��B@F�%�a�x��yd��(YBUf ��A�#�[�Mxi�f�!�$�ݱ)�B5#�7� v�/[��b��<-9k`�G�ju|�J���˒���m�򍠆1,蔧{�!��ǝ���x�72.�8�ֆZ"��6�8,���k�g'B��un%��a�k�!�tQj�6>����`�T����"x��b2�z�FP <x�;���f�?��s�9-��ȸ�K�&�&ռk� ��t5WvB�����L���R�vZ0�p��s>���4�O����+�AjM���������������YG�S�[��U0��3��Č��^���?@�N���ZN1�>5<z�p��n�ޕ%�j�V�(�rcD�oۨx�����w��.b�/�yϰs>����|_��x[yR��9\�j~��2�. �ĲF^��n�-m-c3���D+�35�{J��'/L�3m�lw�<1��S���Q'���q�1X�>$-6��m�y�4���=��T���z��S�ڸ[�E�����qh�[�g�8L /��=�iU���m�U1@��hɢŔP��:ܔ���"fw(�ךȵ�R�ٺ�]W�0rBz~N@�
��s
-��������p�����3��:���V�AO	c��
�B��rw��]�F=fj�W+AӸ�6���r���x��`a���25{�:ޟ�jB1vT]���1)�7��\	b���z=���C�:a��9\�b�ti-hK���y�,
��83a��z�Z�o|�m��p!��~-��`�.��;�N'K;].j�&��
��'2�}���M�|�#Ud~�0��J,O��[�)m��H����j����������J���gT���e��7��K	s̤ȷ�����̭�.��U�p�h��hU`3�.T���l��.�Q	��f^�}a2߶
�_� 6�M'l��[�8�":�,����ib����q=��4Z�&�w�M7�`�j���u�#J#t
I*שEϺ�(8�sO�?���(��"�~}�AB�3!���t.�1�e�K�����~���T���-Z���
�����\2G#*GJV�k��+�%��&@�.o5�?tbF�WaZ���PY�t��`��']d������o�;�c����X��@?�igG�Z��]�֗5�P����L���%�͈���w�B�t�k���סs��oT��?#U6���e�ֱ(5�7�,L�n(�?N2H�����b덢I=8"��S����i&��$0�a����G: ��4�q�޲}�:�E+xwF��k�xynh����1��ʃ�#�iz���#����d���P�~G�+c%f3��D����J�R�6�$����0����9nV^G�be������6�oVK�Y�1�9yo���N[��z]�����8�-o�<��n��� ����L�U��������u�����|��x��X�h�P�X��o��q��cV��E�(я�ʊ�������Gb#��ǲ�����Q(!��.�۩wp�X��L�VnF`Y����,Ay����ay5�;�{�O%�*R���&�e=�����A��Qd�;�۹iĭ�M�og��A�I�{�Y�
�K᭨$������!�+�w�RzﳴS^hu��T}�0�m�����3�ʴ�æ�ƚt��TN�y4�������G��-Jl��:~��K���vr����+�9{z
F�<�v��7�n��5���I�����5A�{RfF�Z�Ё`�����ϋ�������_`��2�A����|t�c�.�m�,K=k�%Ź^ؗ���5X>Ja�^JQ��D�����i43:5����G��%�aZU��0��xҐ��kʫE�^�KE��=���닺6�"�E���a�T�Ή91���! $5/�������ž�Ԗ`�����L�L��l��>ި�W=�ޣd��>����zҝ�4E`ˇ�*צ5O��p5Ǒ�T��xSH�,��qّ<<�xY��cu��Z�m�C~x�r�ɦ3t�ESȒ�쁊��#47PͩR�)����MPI�
�l��_B���k#L�3����L�N��Ж�'D�w�܊BZ��.$�9-uk5x<��#o�Z<<ۦ�K�L�62Wt\�Y=/����$aӪx�~���W���")�b���W`it�Vi,�3�������c�e3�?g�Jm�]�g��$����UBy�?�J����� ߺ�j"���T��E��v�m�1����0�#���%��o�ɫ��.��+)p4����~���h�f:S`�4�h.x}Vw ��b��@?�x�ZUV����,�u�H���
Й�����]u�EXyC�� ޽a���[7����<�x�%z�r���S=��uu�N(B�L��[��8�D�5�-x����6��d��67$�?�No������3�E�ɟ��nFBj�p�i�jzz��ۅt��O\u޺�
c�z�y�Y��Ņ�|�蕄�%fݎ8ќQ��/hq��?���o:H��cc�1sd�6�li�/X�e8���J�܉/���g���J���}����^�׸l!�;�v�O�'�>S
�J
�>���s~��@d�.�֛�w��D�$&d��e̪�����FR�0Aⵉp�}y��݊��ˮӉa7�}#QA����ǟ�mm�E��w� ��n��m>�v���.��[����(q���xLqK�l����J.y<�c��D�˺�[ܬxm��z�A�W&:����h��3�VJ�H=���1�F�P_�ӹ��`1��y�c�'�M��;����M$�5���c
�
A\����!�_Otڦ�uu�Hp��&"�����vƔ���o
����9�C��bUj��,u�՗�_W� �~,�^�Ee��t� {hS�� �P�e�or\�S>�O�K�ڷ6��s�c�zX䪇�5�d0���L��ѥZ�.$K�QS�5p�R��o��M�n�VlipL�i�bTJ�nT���`�d5�y���[P=\�ʼ��7/@�\�����%�"���/�:Lw��A9�l\*�-2=8o�ϙ���:&k^�j�3X8������C����Ee[J�	i��J���S������;\{�Ó2���?+�1�0y�
k���%��Jh��0�'�&"q��^���,�\8n�G�Gw�F�]��?q��z���t�n�w�P[�0�1�z�b���|}��ݏt��ۥ�>zN�R���\��o�-:~�ۚEuBRb�<�5ጥY�G
�aU6�&��&-�����d	��*�w��Iz�t޾K1zKR�-y���~LS�D�!�����1c}br��A��;]!6 Q�%,�yh&��CU��x0,&���"ҁ`/UJ�� :K��˨��C�O��f�O��Es.:��N
�s˓��%�''L���w0eا�6�-�3&�v7�f��ݞ�hW~�A8{�r�s��B��ӛu�x�j١�z�݀�C����>e<N����D}�oqpy$çJQ�
�i �&S+t?n+i"�j�!�����'�r!��Wh��#���)�V��B���5 ��͔%�{r���M��6кW#Q�͇�����r�(�M�?/YV#�dq��7�[3-
$����W��DwV35�s�(~3�4����aՏK��nױ�kG�{���A����_俜{��j\��'=�#R�,�yF�(2���<���dā;CH1%�5�{/� e��y禶
y����4KN45��Z���S�2��P�/��r�D���vx.�3#||��5>��6���O[�M� .���>u�>5�O:ЂI �CZx�N�C�|�F�lB�RN̚�p��!����n�nct=f�.����Y�����A�/~��$=D��OU<W+���	m�r����Bă߀�cL�{n�c�>���`2����Y�"�ܿn��ݣ������i	_<I�{��CPa,�piX���͢�U�ƚ�qr�de��@����Mdh������?@6�Ekn��M�	/	��;���Q8r����tj�k�`�7g��8�yeA�q��>���Nح"�?<U;�\����:��B_�F�gKj�"W��g��рE�N	�]��'�ǟ�k'g6����_)�W_����l�����]�q�����C���Vءoa6�q*k!!څI�I�Â�B�;�������$�ϐ��ʉk���������o������9a�7C6��k"��e�G���sr�򷻊�	D<%o�@qg��$��H{�c~WIwM9T���~��Dz�;1,N�yZ84�F��{��cT�sf5�j�4w+=hRc������ՊŌ�/z�4?#���j����3�GK�r$X�I ��7��492ϸ���N�prxLK���9��u�����֮u��Vf3솟����rcDH��6y��\[��܃>�ǳ�W��ܩG)&�F}H����5�M�b���k	?���M�G'b5|��$G��||�+,��n^�Z��Q.^��w��]ս���������%˳h�<"�_�;����D<u���ƙ�C�bd(��}\�x[�ن���\�p���ܫA�0��w�
���hE%�h�ZK�EǰJ�~O�ć��U�5ql��>�@ �K�S�}���'���c��$�1�k�¾G:v���Ob�����P�5Θ~�u�T���x����Z;^�l%�s��#������Sោ;�`h����fzP=@?}�R�	�Uy��cƣ!j�ʻyd�)���{�C����F1����oɇZ�N�iE]�=�<(��/��˺��0���h�qt�3m��p)��w�g�e�>f�']Y$T�M"6��>|���*Dl��A��b�#��۸�nc�T�u�=J�$ݵ�ʌ���Bv�XT/�l,膜�:)y^j��=2��yhG�޶N�����lVa�����_�pE[:�_�B�t
�#L�6i�w
V��^h}�j��3+��Ni$��	ݒg(h!��B��}�3֦��4N7�vY�ͯW�|/���ʪ�~�)�∣΢����i�)�T�	*���_ӆW5���E���CF�K�)��^��L�b�r�-�}�>��N��d�94�ěnq���\4|�y��</�ܓ]I����@8�my�d�J�3��FY)���T,�ڢ;��W��7����_�g����	8w��v��w��Cms�0i��)�V�Z����K?��כ~Y�t��"]�l��;���J�!�q�f�O�R�r��ϯ��\z����~(8���:и����)B,��?�=<~�a�x�h�����p�p�c8�O<�m2t��,o��|��Wd�(w\��Gl����Loqe��m���E����P���������N�t�Lp���,"�����R�	��p�cY����ì���X�S˥M���a��zD��m�V�S�v�	O��/�(�_].� ��hnD���\LPgK���H[���W�V�����8�T���?'o�l�Q}�EƷ�: ��T������.i�~�t�#��(�%!����A4|���Vϩ
�:g�=cK(�~��������Q)<���n]_����	ó�/��!��YA#iN��~��V�<�'*3/6C
��Es`�C�Ŏ��\��ẔO꼭8KNsy�@��w�l���t��l�����i�����T�@A��ś�"�bQ%t/WG�=i�@݃�_�g-���vYu:��l�F7�rY]
�r�m�];Ï�d |^k�s�M%�Up�����G��6�nB7Uc��P��;_����������`O�Bt�me���ňF?�D��!UJF��7u�%�s���8Z�Nۡ��a���m����F�ÚTJ66,�F]� �N��$&�����m�Y]�b��]DOU�ҘyW��� �'�1��L0�%�Eǟ��h��?=�=d�M��%*1�X�3C���]�Y7ʝ��}?bH�n��Q���~����hӵO���U$?��m��%F/:����ʠ�3����4ܰ{����Ȳ��(f�'B� }�L��sʈҩ1�9/�i�-���6oe��{˽Ak��v��ۃ&��R��@��]X�zA�c��ݹ������`O�鷵,ێ����7DLpk}N�������ξ�Q�G�ֱ�p��R~��}��Ү��ʞ�5*C5�,J1��$p\�vu��G��4�iU�M�I��)�͍=�����n�X��^��<��\XHeHE�z�ob�1��Q�lC> �!Y�N��RE�����
ɆnB����*IcO\��-����ͱ2	�[j��4�:���®#G#A���^O|�ѼV��R�s���f���8�y�W��7�<ϗ�pI��V��kj"c�ʇ/۝���IH��>� �����vn�ɺ�/��d�|��ӽ�b��Ƈ�>�ї������d?�b�vG�r���'�:���Wl�����Ոsz�:���GM��45���{o��<W�
�cm!��R��=;�xoo����(T��w�Ç�����&6@��U��3gx��tm��b��ŷ�XE=��pY6%5�o?�}�h-�e�B=m��:��:Ũ�% �,��OJ�Z����{Y&��@W��{��2����O-��%Q���F���_�v)�\o���'���*]_Z���,�pv~f��X#�e�t�oT�:�:3�3'k�!�C��"1B=l�6�,���崦X��={���y���ٮ^EO�P5/Ud"���ZhI�fz�n���q�Ļ�<1������陵�z=Ӭ�thm����~�RY�ܶFq��u#����~Z3��vh�̓�x`��P���Ty;Y�S�r9���~����[��ۗc���¸8�ԧo�H�k���S8ʯC�c�<��gޙ�OH�Zp���[���0߳��!��N>e��G����h^�w�Qu����n�Ű$����J��;���}Vݗ>^\7W� �T��R�J╽q��/���V��O��3B��
�8j�xa���F���� �$�$/�x�W m��\>P(�	��4���ǳ�|�g�P�ֲt6���ٜ���.����P���a�	����6��T	}���K�b�%�Y\���婫�C��A���#*��O^9�6+����s�n=rzQ�ϼ}�_�o~�r�F��f�D;��:G�q�8���-���\W>�)�"��R%�"s>�D+wa��F�d���R�n�I"�Oi�N1f���?����@�M�y��v��M�񶆰 ��H��k�h�0n�����$�}ck��N��ox����am�˺Y�\L���t�=W~e��%��}u�JaS��E'o�c�p�	K�X^��� ���}�/\�Z�m�9�X�-�^a�uce��M�g�f�����|C(��s{o�'���5��LY�b*4q�l�?��2 ʮ��
Hw��tK�� ݝJ7,��t��tw�twww-��������<w�83s��e�rȉ���z��h��(��]��hQ������6�H?�=�G�$#��BW���н��hU�9�:7�w� �����y]q}5����>G�����5����g3�q�.�%[1��H玩z����Jum���Se��lp���J�F����0`����!�5���(�Xv����?8� �D�#�Y{���f��[i��W�����Z0Z6?��~� 2;ұi3��Y��a-}�-c��l�m��й���|˭G'���9�����	�v�F	��{<m �h>*3J�����a������O�9�=[3��gr���:��ܸ�Y�ɿ�ݧ-���0�,���X�����<P�����.�=,��>�/.�gz�(b�(Pu�K���ڼ�V��Zӗ�^��%q�ʟ���3��ĽA!X��^���99DJ�$���Z�K#\ېw���ل���eA�-��}��կ�D7��3'1D���m�Y�Jp�l�Q�߭�bl3I`�nG�t��E��g�f��bQ��ƘbP���0m4�եd�"�D�~��_!]��Y ^-2&!p�BIJJ��+ݪ�f�K�J�8yp�2n��Y7�+{yޢi�Ll�O� U̬P�O'�ϊ
!˞��M�>��c��K���;��Ib*���O�W���Cܻ��ϸ���n<z�����������_(ᡳ3�7ȯ;2��0V
��~A�S����Ձ���guk����/[��՜�Ä�/�>S�I��B��y&V:��6�	��]����]djuU�w�Y�������$��v�2!9����z��y�1Y
��'[�V�Xp�|�g����e@�J���>lT1�N�P��<��Q�Ȟ��g��:�� .���s%����v+>�B����K��E����	7x�F�"��7�y�����p��-�[��Xcf�� T~���d\8��K������b�l>с%r�/�����A��?t��h�!FL-��^�_OW4�YC��7:XĊu��׷�}W��!�Ť��D���7��[L!B&(3#M�J�p=��ME~?�0t�|7 ���~+�H�j:����C*�f+anA��d��v['�� M������]gM���56H�GM���Z����cR��T�=�����_ߤ��K�uE���0s��5����IP����hED<���W��nx=D��4=H������gm��Akq�FYU�)����~�����4�*�I�h����v{��k{��^G��Oe9z���������]��wP|�rL��8�t�S'���Xp�2N�)	َa�g��b�<M�ߛ�� ;9$|��[��d����>�uSr�^c �Hl`��GN.Z�M�@Y��kX��h��6�-[����P�L�p����_!OXzϥ-�)t��˾�w�<sdԲ�(�u��Tv�IH�z� �Ş|�mu�q1�����oΤ��C���h�FY�ݮ7^["0�N�/̄F����2�� ��=�8B�쇤��B��P]�(�ʉ`����9i/y) y���6pW��"O���{n�ɲ�O�w���}S�w�"�'q��oLY 	��=,[|���z�w{����aD�UR*Lo�a����b���t���ayƘ݄��\�ߵ�q���~�"�'N�V��5{�y2X�X�H�aQ)�������Izjr���(��������5����!x6[��_�ȐBx�����$���tW���Ol�W)�\�d�*�2[?�����"	9�5�	y�.Ŏ�h��]�)��'�'Q&э���&���DK/�~􋽅'���J� �q���lz��V��1gg�3�6S3K},�������ń���r]��,X�6�N�0^Ȍߨw����V���b�<y}."6������<�����y���:��sUo;���	�>x$�3������Z>rcy�M����!�I��d<�?� Rʑ�e$��ɑl��͟�j�����Ќmݣ�(q)�<�,ʛߝh)L�Ua�'`g����x�=�lm�ޮ�.e��.X�>����-���l~��G�g���"&��Es����qE7�e�H_5��2�����`0���a��4�m�d�^�m�u=?��>��6�U�a�Ry�斉��c'e�꒪t����U��.�e���t=�������VH�E|�� �����1�R�5�=@ˌ���wޘim�r���A��Ĺ@K�.c�Ú3tsV����q���o����!��mI�Tj���n5� ]��*M*���I���A�-�����;�y����Oڜ��䖕�v^��������r^�cv�y{�m���;r�<׼�`T7�#��ˌ�� �u[
n}V����h�fY?�p/Dl|l��牣=�<�tm�d���o��[�Bc�v�̒��2�LRT�Z���^�|%�{�Њ�p����[<�b�[{�Z�J4Kn����	`�MZ����V55�0n/NP `���z�����s���~.Z�',����l�4�Sy���x�	�t8������̖������y�_htw��~��'.�gB2T��9����ǱҀ�Z6�+�t�E�����E�ʶ�T�#��ۮ�ތ�X����>��AC�^*s@���i����8c�K�<�Do��N�Wj/&��~)7E\�Գs%c�ik<VT��ʢi����"��d�]! s�:���ȁLo��&�~*�v��o�I\|?3��QA��e]h+v�c����@/���bJ^�lf�&�� ���筎7'��1Np�Ȼ��|}���-�_T�__�{�2���l����ZwȢ>�tpTA@�Ӫ�R���q)�_cC*T��i�|U��w�y���{�_�����6��Q�[K�9f��ʒ����3c�Ey������Hy��,jܮUz��qл��#]�.��Ԋ�����>O�"�O��,e�����T+�p?Ҁ�ƍO�ɼ�;q�N�ɴ�(��L���Eɾ�N#F!��s�y@��/'DDr �[辝�𤳚8Q�nn7��p�D���d��oDǦ=����WG�z\�f�ە�ɏ7?|Q���;̍%L��b�o��sK�f�����m5���ɇ�8�v�S�{�s���aس=QXE��kF�l͍TG[Tb��3V�(hS��rjh��J��o��ݮ_g����Y�R���ؤ�AJ$I� ɜ���)t�v'N4)�>��{��]�4��'���|����674�_�6ť�d��o\��x\� ��$�n���Y��D�q�l�8-����S64��
�K��1�����Zȝ���=_�5f��t`��V��v��Ǭh?TE�*��9Tw۬�%�.���f_e����3*�%��z��#�L5���Z��1�^&��X*sC؅:���L��]�s��ls[T��g"W2FVmBz���O���������J-yQ���� �jnY@}cwL�����x7���j����O�����S���.�\���;1��6���4]5�ϳ\� ���X���T�\������y���:����\{M0Đ�
�W�n���_��G��:�4�e ��$e��Ѥ1�Y��5����(���;���t���գ�a^t��� o��$�-�C��)C,;�уɔ�@�������fW 2�?�,��/{��L�])*�@/J��&1w�5�����*�;�?�o�#��9<2����Y��"�p�s���ïk2����V�?*��q_3=�&S��x�W;�$�y��hI���ϲ�'��$H�5�O ��)E��ayH�p 2ʯ|�j�ϐl� �����\����Os�r�X,��T�<DӇ;a��8 �a�x+�ٗ�y��;	��{�B�za�n9"�_�{���m��(��'&�l~�b~��
l�ym!�r8�n��Uu��	,���ߋ>��i�3"��x�MM��%.=M�|�������XMQª�1�e>@׮���io\Ĵ�|ia���N��$�b6�mVE�
mOP�7�IR�t���kt`t��f�:����r��=�&2U�����$�>'��j�޶�x.��4�N�Z��ϲ��[ I���^��(!����c�_5�P =���yR���o����چ:�P�=�x���y�l�KC��N��i��:y)=�|։IY6Ӹb�(�g���6Sl��a��YUE�X�fK�.�m�}~��*�M�T��|SN�h��t���%��[4��!����8����&/�
��נ��#V¢����T@��~뇅�[�����FT�&\U%���A�b����W�B�E�1O=�U��L�<�S'�"#�}ʌ�k-)�ᢊ���q���&��\�.Ǫ����/!��H�����ゎ��/P�7]�&�\D�8�b��G������Sq�CG�b����'|6������V��#
K�z�����4�Ό���M��8F�$��ҕ�w�x�J� >�K�rq�����v����o څ@�#s��F��_FP��r��ĺ�B׏D��7:e"�
zO%E�C�ܪ�z?f�?�i(T~8��>�9��Ϝ�Qq�r?�m���E��_��;�!�ǹ��/���=�=� (�R�)O��_��a1M�<��;Jt�k�L�
hUc����2=��^�����j4",
�1�����]��_'o��E`)�)��h�U�m}�����8յ�����B;�.�UA��{	�m�i�x�9LoN�����I!c��|X$씀A�?��}�RYp�K�S!;.d��T(}6��..�\4�q��G�Q?�\;��T�m�5���ZPfC.@��!��
�_)��jq��\m���F��4�t,l�.��ܹ��K3SoQ෽��S��YR9-���T�2.h�}�����?g������֓��Eه	3�׿���vm�zW�4��1��|�H�u�	��Nۦ�A.X+��e#e�1�&Pƹ��e����$`��c�\�	D*�b�E�S�h6�7v��sZ������U�% ׄ�a���3~��g+a�D�M�gρ�����-��W�^yL��Ԅ,�9����zm��0�lu)��EYL����Z܊ swXƔ�\���7�J��Y���&�����\�o���*�PW%E�T~�F��$}xI=�Ñ�Lz��m���r�2�B�_�Z������W�`0�P3m�����kA�F�1��i���62_ݧ# Fg�shO�S�KnH�����t�>RUNa����ʨ�a�9E&�0f`���|�v��e�DL,���=�@��Tg���(Fp�Bð�h���H~t�̀ǩ�%r�<�cֶ���GTX�ɛ�.f�X��ѹN�6
@�X�#!Q���ɛH���&8zo�Mp&h�ˤ�o���rx��~�4��Y���CIE�1N��*��(U���Cf�;���I=LdA��,s|A��Y��Sq���G�mn:D�׷�魜��6�:C�:�~x�En����j�k�:�5��il䨾�Op���`�ze�k>��P�]�L1T�_�C��#�J��b��'ȻP�N��Fw?�88�6m����+��(������W~�^2ȧ��&v�_	e讒��bSc�����}��l�?�P�&:��ko��M.F� ��n���= �����s�V�ht�a��G�v�����$��}{��Hx�a�b��kB$�zjk�����v���bх��s���u��S�q�0oۍL��"F`v�
�IPs�(�gC�(-�Y�Us�s��S�'��-����Q��²���㲛Z�9j�3�F��F�'Z��>���U97�m�������ը���-��=l��3���%��o=�y�l�C=_����1�=[g��K�� {��Tf/��w�6 fnf�4#�%`9V�%J��'� �@��g�5�{йw�����擵'��
�z=0sZ̋[uEH#�]��|e.Lb^twg��wK��.ǟ��X��pd�*�$��V���)�0��a{�&h����(��	�-//�NvW����n�^�x�z��T`�`�ߪZ2B�ַQ<<+�-z�l������:�WL�D�t/�B��Eg��j��ls8�0�L�L�����b?���x�'���mW�U�Q<�b+�X���v�o$;`�<2{p��p����6G�G���jʩN2 �me�
��*�l�?�N?���S~�ۤV�����ˣ��mg&gx��9Z?6^�}���6��loc5��(@7�x�d(�e�kl��}g��X�|�۟Y˙΢�̎=��^��n�k�¹c�����0F�|���c��0��@Gu!�G��X��	L�� �H���s��W ��D=2L�����? V�E�s�|<ЧY��}P�~b��\22�Q�+�;��ؒ�AB[W�$�,W�跼�nvxƹ��[�=F��1>WT��f履���ߪF�N����i�i�)<��-�k��������3�}�eO�T�v����_eSFr��%S�U8vy���.��>��Psϯ &��k�6�~"��y���=ȗ	�U$'1?��(4Oo���k.<_��U���gMS"�������d�^�'�QEm�� �a� �Ģ������d�?���T���	�����>V��Q��
q!�ɚ�ݷ.[mu�#�!|��d�.�7ˑ���h��E��0�־i7���9���c����p����~Nϕ7��}��?��!�2�\�Q,�ہ/��=��zU<Voܙ9�j-�:��P`:�G2O�3��"$��,u��GKY��L�8G7�Q�U���ut�/��G[q8�M)k�F��e�f]���[F��;2�恂wG��������	�0��߿��Ð�'U�Hn07�Z�U���#O9�r��k��)�+�[��i$�d.�9'8ۦïNԳ���
I]I(M>$탪B�)��y_��|ۘ�a��nO�WL���6��a�F�:]-��A��ܮ5�b%+��������g��C���Vu%���nk����K2� C0���jk���V`>v���&��2�W&<��O,GyT}*x�!#�
�ĸ!�J�J�[mx�g���c��j�K�,�<���s#�*�u��Fo���}~��D,ڃ���(�41�!�xzy��5(��װ%��~t�8ˋ�!���3��asuSn���y�����HtAԂp����|f"W����2��3��J^����
:��س������c��n(�ޞ�u�7��4i��=K�i�û�S1A�c�CMs�M���S����B�8dl�瀽ڻ�hTx�]���F\1�]9�p�tIL�[ ���y���0ө���c�Rsu~>0:��<^���K5�j�B�U_�N\j��Ƨh��v]zo����MClUOD<r����t3���-m���xZ(G�z@���E2����;�)������	o;�c���iM��_��R~�''5�ZƂ�Ϲ�;����HZ+ =rZfC�Σۯ���:Q56�sTd�KPi��ʽC�\2�2)L
~���>Q'�����Vt3��,��j0e�"53��agm�������\M��fN{�桲_BP��F2��o�GW|FJ�k9,Hu���[�QH�P������;�o����Q;dӦ�qP^�o���ӵ@o�l-@x��!�5��B.Gj6xb�|&2"J�`$�S���n�BaP�i2�lHI{`��F!s�Eq�*g�L�\���������h]n3�
D9��u�s��z!A^�]v+��ҙ���]�d�fY�U�{���;Z�麜/�$��a|ۯ����:?U���]�1�+m�M�l��G�����t��V��9�<�f]O
|������,Kj�| �#��8'ܱ�J#Hid�o���|�0 k�h�t�e�����[��������qo2�pZ�a�N��OL��/F=�<!Z<[�1b	����x.�|�E��4lB3�a%�l�1^��L0kn�됎��\����ں�b�l�SS�Bw+?�n`hoI?�]��r�%��3Be�-�~�S6E{Kﴲ�|�
��Y�kQ�A�rsQ-�zdj��hiB�(�7p�b\���]0�ծ�+&�U{��K��"]����o�t7y�7�;���a`<��KS��e_c���g;��g��o��=����j!����O��U���j��D�p
c_U�cq}l�����1}kn��TJ��fDM<�@U^�׎c}0��~�Uw4�G�2 ����/����
SS�0�m���5����x���z�eT˟��Uv�J�6?�5��W�
����&�(�'���p��Z�������E��l�
���	S�^
����ޒ!��o�F�p��z��q�^(d|���p5u!�1mĮ���S;ǔd�ve�w���ڻ'�"�=3B�z�J#�}T�DJ���N�������B\9�^3���͖������-1NF(�ξL-'gí&2*^!�͞�YIo�p�\����^�������: V��G��4�����t��^'����`�`S�ұQ�c�(�0ϗ��8>�3��0y:�9x}"�In ��W�����Z�s��6�B�>��2��7oR�>� ���[f���Y�MO#����Fo�7T�Ƀ��%7af�X'R,	����I{�̷iC��=ĉ���=�{5�H�m}\�a�?	�Q)�����mm�s��NJx��"��Ժ�۝���cv�_"���:��,�+c���YP�I'
`@qժ�ys�)j�!�{xo��k8��Mq;I|?[�������o&�'[��^PF�p��b
EZPZT��&�5�u�e_YV2�ܻ�tA�\G|��[a��Ag��$�q���-�7�;8D�߆�CjfY�)����e���S�1�ō̜�N|1�{�*A���.iȏ�1�P��_�x:�x�z��W�o��F�{�j�veG3�Z�`��<���
��
6 mU�}��[�^Qͻ�J
�3{3�v�E��֩�I8w���t��K#��Ȳ��Mg�4����u��h�ᝢ�Wj�B��f��ι�"��Q��V�Xy� �:��ߚ�V�&�Zu�.J>�z?77q�K�Є��9H�&) �"sp�Q>��CY�i�ǥ�'�WV =�/c����s��Z��|H9�����ñC�Y��w�w��@��V��0߆��Q����1c��V�a�O���G��3\^^�ck�����
nG�vuҼ�͠~�6w�/��Ƥ�Nm4U�����_e�X� 8�h�h�akѺ���9ִ�<:��o�n<$�M4U�����ȃ��1gV_��8����ց�,mWӘ��7\...W��H���G|>�O?8ap@֌_�qˣ��sZ ���\��G ORR
2�R�_��XwF�7�P��x��3��S�g�9��|&���!�|����]�R����6�&�N��Ŕ��r����x��%y�?�F90�YQ0ML3���`�nx�y�������iq�������%a�9�<'�+?=lܠ�Oɻ=�A̢5�B����{�#,L���m
B1���)�x��X�H,
*��r��[7��3�z�9�hTV�<�27�f�m"�-[�2�V�������C��/eBm�<��_�HB[�)�`�E�T�aT��Ѿ�̼�������@[����Za���lc�Ѽ�h̷c������otO����H-�qD��V��*:v�"�E�o=��C�U������D��~'d�N	o(Zb�\FY���]s#���-4����{���l��;p_fܶZFc�"�Y⯲H���n�Ӧ��s'��gk2 � ��ǻ��jV]j���߈)��L�8~�3���%�Ԟ�q�!��#�*l��:�:ݲ���%�Of_o�x8Ζ]�Y�P�2��1��}UPS"�!w�q�6�HcJ��S�LХR{�Z5��Uv�xi�J��Q�%�s��b�]2ZV�RcU4m�d���m~'���}�Ns]�<�3� �Fc�������{y��sb�])eޮ�a�TZغ�Ȗ���������io�J�\ �J8�5D���`�p�{�E��G�
~����x[�&��WF�]�Wl ���v׋_9���-�۶f��5��M4�E]q����mo�Po���i����N��[|�u���4�H���ww ��Z�9���3q����|J<y�9O{�����;^_�L��+�,��r�'6���Z�iz�U�{m�e?���C��b���?�UyVz�X�\�j||��8�aK��,S��D�x�Ȼ����UxB��|΋��(�����b�h�Un/��b���">�4~�!$%���Rd�cßӲ�&|M�+
����9#�ϭ�4xn��k߾�!
����z�O���l�2sKXINR{%�W|��:_��%�r�ù�Jb���A P��rb�*F�?���
��#�i1���[�}g���J6.K(�讯A�sHt|��˖�3oP�"|�7#\�;�|�xu�=7쑉M#G��6�c��A�5��9���J��he��3�uT�O_�iZ����{�WE_z��/Ҁ�+��9�J� ;�w�B�W%�����XG�#&1�M�h'k���9)�6%>���/��Y��wU�����*�N��P��R�b_��������'�+��6�믨�m�Q�ᷖ6���^�w���0�wˍ�l#6��3�{E��2��O����h����GC�UI��}hs���ͯ1>DJ�ǚqr}>;����:{�G�H���6(��J�|?�.��M*0�jc���D��Z`&GyE�/��Ч��)"�܀�3�O��/N�㭙�\��i$ƥ|��s'c��M�xi�y��c��6�������䄄��3N}A�nM�٪ƪ��d�75�z��S���i�6g�A�,@>
��р/��Y� ��LNȇ�󝝋�1��te��/+���ѯ�`��]~e��ŀT��89���nk�g!G��3��.眣��+���Dx}W��uBڍҀ ��Z-8��~2�|$Ij�\;@�HI����:�_�8�ahs��;[�eT�4ϩ�ڭ����i_�2���({�͙3�`�~��+��IT�l��*爚	O%�c��>�����享u��������j��G\�"kcrk��w[!�'�vU��}�P����2yab�{��2��RhTP*�vb��be"=;h��@Au�ҥ�KQ&��a֑ͬ���*�W�۟����/�߽5��6�����Q���e(�Y���5��*M��ї4;_n��2<��^�6�'��	��9T���h	�9�d�۹��M	;�t6}� k���JI�@f��p�������aｔ����Jڢ}�E���c��`��'I��A��1{�["���Q��3]& �Ƿw2���Xf�\ں#�ۘ<����v�1�5��h{]���k�ʨ��-�ڼK��� 7����PYvOq�m�盕�!�ԫ0�3M�;�-C�-8���2N�3�-V_B_�A�0\�Ҍ���l�c�2�W��ħ{֏U�E���e�@�Mz̅	�: r�`�;�^^�������� Zx��]�E��Svs��H�Ӣ ���y3�+n`��x-��M�E���Ƌ��^��F��2�|^�
����qw��{�gy@�na����byN��k4ZI�64��x�,ئ��� u7���s�vN��X��_q����"#�X+¡��<~�xIok��D��-ld'e��y ��n�Y�M����u`�@��
���G�5ȪNe�q������1�[�����K#��}��߱!!A��gaF���H<�~~�S��v1̈�Gڐ��Q��B�W�:¾�M�xL(�rH�4�
�i��`��
-����<9;T�O�DN�bog�k\�[Vt�Τ�Vc�$��۪��A���H2ĭh�A�H'AD>�\�T����
��I��W���'�����������&��+�~��K������(��6�Oa����&��&t�$bc��
`y�L��K4��;��qk�z�eQ3�_�j�0����4;�G�7����/�LWl�N�j���IHFϭ����a�΂h�Z�o�{*J�l�&����t7���?���i����pP�,.�Xe��vʅm����D��!ɔiqGS0_�W�iJ���uS�R��"E��X���ԓ���)A�q�2���R��l/�@��:u!Fl���dFCgZ��M5���sy(	;���`�3����a(#��g�g�������8�kY$Aݧ��~?~�4ڌ@��W�MA=�Ӷ����)�YS�u��lv�vx�OA�<�H�a�#x��a�X/1�z�_��W6�H�ō\���,��M]K��9�az_"�V��[���n�8Z�^V�@zz:�mfL�܃;��͒9�K2�6a�g��m�cH�]�W�L�9f� I2?�;$Q>�"� 1U�a�.��L����'d\��������ZU��ۑ����欧��B8�0�l�`��0��wYC�-E�`C C0r�����,K�b�"�<�G�"��_�nq;K;��r��������|V�xc$��[r�=C����q����5�����S�~����Z���[�V2��U�i���e'�k7��\��FQ}�����%��N �)�`�톯/�e�xD�|���+ȋ���2u#�_�1��y����;�x��;�l]sXE��N�fK��v�b6�9��q���^��1Z0�_��hS#;⟗M���X���H>#�P���їc��( m� �E��\ ��%��#,�3�����г=X�Z�;��L�НU����2���F��#P����u?T�<�궫�Q��hׅ���Mf�.c�����~̈́_�u���ZǞM7�'/N\>dl~n����HTG�D�9J���q����_����]`��dF�@d섷�+�Ч����Y>߱�gg�uê��-�(�W���i]%W4���=�&�1)IɊ��|f_��m ׇ�w+t����݅��l`1�,���[���ш wM�|͈�%��jo'KDɟf}��鈬:�����M���`�(})�����t��(-qzV]���٥���{���������d���e���՝ȩu��"��V�4i�|aR�\��*��q' �k8t�J�Iׯ�WWri�+�e-t0���]	�$���IG4�"��	�V����|c��~E�J���<b���--��3�����L�9����wE6�yqT~�c����|��	-B��7[3���{��gO
*�A�_]���YL���g0*��n��`��"
�I�����j$is��r�丛��FZ�M2d<�SŎH�}��njF�4e���I��e��O6M}j'�cL6B檣kVض���p�'Z����)�d��$�3�m������v�/���H�X�7���sZ�z'^��4�G�%u[�f%����+Q�]�Me��4����%ό�����cO�牣2���ί>E�$=�P�3���b�z/���K�L5�F���n��(�x��q����y!���.�@�����Xs�IݓP�����DךJ�~L>*Q57���c�̋�u���p3��﵀�z�43Q���r���m^�i7�iH��"���=jO}�t	��6����8>������xb�%[C�5�s�~�s��nq\�0d��K���$C�l�U�'	6�u?�e��x2;�gA�Ȝ��@���N椼I荍S���`%�9�X����z��$�0n�V� c<��>`(N ��#�B'(�3���XksK��uDO�"�cHm�Bӓ�?hi�IՌ�K�x1��g�*�Ұ?�!��y��g濜����#��8�P�	)RuXQ�ۇic	w]���YT�)_A�����&���Ͽ��lH7�Op:T}�ׇ�2q�k�Y�۟��w��} ��bR����ZXXXI�l�,U����k���]��?:���8Uq�ؖ����aV�[����^��\�ޖf��BE�Lz4�T��߈ʶ���=|
��mɗ�k/��'��J�fJ�f�&BX�헦�E��]�vd,Cxo��f�8@�i��Sx�2��A����vh����*&B*�Մx��ɜ"L��'��c�ס���{H4��WJA���a��p>�L�9N��d�[`줯ݚ.}A�x�!�����_N��pԯ�I������7��x[8�^�^`ύ��� B�DV����\�(Ql���I��ߒ���������g��U�0���_�\5_V�7���6u�^"݌e͑*���`|
�$ν=�s3����y���CRi����>���+�f��Ǔ[�8�U�~8�nT̛�2X�pᵿQ��D28|��)���Q�\�����գ1Կ��Ww�1F�5�q|K�����[t�)3'�o��`[N"�Q����%�w����<ӿ��N�neSdڔ��X����۶���--|�9m�"�欮Y�^hA��<�Z�v%��|�m�E|���t��:�5�HD�4z{�)�(>�?�Ȍ��W-g�GQc~_���u+�h�� D+�~Y!!q8��R鋎��s�����HϔG��C�X�,X�&�\�:�5�r2�{�/��N|1���6�7Nw}��n���P9:d�hq4>�D}�d4sa^�J:a�V��1r�d8?X.�ʭ�X����;ȶaUM#��������cYO����I�2DEE/>OfԄ����s�{iB�b�\�����yl
�7�������Ty�q0�����I���%����`I�#\^r��u�AvNǿgD
�����(/I�mME��qiƇ�?s"N�?��.K�5����*S�8�኷�u�B@���4!��X:��E[=�R��O���x([W����}��=��N���Kw<F`�Oȕ�������MY��_��[�c����Q��|���f��o��%L&N�±H��sKH
�����P\����*�떷3&���@�Mj���G��tg�E]	��ҙ���m�F�&���&���]��y�"v=�'?�Ț�뗬���ѧ?gZ�5e�g����8 .1լdk�r��;@���?�S�.>�Y���.;�,ˤ�{���K��ph��_�&�qP%��n&nA�/:���.g��.؝�I�z,��r[b]��Ո��{���>3Q��X�����Z�0G).�fvO�gJ��3s���s�ϡ�d.��2l榔�ӆÜ&�ok���GJ�X/[Z�h�^3~�@��~���x;>G��9J0S^sJ�_�"wj5=t�-=�x]$����Cȩ�t��6-s(��v\?&�&����(��c�X�s���kaK?w0�_�ݨ�ԣOLߪ�vא|����`Z �7X�fI�4R]�U4@!�(uThQí�9x��6{��M12z|(���i�v��1���TM�B��n4CHWSt�8��6�[}��d�\��+.���i��_�H���d�nD���ǳ�c�86H�s�!��9��tw����]Fτ��2S� ��xIF��2��Su�8�K�
�"1;�w�W^���B4�~��-y�y�����vM��]��~���x��3�A�No:�u�����\�N��֌&� ���9SH�?� ����9����s=%4�w���x��H�u	fSV�$cV툑��m�섣��BpW�CV 禕W�>������_$�4FOצ�{�e�LC��&ԕ��k��Ԋ<��sx�Th*�쒤��Vu\�,Š�.���Ȫd�:�Xү��h��xw�B�c�v w��x���42y��?Xl@������f���b���@�wd����.��N�k@�+�J1]O2G���:�8ZE)j9� j��)��k��X,DQ.Q�#J[���[D��x��	�2Z��ǌ�x���(���X�p��D�`�L�hƊW!��5ʎ G������u�Lo��K>�=��HBmِ���Z��}mĶjIB{b���A*އ�\
�r��PB�t�	v��*5��M�5]���}˳�c,tѦ��^�#����\��0�	����.��s�@�J��Dg҇!��	��,�]��Q��1���<;(�m\]�ѷZ_w^�*�
��.$}�ĥ����;������&2K;�/g�u�S�Ik�_x���5, ���|���7����R�E�n�y�6�La��ʔ��dn�tp�z{�m�n�P�[j�^��LGЄ���KoGd|�ٶ�ʶ1Ʃ)��ll��������G}��A��sVF����H�[ݔ�ۀ`�X�?���!�_q|�w��h?b�M����<��^Y������ཬ`/��"�84����k�J�#uE���ر���,!��5)M�/n\�Η�=�n�0�L��2R�E����`�����?�@���\�=as���	��f�K�K������}y��*)v�i�é=�v�i�Yy���G/�>���ŊȌ�T�vB(�G����!�s��B�m�*�ũ	�?��=!\evd.��1���u=��?ܦ�դ�ո�m۶m5�m5�Nl�<�m���ϫ���}�s�=3kf�s��g=��a�T�Y+�ea,z�z|}�7$�5�+�pB�9�F�~�E�@��i|��3�ǂ�dz^����C�R� 	�6LB�wv�V��s�g:��������~<pc�GH,``�����#���o�Ǯs`p�N�E�S��� �A���ƿtQ���~9c�c )U05�}5�×ܕT��Ӣ�n�,E,ڦ�l��޶ax��z�K�Q?4�2��[A�����P+�6��i�vT�7�5X����]��u������I�����`A���[N�W<S��o��"q/�n�J��;��Viǰg���8mp��X�7<��3sOnwi�ZP;��l�8�6h!+�'�YN;R��Q�z~Y��ˀln	�\Hv釕�s�f��n�T�S�&�t���d�+�	�3d��%�n�+���?�Qns�m�r�7B���b$��m�,�6��D�MO/��k�"���޾��E�!��,��r�f(m���~ę�1%CZ.߲��79� �Z���k��L���T5��wC�&��s�l�f	E)���.����wNily��l�����Af��>��P;�!l�N�*$CR�n;���F
wm�)*wr�mNҤm�3�z���
�0FԱ�\���d�(;��7�*�}%�_�Z�\�EfA�O�k`��
�&���e�ܳ��ݨ��2�g���H_Β?��?��-����e/h����z�S��:F97��S��8}`�L$��#Onu^�ћv�$n_�^�!OH�b���!���s�z ������S�'��@��͕�Q�:#�K���MS
j�El`�,��.5�I��
���a�e���	c��ھK̠��ʕ�C����[�Ad�f$L  �(��ƈ�y��z����0��8�AB����5��HR~H���F|���ֶRUIk�4�1���Sr���=3J	M�^q?���IHҀU&�y�b,��`����6����#Y�C�����hځ�s?n6��������O�2|mX���Nyy\Vu��oy�G"Qm:M��rZ�)�P�f����6�qKe���9���:򪢭�w�H��b�|m��l��4ْ�X�vW8�(�#���S�R����6X�X���
RQfB�#E���
��� [�׈Z���?j�2�[e���t ��|Myi���b�5D�BM�<�RCrC�C�E'GIQ��RtF��姾������9rs�2�H�j��݈O�d���_�H
�2�Op�vH�̱���ͭ$������.D�F!��_޳L�3u����|;��QϵJ.dYs����Rs&j�A��i(Ɔ+@ ��bv��ز?�T�$8 >��4ck!$-_�D��0@����U��Bm�hj������3�������"4����nn�-���J��)A����?]��%9g�F���`� �a���ɖ��G?=�2��(�ǫ�(V&�9b�l�i����=��7J$����w_A����������\�T^K��/;*���#_"���f�f�>՝d^Po��EPL��P��Hm�&�V��<qgE���U4��& �tN�>r�����{�m�� ��2?� �g~����M��حo;��+rF�q�)�zgDjr\�R}h4G_��� kTg0�T�B���zf�+W���ь���H�}�Sn�����1�5N�z�[2�&i��S��z�F˸���2��1�`j=���HE��5l���ѥ���&/Z_�]/�����ɧ�/��)��"��X3B��q��4���Q��q�6��J����V���I?9ewj��=�d{�^v�S{��`r����7g$�4���u��Z�G7<-=H�>���J�ps��m$cL:�J�ktm����?�v���yg��o�muhBg!+ϊ���$�B����G�����1��"��������㺫3�/O�˴��q�ؙ���>�i5��7)�L؞���:T$-�����zXD�9�Z!�w;�~;����z�eD
n:�4p��c��5"�A��۔*�ʪQ�
�\��k=�ፏY�{���VX�^1Z��'z>���Į|A3t��-Um/��s#C�+��de�$�xT3�]O;l����AL����y?��������q|�ҳ٧��h�G'�;�Uh��UB�7���B~��F#�.�AX��x}�B��'�� �V���R͘����L�o�\�t��^x���K>D����γ�X�b��w~k�O-�J#]�����7l�M���-t'��A�Ly��[?/�r������� ]5t!W�>�H�3�D	�vx-'Z1"ը���;#��(�Ih@�U%�Q��5tŲ}�0G:�(�D�@KLK�EK��K|Yi�K1�����U%Ij�������
���2�� �?nI׀NwV��7M��W6NV�O�����hA �<$(�8d�˷B���R��&�&�c����Le�ab���\�������a��UD��H�j���yKU-F�D��3k(G�57�$4��d�V��<5J�.T���uݧ}��l% 
h.�n��w��R�"�XԱlluDG�����v��v,)h�����%>�T#+���?�(�䋼Qftj�e6M�XܞЍX�W[�G���%�W�@�lW`-42
�s�"̃�7�0C	]��(�N��7�Sx�qP$m\�\��
���p��K3$��N�~���'a�h{�U6���!
ж�%�*��Z���o�j�A��$*��6;|&B_��\8��������B�B52Q'�?�$��0�[���l�	i�oS�����ǒlQ�:m�8�: 9��[6�*�UE��q��8�`9͑���QZ��W�#������m��<��`��J�?b��U7�:��ǂ�~�@���e9�#zPŲe}�]EM1�9k%*�I�P�!��?��!r������L�Py�d�A�i��*s�\�楔X#�2���ܓgH���gk�	�ݠSk՜ ���X}�����f^\A��v�y�G����"��f$�PC�YG���ɝ5���P���ɝ9�4����b��v��B:yL��`��cّ��i�v�V54Ѩ�s{䴢#��h$	��;�{�j���!.�f*ϯ���W�\�!�,� w���|l~ε&�7d�0B�T�Q��+�t��>�f����
n�v���)D]�ưo��m�D�P�3b����tנ�z<�-N��j��D�C^�(W���I�թ��/��h�[���?��Cxd�Gh�#8>U^�7/�r�%���
����Qh�Ū*-A�V0�R%���NƄ>�{/�M<rS,A�z
W�qnO��E+4�)�L�N1K�x����[��ssȡ	�Z$�d��>Pzsؿ�ҨG��TxO@p�/2�^P�7�0�<��C��`�b�f�M�6e�����m�o�����VKa�#���ʧ�6X�Z���.lk����)���u�hG<���)X6�`��,�e�E�a�B�Js�2�iRZF��=7d,Gi}w�+�'6���s����g��z�ag ,P5mT\ޔ�.����	����J�)I ��=����f_	��5�B&Y*d�ݠ�e�����N�8�/���m@��w�l40����������M뭡�dd�(�`-�����s��+������L�n:�lDk���饔�mdo��q�C�H��^�V��,�@��n�&��g �Ӻ���$���	�Q������ʝ$�h� ��b�}��Hu�2��������ہ*�	u1���r�%�%�V���x�b�P�!,a��"jH84Q�Uf���f��&qO���5r�b/ⅠH��$��UdC�(FH���ʹ��s��|�pϰ��!�� ��<�?D��к�z
��g���d����}EE��ڋS�nv^��"'��R��/�R��:b�4}�w=��A3'=,�C��gC23��\��B�t���qD���¥���&��T�V�<�.�Cyq��1�}�֕[����+)DZ��;��$�_�To�`p�^úSk�ħ�h���Zp�˰8.s_��a��~��D��rY�Q�I���;D�~ ڞ�3H��BTꅰ�ێ2�a�3�笋���*���#���圄�p�[ [��]q&�}@�r8[��P!�D�w���}�}*�R�ߟ���ףʕ:F�%�c���Rn$=Z�y�'�΄��m��ߧ~<i&��B	u�	�	��p�9���ٝ�������!F�THT=[9�� qCen��5�;�.û��71Z]n�=(���QO�`I�D�~T^�R�E�DV�N��[̜��b�G��3��/Z2���;B�^����ծ�e��:��]�o#�����=hޅ ��%.���YA�3�{>e/�ZL��ړk�L��e{*.�,@'X�+�,�f)��*�0:� fP��o,I����n�ujqs��|ffy��rq~t��۔yޮ�r���{��3���&jIĖ' �v��7%W�a����s�6��u���$������.�*�a�XJr+�0��5�w����$�ڢ��H��I���;M�uzgR��-�B	a��8����/�m�m�����c'}VP,Ĵ�S	��B���[����t��NE[+3XB��V�ɠb���
��Ev^�F�i͑�0W9$g&Vd�E�U��=H�_��m5�NM1W����,,���
�T��]�V���G�!��@^[��a��T�CC�董$b���	�P���إH&lU���.�h4�ڭ2�u������Wt��b~E#�c�!��8rC��#�+i���@��ϑ��:oRu����pѡAȉ60�m�Pru$�S�>I�M�1��Ε��C.J�{)�*&3&FAM�I,��Օ�p(��!�A��R9-��8DXq�~{C��L�	��	�$�ymL<��'����۔�^N�m�������lF�E�����G����~�	kP��RM�$�^%\t�Ȕ����b�C����mR�f��2O����⇘���k}q�:,�4&�w���i<����~����&�@� s�]�0���n�A	��/���1a��9������·����F�Q= �W����*���i �q����H��"G���
�^�44��Z�0��<��l-Z:+����E��h|;�1�y�(G����a\?éx�(��:�k"��ujq!Ty��
<v��9���nhj٫s���<����C�eH�(���?�ጷ]w�DI��!A��p���3�8�x�P�wd��º�D��\�yyʨT'akiYTW):�t�o+Q�\�)�����11|��<��RHiִ�{r�<�xm(�$����i�`����n��ϑS�X�?�R�N�%�_����(�c��y�b�Mc�|�$��!�bn���A�V9��Al0I��ͬHnÆ3��H`|9A0�l�/�^��H�blc
0�������]�0~�d1 ����%0��#����P�6���ʎ�ؼ�o�)
%2�gj`��Rd�[c1���I1پ�Dc�_�i�=����Dwk�����Q��.���N�K.�u]�� �~T�ir�۲w�5��p��E�E"���[yړ�Z���ʩ�5b4k�Jw�,0;ੵm��J��ړ��_�簷"��V�ƪ���ԏ�[��s��nu���	^k����ϕ����3&��2��%t-d��x'܂Y�f��幭V�޹HV��[Ȍ��֛���n��N�a�7+Z����0X)2i��������t�D��29���!xm4	�^���-bd������05�V�`.:r�Io}[5���u7�{��=�����7�dn(���������%��-E��3���e����`�Sl����4Ɏ�U�$G�2�����?� @4y��]u��ږ��yr��@(�?y�Az��U T/�.+����k�#.� �rʐKs
|΍���8�!�]s��w��8�EѴ?���f���;L�8�֞(@�J�}��8�o�"�s�u�U��
ϛ*\j 7���k�H�G���B��@|&R]��&;�獥�p2?(���-%�ެ�l:�:'?�k�x�Z+͈ G�ҧ�0?%J�Ԝ
�|ÞBK����P�)�%�"/�k��jH9nD ����z�g�|�X#ݟ4lH+��Rc�Qvz`j��,��mW�v�Q� v�$ �h*t���ͧI,�̝u��N��A2�6��l��o��D;rP�"bLT�.()�|�������Q_F_|��KϽ]p�+�O[�%v���'B����V��%=ska�3����E�6I#a9���㥨���YU�e��o�`�a��p�Y�Ӯ�UB��p�}�0I[�Y#��ɨ�����lP�q���k�+e�,4`'��bd��uJi�Kؿ��_�e˺ns
}�FBgA�ް���AM-�L��CD p���n�*Zr^༞����,�[���V�q�~p��<�]6F��G�F#̍��D����n!����_��n�g�b�m.���F��3͏���h��6�O��gaA���|ND���oP��^ۻ�o�Jw��=���*�Z
Ȟ�
L��BѸ��d����s�l<Y'�	Z��y�����Q�!��h+��z�I��

[geCg�\z�M���Z&ַ<d�lS��G����
!T���qMV����+F�����P� �Rbe�ؿ>��fu\T�۾$�W�G ���Ɩ��ǒ�g�CG<(!o�(@�وNӨ��V�q�D�uun�䑡u}9��8˼�7����@Z�E��'��_1-�CLc7cl�� �	�.��*V�u���Ip���s����G��/�"��,>[��&�l�B����1��"��8��G1������$���1>��1�1rS���xQ��uTP���P�*b;�����S�8�dq����a'-sI��]�a;�A��v�8oa�*N��r|s�	��a2��i�rC����˵��k)���efR%Y֟�l����W�R�d[^B�H~�9ii�#�7	�8v���R�۽�g<�Z{՛��i��.���+��l�댄sY�Ó�X"s�W�^��Z��"ٞM��^���?4J��uk9}&1�
R�Y3Rv?8�B⌤�d�lr\���|��ʒ�\�`�U�frd�6��S�����@�/�Zq�.q��&e�p�{7 N]m��tY� �N�nE4(3�4��'$�@�T�YN�6��e6�_cW}z�����8�$ǽ�YY������g��"��V�w��XZ<��߾k���2	�@f/�m(%C��l�)��jx��V��^}Q��!n�N᫪p(����-kk��[N�����i4��a��+,̞���Ft��Q�px�r�2ҿ�j@C���GLD*� M��?��o��Q��]� ��{%��-\�6�JL��E��^��`Û�jn�L�2��[|<�{ȏ�C��S!H8��_<�}��pӤX���5'Mlb&3�Voh7S�.�,>oS�O�d<iP�%��y]�KUrdE���zt�LTp�mK�<c��[�8�A �����x�Y�cX����8IR���yA;쓖hW什d�	>���uLz� o�eşBG�i��s++�xRRRİ��Q�bwww-���)c���練��iv�@�Ƃ\����,QbGK�O�to�vw&�ޯRlN�������+rh}��5D#�kLd�"$�Ѕ��۝㳁��`_�������J ����T��ꒋ�R{9_*������u��T��,	a��Z��K�?d�YG��������[N�����딃�v	���{�o���ҫ���p��<�}�u/.+��6����X_h�.>%<�ך�M��«���:��w���|�%���8x�6
�e�R���|s��8�|�����j�o5��-�~0�!DQSv��8�����b=g��*�gNy��[{�9���e��n�b��]V�!��h��V0^!�Dҡ��x�ZPP�}��W�[�ps��3�M2���B��R�v.[��5G�*��r�L�Ac�,h_p���P~,�B̢�70�j%�Qex��DI���bQ��d:��O���a�X�����N:���WK`�B�F��Ǎ1�ú-�Ӝ�sa�s�(���N�_���c/��K�W�v��G-�5�3����GxP4R��팿�}�i��m:�H#�x޿uԸN�$8zLr���5,j����E�gu��N_x?p�$Y���8�������`�T��s�q^<�8Of�r�t�>�\�}��������� �=�՝f�g���������E���,��E��nN�oT��^�d_� .|+ +a�UG���!X����B0���pߒ�}�7��0;=<.�Y��:m.n6��x�̆��לgÿ��pڬs����Mb��Od,s�obn{^6�����_��_,I"9M���y�a���)r����'��%�e�4o�r<���^�S����x,%SF��~c�����z[�稏������ՉMe) f��ͬ���6W\FNg *���"�d�J��褳�^�|��=rF3��|�2t�?R$�����.o�v��0/��Cߞ��X�'B�צ(�,��7�d-g3���ܾ@6�=�!�{��q�>��i)Ur�?64�G���px�m������A&��o�����ѸR�Y��"�j�� ~w��6纙`�gn��S�Q�������l��T�磢ٛI�`l{�Nl��C燖�K�W�w�� �z�k������,��G[�ʶk�7�㒢۷�*[���4e��V�;��lxvQZ:��A�[�62¶�*�����b�J� ���B���!f��D�G�|��1IB.�{�V����Bd��<���1�"��i���9.�"0���3��ƽ�3�����'��j.w�ҰS���B��:�C��.>������w2_'%	=��	vk\��o`c��s3^��踝���x	*��xY�0������Q���|�'9#2��8�Wx����Bq�,cY8:�me �{ ks���by��y=B�h������
��F5m]�X�di�1����s�fQ�+Aۮ�,�ؽ�c���ɈvV)����B�n��g1U)��/3�n����͢l.�_L=;6�=D��j�,k�ê��*Ia6��6��޳*�]�̑ldG�۹�*Ys�5��O�]��yn0�9���Af7�~�B��)���ޅ�y��X	('���0�pb@#�i]��J�yp��@U[�y>�1�h%OU���\��T��G���M6qUs���L�l2���a<�K�$)�����έNbXm�Zu��1����l����T2ޔbj����4���D��!~�4����%���C�=�C��q=�n�Z�[���0'�����x�.��������vUaK5�h4Ew"O�;�4��߱y�A2�ה�;Oz�����Y�>~']h��:S���cv)T�Iud�:�*�r���T��2�ګ���0��>�:~�����xO]Ձ�/�n�TI[�QըM��m[��Z{Re�%B�QM;Q���EoL���
vo[W=Y"��+P1��h�42I�[� {���u�o����Wi��rwҝ*~���-�OaIBD��{~�V�t��rZ^a���U�غcM�=}dκ�	�P�:���|0�0�]Mv�ײR�dؽ6>/�{1��S�i�rs��A2������?�/cb)"Qqw��~�-��$~B�}�������/�/����lws
w�����g<��r�`���U���V);]��Q��j���I֯�Co#�x���xdE��>�5�4�M�7�s��F�[������V���iV��2�?�G	�R��6��ERk���=��_E�$�j]�/E �M�wk:n{mz�ˢ�q�Mz	��P6�h>]�3��#�ō�]t
=���)-�q�-B��3����Me���8�i ��bf"�|b�`�iNU+��s�d�Xc�{�n|+}v���͚�44|��J���`�G����6�Ƽ��MP��Yܽ�<���W����z�<�^�4n+w�}dp��f����4똥E�C��x�,SG%� j�SR3�ğJ��n��B߽UR�0�Z �ԾQ%DĴ��q԰G�jE~욕��ڞ{J��A��/��A\�.����$�S m[�+y�cz �3�����I���KW�{�PG�#6�, E��������`k���)Tڒ�8�KC�!*���Si�ڭ��d�]b�
AΤ��{Ғcs|�7vN[5�-l��������e�?�f�ߒya�D��Ս�<t;yLr=��lWL�d��{&v\�F?���^��^��A�7du2���봗�pT*�?Ń�j2�Ȟ ��.'�j��v�A�:�=�����,ծ,�:ĠC��'
�I}�DvBakR�ɮ7��(tQ���̔�'�$a���J@��X]�,GV������_rZ����L��;4�x:dE?��^*H�L�4�3��S	��H��pf�b�tS�^?�|�WO׍?�k��(�;K�P�"*)��t��oi��n����oϩ��v'�&�l�-u�D��v�bv4S �	����$ދ�~	Ѳ'��
��M���W��v�C�k�M۸�co�ݭ?��Mi:{�[�"��e�M�W�8�o�)�(W�H��v�4�����C�L�}���?���+�f�_?���f�������H~7�ny����Ř]�"�.�V��.ٝ~Xh�k�N�w{�J8$�j��f���]�k䄢�����yՓ����̴u�ʋ�2�:�o�S_J�ő��{��ǧKc*�)k���r�չ	�&�q�߄�XѤV�<j�@���u�6��4�c@��w���%*�)AP��C�~��i�D21�f&����h��n�|4u)��Е�9t�G�a�\��lE�^^^b�P�����:M{3�ch���H����CW�į�i����ٳ�2�O�Ǖ���<�u�x�wĊ9�H�����',)��e�A�.�.���;�N�
�1U�Z	F�^�Nl��W������/�-C:�$x4��Zm�%�M�xc�-9 w=d%�GM7_� "��/z���AW!���	=u�|V���5�¨��4�2P㆕u�s�u�m�˗�X�W��{�;�s�k�����>�������<1�W|��A�8���fr¶���"J*s�&�����ΓEK1T3�&�}e�����!�U��~!��V�3�� $���bp9��I��0������K^���q���4~�#�K�n�àOu\v~�t�*-K���TE@�����x�뇮�et���Oh��' EGoZ��>��cl��Z�tѫ��Յ�u�i��UU��A�����-����s5�G��[V�R�{�s`���[z�˹u������1Mm��-<���E�}#��J�R"�SOU4�",�eN�8')�*�P��{��V�M�"e�nZh��(Y�{�~P�L	a�N)R�v��C����t�=.����;ܒ�-T3�zX�ineUh�00�q���$���'8�M���e�~�� �đ��Vז�6"�CU�R��f�O"�������)L��w5����g(vk_��t�ɮ)��yӇ�����x�5��ͻځ��<�Tͺt����$`?��������@�����Z��񫻊
��vJz���ѯ+�����_DfC+���f2I����ec�-���6C���gl�&�ڊ�-G:��ކ�âi��引QV��O��ac��q��ac��'��7�	�B�\�Qv�e,tO����1-��߶Sɴ(�iz߿\0�8��z��@�ՄP^#��13G6U��O4e%+��{4�tÏ|��F��wƌ��;.���QBH�*���(��������ȹ��l�#B����y��
�bP��> �cђ^���Uو�]��Lfur�VS�og��u�ѷ��-�|vf� l�����q��k2�A]���nr��"<�HP�`+`�����zB4L�T�./t;y�����.�.��`�H��_a<�Vph�j,�_��Ą�X�ֈ0V��zM񻜄D��uK��F��l�G{"�
>v����.U�϶���� �`Ͱ$
�*=���NM>W��+5��Z���ܞ]��Jq�*��l/Ѹ,o��P�w��3zI�n����(����z�:-���{p���8?��*v�1��~��3-U��s��[��Il�^�T7�(��w��Bڲ�`�ϰK*4�C�8*Lg���Q�F�6�;�6���֭~���/(( z�o�*��{��o��o	;���&���	��� ���5m�^T��*��F!�W��"�c�C�G�al���!E�T�/^�._K87�v�7���c7�^��y�4�xg��K��&��K�D �fP���x{ ���k��N˙T>U��ǒFPV�8N�,4���� ��q�5�y3�v,�Mݺ�'����e�a�}�鈒�cIy#B�c�U�Q�f(6S��DnFzz7S$_��Z1�\��`P�z�?:�Rd$b���Q]*xV8���oO�kP�ed��s5�tc�qM����q�ktT�q�@��ڑ�m�L�G�3�g�lڦ�\j���}G	�TE�xF!�H��h$�*h��PK�Eշ:�M�aH��YʞFl��_玳�r�Q�!��=P+L}�P�i�fp���Ͷ<O�֠�h��=��(W���"�b�{�	쓡��x��@�LC����s������S���ot�'��Q����t��U3~N�
u�em(n�2]��G&S̮��α#�t����l7�8��i\�647�o,�ч҄�s�m��t�X=�X;f(��4[���qo?'U�P�e<��
������=�$��8x��Kd����z��y��u   �*"��C�ҥ��[��b��Dq�֙�/�K� �X"1�i|٥�m~<E��;���6��bz�hZOk��o����F��j��	�5�?�3"��a����4Q�ʣ
v�s/��4W�<�a���g��N�N?�YWhlD|P:�ϡ�J$��.u�\����1�[ �I�^�{H�h��ec&c.9�=�6O%W�&7�(�$k��X���B�o�M��=\��U�eQ������CL�Oq3�R<Ed���ٮ�����H��Z�ú
��]ǳ�}9�4�%��y;������5k E[�d�B �P��/�����/�8�4�ࢂ�0$�j!��#-g�k�F-��߲���*#dU�3�g�2ކ�i;D�֕b��aX��ؑۘ���~;5�d%��tp��L<u�r���I"t��+��K��_OY��A&/yZ "k��w�>5�d�z^�3�wI����ʳ�q�A|��8�B��J�%�s��|,D�X��-�Y6,SP�7ϩh�>TE������EE����0?Z�������O���}�� Z������`�Z�f�B��K�c6�a	6Gl��m&��K �������G���y^g*R:����`{>����7�t���v��R�FK���]���ņ����I|(����?�Lf�#D7�zaSټ�I���V�'���+������/�[��4h0�/�O		���-�l��1����1��p���g��P.�Eٝ������o�щ�}��z���yJ��J�?�n{�a�K��L��y�Y+��R�9�"�"��m�=��/�_�"t����J�X{hd�_ $a�0��g��x)��)v����a�Uh~���If��K�g��m���4�n@ ?�I'Ċ7� �ՠ�!�d�g`��bQE-q]_�!��Km��̓��m	%rD]�D\F�d�V��	ౝ���s��7t���OU��5rژ������⑿���Δ�����0�\!q5z��IkuB)�A99��nN wkR�iD*�:��	���z�[n�<�hϼ��
�[o`�2�֒�!�_dZ���Y�XD��Y�p��e����X 4I�.Y�^�Bq�nOW�b�*m�'̟��)����~R�2���*b�o��XL.0n'���;�62�$	���E��[�xK�+xj�~#c�ᐶ��Lh��qÞ���m}#�vӶ�k掊�S"�M��X��D�ouH��l�_eT]�m��<��0�^���0��\����4W�ӜG������O��+�O�l`�5��3�޾�-�i����Ο]�ٸ��DX��ѫL��w#|(z��<iHѽl����a�TIA�XlHg�c�n���m��L��#�ϖ�9��߃�9�Å�Sm�m��T�n���뼬,2��t~�X�d����U6���$��}<�Ns������%&�qƨ��.����Ro��RM�+�ܳ	��8��:�8�=u���A0v��S	d���!��*v��d6�K��o{�)��m����B��S�=_�:=�y����y���M|.�Ҝh��2�I@����\�S[��2iD�{�r�a�^YZR��$�"r1��5D~U���#��pXj�-��q9I���l0�	��'�T"�`���t~�3V���/�̭�=�0���ל�_&\:f�j'	�>Cr�p�cr��wN��w�dM�E-�5c�UD�d���{��j�a^� ��L��o��h�K�L�UH"��@��7��$6�� �ǺM監4B�*�4:�5��z���i����0�;���V��^~��m>nE��ZħC�۾Mp=h�Ũ�iޭ�P�K�h�.���Q;�{�F126e��
��A�R�d$��58����3Si�y��N�'��!��������A1��&��z[q'WeY�F�²>D�pp`Xs݉T��\�����LY�ԢT�È��۱�GQj2| �˭5B���yn�/��:R�~V�Zb��fQ	��ŏzd��Z�=�1O��tL�Z{���>��P�X�=�,�j��o��Ρ&Z����Jj�#'���D�Atv�t�i��m���g�+D�s���9��Y6$5@���T�.'}�o�]��n6�ط�?#'bE�g"p*0�A�zI�$�z=�F ���SVEY��Ԝ�ˬ�k<�������,�Y��x�x�l���M��6�Y9����T���-Jj������5�k� �q�D~I!�D��72�eb�R��$C���%c��c"��'TK� Tkq,A�6Ʊ����X��Nz�^x�[X �#V���H�:��ɵ���c�����f%���>/�ͨ��+�I�%Zj�Тj��<�@��PVY~�P��
�^rXs�X���+��>�/�RݗF?�e�,*�s�9^��wkD �xn�[;xb��!���׀.t�s��|Y�p\�����m��~I��p�n{!+ �kW<�F&�\^UF%2�:f.�\$�֙7��?���'���$�k] m�Xi!��Q�vAG��\��dG�<)��3=t�	M.���������0��}|��Y�+���ǥj��j� $d"��O��G��Oq@�&M!A����b���c܂�3����g��ó�Ǥ��dL1�	��N'��[���i�F쉎�������[F��SP�'����`�y^�|$��6u\P3q24δA��z�������P�S��7�Ay�k2�B�h�ι�������S��oQ^�PdNY��q��$��
�.[����:x�`��j�B��Z���5�#�}�>L�].�=��O��VwY������.f|�Qg�e��Q_ʯ�D��4�B&���0ĭ��@V���7�4��g	r��kAtC
=w+Z<���@�UBO�%�]fy�bQi�-з10�Y��4�t۝����"� ���f�G��T>
��ӓ���dɁÀK7@!%m:T"�,v'�k���J��*�g���2i۳�q[�C��RLmh���~�ڋ���vf�ҪID���d� k�������H�iKČb�+�p(T��k,
�[��1��+��"�m����D�ڀ�bI3���j���=��&�)���_m���n���p�fBY�����L���򩢋c՚�xX^���v����Ie�
�L�p��u�UO���;�D2l��c�����&����|Rˆ^�����lɵ�,z�}Ȧs)�a��3j[3I$Ԑ_j݁&����9�Wř�}��GYxb�0�����V���)��7�G߆�b�Ĳ3�
D��q�e��:�kf�u�u�z��'������#�h��Ҕ�"�7�������R�lz`i��G�t,�ǣ}a�[�y��t��g�����������:LsjB�:i�Ngy����#F8<����]�-�=�/��^�}aݣ=��4MLS|<6a��QQ���`�â�)m5Թ�� �ܗl�t��r�(�h<�YT���o[#7CP�	�C%W�N
;��ĝ�z2(�W;5we��i��5���.�Z$[e�f�{�i՘˻��m����C^̐pK}�
H�j��� �Zq�G�	݇	�����Au�$��M9�]��K���x�ea:����:�6��*T"B���?�_]A]:Y-/��f�*�����;0f�4m��m۶m۶m۶1�Ķ�+�ض'��{���������]]�����N�>-U�~����߽�~�F/���$!�=n�hR&���>`�u�@|ǹZ3 e���}!܂�Ņ�*����q��,BI(��ez"�D�f'|z����X�U�p}��q7��I&���$e�pcAH��^��u�����^/��m����ݍ�~��}��uF�B��j��B�vP%�4�+�pRe��3�W8ü�������q�j�8r;v�~�)@��+D�5����8��Cy�xS��qB��n�#�]�pF��C���\��X,(�^�|5�PĶJh4D��/<��@X��Tga�,�HI��6*�e�:r�,�mZ8�w���aD���~�sF<ʄ1���z"9��NE�^��+�#**=�!ϩl�Hi[�j�pk�����p.��9&{��,<���1)SA-���-�O�\0۷=6�ҺP� �V�ɭGPc���:��U��gX�3qc�/�~	]�pR���.~e=E�KZ����=<�@Vp�Dq�S��l.�����G����>��ypMwh�J0���Hez�m�ӕ�S2�|0��oɔ�#NK��"���Y���IV��X���!ۯ�#�H®SƘ6Y�4MK�[rJ�e,cdD�3�Mh��V�Y���R;T�� ��E���Ql�4?����hZ9�E�rZ^E��� t��}�g�"�=.�EX��|{���pv��G�;���gN��q�E�Un	�PXƞ��~a\<v5H�������{/#��/5��=��)V�b΂�{�=���햀����cƖY���0G�*�0��A��yɧ_Ƿ�:�2�{�+�~H��*+z��u�_WW׷.�i̮���q/#$z[�`�n�s��2�1�p|o���X�l��J+u^P��+���6s:n�tţfZN�R�!�m��������x�`��cˡ��Lh���k2��.뉣/*�j�Z�`�g�G.Ճ˴�a�Ғ��z�~�񰀋�ND����b�ͥ;�t]�g�2Ը]��{X`���J�g��X pk�t �!V�g�=�H�oL�z
ɰ7������W��uth!�	�y����iD�߽ ��	�$���3p:�W9�~⮵#[���N����Im���GX�̃���~� e	�w��3�d6T�IL�v�ߓ�SӬ�T�5��)�F�qJ��F����ΠcL310SYG�����!By^{��{aBd������<��W����a�V.@*�]5�<�5��T�'�-{u�S�A9�(�Zf�rn0[�m�-�9|H=�;A�P�f��c�.��a?QyȾO(��:�@	A'S-7����La��w������ ɽޛ���r��8��l�p\)�n�:��X7�D��u D��c8�@;�y>�^�:� ���΋_���z��'�T5�����C�A<!+�*5��;5q{u���4w����<��������m�k؋���.�����LH���7!F����~��e� "���9��]C�7,�ݫ����k�\�0�k�Q^^��4��k	ֶ!Ε��ب�uL%i��)��XA�01�A.�L� �%��E���0%�L���_���T+�]z�.�E��↧�/�xY�7�xe�I9��۝�L/��β�0���2D��/jT��#fm�mDo a�y�ʟ�����L�����J��-U�}ҩ󏫆���&��vu}o6����~��6]�z����z"ܖ@5[��5���M�<ϰ-E���4 D��Ď̓����-�1����'���ޖ�cs6�Y�{FO��a�1�s�S�V?��L�̲aaH'V,Xױ�=�c��cڔ��	�`=�mN�l����z^�{]DM H4D�	��r"*+� *�-�n`�zp�iX��6��s�?�jAbJ�:��ce�i�	���K�N�D�0�׺eu9�ǌ��;�0w�����5��O������Y���(�թ�wST20㰶�m9j��
�����7["!s�FNa��rh�����U^"��[�����E�E���0G$������btG��� d�.�f)�W� ���XB0 ���|ex.�|��#�ɮ�)~�؋�P
�1B�;�P���4`xV4n��O�*�*��>b��:����`l�n�7d�=WH5/�y8�ҋ@�p0ځ�,U��N\�a�U2��uwr5�3%�3��;�?���Y���b���*K��ӹCbɴ$U2�����uGZxh�Z�*�*�PvVC��K�n��RٺՍ%�eo�&���J���X0�V��r��Z>�
8(×!���).���$g\���=.e T������jd$(F�e����gG�WQ�����-W<J���;��l: �+�[�Vm�@@1�^�"�
]����`�~��^h8)]�O�`�����e;�3J�g�-�a�>H���{Ϭ�$n>�OI�~NQ��#��`����N�VN�3������B�|��q�Q�)z���z�ȢLy�E�&������1�9bO������6��f�u�}�{?ϼ	�\�����ƑS��jF'3��Gnm"T���Õ�����ߛR�!��s�����/��Q��j#�u[C�4 \CC�����xDwPw�"e�Q��L ��ٳ-c9+�rZ��>�ww�h��t'�@�o`!�_�]��lm�l�WRY~�2�ݬ��J��� (
$����$�	ƾ�b��=���9�6y �'�{�$�P�����\�V�V���w2�iW{fү����i����{B|ՙWݵEH�A�Q�<�(���υ�	X4i��b��V�7\H�M3V��&����O5���6�rnu�H%q���˔����ї���1+��A����@5�:��wZ�o���ʒ�r;MM0���^��9��{^�����8  $[| �t�5(v�l�,&n�&�%)���a�߻͸���;dxz��z�)	x���.V��*�øj�YgA0�}`�,�v���ƀ'�6�!� ��f���9��Z��~�;��,Ν�+4:�_6�e�������}�qDo#��82���wD���`�r�C$�>
��h. ��z����4���E+���|����+�2K*|�:u3�9�f���)�Z��1g�y&f��n��5�r&q�>_�f��5�W+RKE��u8o����{��Z��|I�P誙CkYV���mKF���(��1��`��ٿl�V�5g�xRs`�^L[ߓR���RyF)��Ie>U
��X�@ U�	i��x�bi��U��jQ�_M �g�-�?�5<7"6��.��W�D������2��a����p�7����ΐ�Ú��cu�WW�����{(lB�y�}U~F�k�բ0-�b7�o�H����`����@�
l3��pҗ��{iw8v��Akd�ް�9�q
\���D�ט6�e�'�t�UD<��RQ�[��G�-@�A�w�Ou4��;;�s����q}{[+�n�
�혂>O&�l�T���eK�_.W�^|��S՞�6������#��	e�
��9jd���z�k-t��M�L��5.�T�d�
�s��:�&lY�5v�$}E�U��C�ƨQ/��Q;|��{~Gy�������1068��]l۾�z(�d�j���uN_ӳfF�t�x�W�{ h9Tg]�	 '���C������m��.sL��������������j�/�D
�I��1l�Û�#?91�T�EqN	��05����jw�'`�BԎ��=�8i��慡��ÿ�Y���e�ղ�� ��WJ�$��)֋�ʒ�\�J�@"�B�J�خ�������cm8�1��N�_�
�z��Z{�;,�sc-���Н�J��1c��`Y�!oa�׫��� $�Ү��u��_^�-����8���ޅ�\����"eh�J��)���ֹV�����q���׮�q���kt N�*���wʻ;����
<��dPҲ�l7 6�U�h���%��e6���^�q`��u���u6Р��u����2���BqT�Sޚ
:���o�pK���D��XӞ2�2��ئ�z��ap�;���	LoC0f-`u�e
 �
�����B��a�ɬ��V �A^�b�s����,|Ap�4f����s��O�/F]���`��5��Z/�L�+��cH�K�D�ݝD���!�-�5��t�-
�F
8p�%��>�����E�(p��?�l�#�+T/�AT��g��������98M���b��v�u��P$KF�>������ɩ����a	/�.�!���P̰�z�+�O��/8Y�>����K���D���ɇG#B���f����o}�ϧt�X܎���2e��>�y8ԟ�x��xgU�"� ) �/4�b��f��	������S���5)���*��Џ_��7����)���e䇫)Ji&ܒ�-��B��DƓa�����P[��温Dm/��m`^���G1���}qt�$ ��pX�6K�X��󈳠����03[����]����TP<�MvV�CK���Xm�T�����Dx��g�q�G,��c�g����z౟O��T�V�����`�+�Af�=N�
���k�����\"�C�i�}p^ʰWx��Z~4?��^�#V@��C4�������w� �x@lfƝid�����zm����2!�m�M	C���u���e7,N&����zd��oO�+���#��Z�1�lEU%(t�)�!_<��oy4i�(z�o��rYGFŃ�����&ewG��6�~��C�E<�~��I�Qx��<�Q��,݌�������O��cs�z���������/��w	=Gq`X�Ǻ�<%���Uh�7�=���jEG>^�e\����F�3H�B����<��;���d���%p�4>mh ���}��ylXWX'b��1�9�vpM�a�N�Q�E��4����2t��:1�2wD߇/��6.�;�)ː�������jb��dad� Q�U(yS�5�u*|X�n��~N^���p����<�{� ������M.nĽD����#˘������ϖ�$�� )��-$��t�տ�I��'��;3�7r"�;�7�CS�^�Y�y�2�k��;gI��t�`�:�.������/ݑ�Y	<�z8����Zu��>�M'�β;f�Cϰ����t�m�v���|Dt�	s�E�iܿ��_���=0���e�M���IJq���PÙ�s�M$'pᭈ�1�iY�'���E<[p��ϟY�	E�����bf�������?��	Z�t�T�3%��$��	�`�nn�,$�(���s��$��E�����;�Ԯr՗�z=w�4m�n�x��.�?�z;��ǎnCbh����Κ�-�+�#��""X��O�K�N�� '�w�jz��|N�`/�G���j���ƣ�������s�q�1�@`n!/qI�2�����:˸���|!��}'k	���(�`��˴3���NȄ_�Wֿ��aH.�
f�u��y�f�k�fgccc�m�~M�f�� ��:�N�	J��wf{��a?M=�1��$ ��FX�V�8� 	k�f@�/C�X���J^lkw+��UA�������(hkݬR1���mj���=��ӕS����+�i��hEmӡt�h4*���o<��=��_l��(k�2)m5����"j7=r��?��ذ��J�5Z���
=s43�Ƀ�adi6(�`�N���T}���?dׇ��O��[E��w�tNgP�Ѥ��/w���fJ1��?E����1ھ�n��6�E�^��%�|-�i	v��
]~Q��c������F�L'Q興��U ���r�:}\/�ݻ�L��'w{\�|~�R"����af�S1+��>�-wq���tN�<�b�ǝ�,,��N/�<��q�E�5���ec�4[='�v��~w](�*l���7v�����W��aV�^����:>歸u4E�E=˺��9��+
��}_�Jw}eHrӡog�(  �[-e��
u\�q�J*>�20�U�Ee�p�*�p��N�7>^,���:���Gۦ��=Gr%v�H����h�"տ�Q����wc�7�m���^V�T�w4C�pkjc��������
=?��6��.c�>�-ܽ��k��^�������tW��5�\{�w޻�[�P� �6]��gN"8�M������L}���gBhhe��0L��ߐ���c^^���g������!Z�V�PE�~S�Tq~.=h�܏z�i� U�6ԧ��g8�0mzM��t�q�lǘ��F�z:Um�9�^H(�����[���	�d�CQ�c��~�l���D
���%�y'tډ�)�A��,m����u��<�G��rZG�T|2�����x��;�A:> `5D�X�z���p��C��aVݥ5u�Ox��2 {X>����6He0Nc-c��/�N���c�Ͷ$������B-��@ES��H�������x(�Bf`C>��!��PD�@��L�=���+�e
����w��[�;b�u�%�
-�D�]ZR�W]�WuO�����M���k:x!��v0�{���2t�� �����{3yF�,׸!˾�Z�sf�5������u�f�l�!�M-;����h*�m�T��\'j(�2L2���r;ﻝ� @hZ�R5|��҂�������+:}:;�����A�l�m{�x��u9��Hm�x�F�?�8�,tΧR��?&�p	��ţ/��]�q��V4t��j��C��`&F�99���5��O�\&ǜ�zo���s�~A^o����{��������6�
�D!2�oI���d�I�����r�'ᇖ�azS��D~��s������b�N���2����j�"�\�����R4(��h�_�Ak����ʕ���<���G��E��,] �� h� B˰���A�����-���5[�+@�T/RH�E�N=�'k�>�u3��OЇv6�6�O�P���x�a��V�����b�YHjy�nK4>J�'�L9��D�n$ ����H�����>���
IGCM1M�����l�������ec��f�����2	�O�Y��TLHP+�mv�5�_b֗�(��{<&�3�A_r�9%H?�~��	 �9?�--�`X�15�ev�#N�R��`�s�.�k��������=�{�Z��Ss�;`&�W�-/�EeB�z�U6��%�l2{�GL]��-"lî���x����Umv�1�hݲp�a4����M#���grcK&���&Y�M�v�e �L:���ݽC!�m��m�G2�Y�gҝ��������K�Z���5%��t�.{�/���i��y*	;slm=5)xpJa�B�2~���D�B"�����W�|6f���fe;���Z7$�
h$>��w�*f$��<�Dwz;=~P���V��m���U
�<�]� �^���-��('��8P���c�^�����2�����q1Y!
���!�,	�t0�b�ɒԯm���g�d�?�̺����1V�Za�Yw����û�>g[|���1YH�y��;�F��a�M�/�h�@���,>\��1.�r�P���%���v��	6O����c�+Y���X��(/a�7���wBLǆH��\�{�@���S�ޖ�=ns��t�$-/�Gź!��R<��#�Gn����n�"|	�9ʹ��e��Ezܿ��cj�m48�����e��-(۝�Uu��1�!���h��:�ڭD�:x"�z:h%SCO�[��U���Je"sd>皩�ʺ��}Z�a����i�1���Zedw�]$�b�y����8(n�"�]+]"g�O^�� ��|d�dA�2���-�d�m�d4�y1�G�ƙ��y�/S�書;0q�$}�݋��WJ'ׯ�B�B����J�o��������[��%"8pX.�%��sn5ĭHݹ���2��v��U����"������|8:ϯޤp{�(F�6���C�������O�0/N�c0��g�^�D�!S��|kl�.b�g�_��mӆ���
��غ!H�˦�ޗE��>�V�EүJ�Y5X���z��� x�jU�6Q�
��Bo��$郴���֝��'`q���m:_{���<�z9+!_H�Ra����L��DKh�~s
L��S��ʑ�i5�JGGG��݇��`�tG�����:n��p8�0�$û���N������b]��2�=�'Pf�AA�hk�".�-��T�rA��!�< � �G�/�a�~���?�d3�&�����W�Jd˳cO���g;�r�	"�!S�+d�M�c1;�r��]�5|�&_����FV�\|���~�i�E[��1�}1��ڇ��,����>?��K��酣L�}�{������G+��F���R���Ҽ���؁�d ��u�窞��=�z�j�������l��A*�F���
�i4��׾��BT�6��[3,�����_�c��Vު��QeGV����jo�̀�k���E-g������A:���Q����
??+Itx~0�!��[���r
��4���m#K��7?���0,t_��I�>S�k0�l0�I�����%_���*��'�0>|=J女j�2�"�
sC��%Sa\!�&�QǺ��#����E�j:���et�9�#�zkɧ�'�(���c,��+��P�m�5�#�o{C�]iP���,��F�0g�x������ݚ�ON�mA"z-�Cm3���B"����B� g��U�m��[��
Ҍ�@J	�l���.��_�哽)H�\(<
P4����~��w�'�����w��Δ�l��<y��PQH��x��R�4�0��<��YT`eQ�4�	qYX�v��7�o��K�K�q)�YH�nն��ӝ��g4��IǞ��.w���<n?��m��)�$^�
�
ٴ�z����	��=�vz���G��|�Ǯ���V���s�k 2h0�k���q���B>����ۡ��&�28k+w�q� j�M���^ൻ^��t�D�=�`va5�F4�6~$���:`��3��a�[��|z�g�O���{"����,�+����&�!����9J-W���m���$���R(���-��^�q����	�56y�O�ofy��E.��(�J�����U�g��)i֫뷢m$g��<�,���Z�M�����6DU"\|�,P�?�}��G��x���S�g@������ܟ�GX�ڴ08� 4yC�Nbi7�N�T���[��i+������T���ɂ�^�zb'�<)٫�bz��1:�X�.�KN��Wͬӗ��q`E�N9�OÔ����7��d4g��.�q�?yc�>�N?�lW�0^�SB$\�5�i��Ի06����_���C�?��a|�*v��*>�@�Z�1Z�/�}�	V�E֤�����0I�s�)ˍ����t4-�?:A��IVA��N��F�yw5�-�? L��r3�vO���2���h�u8T��M��PO��J�Þ2�(��^?!�����T��t��������%E����3
��es���9����o�?�h}�zv�VtcJF�����--a�f�:��L��{�(�+3+����慍��p�����2�IuP�.��^Ii�M��G�@Vm-�k �iT���d��ߘp�i�m�G��=8�6L�ܶr�D�-|h���
�j�&@z���\5r��@{Yċ?�C�3��!�ǎ;��.�	�"�q
e����\�'�Y���帤���7>�9���0'������~�h��y�Ua������AiE1�Q6��+_{���u��y\�R���7��a�G����H!��y�����t@YT 6^FݠPF����眜����w~�l�QO�:TA���w�ݯ
RO'�mi�($C�<R����*�ۙE�kC-DEN#��5�}��0/����0 Υ>� qKT
@5�X���CN��P���S-��A=]Y�!�U�C�l.�5Yr

"�*6�ùTI_��t>�K����C"���2Q���/iz��Z��Ȑo�O�u�Λ��e������6�o}�]�3e�`�a[�"��!v=�s�(>m6?�s�>�:���S�������k�m�(מ��<���g�%i�����ur�s.�?d�E翗8'fE�|i��*|du�E��&ޣ�8,U�׮��#&����Q��c3FN��tȱ���qDB\���H*ޝ�)�Y�td*��\~��d���C��씈����&�vӪ�|d/~�F	Ʀk������c�K��.�5��]��ְ�0s�]�����x���n���-�3�Sk��d�nw`�"з�i%+6�'�B�	~n�]�H����ς�����⛶чYq�b�u���H�L�d�X#�L�]� cTB�~v<.�z�����B���MĒ!�R^��|�L*��$��Ԯ�&��[k?�W�F����Z����*�~��3��#i��;����[�@��H�p#��Bsr�D�������>�?N����MB�̐��Pw��Ÿf%2@���c���|�ύ��4�h�W)s{�l�h�%����b�%�X`b�m�RM��Ó�4�g~6��N	C�<Uv����_Gm/@i�H<��ÿa=YZO��hk�{8�a�Kr�¹�n&%��OVhWuj{{�V]ݪ���PP2��%��]>�5���s�h���
a�~���t��,���,�?�0��ٙ[�sN!���)L^tf�?ܠk#]���?�?:'zS�;��5�K�*h�����$��t���f�M[U��o2�Y)[�|> �<ͭ�y�������l} �����v];4Xs���)@��V�P8鋷��
.\�[�<�o��&��$��ZTg���.s�ʼwҚ^������)�I&�"��I��`�]���`��	�v]U�_����ē$NQ�i����m�3m��O���.2}V)r�u�y���ەgh��O D��x����x�D��8�FiU�2q�g�#��(���� ����2���Nh��tkK��<0�}\R�6��i�GS�r�T��/:"�2z�_u`�(�������$-�C�'�xx�s��A��Ὣ��b~�"}�����c/v ����o�G��`����@��v��� G��d% �&(�����'O$XK�eC��"��'ߝ��$lsS~=I*1.�ЛK(�\Q�&����>~�r&����33�"���?�Z��^K��p���s�O������O
@�Ŏ_2��Ax6�Ȳ�����U<���������:͉�%.���^���YF���o�'6�x����9N]�JsW����!K���N`�T�����Ȫx���AS׮����-�a�JO3��栛aQ~<��]�)1?\(�^r]�@F<�V1���x�}��q���F.�l�9N���_d�m�H�8?�uP�/S����<��QF7�=��J�0����/�B%��V��t޷.ަd�*�t*[�u�������_>j�-��yl��!w�C��95�
n9AV�d��M�\�.�V�.�� ��ή����z���J\�4R����#�W���
'jo;�݄+�p��ݔq^֢�n������_oz[V�9�;'�he���t�����I��ȉ,��<���6-�� NYIY�r�g��,(HT� �ċ�K	���Z!C��W~��q���c�H���W@;S({��ն?ﺿ�@���ɖ��bF���K���&S"�p;#湟[mo��D(T�O�>I�`���"�\5Ԃ���S7�B�v�7�'�ˣ;��^�K�w��"�۪0��.8�m�ſN�sh���he��(i}�؄����E$�P��7�w���nO�9c�؉SC��M�����%,:�\�?�+8!�>B�J�e^��6���u��[��(���M�\0�;��HaJ6�S�?ԯr�}�> �#YrY�.�����l����I���#�f�u��aN��������\�;�����<�M&肑&������h�����H+�O�?��B��T>�FNa�W-��dA�Ѯj8�}�e_�gFn�fw|���dre��p2%u����T�?�KN����E�	�0�.°`A���Z;���L��d)�;�R��ǯ����-x��w{�����g"=(���;���m�� �	g:�Ҭ�&�6!���s�Xi��,�!&�N�6���B��oI�6��>�1���Ӹ"��Z�N�힂�U�H�鹭˓�-ߣ�hԎ���>`��Q���o��#9�6�+���K�r�%bᕔ���*��}*B��� B�L2�t��ޠ�b�{�����ۚ3��s�ʴ�|�_������-+L�L'i%��>�͌�ÄE��H�1����m���%2�4lg�z�w�C�?.(l�9��M�-q�~��=��qc|(����s'�̏zj��9����@D�S}V	1}´���v�Uw�{&\�Gb4z���eu��a�_*=�81>�A=��eH������s�}@���X��9T	�ן��hM��m�k'Q�@�o��:t4��o�P[(/P$�I�@�[�S	>�|�x|�H �7@L�����7	�
:�ѦY� ����dD�"0�R���O2Q�G:
���(�U�?�ȹ\�k���gE�g_D��?�s�-�g&����1�Q��t�>G9EӁO�Њ���ʫf�0��}��x�SO���)��X�������C��T��KaTY���+��-���Ǟtk�/n�B�8��7��266=Mμ/�N�`�5
�ε���5w�[��:u��r۟���53��C��F[�np|�D"=
Y$����~��;���D���v��T��8I�u��� aV	}(�;���5��p��>Dfz�ʙ���DXl�׬n��bv�۵#�p]z�S�"�U�3"Rw�k)��V��  �?�B��o����kT�j��5���Bz���A��͌v���}&}ppj8E�ؿ��C�_��b�z�UaQeI�)��V�0bhYx���Cq�h44������Q��!x1e�xx� �L���.㜬�8�x�HN�՗$%�ws/'��[�n4�s^՜��t	Z���NîC��z�w������M����m�-|�>R�x���r��h.�DP���\�Z�Ŀ��ܺ�����,�H|�Ɇl������*��o��o�E����΃�<�E����~��J鋖��0�BWA}��Z��,��eP豥��.@7,4@���ٶ��#�D�0BvȪ"w�(�1�Ju!��8��?Mz�����%��IPȴ?�˱5��l�#r�#\&q�	9��4*�f�j�2���~���ޡ�~�	?���x8�dM��z�J�ɸj�G�x����/�5ʠ��N��M��X>b�<0?��F�˷��b?�G$!!��(���s}���Q�0���1��9����{ֶF���o�a?顷]c*���IF��I
īM�0Ձ����̟�G?�Gn�;� 2:c:���6��?3��?� ��2W���!�4�P�����¸i�O��J&�%�IaG/�c�uwvsXzO��_W�]
?��\��`2��E8�Ҕ��m�}-�+{+;;1��q-�z��U����� &��׾�o�L�����Ŧ�w�'���}π��ď;���Ycol���}rj�Ma��]�鳒����bڬܹ�<ݒ`6.����7�o����@����d���I!>' G4'iL@��g��z�Q~��0�^Sf�lf>�զ�,Y�t�]�y���2����"q�!T���>"��iv�F`��#.�Xc�_�T%�[���UţI\lȰ��z�I���)�M x<���kf�ݸ���y����1;����}�N�b-�8�O~(e���$;a����t9v��wl`YE���O�p�Kq�`�B�b�Ǜo�}�׀J��g�B��#�e��b<����x���a�?|�x�fY-\�KK�������GrzZA���ĕZ!��ƴ����(߈<�r�Uqv�&j8�O���4^��\A���������0���M�A�,�.|X��p���U1Q廉:�y�̪���-B-��x��g+HO�K'c�����l��eO�x��Z0��� 2+���g�0��WF���-w��ۛ+ۀ�j&.rH>�Ն�|�b�AY�E��\�m�O\6'��[+�am�}G��ӫ3WA~�$��Jߔ	w�k���*��m���jD������b���j�%���j[����qzB�cH��Ȃ`埭���������&���K��׻r�LWN�tK�;�b%�04��9���\6)��id��@�V]��L��<�((��,L,�{�+�i���w�,�fS��+0��/�DT�B����Bi��B�����&���V����Oۃ	Lñms���4�ՓB�B;�<�B4�(�Gc=Y�_�&r��,�ե�i�w0#:�\uJg��B�{����`�	�(OE<����۩%��)pb����^�\���f��j�)]!��Iژ�'na��;іd$�R�i�����r�m��h8!�5�?��5m��� `�k'��o&m�7%<̦&����V����hڔ8�\�^r{�_:OF]+X+32�:�8lH�s��nטvMq�x/��sZ�f�a�vlCK����?LlX����.]�������C[�q���
I��GL��ܓ���\�Z�i[e���@Ivj��--�N�鬜�C�X Z֮�k|T�j�^�.f���)���q�A����R���L���2D>��51���\i���Y�DߤH)���*%]<���>������Ncm�խ7(��Cl�!h٘V����D/��:r��5&v��;6I��9x�UuW[n���r��Yz��݇^�։l����N(����{�5����H濲��߁�B1QX�`��/`��
C������[���g���%B�����G:=��c��l�X'a����ZebDHD~�6��� ԛf�����&s�^ɣ�F�5�l�减!@�6&AT@ZD�\��(J
�<�.I��,����k'���w����)��p ��-���C�lm�n"�nxؑ�t�*
2v]�T��4�̄�N��f���p#?�E�K	�ix9J���G�G%]�mӈ2�~?�^ }Z��,_����q'��/a���RM�>�~~�eg�g��):
!N�UR�YN1�P�đ۱�ަ�
ʅ���>�Y��[��3��oJ����&����m�P�.�ꇬ<�jhi+RgVh�!.�yq�(��6�G4�X�q�Ԥq�0�m��fzl��8�p���\#� >�y�n*�׫>+y8�O+��>;�mb�I��>�ϚXEA�^]�y��۷��pJ�9����q^z%��$��%5nϮy�T[(�Є��C}�ҦZ�Xe2��M�,�tu�{tAq[�a@��~�rbr/#]"��^�ٲV)w����*2��MN���.VR:����)ݯ��{{�Q��R���������klL�˨����Ҋ|�I������B�s\S�J&k�=�T�]4?����FŅ�}�Dc(�lA�1R���9x�͕��1�ᴮi2�#����R���Nф����O��--������W��.��^�@���#����� B.���t�#;���k�?Z��o�W~�vwclx��dY'T�Te\XK�������i�Y�:�]@�I5�9�жA^�W Z�UX�Wi��$��B���� ����8�T�k�L4�)��8�ŭ�?�����	���
6U�9\?�C�Q��3���z!H=ZNK��g(*B]�:@FH���k��H�s!����#X��VBr^+��@��:Q+��fn�K�VU�I���^Tg:�����i�'G?��,Wߝ�b�N2ߕ0�Q�t�lx�q�Z����D�*��8�o)�Y'��2r���M� ګ�uk�7J�1�Ae���E�lKj�.&�,/�OC4F���y.����;��uO/+��0�/X�	��4�yX�Mڑ7 �:n9^q��2P��D��'T�^� R�����y-%� �-�h�Z$'%.�D��.]�d]��[yy��.���,=��a\<X|�플_+0�<}�i�������� J�!�\�eeޝ��y���)e5<_���l!a�F�m�­5К�@�^�C�)�l��;�R���;Zf���Q�O�#�.뚀���?����f�j������ 곁?��T�AG��p�?#�.�%����>@��������1R�Q��!l�)��Iƾ���ĸA����ͺ��ٓ�ev�+���M]Ӭ�C\�$��5l?y���ɮh]S>L��#~퀾-������*N��>Z49@XN�ir;f��0"�Gu�Wt>�����<_B�,��1�k#���6R���k"L�d����ox�YZ��D=7\�/D�/>�8v�G�n���6�>u,��fڑ�3��z�x˴�g4���8vw�{��"Ɨa:ר�v�.v��&p��D��"��&fW�`dIU����I�ÈDKUnm��v]4�~*����([z�tJ�Q��@� ꖡ��8�0NCW9b|��j���T���@`��Ҕණ�;�g�W?�6�2q��ov�9pl����x���4FCuJ��#?�)��ưOk�͛Vq�
�)羒(H�;h�찰��a��V�˅�Xh�$xS+�#xZ}3̱��#MRD�ױ��(���z5z�����˯�;��"��7oX��=��1b�u�ҿ>��4�s=�7�hAE�g�!LÂ��U
�oNi⨑�M�ؾ:3G6�lC�AF߃�&�B%�y���`༖�b�-���,N������C�Ԙ�p�c;
!��,�p�ݩ��R���%�����U*���^9jA-7'�����_��}�"B|���N����.:�����Gs�5?`��%�smZ�R~N�D�a��6�}w� �>�9�r$����4rX�r���]��Z�v-��UU= ��l�D4�b$Jd� p���>	��eQ��i�u]���ĔѮN���39gQ�r�l�E�F9���/�ò@��?Ώe��V�E�hyZ����]W�KFݏ�oM� |��߫���g��i��X���I=w��֘Ll7�b�1<�19�	9;:�g��6�B��M��6���)8:�I��/%aQ�u:X̳iEA��h\��M�2I����
o7�;m�6�`w�-h�F*d]�	���'�+
�!�2�օz���Ӽye[�E��l����9�C˃�*^��`�x�m^���!�ׂ�־��=�E늙sԉ��SBb=���s;��C�2Q^�:l4u��ͱ��Г�UF���,s�\��.a���H*��
�qDk�Ǜ[	�~<�E�ָ�&�|�%�>J/�iW�Pd~5f4��韶M^���%�,�،LUV��B$���?l��&�퇛�އ_����7���p86���ׄ�o���	֗F���ށ6���ؑب�U�	9W��̺(W��AW'��G����K1t.�9��*��B��Q;��$�s�"�"�&v�,�J�"������sp�1;��Sq٨�!_7?�{+|�5��*U�&LϠ[L��f=�s���#W?��p���W��Ϣ�����{ʡ�l�uVGj��G����6�X�aN���Ba�b�C��'��M,x�kx��M6��7Pm�E�Mv���`<��d�x�9��V�,��Cw��#�A��X�R�WJ%t�rx�jmH�^�՘J{#ћr������9Kk@h�8W�W�o�vD�~��p�E���s�T���Y���3�\�B���v�iF��:�Mn�������?�CX�0�}�y���S�e�\
��%��s�3Q�JjS���j��8m���h��˟BX("Ŀ|4��Ig�v��k�9W��u��ж)����Y�ZÀ�8:j�ڹ��#p��nP��·;I���G�� �a��m/�!91���/�"˅�b�G���8�ф\TO�/�<V),��:�s�}O���O�*�V���ɊU4DA�����|��e 5��D�O*L��L� ��y8"	�s�~��^�$�y���s����1t�f�꼻����'��vO�4x�:eVݻ�����F��y��E4��N�8��Hb=R�5���tC�&a��AUO��C-S'w��:��x��BD�sN�0mKE�p	a�j�n!Hc4��j����`�i�հʠ�8����*����(���8�.�V��J^�e�P"�ĉ�|2���h.R�ddO><�Vt-#W��:#�:�x皠��I0p�Ǝ�s���&\����rq��'�;�Dte��+��!3i}"��sX���9���v��V��\"I�82��s@�݄$��B}�v�Q(Hi=�>d+q���L���ﺔ^2R-w����p���1��{~���)X�J��BXr\� ? ����U��䶠F�gSc�_�=���_r�-Î҅���Y�	Z�Th����-r>�J권z�x�����ޒ���� �nd���(|
�r�T�U̙7m�UDa����N4HD�$܋��B4x%*K��k}&9K��ng��� 1���E!
s���a��d�~1�T#xn��V�q����\��zSQ��R��8���D�BZV��^B-!;0�>ۃA¡�D��7�Uǩ�����}^��M�\mvqǉ�~��涢��]�tgb�M۱��XD�^-hh(�s�+[��g�|ڞ��`� �,�4�)|�D�]�v�_��x���W��a������_�q�l^	K�{y0]{��1��E�7@�l#%[��f��@Eq�C����2���c��B�C"�l˶Q������^K��ҺRƼy�h/w�/@ǉ��T��nA�~�T�o�崞�q O'a�Jx�I�>vFj1���B��Osh����MQ���Q6>�v0N�í�D�e�����;cЊ%d>�5�Hh^֤ [���i�\0Wm�r�͛��ɯҘR��K!���Ày����sox��f\�C����Pq�0�'�Ј<JQ�k*�2���������~��^y_
l}K�����Ŋ}L��󙹨�19GB?���S��ih�S��0mWG�/k!�{ç��I\|8m&f̜�����g�M]t]>����-�t���a�k`�A}���~�㤞_KO���%�:�`a�'(�ա��\[>��*
��s��F#	�ۮ8��3>��K^��%ر�ީ�.:��,���j>�HP;�E��EX���&��Bb�PU�y����i��fVC	r���̙�0��xi���8C�S�k~IYs���n0�n8+��U�D���:&�m��FY�E�P&�Xѱ�F��痊� T!�����u-�-���/N�Aĸ�e8�j@��ʁp-�4�+�ӥ���y%בI��v�ZkT~���}��^14�s�N?���̹����x���xmrGT����6dѧ��p6�`uЂ�+�R�j}qIpǑߪ	o*��h!��	�N��к���h��Xep#���p��Q�8�o���fĚ4�GT	Q�[4 8�!�-���zj�B�B���[n�)��/��s ��_��%��k����q���*y^X��賰��+��٨Tj��J����eXܯ�2?�gG<��U����p�ؔ�0�L+�VyZ�^Ip�bfX��$*�^'��C�G99�%L�p6&O��kn{Z�f-�O��Bɭ�_�<������v^�[��<�i 	��4�q���������U���m�<ٌ�Gn�(d��t�~μ�VL��*>��uK���Ht��e�	Pt��ɉW-���o����ָ�������Un?6m��3e*F��uZ�[.�_�[�^�҄�Ս5��?������Xs�!��CJ�s�]G�'�*��~� ��XS�k���q�f9F��7]y$~v�u�D�K���q�i���l��5b�4>��I�Ҽ���Z_l�v�Uc��\�v�)m$��$������w>�ݏ�E}�v1Y��Hs�q���Y�Yï���2V�����z=��9�<�\�
J�C�=�HqP�R�^	z2�͸����Q��V"��������� �4� B��Tkmh(�G{{���e}���>�]�	P���/C���3��_a����� �!qn9�n�$���m��G��[0d�]$|�q�9��\�ˠE����v	~�)����q��n������_��M%r�3a��I<���Ud9W/�b4ݚ��h�O����
#uItT��g���x��K�[������G&�U瞸�[k(��|D1MG���H�pU\>%��tC�T�nJ�Rb��Of��.ん�ž,. �g�%�͝W��5\�3�KꄏT8G��-W���a@s�A��H�i�fk�,o�?���/|�i�c.���߅]�QA�ܿ�8h7��
�s�7���Y�(/ �ld�Vh�\�Va�i��ŵp��?�A��ElE�ʨ9��S�$A"�=4O�6O̡�P-��'���"Ӳz�Ĕ]TQ�ֆ�?ι��z_�����������8p�-����h���g�����z{AD�U�}���8��*I'��!��p�!8��[T(�����W�s���R=�Tf�FQm�����K�c��r4�� ����{�� ,"ėn:��Q�����?�
��4)��Ļ�5�_5r���>��!��Vh1q�A��U}R��o ^�.?���ԫ�jY�rX;�,*e$	l�	A�N�܄����I�<�p�L�����~տ;װ=��{���E��Շ�F�A7r�Y��z�z�;��rH-ș��-�T�������p��� |�^n��0��d�K뀎 �ILhd�����r�NO�#dY�"	�8k%g���
q�9A��B�x�<�y�M*��3�ŀ�6\�?!� a�9�Z
�6;�i�(&�qw�J%\s����i�dN�d07_�+�V�9��zZ��$�3��*��p�Aͅ�Ӹ#���蠒�a�{�8�ռ�u�/�����3�����C���CwE���F� ���1��E��?ǵUtX���a5���+�jhnvp�Y���ȁ�7��G���kD��U�H��	�i��#2�kh�33U�Hh%�~��������/6"ĻF�\�w?��8d@q#�x�ӠGI�*Ъԣ(�+
K�ONk��)	�-6^/M�qo���V"��EUG?rPT�[YG1�z�����Ri�*�ϙ3�U/�DkË�>��<�TW���n�V#�������vMe�\L'�Eõ���O�����Z5$;uH ���_p(�<�F�-,l/��qZJ���#CU�7�����-�lr�I�$-2��*<U3Z��?_�]��ƝsU�=O�s��~;m���ݘ���[I�$q��"S�h��m���pM�z��}p�E� �v����Ah����՝$�u�U�9\W#XEC9�q�#�r�������������Թ8���p��������cr纗��ުҵlÂ��cv3�P;y��59��:N����u��9B�z�(����-7]��N~,���gy�Xd��IV��7�a��JWs2=\��؈��
|x�y}�W�r�ޖ�F\�9�UDn@9)Y��{�K��q+�6my��7���w��Z}]�b�������&G�[�uV�U�o�W�)y�!���B_���Y����ݤ�B�����h�y�C<3�j\t�O��jP+��D�#��
\��P�i��j���$@rz���G�\#}ƅE����}6��~L�����i4�:lbn���A����c�8g�%̘5G�{���
��nl<�|l�t����܂j櫖L,��{>�dqğ���������&��H����2/_�I���-4�r�j�,���P���fo�s�VN��x�) Mm����c}��FZ^���wխOb�?CSK!��yj�`���!���V�S�lMUVOC��a����i�u��3oJ}��	�J8���(�ZǱT9�z��������IY�0mZ�I��i'�sÿPI�Q�!�u��m�K����N�[���$�ȩ1��F���J#�Tڛu����P3��5�$�͸��?G��/ҟ�k�[���V@R��i���|J�)�Ua���3R���,0�q��-[�˹�S.�;�9x{l��z�H�� �pB�+Ts��8!a�թ3��>Jf�
[�x�հ����k˪",�z��~�`&5h�I´Hs�����l���|�LvdZ��5��1\������b�f�s�Y������ [kA���I�z�r���N��{�	n"f͕n5���t����ƫ�J��2��2?E���U��j����h��dK�=1	����
E_��G�z~�>Xg���jm$ ]xܒ5	�y�j+2膥���0Gq�c�o�Ǟ~S�w�x���?��M¢�d�@�,�UX:��׸�,w��D�w�(�R��ڞxf"���C�R��!�t�s���m��U����̒�9��ZCCj�vh�a�1�aB��c�^�%�S𫃷��<a��Kҍ���CϊH�q�r��p�����-眂zS��k�����G����o{S?���%�5M-M�[)�Vj�� �U๽�z$ɳ q� L��x��� B\�_��]~����WB{�l�Q�f���BC�F�Dx���8�A5���&ি=�e1(��3�xG���4��jJ��I%�$�:��(!���|\|�8踫�^��	|��]HU�Ϳ�:�����=���X��4,)���n�Ǟ}����r�E���#���t1w�\�A��ň����^�.��aME��pv�(u&,x���л�k��������A98��%�%�y.���%G�æn�ϛt�]��M͆�!�t��m�i���.=�o�����1���a�rj�E��dU�DD1-ږ��GËc��շ�CX:��ÍP�RX������	;�:c:��d��U�5�����Ƨ�,ù���y� ���� �����l$����TlBf���Cw=8�������?�.!���߱���o�Ĩ�d3�j)�����2��<���r�n���xw>��eߛ���w�A��Ӷ��؄�V�<,��8�	�1��� �!�'�#\<�Q�s���Ek
�Q��z#	mn3Y���W��B�d?m�������Ij_V�����~}؎1|u��
��i�L�C"X����ǩOkk	�����qc���q�#���m�w�GJ~b�c̨�j2M�^�UU���q��;�X]R�&���u���$�~��A�ʈ_z����i3fOZig��}���y����w�\'�6j����=	�̆��8��`�_]�배�e��TT#3P�͇��Вzz��ķBC	�Jo��.��,�#��+S��r��O��%#@Q�P��+O,z	(ǀϡ�Z+lZ�K��< E�f��Kȭ�l/�n��jH�PA5�I���z���|%էV��!4y��ţO��;~y�8K�^8��$�|��y�:�S��ix��w%Hhn��\Ps�uW� �7�{{���FMjQM|Q!�Ɏ:��qU�_7Q��p�#O��祈�:�Op٨��#sl<|%��N␿�H6��ؠ�Њ��'�`���ָ���r0%,��|��_���r-�-��k"�H�K5IJ��-�J�	����hy���gN����{�e�P�Ad.=x}��g���]>t��g-IZ55���3*��n�İ��D�J�q�7[M��
���"{�Mx�c���W�B���^r�^(�r��Hr�i��H�gZ�=��A�mr�-T��<��^����������w1h�A�n�es�h-�����;�۱�E��&nv��s����J�d�7_r<?q���Y($�<F�ۈ4&	T3M辏�*bܛ㖿��\�!������>�1b�i�Mș�`Ҝ�gܺɡ��W护�B��/<��|+���嚳�א������X��=�kH�8O��}H�V���S1��)�UD!�_�8�����J/�� zFs 	��ʐ�U��M�:�5 �kЄ��贽��������p0��W�jcТy���7\�:���{�"�L��Z2�B~�@��Y4��od�E����jA���>��'�eS A�K�å����g����փV���A����0�NG�΁��������Ĺ�O�']0Z��%��� G{>l�C�8��8�A�i�J<�Zk*�ƘS�p�e�ay�+D�p�0�#�X���,FC���JYU�傀y���戹Hݏ2��ޙ	��CB��p����3Um�[ٞ�0�M�WH&�a��-�0_���9?�/}������aC�!�ˀS�a���ˍ���i	\��(z�1�e}�u�XQET�4���ɱw�*�ʵ8�*#an�s�JLEI;&}P��w?�\���g_|/����ѻ!�Ev��J�r=ZK޸����H�~���hV��p�N�Wmn�Eӱ�ZP�a��KNa*��F򋪴�Us�*�����/�K^�[;�%F���g�{����{�2�����zf�%Z�i��'��{頻!V_�7v�f|z��/U�~ -f�4������m�Q�P��(�-(5�m��}�(,�� ե�����A�]��p�)$g)KR$i�D��9f���%���ݰߑ�6O�pۥG¶S�| �ITXm�����Дn���f�ԋn\���^N��ݸ�cQ�jG����3���ކBҨq���q�eG���г������G�4���Tj@���[I<q6/o踰Uw��/�g��g�֏��M��H���لa�y"�?���iD�gp����g��ξ���������a�51t��t�c䙥��bуI:YW���}D�ڏ�p�J���ԟך����1��K>��%D�/}�)��;ힾw^���<8}iR�:�0�'�Γp	K�:)���o��?�
'��3Z!,>�_<x`3��F.���P�yg�D���i�-�RĦ�g�N��[�%����y �����j��ʌ��v<�o�%$�m�2�C4��j��B�\h$�`��+	�	]�i�X�]��0 g0AHs�i;���Ov{���O��{mK�)�˧M$�uOՀ�fVZ=wT!�B!�}-�B��b	��!�TQtm��$$B��m��j�
��ShEME_t�ٕ��c����[G	D�l&�?�t5���M�G@��,��q������q��۩N:F�)A�G�L�#M��"9"45�C[��8��r9��l�1g��(���%���Ed�~=���&N����ڃ����eTM	q��T�0���l�\7��E��T�i�&�c�9�!
E5r�t���K�@B���+z��sc\��e�B�W��?œ/��-F��4hS�ߖi�����%>�̣*=�㜓~����~�l�#|����@b4�%D6	qr�R�ʠ��ު�m^	�f��I���'w���ȳoaӑ�`�����%����-j	,��"��.���ʳ�1���g³�N: y�C7H�Ӛ��/��:�)WM�p]/�1���{l��͏��Y���4�/°�����]g��X�H�����G����?����!�"��Ƃ�KO�9]/Q5DC�ޣ=׹�]oI�H�tW�r�ķ�R��Wf��`��L�t<Y��t�.#B��%��3.=���]���VM���8�y2��Eۄ%$6ai1��(�9n��0��� R��Q��7\��EL�/��Xȳz
E��X�`�y �؄Q���]�+nz��hCh���T���sSS=O��	.�OP�5�#=�E���&0ԉK�W�i�j��'[�ł�]�E�lg^�p���<��{��'@����Z˸O��ۢV��G!Z������fY���bRrɁ'/�O�u�S��3�-��9�'�bO�F���ne-9��}`N?�@Z_Rh$��,�5�P�u�@�su�8�F��\�ń+��p������QC�W=�^�hlq�pME�A�N�D�����m��r<��KF����	xZ*���(�}��_|��7?���&��F�i�j������K�f�Z�BIC�x���N�']x�,h_ �(r��&�ջ��vZ�,�&�uy�����Z�x�#L�2�>����b���Q��������r��<!��2�`��Gb�=/A�yl5rU��<ph� E�F��Ӧi�����"�${I���2�7>��u����@�q²�omDH��vt��i!��du<��=�?{�h38��j���"��v�\�(h�pH��^O�4�[Z˄I31i�4_mED�
�o�e�(����]�>@�C��O�%����=�?��Z�[�Mu�F[�|�<d)G��\����*�LXrr�Q6��Q,μ��'!m��@�RC����)m�?���l�֚�[�
�b�wg~8WMg.9�]'&��Z@X���dH"kX�1�������Iձ��I�V��Vn#�M"T�����J�Q�pm������n{���[�~�źВ��D-�������u���&ݳ�͖k�/��,�=]3q��[�Ou4�sҮ���	8��q��L�<��BwK����]�����K�C�(s������ҬH*D�%4��Pp#�ώx����~�,س��v�">C��?�h�X�TA�Y��7J��)���ItGx�x�/`�?VsCL�(��k��m4�D&�����_�ߜs/�oY8��V:6�"�J�>�(4�>]����"�/��,,!	y=i�W�N������Mzu.t)!B��%���G�7��F��B\�dDj�,��U3�4�fN �D�%4�)�&����94SG��y�������� s��� �0t��� I`�ñ�c���1эû��q�����7����!�Ͻ�Fn��C�9��[2�s��8����<8NVlq0s~ ��P�sxEi� �a;b��6V�,@iЊ$Q����a�}�T��!ޚ�6X�zVo��6�[	,CٌnVItXh.�t��#�b�I�����ڑ;��BYFs��r�-�P�j�S���X���k��?�ԙ��
%D&���Mv3��-��N���	/6�+�&_&������믄����,�Q���}��\��P�]m%�a��胥��*�6���9]�qm����� ����ǟ�X@��b���K4ۧ�hlXb4j�%1��i;1$����A�Q,i�f�����9��̗������s�ٙ��e�����<�9�9�2�D��凭j�'���_��oyih��;BFĻ�`�x��[���(��/�B����u�a�<�#PVq��W�H���c��P_���9 K�>���.E6-��S_@L�P������_D�h��=���0i�I�k.1�l9�q��ći��F��rC<��[�P;X{h?����ǆ�L�B�r&�)�X_�����Sѓ�{��w?��J� �x-� x���/��Q(0|h̘9j[n�نB6��`k�䡕̄s_�k��IBD��)��gaH�M�^�RP,o9�e�x�(���D���w����+�!�:�{�c~E��Y8�tξd'���%�
y�,�x���W
`��8J-��)̠�OCF¿sdD�����>8����{`u_3Ir~@�Q W��9÷��h2��0-��۱4�Zې�������߄���o�	����N���3���<n{h
z6�;s�6�ЧQ�������d�N��CWM$Q��w�
���T�`�=�&*��bg"ԄG�$2��s����0�c�t<;�#���]`��B����⣝b����EF�kr��I���X�PI�-yq�j�,k���?����Ǧᠽ�A(�<��E0,*F�G�!���� �cb�Qឿ��+�����ׇ°<��A��"J�2�8��u��'�C�zHh�ꆎ��1�e�w��,�}62|�Ȉ��.�{�/�<9��~6�D��K~�(X�$;`ZUȾ{ՐA�����r�T���k������ޖ�0�����Tʊ��I�W&�>_T�����i�F���aa��<����)�i���`Q0E�.�N�kL3Gl0F�Q@�ˑ.�b�u�*��A�BSޜY5N��?�5���G>_A�R���4E����Y-�#(��T�ѷ���>i,�'�>t]��Ę�?�S�"���x�WX{�`b�8�z��V(t�8v�D���I�L��w����F�L-ܙ�7x��O�!	ۡ�6�|oœL��y��j�|���}��V*��$;ml,���f����]6�Uz��Ȳ�]���X2{^�^�`�]�2��S.�LU(~Zs��[�P5�a ��a�-�"ؖ!Bҫ���Cq�e"smd���{��!�h� ����r}:g>j�����/��V�1Mx����S�T+�r��`a�8��M�]�	����t%���jI� pI)�65�Jz7֣������=��~���鋕Gs��t�.�PJ��#PO����	����#R��$Q�DF��H����_��Q�$�̜���|)2��|?�Ϫ�T�VbE�o��e��/je'��������*�(�FTh�ᢾ�A�V&����
xlkD���ۨ�m��Y���HXE���	o�4�.I_�]���`���v�KFl����ꬍu�p�*��+�8 4�8�R�W�����|΄\�4�<��!pꑻ��;_�y�뺼N�P �����$ᝣ�:?��苚�[�N��3�w���|έ��b�%��cgx�+�H�<�n̈x��wZ���Ô8���1)7�'W 2^B��7&O�� �^{�{��r�M�S2�r��J�^�d/y"�-���ѷW���0yN6��[�t�\i�z���6cN��&x��y�7�i�x�۴~�
�*�ߡ=�����/�X�Zۂ�L�q�NX{p��8���y"�����\SYM�*"Ѡ�T���x�`������E�Z߽����ӻةe��.BFĿ_�r��-��<�w��?.���9��YƗ��!}�r9��Y�-�:9[RC��Ců�su�-�l�����L���0�	�E
B�G�*�"[�2Ҁ)�Է�V�	��ͭh�'rt�PB�M<�,� ����"�����⭏�#C����*4"�Q� Jt��M-@�B���PC[[+�^Z;"K��V �|s�1o�7��wf>MՔc ����g_eD�0tp_9�D�
��
�l�"!�Xܐ[�-kF\CL�w�P;�}Ä���ۑ3x��8j���aˉ|pU�D���~��F�c��y��D�m��/ o�,�HX53���U�H"Ī.m��K�-%X���0s_�������}���.EFĿ,���W���[��ڻ��ݤ �HV&mƼ)�C�,G�^�@��]�v��
m49I>�:l�[Kxe�g5ۃջW=݋"""�/
2:�8������o�u<�琲�(����g\N1�jB��@�~��=Yb�:�,ڵۑ�vb9���/{��-A��z���I�;�i)1�п�������1x`�΀���w�n�c15^����kO��RiCN#"�x�mK�\���k��x>]!�*s����7�������ˇ56Â����^�}�� AQ�r�rE������{��i��{�޲�����ǯ��k��#6\�W�224�"���i��f?�aq�-�ɪ�g��uڏy�(P,`j����
�:=UX��R�/��!.�3?_Z�d|큽��*���t�J�
B�2�����E�BC���~�AD�I���iBO|�?�2�6�5���".<'�v@$##$
��kG�a֗m�~� ���Y���	�Ԙ��B�
6ڄG�������Tȳ�D8�*Z$�������k����9l�AfK�G��r����S��P��a�൷���$|��^8������Ss\�O�,��Ēj�1'�h��H�w��"��;�� 1��R�s��=D_�i[m�.DF�W(�Ǵ[�}r�'������t%1�<�8�i(r�a�d7�5rn^����Mp�)���3�&��j��7�d�B!O����SӖv
����Qk��0����5��7M~��d�t�K����N�����Ϝ�s=��f)��d�����"3�)�j��C��@���В�1;�#V&N����/����������a��}��Z��+T��~q  ��{F���� �)�;�(Q��7���$Z�o!�*5�Ȉ��/�%��7o�������r���m9�#^؆��X��P�AL�o۰�����J���)��鳍�4'���z�����x)���|̈́�Ʌ�4b�Tj�G�\�,W�EGۼ�y		8u�e�*��^�u2@���[��o�e��aP{���ˑ�V4E�&�v#�	�A��W�zd�����P�y�>����*U�K���/|pŇU��w�*�G�qby���9І��A��Yb��jCKJ��upyl^���:p��≯~1��fOFZ������[}�����M|y���	ԤW��jF�Uz�KE� (:}�NW,&d����b��W�M�B������#p��wה��C�h���C�bZ1�U�fpϐ���d����OWse��&����
����F:U���L��C�c&�(��xy�H�R_xg������
�ZAZQŶa�ZHm$!_��+*�dFܯ�
�����C�T�P���ȷ9�F-�W�5��k���}��"�D��fpr*��R&����������H������^�(�y�ʿ=��³�['ƒ!y�T�e�6f�ͧ�-��P2|{�hEW�CC��Ҧc d�%�k&�i��_��_3;��R��+�^�t����d�'�L :��gI�.�D�?O]X�Օ�"f�,�K2����O��rV�E-����_�!���f�A��e-
ܐ��X(��f�K����	�IޠW[��{C��W?���}fR߽wq��(N+J&0i{�>IF�U ��*��%�x]�-��Cϗ�B��3�����\Mdƹ<�ga��]~%%�r0�q3q�x�t�nWTQ2d��,C,�Z%^����1eyz'�5��1���k��"i�O�?_��>�˵;���J��Γ�>����ÏM�����O���������fj������w����E��^��""�e�(	37ۥ�C#15��s�5��/���jo��jFF�W?��|��N}r�]�޵�6�/a �����lZE�D�}�!,˂�+�<q������;m���[���~=mm%r���~�� IIT)��
�h�����%���o�ז��'�����PhmmG���V����g�G,t���$�7�}�*�a��@��p|������ �<�"(Ԡ�%� ����Vt�������p�>�c�mG������~����1�+�13t�r[Y���?AO� ���{DFĻ*�������e�ky~y=MU�L�̭�G|U 8�K;��� ���f�Pun�R����:�a�A�cޒfL�6=�-e�	g�ih(����,���>^�~[k�,��D\H�7�'(=�62���2�m� �+g� �dv��XV�q�f���*�JG�zzP��F��Ғ�A�\�i��\^���8��uQ����6�Z�7�\��9�!�x�̅��O,�ź����Q?��H�t[๪]h��UH\�vg�u�cГ�G�_t��>h���}����t���fuk�X�#݌�dI���S�0��kϙ�7В�/� @�X�!Okg�E=����!�!~=f_,�f}�s�d�.\�@	a'�اk���={�@D��|���ڱ:��]oAIbZdWV%t?
� :��AA�����P��p	�[{0,�������i����("4"�J"��u��k�`�l��@;��lDdW�:��"��v��d�|��È��I����D�%ɲt���=��S{�ٹԖ��߄ب��5�"������4�{�Y.=�a�%��6�	g�3��/h�r�,��H��%�H���������vx�?[N�Bfl�����ks��i_x�b7BFĻd����{a�=��/�4�ITg��"��e��ڑ��eY�'<h�
d=�>��T�0M1m�����o��a'_+��{"/ik�(�o'x��m�鈮ۚ��_Oמ�� �t�~p�05YR)���b���60A3h?�� ��}ږ9Z2�@GO{:�6�����!��+�WO�}�I��1�2d�̞�6�`}�A$ER�-:#�#�Ⳳ�li��5Pk��Oo���i%D�����.c�c�89,"�s����8���S��^�X�Д��#ސX��G���x��W�~���92�6dD��A �~}�-}o����;�~��*:D� V@���n8΁�T�Ԍ�BA��ا���4�(�H��;�T����=2LX�\JG�Pp��+�W^ 	�������f�X{ؚ�K!켆6"W�,�M�bY���G��ϿF��������6���7�B�C���XST��5�g�P,%	���	�TΖ�
*fdD�V0�˅�w� ���g}6U�h�`?KdS��1h��%\���#2���!ha]֯1�Fh/�,D�cE��\1���c�	5>jO��k �&�h䶊����r,��;�_|�c�m����~��{������5���F��%�&EL��1q9�9�H��"��<܊�2�lSQA�Ѐ��=	G�z]���[<)��O�W8B99N�!��#7_���4��XgH�*�M �#����a7u�'�EJ�XdXK��C3xo��k�Z�ZU�D�uZ#q��`gǭ���7g�����v�b����IµA�N%��_m�e=�Xd��X��a��Ri���<�����8:�������&̜����.E�zrX��
���!�:6�EN�Pm�m=/S�$�αG�28I�H�dD�K%(�;"�h�� ���翽������g�W�a�"#�����p֒���]����C�H8q�����RaV$����4�#u2���4��gݲ��{�/)w]��-�}�w�;G�rC�*Rw)8v= o��ىkH
�`E��:C�B-���V����S`�a`@3�u�x� +��\=a�cᒌX�
��`U�D�	)t,'h�o�ʆ�u�h��x��x�ߕ�7��˳߼o�*�R��X���:���<b��_c��v躃�w�j�<��3^#���9�\l��0|2w�����ts�&�Vm�V�y��7o!�b�Q��Cs�P�=	L���(4jE$\��m���w%t3A���h��f��Ͼ����ůї�!kn]�Ȉx����:���������+��:��I"��T�6�4Q�x���~�ò5��E,�Y�>}���w��kN�1��=�5*x��9�f�5� `��/W�������k�ǉG=}��!m��r=D���@Q�ȷ&����8��Gk) jq�`��V���p	�M
�)<q�+%D�P`h*F���)��M������E�3Έ���˯�@���a9ZK��;��u+*��z$m�Xw���r+V��b�P�~@�[�C�x����uCKL96�c�wߟӣn	�w]u�<t �:�_��c>��ٺ��u�����؏�ʉ�O���s_�L��I�Վ��w_,�y�/���5�>���~�W.�i�8z�I�2|;p��6�F^�ƕ/֣yY+]�C�,W���p̙7��]�Ͼ8[l�x�����+g��q>g`����Oѓ�Y�u����R��;D�"�8���G�S��"0e�{�I�R���[�0q�<d;"��3�"k�9��}X�.W�Dd}�M�䫞]n;|P/4֥*زM��1ْϕ�x%����������x�m3��B���N]1����4#��V�s��5v�j8�/`?�<�|J�%�\�O{��2��Ԅ�=ƿ�_��k����Kq%����&'�2z�����`��KP�(�3λ�A��)��Rd�Ȉx���K,�<5y��{�Öy�P��-)<�yy�RV�d'��.*������'�R�g�	�-v��U WTq��18��[z���9�k��V����;�<p۱�&�a�����G�3|�GѲ�W�irv��w�u��DO0a�d�-���Lq�62{�&6���2V/�ˠ�:4��^;m�O�y�G˶�� g�bmyi�T|&"��-A~j�;��dGW5��&N�N[�n�1LS�1:ub!`�:|�c�7>��=w�l����v(I��+!���I��C��'3�>���=G􎫉�'���l�"C��*�F-ȇ|=D�.Wo�Z��m�_�t�¥�c�*�g%�����hf�_���-Gna�Q�Q�M7�8�e�󩪙�f�w��3+�,��C�cS���<4ۃN���i�?�ν��w�@�h�,4&m�m.+?�t"�m���c�M��lpO���u�� K�dWBW)x r�Yq��-8���q><|���Θ�𯱸5 �!T
�3��`p<�}A�'*�,��v9���RO.��u�����AX�T�"�=�L��O��6��۲`��0w~��F��zG[�5��!�5�U#���D�`�MBː$�p�<��f�7�`*�`j�!WD=��Ҧ��Wp�eG�hZ�n�r�VȘ\� �|�	�@Q�I��++,Kj�(<"������[�.(So���H3�=� �������1��7���/';��7���m��;0�����)�ԤXWS�:���18��[ ��W2�|���pҡ��u���PG�a�)=�@��豎��쎱����>^����B!�HW&�2���2{�Q ��|EL����T�*��g�V�������Zg��a"!;Q�W\I�`���c��>4����l/��dD��b�B9� PI�x*�s��p��x�շ�ؿ����a֜yXg�"S�k��J:�,���N�(@]��9�=�>z�J���{I�����"�xRg6�R�%l������4S�`��?�>�&�{f��]	]S(TQ��V*⬓m�����U*e/p�<���=Jo�R�����!#�ՁV��&_w��N>b���$\���m�Zі���w%¸�B#=�P.�B��ލ&�9�H���;��������؃v�f:`AM.��R�Jœ��N�S�^;o=&"��%��]v�D�����prf��md��Pf�ӆ�1��g�������;^���� �S5�D�YqA�u$��jF~��Fn��z g�ƝF'��x0�\J��D(B�`@��U��"n}�e�Dr��?��o��9\�����f5VM��+M�`�2ˀ��k���x$�l/�o=j�Ӱ�j"ף���a���q�2<��&�y�#T3�Z毗�~����)*2t���(��q�p���M��&�����&L"sd��l�j7DFī_N|�I���l�C�5����4tE0s�xx��OYh��^AC}������5q텇㗿��j�Ί/i.�O�:p�M]Ι,4�d�)T�Q0�෿��x���t�f�v��}7E�<4ႍI�@��H�D�%�6�KQ#��l̚�j^�ka�y���
"
|������DBCDa��b/��������Rg�'�K�O:bE��u°�~D�v����t���C�{�+>ܰ��*3�
��oCB�3Q5�%�c e�*���G�(�}���f������
�ӏٍ��3ܱ���!�]Uc�+B�v9��'��El+�[�Ρ�5����@,��o�B�xx�"���nr�c�D�UZ[�xx����e���Ƨ��_"C�DFī\N��c��������E�b(z��ѥ0�:���Bє�����q�y��K�R2�෗ݏ��>����k��&Jn�����6y�!\
$�6[O�z�{��K�B%֤����@C MW��)L\:�#6;V��d6��?@�	3������$�:i�E�I�&�X����14�P����v����:z
8�ݖ?�����B(1O���K	B����(&Ê4��6>���?�f
�g"�U�\�w�oĬ�`:Px�vE�w��<�6z
����)�ښ��D>o�b�M(���kȫ6*�/ۡν�^�jk�\s�Aִ�R�b�!d9~���mp�(��S�t�"D����x�yiIz&&�M�����L<��7����#�&5����3"ޕ�rK5� �*,�z��P5`��F\q�h�����Ѕ&h)��6���.XJ}E�rm�h�,eg�����NT;�<�����x��OB� �Kk#"XI�87E���ϱ��ݏOˈEM#��w��F1��/-(�����D�s�J;t`�cp��oA�����C�S��Wd?x�ƒ���#�)ڶ
?��'&�xw2�2���[�w�]`r��Bm:+q���=�TyBID�!�BQ��/<�Ǹh�U����rژ���*+ȋ@3,�'���ת�\J�!QĲ�����z���a�^}�D8�>h�T��z2�ѕ`�+�G�����xE׋A�:sF���K�-oٜ���B���3|����g��t1����e�K�����l.��Hx	y� ����f/\y��8��:2�������y��--m�su�,]�)P�T��	E+Ӧ��W��9�����TՆJ�����F`�͇�ko�i����J�L��I,ئ�2���ޞ��;h��]����O����lG�d�5W���H�'҃Q�au��T�p����תv�W��N�fN��� "reBc"A�3�\�·��	�d��A��7��;o�"����͖_���&d?<�=p��66�p0�s<<�-��Z�̀ߜ�7��ҡ��A>�s�(1Ӂ���D����;ը�{���폡k�*���2�D��A��L����2-
(5/A���R�����W?��L-��##p��k�~���m8l���=��B�.����B>��!��AQ#�C
6=�ZfʑVk�a��F㬋�:w���_�U-��P	8p"�>g�˭�l��S�������{n�G�0X�r�5�����vCTYJ�`^�����9r�J"O�'Q�QU	���)d�����7p�>#�ly˶~�����B.2���#�L��)>���ϘM�U��h���6�=w=�`�xQ��%��J!"T�/�1��A�����Ӑ!�[��6���-RS�ӱf���A3Uh\}�8�Ga��s0wᲪ�#a{9p����F�a�
�mm���^�oE(C3�TP�-���G5��s�оCa$.���vU�k"42*ޕ�X��`��J�]��WK�<���\�΂6�yh7GFī\���W=����Ϩ�o/�QQ�}4݁�ñM
���Ҍ���Ⱥ���"mRwD�r
#g�bT���b O���>\s�h�qIu���
9��1�c��L�E��T��m�3}*D�Q�@��z��p���ዯ�`��˪�\(�]�Eg��SFR"�QC�D�C߅i�8���)f�eV<��q«�Ha��n�w2�;lw��/�C�u*��0�%T��x�'ρ���#v��seV�Z��'شѝ����r"݇c��<}&7��AX���"_�q�Ƶw=�,���	^/M}{�64�#���0��o�D�\MV���EB��4���p�Y����i������C������'h��-	Q��-**��_��6T�{�X�����~}�Q���R %D�-�[&�3����>��;�x,�j�v�&�R���������z�1�V�߯�^�CFī����_9�7W����?�-�p���>�	9z����M�.�ʁE~�G��������#p�%w#�"���`޼v�������i�#��O�ª��(�����q���g�U��-�!����з���%Kѫ�3	90�<�0�>j"J*rΫ����{&!C�����O0z�=Q��^�r\��)���1�+%�9���@�(�*n��w���Ū�3db?Qq�O${��/(�uQ����8&"N��֊���t�}�ղ���gȐae�x�d��fS�q�9r�m��"��
r�<|�lS��b��.�ϻ��+�=QU�&����9�81����£�ܫ��dx�{C��u��ª�0���X�R]:Z�׻���1��d��]�����"��)�ǭ������"��/�����O��Y�����U2"^�h&�5��g�}��CU�e`§����l0!BS��ebn]	�z0��B�r;4GA�&W��S�u�2���AD'~s��x��s�+�hm[
�鍐'�s���k�r��R[�\���q�uO�Otۃ��yz��8
��QVѫ�*A3�ź|�B&�e�&\�)�r��ݘe�2��s�8�s�q�� Ǡh;���Z<���JR�d?�K8uw^}�;�V��趇WL*����Ǡ>��u[Q_$�T��|���H������% r��:���!+���`{9��[p+����]Ψj�����u�9֋��e0�hA����ʣ��3o���nj.r����ܓAA�%�l��#oX���XF��ި�C�Q�<x8�;�ƿ(�C��MkBOJ�̞.��h2�,���9�=q�$j�/{����e�J�֌U���W?f=�������{�M�-"�
"WQ5a��TTd$�k�3Q����6�4K�Ё���W�q�PDq�}O�g�:9h\p�D=N���\.Mr\QC>�oO��r�x~�G�n�{?�_�u(��H�J�Id�Ȓaip��׀IQ���#'tma|��b,m�!ÿBB���3�b�6�BDm�FD�w�E�\ZGZ(�k��=�5�㦫��������c_��-6�_��#��2<"�R��c�B�|=*e�XTL��F~&�t�^�2Gfh2&��_�����a�����0̢Tgb�����!נ����&7t�5'��?݇/�w��+&��n�.ƌ��l���iB�5g-�أ�i�Udu�*J�t��q��S���*�%��Qpͅ���"��	I3t�@2Iƙ��:$<f�?�6���O���4��2T2"^����W\���C~�Z��ػY������Y��x�TCCM���	O��eh<�,�t�@�F�^z$N�ݝ��D�ܳ��������bКy��$��x��צiȒZ>ɷ��ǮC���G�5��p��S)��.х��������Y�k����r g�#1d6�4��)G�hzH��O���c��'ÿE��w��6d��'!bD��B?���v�����\>���7'��ǿ��_�����w���tw�^+���b�(�|��$'I�,�4U"����D.���۟C7��2�F0�>��p�e' ���T�Vد�uE_7��'�}��c�;͈p��G��{^�s�}�m����m�~4
�hC�s�5�|���5G��u#�	�@Q�P[a8u�=w1�?�>��^R�I��`,��x�=gA��g�2(����w���3���t��W.���ӗ�CV�^uȈx�@m��|��w?x����-ٰή/�>{�*C�AcQ/
DC!��AWmz� �*t�Y���<g\tJ���d�E����]��OǣO�zD~Z���8o�IAF�u�Gq/yj���!����j��8������X=+g��N>j/��p�£߄�/*=n� /&�d�XE���r&}=����(���n�@��+2�6pi��݅�ǎA��!��8�t�P�j�UI1������7���]u���`�0\��Vs�"�.�Ձ�n?D���<+A{�+�^�\�<�+WxN�!�1JLvo��mN��NTO�O��>�<�q����=�Z29ۧ ��"��#�"~��'G�<�Dt�;r6\ ��<a����/ב������ލ��6���R9D}!�
ٹE,\���⯤:�X�P� ����X�{�I�Mc/=�f�Hyx�ͣ�NC�����HA$c0��l���Z����'�s�]dW|�ۂU����4S@����xb�S�گN+k�b$1��Ⱥx�<)��E1dY�'��=獓���4u���	���oAs[��cU^1'��&�z����8�#���|��'�p]7`�,�n󛑣�_��}m�z����I���d���y��{�۶�q�����
��Ce%t��e�&�e���:!�@YD�ځ?��l��d�"���$����v�/�'��OC�M�{,Lť�\���y���P���%l�a_<0������+!O�M�=G����#���=P�#�a¶uy}Q!J"�r�JDd#����s�L+G2{����xn����8l���,B�?�rl��ijp�e��$���X[o67��<^�:�{�Xb�r�n㈃w";ue�^g_9w�(�5�5U������0���$T�/λ�*yy�U�q��A�Y�"�_am�P������WP��d�oq�ű�e9�+(U�_�:~���	��«�9`kmy��O�����w9�N���u���it)�؅�;B��!����[�����cY����c������f��;0^;��qx��12�%R<W�ҙ�~����H,E]C9萮_��"q��8���1��xe�G]�sX��ƃp�{����Ѓ��ð
��`(�J�'��Gl6B���B��:c������+�Y��� �����8�]`�gu�2T�HDP�E��*�����mBd���q9��j��ѻ��v���<��f�������m7[�<bg��5�HD Ŵ�*6�1��^3X""UJ�-���-?�~��������7s!�{���&"���+ۺ4]��L�5g=��.�򘈮���(��S����o���L�����ſ���8�g?���P�
���F"E=YTĶb4�Yއ���OZ�>�e�6'�}�}�p�h��c�Ň"�7�׆�� f}����cF@{��M��R$b��#Ά���뢵�uћo}4��I��Qe</<���Y`C|�o�O����������]n}��I�´T�%���y8Z���� R,)f�����\��*݉R�O$�;��[�p�q8����{��p���קp��P��r�����y2Pt�AD�.��Y��ђ�\"�:r;���q��I���l|��݊�����6����$�YD����׃o>�.�%U1d��=�ߝ�3c��#2L�6}&��ob63<��o}~��h�]��5�� 
Ц��U��-Q�A�5� �m�셈G��ç�8���%8���ԣM�r��d/s��F�.Q��n��8��8�kh#&r�Dd�,tA�_��L�\ݦ=��p����f�>N���^������kZ47<4E���[mBk�#��&��<��$��!�ъ�T!G�1)���L_"�������'a��s���6��Woa�M~�cF�Ava�\B˹ٚŇd�ZB1�"kc��K�U��o���P��Ki���=���[Y�z�~��K���j��������Hx�ç�%��S9T?BR�J_,^��5��� �e:2^�Ȉx��Q���W?�p�5��E��w�,S� ��1�&�.H�o�$C�!U��y㬨�S�a������m�bA�38�����j��8��}Pp4$~3*-y�������ƀ�pS����5�����m�~v�8�';a��f<��T̚��T���D��%�U41|H?�6jSl2b
|"8�eV�� ɴ(H�)�K�� ¥�.$Rns&��I�ERZl!��/V,���'w�K�8[�o�z�7`�������SZ�E<L�|��޲,=QJ���141��DvcV�.�p�O��	GY���<��t̜� �[��z}r.�o��aC��ߞ[a�֔�ݖn�\U�*̵E�	���(c �P�=�*4���b���D<��r$÷��+�x�k�[E\��:h�!�+0"�e��T�5���0�ǁ �*�Ug�ģv�Ϗ�3?[�'����>_�e��_�N\z޿������}w���%3�,������w�xr Q%O��ף�U��kA�`�-���i�'|���qw�Ǵ����C�M9\v��PY�&km\�ȩE9�/$���0�5;l��_=�O�>L_~	�zdD�g��ۦ�������1�m�e��RWm,���/�nG�Xd�BHNBa撡�`�����*䩦f
d.;�H\{�x��y���`i껟c��q��C�mX��DDzQ�n!��>|
���A������U��������.��cz��������p|�e�m�p�R���+����0lP��x���]�>�۰!�v9nL4���q&/9�ͽ�@���ɫ�PtG:55��[�WMLx�=���䌄gXe0����S�tY;�>|ԫKP*��^"׎T����:�2�Ui͆�L"!Z�re4��2<l4���;}���^�5w�|w�Ehi-�cŤ�t��N�Mcc�� l��0l8����(����]��~��G�i?8ك/�T,2��m|xH��V`�k���˒�p�}���Wgf�#V�玽�E��Q�{��ґ_Dxy�dx�MG
���JDv��/e=�2��>�ub���c�!�X��´my����E��9�l�<���DdwI������E�3�/��t8��%&�U����-�p��=@1���U"Nլ�<$	�L
r�����ߔ��	�����̞���F��+��x(~w��p�et}v6ug5#�i�[�l�s�B��Ϲ�����2��܊U����\,�jIi�w<����;��m�o$*3b�a�A���C��\f��F"���9νɲ؎��c�����������j��ͤ������kO��'@�Q��#�$[�D�X)��%�,��K�G��2!��Bd����@AК{lB�&���L=��Q6in�@+r��b��w@㹚��ǐ%���0����\ѐ+���K��u�[DL(L�}W]7�ޙ��2|W`����1i�'������.���u=�IF��m����3��0T#�C7T)�h)g%�KvH]��=d�z��$�LL8��">L�y�,pڍ�w�ko)�'/�ܹ�\#ZD�W����"�7�'X�$��g���;Z�~5��>��ѧ�C���d���\�&��?�y�<�_^�~��3bI|5̀e�R�C ��y��K�~T"�E9�R�x=����\l2<���A�yS���X�_4I�c�E�ׅ$�L��op�P������o�K޹��'��<��`�l��Qa{�\�X��s7�a�	�U���8`���}UxT)g�-dX}�-�g"�V*I���|��y�Z'ӗ��6������x��Oدi�=v�x�D���S�M�ձ,����t5
yrʾ67�����]�ɹs��A{m��MM���纽��n�#O�W_����HR3Lǐ=�,P��l�zY��sa�:�����@u�xDR�&"�}���I:��R1(�&ܓ�`�D�yff,�q
���6�H�RО���U���֔D@
�ͭe4���m�.{/rp�/ǢZ�����Jn���v�^|�?����Ϧ`"`�L�<�C��m+'gu'qZ&�\*N�5�2��}�&ۖ�J�IH;
E��UNڀ��,qgb�廚��c�(�ǜ*V��� �
���P��a ����6�^R��9��5���ⴱ2;����?���N�3n��h4�LZ�6���1���W�Z\1��/b��C����#�!�/l"��-d��⦂���?��p�J(�?��I'��#dr�E�\�.�o���.�LӸ��%� �%����=G�T:�����%�u�mU�_��9fOl��`���U塆p_>2�F�(���#/j_���������EV��c��V����S�2���Fj	�QYDD�^ڛ�u�t)X֗*�&
jYuܱly��D<o�0j�A���`�s��n�rU�>�#����-�ۘ�@�
J(���T���Y16ȹ+R��T^�������d8��o�2�HU\vM�l��5d���t���}��Ll9�=6�$�:�{IVx��F��'���h-���,4W|<�k\��2O�����Q�<�f�z���a�u���ՔPD�S�[����\����nK�&�a;�I���X �!� �$��؋8oå�Ҧb�#�4u�w�dѤ��Gf�� �t��4)8�{+W��&�>y�Gw׋���}��P��=�سn�E�����0S?A�g��9���ds�ةgR"�R��<���b������_G�p�EF9��}���{���F�=D��
C�d�����N��Hrq5:�r9I��q��U�:x⹩���Q`�}��~���u�IH�c��]�h2D!*Ȱ�@�t\.�[��o�q��Sn��f��w�x�a�"#�=l��/����rr�N�Z.r��A0ӱT��/O�eƊ��Q`���ڴ(`�p����C�1��Ʃ�����7b���'��)�ᒳ���|��]C#�L[g�ܠ�R\A��DB�;��<�`�~� &��8��S�PГĨ�,a,���S*N+I~��~#H�~C��y=k��#@�D8X�Zs
coyo~�EF'2|��������3p���1)��U�%�ɹ�\Ӟl����DK�Z�aݰ��(r�0��$�g$(CM̎�6	�3)�H��B�$;0Q(����9�q%N��)�W�D���ˤa"GC���.�^yf}ޒ�K����.���jD?�}�R�-
��C3UZ穆C�1f}��GB��q��&g�sKG��n%�/��}ĉ������B��qƛ�g�\$�.��'[
��&��)����
6�m�	.�������j ߎ.=u��"����gyK���n�)dX�H<����^����mȉ�z2"^�0��u�Mk\w��u��l�e6|b�w��f�:�V^v�\�F�Ĺ�M$1TN��݁I���&�]}�>�ƪ��~��ǉ�\��w�#�:g�/���2#ĺ��cR��P��3"LB��@�\�|8�s�9��A����T`��C����Y��"��^0�"���R\��ʽ����]��/���7���.n~p"��l�gX=���%8�?c�������4�Zm�P�$�|�%3ކ"{X�0�����3Ua �]�k;u"��b{I�nuYg���U�xLe��iH�ؤ�N���3�����A�� �"���x�ɸ��7�LeX�]z�_��ƘCFa����u�η�6.�$]�z����rn��>qA�m��:ҿ0�}��xZ5��q��Τ\��*���u���EvV&�m�%�\��R�-�`XL��롗���"���$�ƫ�D}����O�Oa�=��e����CVx���u��]��l	�Ȉx�`�6�%�������3�pS��IH$ч���%R��q��^;R,%÷G$k�ى�������;|�6��%�b���ۯ<G�yC��t�̣/~��^�?9p[�Ƕ�����'���p�2ې�6��2M�F$"����L"4&�)9��s&�,��(T:Uf,��~�,����&�� u�fy��2a��
bM�����SO��-Ȑau���ާ�c��w¾��p:b��i鴦�.X|*�S�����+F�$�[�?QK����X�q*J�9r�R��d=�ӲsE��^�azeDDD"��؈'&������Hf�R��>�տ=0	O�2����[�C��.�uE��D ��Ƀ��KLݠeK>V�#C;ES��Ȳ�N����:J�=J�t�3����r)� �J���Z�t�b�����������:����\؛�q�I(濠kl�1��Gⴟ�&�qF»Q��r(�Uz�A1��OMt�Pι�5�&�[� C�DF�k�͞��W/��蔆��x�~!JM����R �<2~�Y���Д`�,2VI��2t8�fa3��=غ�Ƽ�;Ǟ�ν���q����M�}��}��A?��R��P0L%&]c�ʵ��L� 1YZ���g>�mS:zaUI8r�:�I���=�<���V�EZ�D�5GE *еzL��&Lz��-B5Td�-,jvq�����g������� �C�Q�尿��A�$���P�,J�c�%%��;�6�H���4��ZDD��G���D�U��#�E�
x�ix��X��I���ҵ��������k�w���˨MP�ڑWڥ��m��i<�ۑ�[���_x�����y�/�М���l�t�V�yB����#F����u��������QMEV9��͗���Q���~8��C1g���+�ዅB���xlڳ�?w�m62q��������������i���(�mp���=�|ʫ�90�HjRԧ�g%���*���,� �BD�N`R�p�'����Ƅ)����H@���'�ၧ�aב�c�-�b�u~ �؀(�dƛqT)XEA �f��"p�@,�e�B��h-��LpY��19�e����
XN����4��ܥx�x��7��RE�Q�w���]E���3s�+��N��J�@��""RD����'���"Ho�;R!�Fh!	���!H��ʭs盹�A��P)a����۽���;���9烖6���4ܦǁ{���QC0r��z�srh#UfaɁc[�����=��T�"��y�l^S!�G����[���U;�弨T=LQ,�������w,�ęs�'��ٻ��]�D�����o��+�8p�-�Ϙ�1�_$�D�T�~K��1�M��T����}aK拺EU�I�2�2������쑖^�A�	����K0��E��Ԝ|a�����#p��{��ڶVM.�PлSI㊾���^�Q�$��IK�k�4���Wק�JI�ѐ�}��m��t�ċ�:x��>��N*�^�ע&�k���'��~^���u%\m��Շ2Փ���|�X����4B��L�b�xԞ9bm\z�Y�>�_�L��j>�<��M1|X#��fS4�b�h����<���ݾ=u=��IlR��ȃ4
��h���F��>ﾻ�>�
*��+���D�nT�[?v�sxp"��!�l���4a��7��Sc�D��Y����τ�#�<����U��kO�գ(�B����`<��,,\Ԇ�����;=-Dwb� Ο�����h(���-���&l3jc�&�<Z�D��Zn_�(�G�y~L-�j��\f����.�<�2�;�L�;�ӊq�g�H��(��"�)ڏ�m���V�N_؞�o��/&�ש��^���a#�#Lxmޒ��/���+��s`:�=�#����o��+|��U��Ⱙ��Z��v
����Z�� V/��k�^�W.#��<�.I�s��7m�"2;n��+���B�D2�My�%��g���}vXÆ4a`�2��K�׷�����}�)�#z4J47W�lY+�C����`q3^xe-i��7ѣ�:2���Ky��	h,a�-���5����o��W?;,��{;fG�=�JU?+-hn�`q�\,z���}Z�q����!z�Nn�%���;�ޓ���l�6jD��"�4�g����c_</Ο����`yK�J5ż�V����u��NB�{n���yg�����
�7_��D�z�`@t��eX��sZ����GϜ���.�o�
��cM�
�N����W���<�!���-�W���"�.����V�$΋3%a f�q*�BC�<���wj��0\��o��s�n���'���n���#O�w���#P�(��*R���������7�C��Gb�	��=�UL�U�p���Ms�)�뺰���+��h��$2SP�T{7��MZ~ST��v&
��&m�j}E�3�<�����z� ��{$�{/�o֢h�/~s���:�O��ij|����a�)�_�p��+�Z��Y��T*�{�R	2�q�hŰA��c��K������{w�����տ�� z3��P��,�����߈�u�4�ӿ���8�y�j�� �/������$�6�$ީȰ���DH_����h|r}�Z��"H���o}�ޱ������m;^7�(|=qK��:F��$2��e��e���<�jj���?�e�j��l����?;��3{j.@�6AA�=�l����j^�k���<�B����H�\�����i�2E������G&�9iμeS��� z$�	�)<������l?j���{�Jyl���8K�ӣ�T������I����q�v\<߻����˻B�7���c�q���L��D*8���#��q���AAD��o����VR��
B�ÁJڋ�9�!	M�6A"���I8��45[+(5�k+s`3�*��g�]<�·��
馐�)�e�'fV~����i�O��l�~_���n�G��4�y�g3����S���a6��i�X�0n�W�o�u�d,�[m�����.�����ww	������!�� �,N�,�z�����������[e�,��������P'E��G�ݰ�ʰ;<ā�ܺH7ڌ ����,�Sʁ�ft)Q�m���4Z���U��$�H�"��\�+�X��y�����;����=��^�*���r\��)ǯ��=ݼ�f�!�Չ�촸����q��R��L�Ϸ��-���Ŋ�POy�c��=Ӵ�k��v%�^�Wi��HY�"�0]j���~:p����#y�c��G�j����o�B�dyf.q-�ޙdC���o[ٝg�nf���ܤ��^B��&�L_���Bkv�C�?���@^��Յ��;�`�! �Fm��mtFji)�`� ���s'Qu�F��f��R��D���� ��a!�#�'�$����J�e�{�7�:8�}Q�t��L �Zu�����7v�F?�J���9�����g/���zE�HO�R�����ټ"m�8���,���!��Sq]��a�+�ۉ`��,l��GxJ����T
�ыן�A.�&��im�0��"ö��a��TV$2�!����2���n(���L�}O���oD�C���� 8�t�b�V�_'�ȸ��2B#��	 �)v��40� �Fw��BS�O��;8 �n\ʭ�O�+{g���
�$�ε�T�yƻ��;����@���?��Mn8\���.�|���ЛҀ�� �aj�R�|C�qwI�*��A����j!fN>�#�*b��^�S��߮�^�Ǒ�9nA\b��)_:�4fJ#�ԧ����6���]����OH�1|}�Q!�"�u3��+�����2��&��w���Ͱw�;ie~H�yݣ���a���狾�N�b���5m�O۪��x�NT3A�i��2�
sCҜ��DĲ�����9|��vz�E(c��O'`>�1C��B7<���l'�$�*ԧ�G{x�_��}$��c��������6�>�}]&)�=N�+˿}��zr7I Y���{L�y!�ɀ���L�٘��3�k��I���0�S�u�U_Q�����/~;;V��B��A��w�@Hl�#��㏌�ye)�^���j�WQf�F�n+��/�U��Ns9~]8��y�e���0���Iث�a{ʠ����~~^�䴻lA����o�@&g9R}�����*t��0����cP� S��5 �1���}��	$���69<#�2E}�`��+8���DX��[���3����8o|�g���0��7q
^M�"��T5����
��l�Xˀ�|O��S<�vBGY�bV�cL~� r�Hq=��q�O���D���6�0;ZZ�#��v��P�TE/�n� P�x]�������8of���|��{��%PiU����a�}K���,
Vǵ���Ԃ�chu�3���S�A��A+��ŭ��^�?���|��w��ȓ0ˡ�p��6q5��� DS��_����L�3B _����<���]r��"y_H�K��� �ߞ��ӟ����Y�N��n�v{
�����܅���4�����}i��p�̱�^�� �����4�@���](����0�f��k-$�A�aI(g��h��d��u�������J�6>O���Q2�~�u࿛o^0"�����F�gcj�E�i4?F���V!Z-�QG��oK��i�d�'(���ɞR�b@$�/��DcDLfD���w��L)�QOq�P`h0�J 	r&��JՓ���4�k��_�5�]=���+f�bn�`c_Ȱc�_cM����E�}�_�~��1�h�h����_-�B�ƛ�GC�u��JbT�H���	�
LwW�z���WX25��	e�&!�jX;YG6;��D
�,���Oӣ���5L�[sD)�|��{����%	�<`v&�B�o�vZI��b�'�$�G���uf�1�0q��"ʻX@t�a5�N<�v��?o�K�0�jnf�ɩGf�zc|��/�4�a�p��U�BeD���ʗ�)�s̨�7��b_��A8�7�(��2±2��/��9�����؃yq%�����f�v�^���Mv~����"|�AW���a��r\��D���B��K�Y[rE<w��\N�mxؾ]�;sHS��.�M�����E��)�=���DL݊�&砢�RY��6� @ 6��wy��H̗l?��vt8��}�=[On��<�"{�����s�u��v�JT��}ŗ霢��"��d��B_ Zu<���S!��2zB�|�o{;zj��5r�_�5�]�Ak�y��j, r�,�,GH�q�Im3�����T+*����"&a����7�-���P��r�8ʔ�C�����J��Y���A���0�軐�]o���p�=��wi��=���Fܙ8A�VëԻ�}����k�!����7���a�ݍ��c������88+�gٲa<<2u@��B������B�;)t��z��36ʬ\żJ��L�|D���MyO�%!����VwO�E�rTP�����o0�Ǵlz���xB'�K�]��ud�~�	̲��ڏ����͵�;���Wˢ����i�O�O��Z��Ē��j�O��h���O�i��q����˲p��*\���?@��j0b:H-.DqJ����������9��5!� 	��h|����a�W""�1�N�������3�KN��JP���?K��ox�w8��q�P���^��W#����F�rJ=� �"ƂɑW���@b�t��t?�-�\�]O����˦��V��	sg�@�x�+�ǧ� �%���S7L��4��8�:���f�v%(=0Q<����86��VtV4~(Y�OԘ	� ��?����ׄ���l�40�i/=P9k:���C��2�	]N�d%�\���i�_���yp�D#�y>�vcuV�G���qrT�1NI��,������詪BK�-{-1ZoB�H��]�ܶB��l�"w���
�!���|5�����a��w�$Ҁ���_�Zx��Q��A��f��Tx��u\P��v�s8&cB;�-�w	K������yh|���:w=��8����(kvUQz��{_�\L����]TŮ���-��&�܃qS�8��o]��vD)�1xo��˦54պ"�ȸ'pۃ�H[��'�/���%En�L��6-&� ���ϡ!h1yB�M���)�4B��͵�l1�y��j�eݶG�[P���I+�%��NK1A��	lP�M�&�O���n��"��Eڄb�8��vl�6�f�= �}:"��!\���Q)�f��y� <O=����H�O�����S��/^��y��d�e[Ql��K�^�;��^�Z����2��iΡ��0J^a�-�[,5�_��E>E���σK=��c4֕��k=�)�I���9���B����Q(����#�N��c����8bY�{t~�"U�i �՚�R�7��m>׊�*mmk˲��rW�՝�����K\EO{��,|��1=/CH�&���P2�A8�\(_�&����~��sݗ�#����<�5ܒ�V���T������ C;����&�=�j���ha�#	xj8����t��~[7�Dhj�/�1�����_!��ɋ���6[ӂ@;#>�(�c¹�1����� �z�����j��kŐ��n�Y7!����"����w����|s�Ӧ��u����šW����N4|~l+	�l�s��6#!�ì��'��o.zx4&l'[���\�c2+�!Z���V�3�j~
�7�%G�(��B�=��(Qf�n�Ɩ�rJ ׇT�֮`��l����=,&il��\�4�Rd�g������	� �Ʉ�H���@"�ͪ�f�^`d����~���C�;��5�#�������9�}/���t|�:���G�۞ľ�ܼ�uv�_Xfb��t)$�D�%������M���V~4!v��� �g`g��F�t��<�|�4�b�v2F��ᅬ �̗�D�E��t�j�UJ������8�����A�yp%�Sj��8��{`�m+
F�ش�xnIB���7� R����Ux"~"xޙg��L⎗�CQjV1BǏ��"f�Hh�5E��>/���u$��KWU%�)��v�|T��I�
Fx�2��`���c���6ylS�6v�XG�E� e{O�x{��Iߋ�
�щY&V9}�f�Ei0�VF������Ù�v����%��g�e���m���v}HEN�24c;<�M&5��0e���_��ⲱ��JU�斪��P�8���.}�6�<��W��~KUK�����l��JP)];�*�`�ػ^�Q�/:)ۺի����ʟ.�T��҉%[%�P�"Ew��p�}9�V�{���4D�. |�ɑr���M~x����)^h����!�J]�����-�'��c�V+P��$�8�٬������KN�p|��t]�g3f掄şR����v�
�A �}sY�����$�̞���I�[�������ď��tز�A�Q.���U�t�l���'d>p�y�!6g���<N0�6���Bv�\6:�q��ƽ}��%J��X��9�l�����fF��c��#Kݬ~O0�5�%��:���}~��:�s�}���[�^��Q��������������>�E�%���B�H�N�k��ͱ��]��=ӄ(�G���p(=�S�^j�,*��EJ�*��BM���o��_A�I��$�|���r~ǥApxr�g���ޱ`�I�o�V^�r~��)��ڭ��?>��Q�U�����ՠ�.������F#�v��&�n����>���S���C���M������}S���SQ�! Lk��k݅���2���Nh��o7��oH.�%�7������*�E�O�P�
�b�v=�t*�d8
D������Dƀ�i2��#��o�.y����qԀpV�)��"�sv͗�~U�9��J{��.��'�R`D��
Y
�L��f�9�/� �������e�Of��	?�.'<"��e���p�5`���W��ҵ�����c�ԃ"R�fx�|HE�h;u������	���EI�@��	уL߬�$�wԔ`��]�
Ʊ·�b��~7���Z'�R������{dI,F���e��� �7���~{X� ��@^$��حl2�0Qj���g%/�y�.�$��;�[�Dٯ�F��$2�x�K�U��^v�B7$J.?����O��ˬ$�.V�F�������	V\V����ӳ�1�n�*I�i4�b U��|[>޻�C�/w�������^`����vQ�
�	#�IJ�\Vw9�{���x���X|�\�4@A�j6�����Q���bR2�xn�#�R�WB�����T����������?�:���z�<�GO/��t\Ii#o0�RDչ�	
8ȫ�RQ�������x���g�X����k��-E�<����v�͎y�r�\��nؼ|�$9��'AS��|���>O��Oc�a�c���ѡ��X��u��I9�B��c�m���j�u���*��(=�\���e��*�uu 
X��d����܅\ɚXZW.-u]NL�Z��~,���˚a[ ��!�wQH����U	ͮ<\!�M1̺`��09̝u��d���m�fє\����������h"�9��[X�؞KuG�y�7�<�c`��5gO)%��m��@��瞉V���u�٦�t,�-}S����F�}���i�m�q^ѡ���wT�Ɲ�O�w�(�n�
�ƭTǉ��ETz�䖀�JIP&$qz�M:t(�R�+�.��vmV�:�����, Bţ������+[?E���l]h��T�y��R�P �d� �c�H��C��7�=�|��cy��RE��d�����Zq('��c�.m��P`�L��pYP�3�q�=�G���͓���?o1�[��tY�ٓqW�w�ERC��c�V�[��.R]�5/��|�_Va~b��t�	�.
���>J1��E�����["�
�������YXz�SZ}��8x؇9W��To}����O���Del�KB���flD��5L�/V(RX�ߎK�Gv�4p���Hg����~d����%-ZpܤT�B�j�V�^&�6r�L��O]�g` )";R�r`!"���=���O����7��ƪ�A�G���x�0Cb�������q�o��)�����r�1\�c�����mx>����qN*R*�m�[kt=,�D]f�o�t7�b:���_���:O1}�^�V�'��8�r�v�;�b�����t&��E�JO�B��ۇ'6Ĳ����%G^ݬy�g���,��p�K�(�m��p�~�ӗ��e��i�h��Y�6b)�1�?��Mk�[K�2C���Lb����b!��+��QmUE�F� �
�׿F>{�G���?���bl�p��u�?r��B�&��hKv����o���i�ƃ���5l}�E�!��p�����18����age���?�Z�H��W��2+�4i������8��ln�������<�}�ř���j������a��J.��i��8���CWOW���3[j���Bin���%��W�l�GQ��Иz\�����B��;�� U�@�����V��fKʤ��i������ʵJrU+�x���\�֋=0�i��?���;����@C�
J%�Y+a��Y� �M!ҢL1�o�� `�wuk������g������Me!V-z�S�N�&Y Y�V������#�d�Ȍ���z3�4�Ø*�(�s����y<b1+�Z@K R���m���x|��RR&Kv���i��m��a�!Kp�I�}���d���j�N~�ˮǯ`�M>�i��	%�RU4*1BO��cD<B�v����J��dkǐ�± ř�rd0��'���˻��ߌ��LJ��h�?U_��,HC1�>��V��%�U�v�q��k�@ڵV��qt5�~�w>Т� �����)���֨d���a����^o�8�g�+��n�Cb����a���+��w@����f'�"����� ��Vӝ�{Y39��ں�`5�
���z]i~�`ye5T�t#w�W�؁l�L�[��3'��>x��Y%,A�"�l�!��"�K� ����AoȉP�j����v6"Y�X��)��B�P�	jg����{��B�t��+��^������-�4^4�;�w���c�c�_�)�6B'ڝ-�
��{�<ҏ,���N+���m�b�y�������E�I���c�ὐ�������-�r5���L��q��~��ݶ�؉*:�d���N}������U-u�)�Ä�P>�c�^�l��`.�)y(ߜ���#�1�rR��ظ��D� ��l�����_q��'��i�x�?=�x�ҡ=��BdQ�I�NZ�9qi����?�K�y~�X���{d��G�5asL��K��Bi ]�[5�U7Gouh��Rz1��[�Զ��چK�];��ª��{�!�5���#8ÓI�I�yf�T�v_Ȉ�U����O6.H��E�*qw*� ���5@
fy�ב��*�>����h�����E&��s].m����� l����sϑ[w{�%��GZ(�0���x�f��8SXZA?�׮�ҹ�IY���2����"���itP�-��1E�aJ�ER��L-Ac�i
��lT�t�M���1��3�9��T�ة��&��輧B�wbV�T�>�y�(��Ӭ����aJO.Ŗ��� [��wi�Z
ͮPD�����CI1�F�JY������!�]�p��!�%�V1-�Fo���?�I�E�zc$�����\�#��	nq�^s�j�G�Ң���:�v����+���}����'�9��k�h��C���Q�݇���^�G_;��;5������=�ޡ����:V�D"�z��W���1�0l�+�5��5����<?�i`��'�kM���;��\�⅑�s�>�~-��2sdJi�wF����n�sW���ЊN�l������Rx�2�n�1�$���k����tD���r�+#�9}��4�=ο1��Y��nk�]Vr�����2H�ڤ��$r��-�"�[�b_X���[���V'Z���t���uϣ�m���n㲫�h�����2̤k9��m����H��V��_B�gGK��~�Ġb�����M�$f$��Yl$U�����D�$����cU��k�x���?�@�_v�Tl/��-S�{5C7:^R�nF񾄡��
\�:j'%Ҕ��F��M�����K07�c5pK��d�G���<��d[uI�#�i��0q��>��{_ܩWd��"�T�l߷���(�OM��]@�x�]SӚ|�o]�b%�w��d��긪�X��:�l&�?�{W�E��^��'7�4�	�!�|:+�z.*��o誶�o����,.�H� 6����<=�F�̚:�ܬ�cy(��bg�bs�g���a�(h�A������zb�&t��ē.>�\{s�C{���d=�s�b"�3Yc�jׄ�"�~-rS���OW7e�o=�;Se!�;[ꇗ�-� ύh��WE��<<��q}H�t�&ӇU��*<yG��ny�-�8Apf*���)_���M�V�̷)������c	�:��v�[z�&���g{E��RS2],����2�N�6�	G$��8�R��/��Wxo�}�f�j��
��J�"�`����h��ѵ�i7��%�;���G�3�Yt��Ys3������}z5���+�ܙ�wa�>%�� }��
�Q+i�����𴭕����rk=S��m�q�+�i��Φw��A���Z��W{�ڡ#J�?�9��Z�I� M���@�nY�������+���n��l'"�!�C,e�nT�{��eP��}�W_���B!��3Ee�~4�4���Ჷ�lO���7�f�}p���I�
�V�׷���.c��,�0�}�{"�u���vf!�"uu� �,zU�]1Mh��`a����27K0�B�G�`vc/1��b�_e��3�b�]u���4������ҧ%��T�s_��	�(f:TƎ5JHaZY��������f�jZ�ۛ:��7Z�i�Dh&����e}��VŮ�\+,���0��.�k�����^2^��<��1��vt��O˅p`����;�������:T����+=q:�8��m��Rkl����p[fJ��Ǉ^ޏ>��������0�Y���	F]��e[:�m2#��"�Ń��n��x��A��?���2@�k����r{�O�-���"D�XOr�=���⊿<gr��~I�k�&�T�H xoN��0Jv�x��H�~V.&o�pCzP�M(�_����%�w�`�����r��ȤbA�\����6\���k���Z��A�&��Y�������]�Lx���}�����
��[oQ�D�]����ԉ�E�|��Y���Q�̋A� ��0s��6�� I�~��p�Zd��i42mR����ui�c1~�bր�nl80��:��#z�U�~�k�ajy`�7^[�l��~9�͡��G��x/�资|��[��w[vc@;.(WO�f������Z���A�p��i�R����JC�N),Q�|!�����]���M��r��@��f��f{,_�g!��{K��ϗ�z�.G�������kƌ��Z��`��ES/��L������r� �K#�X:D#J9�+��B6�&.���Jy��ʧ�c���M��l@�it�	��<�~�~SB+
L�Я#�+ ����#�,g�X�k��M zh����}D"}T-����'�)��,�o��g]߉�O7	G��a
5�+�0��7ᐁ	�������:6��ǰR3�j�eɌchG.�	KԐ��5-��n�P9H�::niBY%��ps�e��`䳚�kۭ�$����o�F|	�x�R5�pˏ=��M� �Vf�N>���{G[i�4z��r�#_X���[��G�.٨���0����b��y��q�~Hlj���Y�yo��~V10�� �/N�49x�ޗ�L�^���=�,�M����c��D��YmR������z@��cQ����&�U:d��֣�H˳�����ǋJ�:�#hu����OL�&CmF����������{@��l����uE�f�v�Ԧ xt(y��@N�Ji�rj�-��`Z��fſC�|���nyg��ı�$V�}N��s��F�d�(�٥�tX�R��'f+�ʳn������T24i�%����P��o�[ɋ�0ML,����<����)t���QFvy����UCR�+�N]ƥ�.���)Q"�U���"�M2�P���/id��z��b00~~��xJm��`�#A���uy9��|��y>޷g�����.�� ul�JJ}�.�J��
�0"���;���a�:���>h���U	ᓺ��*����H�Y��c�	�{���܁���?3.�FG{>�y� }��;��;����z�d3
q���Řė���Ãy/.�v�M9�
A�I�������EE�\MI3�)H������'ɡ�E���O�/;�%�ϷA����YQ��i�G8���B� .�q3SU�G����F� �KХ���o��<�ZL�:��K�Q���~O8�oC���PI��ǉw:�����ɒ7zIf|LX��y)��G�#E�H����b�)��_�f� ��
V0�H�Q�WUt=_����f �@�ۮS�l�߱�����4�h�L�~]�[m-�P��yߘ�)�������Y��-v�A�*�&�(���6O��fh�ΐe�`nA'�/.��	݆����Z�텉�ב<bݤ(�mN�x��V�'(�'�� M~
�/����샺�q����m(� >\����l��J�To����n�wt�0"A��j��q�~DE?-AU��<��:�i��@Ԇ�l}�l����o�D�w��D�mu��UrXh�&��$���V�yP��\����R����5�~��~q+<���)�g/Ͽ�	67��s�L�mT�m�4�_V`1\8�7;O���RI�˶�"����qiR#����2,�a��g�ꏛ ܝ���÷�Ǭ��D"�6<�q�K�wD�>�}�i>������*����A2^���F�{iҰ���] Ó�����m�窈��j
!h�344�u�2KڏN�bz�L�F��o���lry@(@X@����t�i__L�?餒���Z�,J���z0�P���M(�����p�w�KiT����֤����$��X��s;ݐ���_oZ��k�j6�uwCk�))�!��x�cв=r���V���X"����ݓ?�V��&l�m�_�a�K��(#Wd�V�.;�S��[�q@"��~U_[V������ݰ͒&t�^��	�/�-s �h��L8���Ǒ�����e�em��X����2�؁h�������f���L�͐2V4hm�n������V"3Jl��y����Sʆ:�r��G��'Fg9�#�+\�S�+�����w�C]��H|FQ����jz9&�~�`N�.�������/���Nư������k�NU�c��1�p5�v��)����烳��i$b#�����L�츦����`��t����L�c��u>�:���%*���yy�]��X�^�O����ȢU�a�Қj[���o[C����q�׬�+��%�=dZ���I�?C�4�/e�4����n8,y��O�stf���)�c�wUlb����r9 �x�`n�m��'��۶���T6�D�)�CMz:(������!8Z���"��ʒ�)�7� kfg�,(�r����~�Mn�K���~��ʖp��ݥy�>�
����qP���Kt���=�.K�ȩ^���|~�ٶzܝ��l~l !���?�/�%m,���6��Z!�_��iU�n��F{��V��TN,�M]��F��9�F�CˤG_5������>wO��^&��e~��=�C�]2iMC�S	Q�f��ޭ>�jAS=�(�f.VQ�0�E�_Z,-V� !A��x6h�`�(d���*s6?���qM��4�/�SM����o���?����vx{��O�ɛ=�|~ه�m�O&��@lg Ǫ�?�j]�L����+�K«��򑜺�kw�p����l���P���fq�w'������}^/c}��E�F���w�ނ�CQ���]B�-+��������
L����t�.c?�d,�˽�LpunF�BuxH�q{�*'���6�4��tZ�i��in�.ܺ�sJ4�#���C;MF�SYHxm�{^�N2���E�l[k{T��	r#"��3���L��!I��|����k���[!�$3�;���!=V�!1p\0��
E�%�<났lAo2�"���H*�zg�_tU��~V&�-l�-{Î�M�:s�R%�ѡ�R��Z�b%�0KA�T����C�ȳ�3P�ޞ���%7-2��F�>����}W �I:t�����ߵ!�k��E���?�a�=�@P�&�e�c��eڐ�Y�)����PSsz���!#-uR�i� <�;�"FFn��膏�e�#��ҏ:
j�ϔr>�� [ ���囐��o�#�.N?�Ӽk��*���CW�p�t��[=��SB����VM���e-�G���Pf]��C�PYͰ]M%v�L:�~Q
,G;��˄���|�ވ�쑭(a���$�=��Kf:�n��eyYs��B%�^���w��0�i4�����^����^,V��γ\��
g�<��T�il��.�V;Y#9m!��$W�t�So�A e��G��J��c�*�Z��M��]�����uQ�?����Ӽ;biS+�,�/J��Ɛ��$Ԥ�e��U�!#���kJ!
�+"�?ЬP���n�'|b��@�(niχ���YuCy\\��;pU�$U�5XV�u#N��^\ L����N
��� g���jꡨ�.��a _�ȿ*��6���|YF{�5�KTۙd@w�v�Ź�>��*=�˻`� }Q1f��L���}��Uuo��҅t���sQ+� �_��M��ձ4�q���6�t3ޗ���n�6g;C|g;50��A !Zn�*��o�Iٵ�J���cm��Gڹɜs�!�l$4���0S���ꥰs���g��V�2� I[� �;z6]��T9��
�A6 ��Z�k��+u���i��1��܅3�w����,ZMjlW^��wc"�b�'-N����%��$��,ʆ<w�#hpf�9 D�O�x���\����_�ّfVl5sqxpW�縟�����?H��'&2fn��(s�4�FU7��7���:��?�/u)��nO��7f�;�L�����0t�� v����ô<ol����}��˔W�JkI�\��l��~�)o���_VA�y�Y�+�E)F��%B��ᅼq�:��,�-�4�� ���b�5u?�p���-ьgZD�+����A�K.��;%�-e�?���9W��P4���6y\�� �L~D
' �)M"9X��Έ� ���,��v��i���N>@�h�j�e�>3>�����|�[ӥXND��������檞����*���l��rj��:�UI����&�6��s֟@̙N���|�7��N�.Ⱦ�(��rfɪ����(}ȶ8�WA�)���}�<�?W��Y��g����lY��8�J��#�m�d"�_��U?n�����b�m�VO6�b�ଇ)��K2��~�7.�=T	�N��S�˥��*�\ND������n���/��;@��|�=��p�,��)R�G�|l閨���;�hČE�t��M��ǩE5eH�����Lْ�=��VK������XX��;e�=�j�:��SQ�<x}�1��Ļ�4��K[ �s�z~azӶQ��A#�i�$Ek�������W)��<�)q`�.ߤLta�l5l��W<oF�,/��$q	N/5�;$�ש�����eܬ������{�e���x�KN���̤=Պ�j~}ע�m�����s+�����Y�+T��[	���*r�2��B�
ҏ�q��`���v<�"H�R��DO�]'���G�B�Ⓑ|�)�Cb?��v�i��8�ݱͼ8�|�����\6�4<��lUR�q����$
����ڄf"LU����I�H�ܥ�	���;~`\ɓ�[�c<�v�:�ɜ�ov���1��$k�yE�ny��n�F�w���yŢm�u�xr�d���	����;�)_�.l��M����*�aR�}8���?.1�P%�V���b� �wH��)��=�d�e�@dEy/E��/���%�~T�b���H��ÅQ\�8��
_�?�X%\$�p&Xc�gD�0[ʫ'9U���L��!?>��A��ĕm����y�i�C�x��oA9��R��Ӣ)�E�U�/�G����,�O��A�p��^�����Tk;*VLh���3��	�U���[��Ղ)-��芏�3d�%��lsˊ+H��K�s��,�[���G�+�.�\ì.2��lx�-��k����u _����<�r3���r�����ܤ��W9���څ�,�L�B۠X��{�����3p׌JL5��DdU�D3�ǐ�)�q���83�Kt�ɫ _�Tyz��)����9ò�RR�<ڤ���tj�j�|�»�r���+�[M�/BD�'���Vj����8u�7>ϼ�6R.[�͑U�bI��H�'o���L�M�
Tk�F���	��(rH�L	࣎߳:�3��u���z��2L[t�0l,��k�(h���ͭ��?�σp��P���%V�|$1s��ܒ���-T�눟��8��V��6��&��'^�C�LI�>-�(�f����-����W=�#�A�{'���ͪ�G�_g�raꙈtd~g�:�m�n�dP������R
#�|����ڗ=ԗ�K�m8+�{��x���ɿ��1����9���>��"���c#z8X��A|:0�^J�7���/=���#�H���I�ˊ����O�P�P�\���##,��lT�W2�*%�a��؂��>j�'�^۷������*�!x��X��Е:�|�·6ㇷ6A����~!o32�][nc�W���3����%�~�W��jl�e�Nf�Z�X:gp��6|zW���A��y�{�)��}-�؈��&��m�vMT ����8xa\j�c���3�j�hk�+�E$�#_���H9���^
h��I�n�_�k`��̓�~�Ǖ�ٺ���g!�P�'OT�iVD���g(�"�1��t��c/�ѳ��-�X���Rg��'(ޖ�^:A���ڜfu���О������/��d���<���b�p�7�U�{���q>�moF�~W�mS�����h��K�!fs�:]��SW��/FǨ�f7M���a��k�t�����0�����yr>����}yW� 3���3��΢ӑ/_����Jv�$;�Z��kd��9�ٯ�ɣ�������
3/��)���ІQRR��r�sٌ��T�k���Y����,�U��%ž㤑��	���E&}���=���V�%�U'l`��R3"�2�+������c��1v��;Jī�ho�a�����4(V�*sP�۷}K��yhmw�f|��A�[������G����=7�$r+��~��Q����Y����(�W$�Q��bńg�]��%.{�f��ӷ�_fA�0��:ۘš�=��^�˩3�t	�eYs��Z�PM�
���Z;�]^y����T/�q���7�������u�\�hȫ$�@�h���������˅weX���	G���/���s9���e�u�n����P���J'���Hk0���𴳻d���O��я��O������Ā�d+�C�s�ե���t�J(9�un�~���/�q�V�P�{���~�*�C0��jUU�z�u�b0'�e�lyxA�Q�	��5d6M�~c�u{��E��e����NC!'o~X�ǳz�Ze}w�U?;��֏�xE Ї�?�J2h���g����g_y�Kٲ1�.���io�!9ٺ�����=�1VJ�W3�2^�ߒ%��/T���= �M(Q ��'��`��^�_�+�=Ae=�g�i� ��ChUhQb���a}!e��Ka���L����e><���������(\*�F|�ͤ{S��@��̫ �ͳ4�~�L��Zo	x���m�� �g��N^��ADQƹw�d7v0q�n���4���Ϥ�re�8��_�����E���Eѡd�`GU����iG�h<]��
�_�[OZ�@1ݞS(��B�tKwA��ə�ԑ��A�3��u��DR\�,�m���j6���{s�v��23�l�(�if�uD�4����f�_����v���i����g&� ��u��z�C�>�u�y�_)W����DD@	AB�C	�F��Ke��t�#�i�Q�f H���{��l������v]۳��}�s���5Ǳ-�'Z�-p��������"������\3��wy�o����ṙ�lM���#��q�6�1Z��	�ǔQ��ɝN�P�J3��ȸm�d-3A���J:���)f5;km}���l�K �'���?�Q0�싞i7�	o�
������弽�m;r9>�;B]��<��t-��*����W�ˬ��	i-������k8"�^�h����t�0c�/�3�Rd���\
��x���J%���텺]�f�ńh���p�T1p��G������u�IN§\��*�7cu��q�jq\i̒�eQp�1��M����xJs(�	�tpt2۽�XH/�3&:����c�x���i�v�l�^�A���W<%3�r�ۧ�ՖL�vJS^Q�T�LO#�N�G�W��W���)HF���_	S���=�kp��8��^��r�.���ch��WPI�켓�C��x�{��:/�MH�斄j�э�,z.�^įA�6�F�f����B-)"a��s�I��F/}��(�|��(�-��u��q?Y�Q�Đe���AB��]O��C�5Z/UpiO
���eૼ]"�Z��S\��Ќ�u�==���n#~������lY�)��S��l���������"7?^���K�^4����,�L:J�o����av��
��  ���!���'	�Y��`�5�5����b�/�i�+�"�A_�w�+����>����~K�&����?~��u�k��nwo��!}��9 �9.�4y\��8��sV{jR�j�hr����7'�{?\Г	 �z6�9��z��(�_�2vi#�"��Ƣ����w�>��Op��?۰v�6�󵚊���G¨�x�煙�2d�ڗ��C�xm��.�����Ȉ��������ɭf�78ʈ&X� ��9�)�yI��	�+i����I��Vu�Ɏ�I��K�SG}�CaO)v�/_cOtxU;	ڈ?み�Ty-V���^Y����qE��'�ٿ&%�c�|����wIJ��%��ޅ�]�&M	�0�zū䅡�d~����s�5ǻP�%�sa.�'@��7����bI=� ��GP���ˇ�PN�s}M��IXk�9������&#^0���g�D�Mn�t�/����LbF��lw����0���I�I*F������Z�g��v�>�=�l\[�ȡ���%��7�t,�/\��pG��� �\�<�zhjd*�/��bԘ2�!���g9�'���*���.@1�7��ugdk�B���O��QY���:�y�>��?���
��y�������s�v;k��"v7��������\j{��8�{}b<�\6�"k��XK܊����a�gk�Du�<�Ŕ]�$ �:��_�	{�L�1mm�L��'Ɔ7����0+��R��R?�)v���ײ�X�a_`�7\._r=���V����'��� �@���s�|�!!
��. y��SN��nchF�he0�-���WjrΡ�R�_�[i	
�Zp	6��t܂;���_�ӻ��s��
���9|lW�H=A��T�-��<$���}�:�2���R�d�O&^꼸;�l�=�F)���zH�e��'�"���M�N�\7�V��9&+E�tf�@7��L=������/��\���.�F�HC���7I+�r<��P���dLRY����|;!�,�y��<aw!FMkL��<����𢎢/��~��$��]O�Z$Bv�y1�mi�l�i�([l�5���X ���&M����{����-ӠqK��߶)�4���������	��N�>T��Q�F$�R��qm&�	v���_M�V;8��z]Vf��x�c�B�X�'�B�~o�؛W̟�������Z^���
Xپ��Z~`�!�SPw,U�}�F��|g}/���``�'i�Q� �
u���aI�,��v&z/x��j ����Bj�chJ��ha;S����9��U�gz2�q�bD刃�l��0yy ��M�<ڈS��~���}�Z��-��.�8����+�Y��9��]W�p����0��c�As~����_!��.��*fZO8��ӟ|���~;S^��W�)�ez�Fj	���r�&�����;��M0pvJ6�l��4�Gk�����8xo���vL\M��HV���V�+]�C���3]�â^Z�+x��il���T��4�?�}� �(4?��nZ~�l���ut�e^��_R4��T�oR�8N����쮱2)H�DR����p 䇖���o��@�$������J��2Q'����Qy�>���g�0M�� �s89�a�+_��|�)V���Q1 �#`,+�Z��*R���g�U�`rn��Y�̮֠�&`���b�V�Ɇ��ɴ>�D��YӾ�R���zc45WBS"��S�2O ?�B�T�
�9ة�ˌ�u���\�Og����or6Z�Vo�0Z�f6O
.���c�?�&|���\�py,�3~u�s�51ߠu�9��mEO9�8�N��V�������5¶;5u\��V��ҋJg�^K8� u�^Ó8��>6ݤ^o�h��'�'<2>?��<�lZ_��/kǍn�;_�x��y]}왎�Oi�v��<]�2K��jb����#�O!τ�5��z9�Ѽ����T�c"�_��X�{���A �"�36�1��-Vaٷ|�Fh������;5�}��?��5����ad+;�r�n�W����e����a�	�#�n��O�원!z���hL�J{��& �y�Q��7x�P_XV�}M��"��{�+ڿ�A0g�O1����p��5㩘~��s�2�hBr�ə�[m�7+°�(:%�g! �Bk�dV�z7<�:�l�ڟ��Y�^1�m��Ŝq��)b�z�9B�W	?\lkd	e/'����N!�f�?\�>�M�A�&���G�WE���
ו��b7��#w�h~�25!�t8G�H_��a�u��`��I���e Q���ٚ��ӧ���ءփ�	� �F��w�e�m��EYd�/��N���=Ax���3����_2܂��hӸ&�;�UUY���s�A����C,�ѹc.�����ş�d��k�zRj&ڜ���'.��'�y"���0;��?/w� ���"�֌r�a?k�zi�{!����?���򧌜7�y��r�ot@4x��4�1�9�6��1�љ�n���'g<��Ȏq5��#�Z����JW���!��[ʨ��V7�q?��vMC��ܠ��M�����3��r����qj1O4�B�3UrPT�#�7��Uj��:�����l4y�uW�H�W���E���塸�A��񥨏N.���wfw�B]���1)�����.,g�Xо��Ry<�A������Ga~яnZ�k]H/�9Rw�51�R-8E�#3ţNN�SY�:�+���$���}����K-<LJ�FS�����3�21�F����3���[�o,����=2�q%�mقE6=xj�3���`QD�w	��0v�<U��m�~�[��6�e{m�����Lur�H�7<u'�爠�|P��)����=A-��_�ډ��!6EO8�Q�I�%s�	u���d����z���=�����9��s'��j'��<1OX�/��+�5����F�V"�x7����l�h�/��*d\C뿼��Q���0wE<>/V3	$��e�X��������Y�ۦ1�"��I
�S+~����C�E���=��}���ov��,'�FYI�ƃ7/@�W ��F�0u
�ܵ���bA5\U���@��7`EoO'���3Ž�S&,%�m����A��?bqt�� �J,%dE8$?���"�)
�/���CyP�k�5���c�}���ѮtH������a�`�4c�d�4�e���-���n�Ή�W�j�@�-��U�]���ci���w�T[1k�!Z��.�q��9��(�W��Z�W�߿��'�z�����?��w�Y$)��61k�MAs~��ч�=�t#�ĥ[K|% ����1����=��cg����d�L]AǙa�`+jȽA�Hb��Na�P�!�Hg�ڟ������u�Yx~��2WNՎ���� ���f�0M��<�hxMb ~>*��]U���{_N|.`4|��s�o;�&�k�VH]o����H��ۡ���#ePF`��3/�ƀ]Q�O�/��ăv�N���òr��f���h���Lv��@֣ܯ��i%�M�uٍo@�i�&d���l�;\�5��Υ\�=���҈�;^�[?�g�z6 �����&�S��9����}�%b�����S��n�U��ņ$�����QcӲq�U�;r��ɹc�ȓ'ߗ�)���1%��I��T��JO&<o�<+<Av�Jv�5�����-��ƚ3_�� �C�1?���i�uc>�ׁ���f ��DZ�	>5�,��h�Ɂ�(j<@��}|M���*o��։N@K�UWbS���T��sX2W�K�M�cPU��l��`�q��;�Z���S��䭁�t�S��x/͠��p�<�ou�?G<�=��;����g��.��و7���ڗ�/�K4����ȩ�渵�樶a���_7�W{QFZ뾳��W^�/��f��t���Բ�f9��z[���D���8�e-C�m6���{~�~�r��B����ͽ3�����.F`a0�'��ɨ�J���Mo���l򇱥j<Zj֮n���u�z��T��p����X�T¯�#]�#�?��X\��N{�.�7�͡]��gg|��?�>����j% �F���˭%�pS5<�,��ř`0�Wߛ1����^Zlsu� M$��w�iH�����x����w�L�t�f_vB�% ]ӛ���g9��1V�p�dM��f�lC���㵓q�Y�Z��h"�7�t߸�
Z��%ގ�]UZT���t�r�b����g�7L���7�8r��$�O�y��t�$��_���m �`~��n4*R(�s�o7z�<��((�J9��h��]]��V+�k�Q�.��ͮ�T�fji�pҹSk�	�Zi@C'��d�/$c�P!+:�}$��d(s�hd���+��?��%R[Y���P9x�+V?=��]]�Ѕ����9��v�t�5�(�*��c�yK�Cu��{��y�6�V�Rw��r:b�u���^�q�}Y��q�-S�?�������R�t�GX]׸�Gl�Ei�ͯ���5C`��|9^'f����ôC.��\��	���G?����dG���B�M�U�d��3��&3�Q3�	R"7�OZ<�X� .���G���}=�;aN�O��5��m�����4@«"���w����'�;����g�Oj�+�Qk���=^��}Q�N�Z����n��q���쪕��f:�(���Y���t��c��ƫ1-.^��5I�S�g�s�?+�*��H�3�2�	Ok��z�����n����-��W0Hm���#x�s��,ݞ�P:6�'/n��$�d��qR]��\k���碞!f��v5�9m�a�M?C�RH���F����Ϻ?Q�FLff����3fW����@ְT����K�LM3�Lo�׭p�!2�N�lQ�e/����Yit��	9_�2��"׬�rkz���]و��!�W07�q��$���9w3�jl��m�4x�#M�r���+�X���ȯӂ#o}l��H��8�y�\1{����h�ּ���t(Urq[Y�F�T�ɪ���g����"e�	��i�T��6u۟J}t��亴+~	�rS��ʪY�~K��UZx�E���O���<�#��M/�ýˌ�m7��� ���z�f���&���#D������՟-�Q?�����.]����b�%�Ծr�l��{�Uc<'^���&�e���\f�W�pLK��Ҕ#.}� �B	b��l��B+ƴ-33��v��T���1��xx�����B��.`q���*����;�4sWy��Agy�5E:iǰt~�é��Li���>\��Dˬς�q��ͽ.�U��-�,����q(}Q6��X����,Eٶu�<G��/4��W`�k	]YD��~њ�L��$��1z��w!x�ǌW���E�KX\�n]*6C@q���S���|7TR����c;/�پ>����h������y����L6�v�m'��O �ׂ�)x��D{�͹RZ�N�Qi�d\��7������i|�,�j�î�F��3�����,w���5:��W0�|-�p��|�O?���.���8~�ő����L�HI�BdT�`�,F`�Dޑ>ў�9�����U��ݩ[�<�s��c�h�;W��U#>�q���C�����v��5e���|`��Ϣ �?�<�W��'���Y�m'�bՑ*s�g��"Y$�Bv��Ͼ����������1��E�������tyS��B��o�:Q`���ώ�Dg�\�NܡG%j�S��u,�Q�P[�< ��Ï߶^��ڢ1i���-q$py~�����*=�q�o��p�N�8}��#ہ2kae�]��qTH�^n){��j������w=��,����b����b-K&���G	ų�cX��N��pv�|p�����.TL��s��=���^�B����&kb���
�4���MK���9���HJ�m�E>�����z#�==�[���W�.��h#ѷ�t 2":�}6��,"�ۍu����؍�XL��Y6�ɭ�.���?���8&��[Hp�W?pS�d1��^�k�:��ap �	O7��$(	e��Y*���k#"��+���u႒�ZL�T+�}�ڐFʓ���ְ^�M���-�[��_��6}v<8�\B��j�gM�b�t�*hI�g-SL˃�2o���@��"4i�(��9]Cųۀ�#~F s��Ŵ�I���m�Zϻ�����G�u��h3�!���u�_��I:���;-	>��N�"��y����~�{zMv��$OQ1�C
�F��g|]~�B(��%}���MYu��R}'�|��j4���������$�r�c@��qK�F�������	�J�Ꞣ���+Rq�O�o���������>EO-��!�ٯe���v��h3�w!�
^���T}��y�w�^��c,Z�&o��ڏt�n׾��7F��e{�`O]E���c?D����e-��>RL�y���6,͊SB+I�Fl�O��/u�qU���"���Ϯ>9�M߲��)�i��l��7���a�^�G2���)�'��G/���u�����0�H��ũM7O)&-�j�^�#�g���h���<ٰRqgţo�V9��3�a�w�C��sJ�2���	���[�=�u��3*��Wϗ.�j�c��Xz�{�|8`��:��)r� Ȃ7��������g�}}!�&2������YJ;1��.���p�kz�����y�%B�a���;�ĭ=�HeP�,��{]QE뜴�s�p�[[ �_<�ʩ��)I=/4Cg<a*`Q�+��,�%�v�"�z��7��V��E	 ��F�����K�~�$�H7`e�q�M;6h9�df��{��
����nE0�A�h��դ�9�v��N�t<4C>�h䍸��>-��	4�B��f�r�_�i#~V�@�?���o����`3�X�Ξ�te�͐J{n�ڔ���(P7#��8��Z6���$k7��	-�%���xG�=�5l����8vPP�l�ۓJ�c+��Ǻg�F�{W5���z\�]b���H�e�����E�>��ݯ����qI�s#:ul��Ϋ�m~"���zL�0��UU��Xn]�U�M�b'UF��M_���ٽ����.L$��y�X<Mq3p��I��$o�)�^ʌ��A��� �D��h��@�Bqd��6-����>�?HL?[47:�G--�.��	 �Ю�$�� W�6���R,vL��<�6�nGU>�����vkt1Q�0���S�E0�Iy'I"�����:Pm��D��sFn9"0C8NB4Y3ɓ��|�b����עY�ݻ}o�SEӤ���ФҨ������]�P��e���g]�7ۯ~]ʾ1}FA��D�����g9WE��]��B�u'��~�N�i�8o1Z���Tv��W��p�.Wʃ\�1kGo�&O�/;O�^����>�׭f{��~����ޅ�~~-)H�:R�g���;�o@��F�m���R����.����_aLH�QZ�)}J�u�K�Àl�ƙf�,�Z�e�Qȃ"�TIj��!����a�Q�;����z!���{�7���ɩD.�J����,��쀧v�S�e?����oZf�C��V0�*�Lڬ�;�I�;���;v���BS�M�z��������.c�d9�c͊�~��h������ U�f�Ze�|n��ȇ�һH�o�n뮵�H����_���o��b���11��-ǲ���{�5����Ѥ��S�3Ł|M���0nÕ���]���U�9�{a�ȅyu�Ȯ��7��-J���.��o��	s��p�1�*����~�_�ȍ�1fQ���Eh2�M�f�_odk�$����_X'��H�D�]$�û���m��U;Oc�m�)��otAK�^��.���j[y<��&{zN�-]W������^�t3�|�|Bۅt��k�g�SG����Oߟ�r�G�&��>y��SrP1�+?jg�V���ii�H*�3�2i��N���vt�]0T��]���4t_Q'���2r:姇:�O���oI�tR�:��.y�m;wQB�Vnr��D�2�_/�V\�o.~����G|� ��r��ȿ��nA�US��sG/s��ן�<���_$�����v���8�27$`?d�Λ_��Gh���2W�2`�KG���>���	Kى��D�䉶.ǐ@,7�8�FV�k��#i4���h�Nt�W���T�^��JC@��=bGb̂��ؽ�[�.w<�ek��溰�+~Id����IZE�^��B�!���͔FM%y��5�g*&������~�����lrY]����^l�6�Ɉb�dGk5�*�����㣉íc�Rf�c�uC3���f�`H�T9�q����t�4��<�x l���id�j�Iܞ�P����AC���pE��I��I��߉\.�\��H�,��y�c���5�ET5E��Y�%�jg�k����"��9��i�TH��<����>��Q�ɾ��yw��n�}Q�`�����,�H"�n*^ߩ������ޕ\<�B�wݾ7m3'���D߿��a�Ĝ�ssV�0_��\�jhƙ)i0�/ �|�,�p���C��5k��_�B>%؄dL훛�z�p1��4���e��l0��oٜ�)쟒�P]>�3H�U�b_9�t��	"�^|��WS�*�ij���+a;��d��mB|+��7�0���]�><�[�9�����Ʉ�
�"',��l�U����}?�l9)c��-a���в�|�\3��ޒI�,r�^�N�b ��l����p��v�����ֱZ����l[�z}#1��3��$��{�*+p
Ik��W^�+�ſ�*���g���Ji���{���쇲_k$XV��*�=8n�i�y�B�+��v��Zw$�����/�B�&&��1M�	�-����pk��N�O|�5IH��`z��j.e\ہ��>�!��I��7�ۊ�+%�'��1f���SAj)�y��
�%g��i�YAP�Y�V�ꈈ��U��{ �`m��H2v�H����E��~�X>$垚��}�?1����"m'g9��W5����k���/���F��Lnl�N�.$Px�W��cM*Y�.�xQ������6ыq���P^6o�� Ěߩ���e^~?�����m
dX�)/�5��P��H�wL����ކڬ#:�2�����i�IG9��|��>!S�yX��C	%���N�coŇ�� ���zm]����%�4�@����474�e�IK���B����j�	CG��R��v~����1���t1�[dh*����`�(#q۞��k����m�8��0�*�j}���/Խ߃ܠ��o��'N��^�'Mt~[~)��Mn�|�%�A��b}�}��`>����?[jp�X��4sD�S����k�yk_?f�����C�hi��21�i�Sœ�RV��l񔖾ᢨt�<W�V��l�Ԡ��:�B��|���/y�|��G4^19�){TO�\e��|�1����ټ*Jo>���i�,Vd�7ަ�%3�����=�!��l���c�PYV��Ü�s��h��O0�d��ʖ�@�d��(]s�'b��]�����S�/h���^f��$���xK9����҇�O�o&����y.t�XG#}% �8����,�2����T���$g2��-ˉ5&"���'"t%�b���0�>���7
� *��}���)�޵��Z���:�ɅQ����b���|�A��"=9�������C���'�����)��Z\�8X�ױ���4�D�Y��b2pK��ۏg��=_
,׸s��<����H���Ά�	7�VC#�����S�{[�j6�x��3~u��*����k��js����N�#O��~�t]��N[������H'hL�F��4:;)���(���~��]���)�@;~��ͽv|Z׿��:���zJ���\�1^����,�}�Y�����>�z}w�h����(V���Ǹ�6y�ZCEG�h�� PK   vOX	�\  \  /   images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.png�W�W��%����K`鮥;%����n��I�EV� !݋�t�>��;�̝{��qft�U𰩱  ���"��:��&�ߔ���'X^���  ���q1��w��S2���t���y�s�p��z����T�|M ��)���YfO�����~qv��ّ��v�C�m��� 91��3�,.���3��2м�P%sVOV����$�\09�U,��Ka�����fv�6{{l����c}uu�ڻ����\"�4����h�v�Y�!^����!7�)�Nʑ��[��������y�B�{rrr/[��q�$�|g�Q\P\�_��m����?���Z�|�}�X__�-��pM���������O{uNF����0M8�W-�Դ��۱�茀��4�7�/c���'ˎ�{ƀ������ka��r-�v����}|/}||4�y}>~�w�R1)d�-�uYvW��������kkkW�O��V.nn�� ��|'��I����K$A~���:���0/�j�ڍ>�^�,��ۛ���x��krΖ[�2��������I����}b�t�#���3jL�Tp�f���%�M��&g>���h����Ŝ#)}V�c}pr`�A�W�rm('���� � ���0���7, ZB��{����p_�u~�>55��ŗ�L7u��aMH����euU�򢻋�@q19n�ViFq�{$'��Q2��SGv�< ���Z3?d(9_�S���'���Jߧ�kc���h���dNF��1�;U{�K�����B�~�o��JL��S�d���b��*��+f`uy��[!s^���w����%]�sCã�~�����������x� �r�fr+�T�^����>uMֵ�컁1t���!��Y*��%p�fWD�����Auu�]��E�R999�e���R���M뭡��'�i�=N�#U�LԾ��<�ۯ���g~��d,x�>�-�&Inv]_���]����*V �|�������B��.{��,s5��D���#��Y�]��f�h,�2�@������?@=Y-���犸��{ǦvFϵ{�����eI��<�T�ۮ�?�=����#D@c]�!��Wg�>6���g�T��Tnƻ;� x��ú�(���F�����.Y����֞N�;=��U�v#�Q�EA��� ���o����T�����<�]Ц���P�U�X殎1��ٽ���ş��z��ɿ�eN�]�jGs���\{{�0W�5(���f��,4��S*��A� sIh��Nw2�J�l�ਜ਼��X�2h��3x��%Ǩ�j�L����	!Y�@�G�s��*�l���#�ie�	IM�f�� �����W��D�����<;a�+~"�
z��;B�t�U�ť�&֗ff�1ɭ�}q��2JZ����vj�6q�^ c�Ì�M���(�0E�⇥�<���-��~ �*�塈(-�?���Ć��$??���q�yr!Y��:�	�7�M��m��;e |F]Z0�u��Ӿj\pW()I�+)�F�8epr/a'?�޳����]_А��Y�5�����ff��Eig������G��i�	��7?���y���yVq�]�x����
��1�fs�(�/�s��l�R:-���^(��6?�s���N?���eu�-�&�i�czkH��Q]��"uj�Fz�0��a��5�f�H�EK���c/I{k`��pG��ߥ=n��[����ڥ.w�p�a�a*h4�Vb%F�J�觍��vgc����<n�����a��eG����U���A�5��֊	w)��~��+����i�f��uaΚ�¯��k����[ ��陙�.`ra�AlqC�h����6�S��'i���nSo�'�$���ٹ����WKF~�!��%�0d\��Em�O]䃍��+��qLi�\���k>
;|P��&�Q6P40L:G����J7>0�e+��f�Ԡ���,��{*�$��Q��$h��#��~�i��*	:�R=�0O�!�������d�!8�۠( 4����U��-�l*�L�� ����\���ch�*���bh�J؆*�m K�1��JM;���s��¢k=�{�5���l^6�&cW4|Y}}wl��j�i{�y������Q�S
�	�Jk����rl(@�%ݴ'm�ڕm~�����=�tLV��%0#)��{C��@Z3��h`��[�0$/x�t ��g�?�H�!�B�tV�+61��BG�nna�R���o�^2�J����+�Oic6|������$��,�8`��~K��	K������儃��{(������v�>�)�����'�ςE�\���udJ�HG����5�ؑ\J�M���M����D[���#y���� طt.����Z������C�+[�H�����nK!IG~\���@�#.f[��=�-�#�=	�k�T����B-�m�7��p�������'��9BL�[Xvل��Ԥ0��L�;,K��Rd�n��5���,�J2^�A�+*RR�����g���U�)��ݗU4�����s�c������Fۦ`e�m6vX�t����V��X7��������F�M���1��7?tK�z+~>�\�鑵z���.���il0Ͷ��z�����o�j���W�)���d6p�n��X�����5D���'�((���W�_��r�wu�5��b��ߏ�7{4����۔iA2�x	O��o�ͩr�Alȅ��o��)�?�P���/J��(��)>�-��qQ֒7�������q��a$��7�N#&msܪ��/pѱ3���H굪F�H%n�58��G̮��*�'B�87�����%n�p!=ExC���'�'�F�+�,�2���(w�Q���Y�� Y�XO�Y;�2�����dI/#|�%��z�0%%��=J������8��]�@y�? gnd�ns��O���kI�dv�E���E�/%����@���q�L}@N?:D���,lJ�#˩��fh7zC���[��K�1Æ�5��Y��5�UEd��{V �8�f͙��:P�h9_���%\�}����7�E�P�E���E��1D;I�8}��rO�C��\�&�Z������8{3ͭ�M&ވ
 p�����4�BtuP'^
��/�Q���[�$���%��U7��Ĕ����v�����Z���*�\�W�U���gj���=}���D�hR#��E0��fi�ۑ��>5eY���3viܵ�e�����hA�v\z��7���r؇�ҭM�iPP6ֳ}��=����u����!x/�E�`�%��c�<���,G��
7Ŵl3���}S�A�:1��	�p�����_�ð5=߉|Xj�W-G4�Ҧ4�����[�8���UP@����m}M*�Q�CQ�{�nK+hb�M��զ�Z{m���JM�W���1���7����h��PO��)�y�~�6�{�$U��F 3��U_���h �=�������l_G�R*�MF)'<���H�~V��BI��vp�66.�+up�nf�p�y��ˬ�������%��#Ҿ��� *b?0r�p )�ʮ_FCg�^�u�NkRa�lI5�x@�	Ub?)�Y�����𷌌z�|�<04�'�m�r%h?�c�;�_O��Q��I�F��bW��9`&aL�8�S�I)�P��M�~3���Kx����ދ���2���qc��)v���4Z�p�o��I��	�jk���4��V����V6��2@:\WD�5F%�D��o��پM��g�\�!��@�����[�Qxa��F]����/���mA�zl tG[r,?ɳ��h|f�C�f�xgW���tg���	Q�!� ����<�2���
��S�����uʫ�H�1c ��$7ے�]9iJ%��K��x|H��?�u�R��䥏�~�ꄍ������p..�Y�ܬ�ܨpS{�!N����� ^g5K��;U�|0�.~\�p��Y-8/�ة�{^|�1��жٟ�Z:k�2rc���yrS���\�M�A�ǭu��w{ۗ�)���濆���w��Xw�/��}��6�'�Z
��b�!�|��լ8#��;�o7���i��I[�P}����Ę�-���;ɵ��,�E.r���aUț��j���}9$���LZ��N�����Sw�웩N^7+Q�ZrDoo�n&���.G1`��8C�
�v�Rl~Yk���J?:>F JM=߹5���%��'ב�pB�U����V��Q���&3��]M}��L�؁����Ц@q%���v���ߵ�y$Ϥ w� ��?��unin��}�[C�y���a	t³�{�}�^���T�U74L-��9�U#��!`ƕ4:� fPpF����v�N��z$9�;q9���cO����{�m?Z۬.j���Fw�*�6��k ��A�R  ��N�2Ͱmz�����B�?7&&��g�Q7��p�%Q�p��*��۹M�[.ԉ�xKK�s�4����e��".�1* �0A�Yc2�PH(i6D�w�`bQ eZ�:�tb�y9%<�	, �b�����C��+�a���&ղ����;[K�������`����E	�sy֝�w��E��W���������̃VެGG�S��tך��X�����،�����)�U�<��x���~�ݹ�l��{Sj�w�)�ƺ�a���k������y`eQ΁r^��;J��r�2m�慗B�OQ9%$�&Yj���C��̪0�[�E�^l�k��Y���/'�O@mILdw��h�7�܉2���c��_q�������1c����~��#nY�JB��g&jfE�rP+�" bzC�Øp��x]�U��� �I�����gN�@X�5`/9�䊌,�&��>�<p��s�ǆ���zu�k@���9N�v�o��=�	��y�Z�k�.�>Q���+	�R��igF�̚��T�Ǟ	����<D��7w���vUk��ٔ����*�'��'L�.��-�� q[PV���eOǻ�W�q˒0P������sۢ�V�SY�n"�T�N4@�y�M�ܟi��{f�=E�}|��_��#��2����W/4oT���=B�`H�֙�ɚ��JS:Ed�!e�%`��n���q�v\.��p�p��]�l�(��"�J\𘵾V�v�m��g�B5>�w�'�%� ^p
q�nބx��+��>�f������k�Wj��|��j���o��_�ʈ{K`"��vZ�,�[����=*w��Y�R������i���
��[˵��ж����,�"8�s/�(a���M��;�?Zr7(l��U� � 5<��N5�?�Zxn���~Rx�$}I,�OYQ(���8�-�z^��-$�W������0cg���Z�	ȋ�)��R�dA=͸���z������Y�\�+zl���y��8Ϻ�q�=�����6:8m�R��N���`-�J|�����,��!V#>N��Oq�g_�"t�uU���hX7o�m�i�Rr,L��z�->�#8ÀU�#�	6�s���Q69��&��w~�4�~���VC���� "�����y\U��j(�S�����Σ�Z�X�k�O	�!�$�~Q��X5�fѐ���,�4�#u]�1N�.8F=�Пux���|���(��:'�/C��[<�AVĐ!�j����˧��1���:�
�]�}1��L9�?eۼ2K����l�vr:��{��_�3I�p��P���fۼ	O����(a����w��r������̒I|=�����|K���'wJ1OU�#�AT?�^
q.b���\�kr���͸洘�%�Ct3˨��A�|ؕ��`�� �~�Τ$�-�'[
iXS���J;c�wso�H�=�
�w�HKP�~�^:=�!���B��3'�z��G����Oʑ=<!?]`;
�6�������H�&��5U��,/���P�}��մڢ
3V���\[@�e	O��i̝�KBm]�V9�}22�)�u1z��I���B66)X&�ր��1n ���Ph�ĉ��ۘ���BG�AAa��S}}ɯ�*��I��z���C�;i�F�DV�O�	�GV6F�2<��v�����'�/qK�E(�Wኬ��b>��Jbd<���T<�VJJJis]]p�R���SM����3�rW�����BF���7��!�����x����!w@=l̺�㮌c��*3��ڂ�L�/��"U`�*_�!��?��^�S?�z���I�^E��[�ןb��R�G#��ݎ�]���z@�������]ϣ[Cگ,��j=���j����4ݗ=��ڱ��Tu�:$sy�ab���0d��1�L ����G����5�>9�iزiK�VFQ�f���u��?FSS���X^s��Ja:���?QY�����]ǁ�%��[����n�t���>cd�n���5��e�#n�{~co׼�X�LJ���%��2���W�`�ee*���K0Ȭ��RX}	y�q��/����(���L.,~�{�r�*�Ţh�H@n=w�-�˄M�8�sũ
�Z�1����sqw��5?�mVYuz>��7P\�?5�*l���R���"�<=�j�"���3��ՙ����-$ ����I�7n���b���1g$���i�����9���L/��q�#������&�FFJz3�U(SR�S��y�.��@*�'Q1���X]�./��f*�����'��$::��Q}kY�u!>K��~�K��z6x��0晀k�˻:ݴ�+#x+A�`w7�s�dm��q/ɵ����\�ig �ִZ�$���H)���Hd�g��u��#�.����[S"��u:�
8��k5Б�~�(4�}��iM#�����32y5r�`K���\c���׍���g,�d���qJ(�HDKR�Wuk�WY�
�ym�fg�ؒǽ2SI)W����qȮԒ����+�ϡ�36ZB�!B��V�	�(�dϓ�S�,�g�����g�Ih�Hx��Ȟ��|�b��.8x������+\b��O�	������_�K9f�Ð��n��T-�w�s�Ǻ�奯O�F�e3^�����"X���/)7�z
l�50v^���f� �T��剡��O�Z�'�jJڊM�6Q�PK   vOX�R�{� �� /   images/8b783ee3-b9bb-4285-aa49-cf7c99b593a7.pngL\TU[׽tws���n�A:����ݩH*!� ��P@D�S���������qgǊ���{A�kU9TRT�� /�!,�@�JȈ�'(�.��7x7I-d��C��z��E^���z�����>$q��s�t�r�2s}����u�w�0sy���j�y(B
Q��_iyg�/z�i�y@:u;Y�F�FA�� 6Ca�b�E�
��1 �l&h4�'oh��u4���M��yM�Oڒ�~��wic�7g��}��æ�ͳ�6��v�?�GTĶ�傢��䙝��������;[�W�L8���zg��$�=U�9wL�e��	�6�H�E�epd��ӏ���̓���p�����e��3�mLaׅHk�887�}� iii�Rn!�:縩;���ƹ�;;*�^�p&
x|>Y�"Q�М2X��a�`2'�1��L]V�<u���aAa�d�G���O���'�*r!>�YU�4��<���f��}Ree�v�vW#,H�P��
�m���C{�ͶPr��5.b�#<��g*�R\�||*T\uܨ��A6 u�����2X��J4��-J��i���oP��H�|�hZ��ݢ��y�C� �����i�)As�x����������ȫ��T (󺴔��H��J�/�5_U}��:����U��P������Ոy��	�$��E��g�Ϭ�����}���Gܤ�f<w�k�ԍMaP
� |Bq� � m�|5�j�S]���W#���ي�a�d�/Г��+�k`���w�A�Ze���<B50�pI�T��o�`;166��֢@�%���s��DK9���Ң��~r��t�$ m+I�(P-�ewt}�g�Ҙv%��O�n,��|m�n˺��.�:[�}{M��=gwL��,�9�L�?�qi��(��.�P"�'�N�#2�[4.Ab�(���~tol���0�'�+&�SE��ޤ�Fuc�_�A�O"C/[���u�l�=!B?���L(h�8 [�m$x����E�|gW4�}����nR�zYb$�''5�*���JZ��U7l��k}'I�8 4U��J�IIs~56����[��h�f��toP�5��|V�g�%2<�u(:�MJS�۬�;�8��PX.
�P�ɍ������1��=��{5��>[�۠�u���r�@�'oɟ'w�°i���5�+��cZ#��<��8X���5�ˊ���$&��U��3hȃ���$�!�dx0��LS����4N�I� ұ��_5>�
�hhJ��S�������XA	�ލ%S����h�[�o�(�_Q���¿cW�/�������G#H"`WvP7�Fb�ޱ(�%�����"�=�vg��9�����;a����$^�gt����'��D�`,���H������7�8�I���`�z��'�#�y�6!����|�o��~�C�7[�o���$wJ�P��E�KPډ
��>t��.�1ʯt����s�%��VL��Á�Io�UL�T�S։����W�-I��ӝ ˜�띚g�쐶g�����7O�pLҎ���d�3KYLz2�`�H�T�мn!�e� �`�~��/����^��n����ކAv��]g�͏��t��q�`�=��T�>�Ҽ�>��-P5��\�?oOǖC-ڙ1a�D�0Ы����u*ƶ�ӡX�5�����Dk�k����HTb��J|4����v�a�@��
��tO��"�d�B�/�$)�h,0�O;ӱ޳N���v��T/�x���x�̙:������$�Խ�dI�O�o$s����0e�MW��#�`�g/��a�H�#�g�A,t��\����'�,�����8L��>`���ڟ��W[q�d����VU�ӑ��I{��n*'�s��	ۂo��G�/�"&�.b����1����Kz%���s)n��Aցl$��˕u�Y~�]A/����7#˥.iJ�z���rhurء��o�F��(1o����Ud�
Sz���Ua=Sz]϶D;��#�VEW���Tc:������:C��Y��z(ӕe$�D�X�r������3!��0�ɥm��I?G��a�nk�ld^����+AqG*�!�����IĬa��k�lp�W:XȔ���δK�	�T$��U�*x����Xf0KN�E%@J��@~��<:@���K;��Z��);�ߐJ����2�I�5Y�/��7>н��A���t��*�ޢ1�G�"�1�b� ��BϦH�9�|>�r�Tb�E��?�O����%��Ku�&kេ'Az9Qx�m2���s����r���~j�Hdp���)��s!ʇ�X=���J�?��(�[�ک��o��Q�����q�RO��o[������y���-8�D�f�8` ��J+����f���v����uѩ�4b��j�: ���0�[��>��6�D��B|j����B�bt_�ƿC���Ü$�|�l��++�;�Y��As9:b���w�f9E6l�C9U�Y8Hd��� J�u��;��m��+><I��L�0ld�]!�9s\d�����Rŗߚ@ rU�9�P�N$�\� �Bu��7&/�a�Ru��4�v�����z���~����zu��"tR\��3�l<�c;�w��T����	�?�h����z�$�%mk��uࡥ��.���;Ji$S�H����ɸp�=�ӽ�O�3�Xl�+���h�)�>����*���o%x�`aHy3��#S��BQ�J��/� ���'���)f�sF���2�!0�i�B��.��mZ����/Sw�9ݬ��M���ӐWPJΎ��u����wݶs�g������E;*zP�)��.g��A=s��&T/�"�x&@<z�I�/��x��p�а$�;��פ��W["t���Lm\��R���-+G���(��$��B��w�B��>W>�i5� [Y��Y�3HE�g�����e=ȉ�Z�G��(�S�(�;�ǘ�d�vl�� ��>�v�a{��Ν݋x��ȳ��q	kG@\'�Q�&�H1�NM�C�ε��Q�7��{�@>�鐿1F)��y�3�y$2���U��-k������@�d'`�R�V�,���YTƔ�re���bb&�9~�+�K����85���uJ��kӵIz���j_`!j��)�wrn,��'ש�՞KD�H�^l��hN�b�+�\�j���I >��Ҹ��ȣ�aH�e�/M���8��S{)/LVM���dV���TD�5�f*���k<���zIBi�hɤ�K�bq��a��֜���S$�BVa�C$GZq&�;(��"�3~:���m�0�^w�x�ۡk�r<�C�Oٔ�!������8v��A�ϳ�v%���DK���
�؏�9�c$���vf��Xr�����b���R�2Z����I��2CI��;%�*w[<Pr:9R5-ƈ^e���w|rH�����LM�w�<n��Y#T5�-��Bq�j���O�c���mƪbu,]����Z��F�X�}w�Ww���Lk��Aq�����oK���?�/>O��pP/�L�G�L�+(�c�Ky�}V�~��'u^��
��1n�ٗ0�ì���gS$����.�)��̆4~�AF���zo��Q�g���ia�w���{�!?�mDn����=W>,6��U����/�������k?q�"
Z�q�����E��
�!8��_�e���k�9aq1���$�!&� �n�PJL=�%�T�\2k�Ѓ�3g�Z��Tx�
�H%�q�~�t������(��=.f��ޯ��EŤ7���~y�����?� �[����'Y?V\��V��Շm@�&��
Ԓ�k[\��ϫc�1�����{��F6�rv��� ��m�!IW@^~� �&�#�A�	&	�f0��z����nW3�DJ�S�_��l���s�t��Rg��J�cej��iEC��)�sف/�IdxQ}<�f'q6y����:W�YME��Д��7zZ���T���l�0ܒQ��{�| ��3�pnJ��5=5ðP�"�<Hr�/S�x�Py�s����Ëԣ�����Z,]�I��<���m0H�nzk�/_&��+��-��Z3��̴�Ma���l�qXD\�����`y�K1:�×B1�����I�ԶC��S��꜑S9H�
c��[o��o��FDx���~r@YI�Z$"RQ���A�V����3�O6#P���gj;��m�X�$Z9NO�J�|�����A�Z���l�S�� ;�WS�v����)���ybg�$���z��}\6��^��������
 �@&���v����I?�$�M�gu�B������T��12S��p�x,%W%�7'����]�J�����@Ħ���g����Q�� g����r?���/1:���ǚCՉz0y�?���O����!i)r<ط���Oz�cT���]Gt�oA�2�����s� ~(hW�4֓�_h(%���[e��t�2�X�^�t��K'R8�����@´�&���(�C�֝�o��}�����[��$̀IX��S\��'�`��V{���|�������Tw�ev����Ϊ̺ͭG�\19�ʝ pm(ʃ�;�yL;��F������ 
^�e�_OG2�lo�����e�]Y''Ї{���+��f��CN��HU��{_������Li &B��b�=<�[��j�Nj���ྱ�L�:�5����U�f�\:]�{[`âVC��j/r�+i��9m�{w~�:u�?Sy�B����_qv����X� ����H>eeVN\�|���)�L}�4e-)UP��S �Ψ��;��@�C�2�������q	�t2���=�H�@���9�;��x���=�/�����+/����aQ=�d����y�Z�'E���<���*%��Bϟ-ڙ�{��Қ�h�_K;�UE?�;���`�PG����6Y�={.w����b�Kq�ׯ�N���e݊�VD]�ßW+��G<����*O��������D9��0�	�fɳYK�_kLF������ȫlz&n��~�U_U'^z�M����LV�5�P�����d��ԿJG�?1Ǵ�����<�r���\����vb1��G�x�(��]O��>�zMWA��:y���p���>�b0��u��f �o <R�Y}|"�+QƜ�K�"kT��<R��aQs�f��FI%EЄ��mߌY��i�w�|�w6��96����Ar?^ͭ��Ŋ�|w�;��4�{׊�vu��aDL���{b�Ij*	�j�`q	�%������]�:deNR
��\�K1<0-]�p/�U' .p�%+����z i]�2vL��C'��fc���'=x��E�R��]��W��Q�j
����k�%3&S1kx#of#,�|bߗ�	�n����!�0,.?�HT������0�� ������e����z�<.��S{_$8,�Q�/&jg��R��&<��j�B���"%���[k�%���%1y�l�J�	��g�3%Ú���l�
&���Q,޵�u�7��n&�@�\~�fj��D1a��J��6��m�I%,J��_*�Й��v��
�3)��v�/�/��S�m�i��+��H���A�����8���dT�櫚��5(�q�n���H�T���=غ����6=9p��3�2�"��T�k}�cK;�eg?�w�p<0�ğبG �AW��*>w����O�x��H �F��ăآ�q��k%��4��)��!��q� S���6�Ro�ӓ-u���L�P@������e�hCK�����ݚ/PB���z,m����̈́*��v���pQ���!ʙ��@��ֶ�N΅���^i�Vs}��&�O��JT|:*����W���7_�ݯ>5]�����W�`x��v��<��Z/`� ����N��=�?�UN��J�!f@O��fR&�_����?���v��ƩJ
xu�>�V/���6�RH����)[؎? �� z���N�6��T��h:Z��0c ���FL9�w+�X(�L� ώ.B����(2R�����)��
)�wi�"���r;�S���)��2@�)7�P�gꥇ�Q��bߥƶ���Hp-�RBt(-P�?⺁4A�����5ȝ]�W�V�X�����)?���6eR�x�	`�0ת{R��:6��Q��h8 )�Z[�u�.�R�\ڽԘ$M-����8�n�?�mrӽtu�:۞�b�Ą����y�ϷQ��l�m$Ag�+^i�:f$�����UGq�����"�K�M��Zo�>�[�����^�Yj�!�����i�	[��>!�&�������W�>C�ĴtK0�c�"]�:�t��ņ�;��.V�$�
ߩ��y��.�k8�>��5�Ǖ��^d���8�H���:�j[��1���j��3�ߘh^/4<}�'_+�8?l�
HLʃ]��F�/y	[I;}�q�{s"��|��1Ak}���7����ך��Kg���Z��?���w�4��6Ț�V��m6'p��0���Ǩ��X"���qj��4,m��즚���t�Xr�zc�'�C_�#��t����B���Cv&ڍ��l���2�}��1�L��^��0<�;��w�.wg&�cY�\T,���Bp[��Ro=����3���{|X�J*۸^b_��U>���ҙ
w�w�/����UL�i�(�p���ܣ�c�7������a�7Sr�6�pv���*��9�|(/��M^����� �rHK���Z�Zǹ�W��	�u�R����Ul��NU�U�����mkd��)�S����T���j�X������DIc���ËcqPlxD�<�q�#��?:#���[W�Wc�JC��(�4�"V�ҡS[- 8[�w����m��p���;[���6���Џ@[���ε�R�Yl�hH�X��~*�y�D[�}+�K�@1��<�1A������A�3z7�M�3u�z�_֏"ӊ$NI��#n��qBM\�)�\QLw�G��E�k�-
��I����8i��ѡm�99C�'�r���K`
>!L���`	`�l�rZ�,;�t���0�o�5��z���!���y.!�*G��Et�&��8^��2z�m��6��.��^<�B[�Knv.��I�8e�]�- B�M� ��eN�����[��g�ܕvf-Dj�[��j��`E�OM]6�!9w�l�l�����	�y��E������'��}p����>��8$�B����wv�b3����\�E����<~N�� ��wA7G��G[��wE�N/�TQ�q,=i~퇀�mv�R�t��T�:0_n�gR���
,��+����1"X\����-^�CU�]#a6>�l�1�d��ne�|]J��>��i�na�)g��qy'�b
�%]���M��0�(����_�ǎ{ɳ�i�e�v7���ڞ1v�э���|�)�M� ��'�̚tR_4��pQ!����������1:E�h°��q��.%&�!����E����<�H�u5+�Ķ@���"��ͨ��zW9I�QV��������VwxvI�w��e ��"�ęյ����
U������l:T�Խ+]�NU�'i���s��ms��N}^����ķY�udi�����������%@h���r�wM>5����
��*~�
�o�E:����	ã{I��G�&�I�t��"�&��Jq_/�����	$,wx̰bI4d,�#۽ҐG�1��D��
�9$T���c�ڑ{N�Ͽ�%��ݤJi������ز��V���=�F\�=X�	�� �?n1�Ƚ���f�6p�K�z>^VR΅�
c��r]m׋��j����VI�����B��z*��2�FAl�_f�G�;|�,�p�vr2J؊!�K�q���Ā䰷*\�X��ɝI��v��y�����g�倫�u�WQc��7�U����?�)o�����`���� ��fdf��������w����[��*�����+������.�\2_/��l����Ɣ��]�3��VG��rH��P�ۊ���D��P�Q=N5m���}��������h7��6��G�l��p��=Z
sDj[���K��t�v�����H���b5�ꭹ�V���1��EV_	�GF(���LŸ�Vlƪ_F���Hlz�ϙȿ�6[]V��������^���x��kQ���Z��-|'(?�F0���.��ar9ғ��Po7���"��oԢ�8���Q�r�m*uE~�����.dvQ�������xJq�����PO�G�W� (���?@��S����K��j�����J��r����ؐ~y<����FNӊ����`T3��Y�YDD�Ҵr&��w8�>��ì\��-{�"�i;*Ew=�Ll,s롌n�c:ѮZ%[�Ni%�|�2�=^P�M�B��3NV��N�#\{��O.����_%{lS.�Zf�*cs2J��$Gڥ}m����B|Τh������0�U+�(�Yd��ٰ������ڥ(����D�Ñ0ġ��~zj��m/a5�����0a�lxW��`\��d&��\�x\O<Ό.8Z�a�خ�^
��KY����󗾻frF�l����L�[l�Z�S*μB��u.&�ts�Ka�d�/��"�=Ƚa$u�Ll��؞��J#�˾�?���G��LFa�Mj1��	�ؙW�Y�%�#��a��ʃ3r��xn�;͇�HoX �&�*�E�ӌ�Y��K�K����r�� ���gip�/��
� 覜�"��6�ǋ�9��$�P�1�d},�K�[,i�#�������a�����*���aBY[
����H���G�ޞ�i|��pWL�#��~���V��d�SwL�O���$q�D`W�?5��"�k�Ǔ%t!�7�ƓF�*�yY2�ȍ�XQ�"�_�J]�sBN���&�<j~�(�̺�X�5mR�z%�q��ci}��y������g�g5���;����G`	j���B$��t�p-�(�S�I,�w�g��.n(�.K;jO�=�J����?d6Q�D�5׭B�#YO���h�]Ri貲�I�w���m�ꧏ!?���j�m-��cVܘ��d��M������Ov��:�N4i�ք����:��U���H,!Ԭ�t�}�f��1���'V�<�ӽy�,��vy":�E}�'3o�\���(���=�·�D�0�D������uǽ�Rf��R�`�Ȗx,��t�v������8��ÃK��	�ek�/�,"���V~��R"���bT+������Y=�h����C�z��&{sZ�-ZE�+߄�����UH�lZsQ��R�| OC��Z�'�ڑYO?�m�ז��bNo�@=�)]��x�)G�#�:�ܓw��Q
�S��o�B�eI���q�'��vV4d�}���][�L4�H�]�ݧ�-���ޣ\��>!Lx��c�����ɡ*FJ]�LH���H�A�c���m\$�mGZE�P��� �z��miXV⤛.)�4�&t�%;�z�٨������ƽ:l����P,ϩ���KS/��ӻDsq
х��E�0��K���ș,����4o�n����:GGU�-���p�HL���'�Ƨ?�%DQ���������N�E-�zx���ё��AO�ZW�`�:��uVn�|�f���������͜����qↂ�u����!�
?��G+��/��5�|��^կP��-|d�.t@4�%#E�f�>[3��ϕ��n% ���u*m�'["�b�b����F���aiHv�R+���>3v�#q�?�[6����}�9Z��<��gx���ó�cގ
|�="��?v4N���?>�8x��TT�$i°�ܦ�LQ9Tn��*~��[��SaKk~\�'�<�/=��7�D�q-�i>�R��fA�yq���w�,?�<���M7-͖�
	L.�Vc���GI�Zc�)�-R{OE�N%�5����vK>�~���}]2Zfװ���ҁI��Er�p;��f�j:��S˸	��Q����Х�b���?5{K��� q�c(L�İ����{(@�٠��
�oӳ�a!��ng�=�UftH"��������Q����f� <��q󀯦����7��c����vTWtu>���m�>(��.P��aO������+z� �q <2޳�-zA!3)��ײ���-!�%�-}�D�*�z�s�yݢ�f�f�$a��Od��t��_B-����˵�S�@���f�o���������s��Ct����B�8�*_�M`'x)iԴ0(62^����WEX���1�z�c�O�[�2r�~�ʔ�/��v�ϳ�ҙ���oH��-����d�WA�6�h26�c��b��.D��`�p�E'C&���2�( ��j��nt>�u��ʢѓ�E#�� 0�$W��FDn�K�#a�E*z����#�o)��T��R-0��7^��IJ�}���zCݤ�_�~i�I��9��C)�<}	 �z���ś���?^����W3��e����N
�����UO8���܈r�]vk��,�7;g��H��H��Z�m��с�ް����8M��`�Ȋb�ۃ�7]������\��a�6j7��S\���0z��>IU��=�>w�=�jq�/�䔌��]�P�q�;���XA1X�A]ϭ@<�/b�5����z�C_>�v����@d.�����m�I+�a|v��m���A�sӎ�{���Yf�k��%����/+�5��Wë���гܾ�;w}q�r��,Z����+������)}X�h8���q�>�0K����~� W%�}���z
)��,��FM��u���A���<������'���AH�ɋ�����N��ɗ�"h������U�������=m��/��� 9��>M�ru�8�O:}��>Q�p+҄���Lr�f�H<ߍ�����9�����v�dfӁ]n,D�;�K�ͭ��մQ��T ���<��F���o�'�/��/6��m�֧���gd� If�wYV�=�	m6��-|ߟa�+l:z�ɩG�$�~��잒Õ	�|��=�L���vMh�۔G�Vg�C%���Z���\�	
A�'���G��� +����~LQ����_ok�'�R3�Pғ�!�B'2���l/1E�d���C��m@�I��$�8�sW�Mm�k���˞�O��O*`��FJ�D�����ۯ��D�����s���!2�W���w���5��u`�<{��$BV)
c��B~�^jgO:Ns�{BXkot�|G�b�R�eMT|Iծ�اp�*�x�3�k����{��t[������o�/92�{
�������ƅ{$���4���<�������c[;�|R(�B���uC�3$�Z��T�kD��u{,;��eT۸Ҵ�,��E&_�ZMk�Sm8d�O?*�v��v���e��p��Ln��K�a+:��m�#�}�ʆ�o�t��_��R]��-�-���De�YV�U��aG/����s�3%j���d8�M%�Lp���	�wQv`�7��d\�IYA3�[@��ߓ�����c��~D�����qFb���sHE��q�l��
���U�b\7y||��̰g��J-��-�X�ꐣEV�*��S��YN�3#!;x�.��-�!0�V_��>�\~v��M���@o�ML��e���C�M*�l]Ł��� ������:*Sbpx��,�d���~;9�q2�׷���Y���[j��U�i/��?�ا&�X�wL�Qfu�8�����B���D��\[n����
{$�MT3d}��l,]��,fH�+����b�Ռu���\�u��܇�0U@Vbi㛍"�{��q璯���#�L>]�6�`�t>�j���UO|l'�?��� �`Lep�����*yz�넰B2Gt��LF�v��'�x�`����*S�b$(��;e���>�������q�]AVxsp���5�����`��՚аjW�Mr��?�>����$�2���K��O�U��RZn�������{�7:�,���~}��,&����E=�mSR|�X�S���d$z�nϣ��忔�ͫ׏>�����bKF�$XS�[AQ>���W�2A
�$��(0t��k�/��	�2�?��Y��u)�k*�%����gљ�6P�"�J��2 ��w�*æ'��v�V�<p��2-||$z��T~!$�������s;��Q��0נ�7g��_#_�x��̸���U#���zH?�5��}������7i��0���
�q;7��5�l��>w��v2�֋&�7�w�r%��Sm O3�D�(��hI$H8vL���=a��7!�@P5��7�_�<z\1��X��!�Z�}����]�γSM��K
P�e��M�a��2�p�z@*�9F9����=�r�!�W���ʥc���L� �RL��=@z#߈W��Qe���H�YK_t8��j'\�����22s�5Cj������9�%8<}�ܴ�:�M��2R��bK�b�������?�W���{�s���o�u����ګ�&T�q�b
����J$$]X/�eljm�[O�����!��N~|� hj:�!+��;���D���^`�Ho���$� ?���N��kV��xK��m��g��$���Sc	L؟,�Eb�b����@��W;�K�K}�O�W�4�Ҝ���<��r���R�+�J~��^�����Eq�� J5z�z�~�Ӿ����nMHe*�V�E{�cX�=���`n�7s�G,C&�P�!��Vx�	
�ՠ����������t<�9��K�ˇy�e�sч<Ư~������B(@�-.gS�$�����̡!����	�De�e5�Q눅�������v莛�� sq�\��wt�^֨m�tx������3�r��6�߿G�~�/��t�Z8=��1f����\t4�SUg������Qj�.'+mד��Q�~��!v�Ult+�g�d����#��mEe��i5�M�NtWKݢ�1^\��%��26�֬�(��3a��:_���B����he{��k)���U����Ä������x����Tx�#�/��7ɣ�ކ�w!Gf* 丵�����7�[U>�;P>�:�{�xsb��Wq�5#*�΄սW��?�TS����-^���?wi}X�n6�҅��pi�nO�"<|�`�)
ԯ�2�p���ORy�-��1:ʭm�����b����!��ug�����k�L�v�w�Ӯe���u�F��R8�䕒��ռ��"Sa��ˋ���.	6�8i�mZ_� _���[U�P�~'����I#���)Ux[µ͇�t����k�~���һ�n���>�Ȧ̧���������?]�?t�V�Fy��Q��m��	*�y��|��� �N��;�C�>����N��~+ձ��m	��n'r?����e-Fo��AG�����_����.,F����Ϟ�ԉ�Q.Et�S으y�$"_P��[����Ec״zy�<���w��s͟�Ė�٤k��kt��n\k�1>��=!�Gr����@�g<  �ɸ2���q@<ȹ���y`��I&�q���r����D�����s=]��4Hl4��_��&|���~�9ƕy�<Ϻ'��|p��و����d>$���Q��Цȭߓ٤�m�mU�;��'k��-0Eu/��)��z�� å/il�wx=��j*I�8x_!����v���6BJ���i��� �Uذ}B�dE*�k�ַ���$���v)�z��P_t�m���"yl�*��iK��T������G$�O}6n�F���W��"jn�x'pη�s7�R���{�jٝ��n�랏R�&j�}���v�	Χ9��]��ܶ�\����+G&����r�(��[�_��}��B�C�~G�98����L����d)ꙶ}֌�����7D>e��0�L��p.ՠ��m�@v�3�8�	�} ��yZ��R;����u��ܿR�LQ��=�s��աW�^��1��r!=�������r|��~}��^���$A��n�Z��u���C�@q�r���Wr-kc�NG��6�Eyö����
�.�~8�	�e�W���GW�Q�����(�^�y�D�������>5^N�^,&����Q�]v��^����4�����P��:��d}p����&1wb�N����Z)5�ƹ}�(v���&'	ݢ�.P|h�6���6 , �W���<-�w
���ћ���Uv2�u�'�\���-ܳh~�u�ױ����2~�&_]�W�]��'�N���cL���
[��9�4$=��!�?��h�2|�u9K+�R4"�����(X���?c�}�QHE�ڮ�����{�a�H@}��|�X�K��!���L�4�8�����̍��ݞ�]y����)S��G�ڨ���E��s����shݩ�ɢ^FZ@�O	�Av�c'C�U��H����z���E��~�?k�w�:K�F6�A pYo3�fv�/Ic����� g�+O��O�T�@�ʎ����g矩vw�����'��#���9!45�.W�M��~��.�F��e,��i��i/l���� l|�"�8��f���{��:���Ϊ��o�ǫ����7�,@� �7���Ƹ}�LߣM1�ҷ_��@���co&�K��g�^6zu�5�/@�g(����[L��9��^��!qQ9������X�Ҭ��AN9���*Qz�Oy!�/El �"(@]��⹗���y�"����iߢ������T�'�Д���y��wh�q��������}�r�V��=��.w= �o��Ap�W�B��}>��	���?��Y�(�P�F��t;��Z�H~_�u��T�:Q�Lc����Aރ���힂�	����,8�_���z��O�.��DWqe��Ӭ�����M�b���P��@�����+aq.�Q�,�eS�� ��d�K��:�ș<�"�J対��\�ģK\���9�KBÁ�`���#�[�����$��:�v����b��6�����M|U��֧�p��Q0I�ɓa.�K�m�63&�u���k�zϫg����h4վNi���1��pG@��'��h��w����FR�G���&k	��C�Ǵ{R1���?"}ݢ��ױW��s�#{v�������^���YX"�L�}����|�,���4�$���S����*��'QR���_��^x���D�wD��WCp�Z��s����\x���� a��ǓS��:d1����yt���q���z�b����f7@9��e1>x�����eb��'�;:Ľ������^��M�A>B�&���\��^0A׵>+D������=h��U�x�M�������?��8�|_]���`�"[����ѷ+�w'3�H��p ���#E�Lۤ���=��;L����0߄ˬ����4:�s��|�|	�;���9wM߱��0�(�j��G_I�����M ��&�Y�7����a��4�	.m"�u�B��Z�� b��A^��͋���R8� 9l"1H&��˔6�կ�2�d�Ef,4O���J/b�y��Ԃ��=M��2_=X$>�����ƣ؊�몍E�kw�U~U�=��~}��P�'&���_��\xь�*�P�������~.\譩9W�؎r2�Q��_�h�IYs���/�j��#����]�3./��ͽM�ފQ��o��zUhc��qI?�#��r�5�~�x����(a�`N�ц��Xa,8�R���R)�r�d�y�xS��Ǯ�ߌ/�~-"�	�<m�O���ʬ��v�yģ�k�5z�^�0�4�Ni�v����[���sn��_v�v%7g���<_e/�]�G ��m����ۊ/�@��T�*4�3���$�ɝ4[�����iJ�oҌ$թ
G�5*J�ʾ�㚺"�vJ���_v�N��%B@.S�ۥ�]|cĳ����Ʋ8��ϧ����]�Y��C���9��7�8K�\��Pk�+��O��Y�*h6N���>.��%4���;x}&wrkx�_��&��?>����߭�+�;l��N���H�|	3�1c�GG$��&
�@��>O�.�A�Xh�3H-��v����E9ydi�%����蝈��Qv(��p��aS�xƯ�W	�FZ�ݰt�,;�>�f��{�?m&��a�P%g����y�����՜5�^���,��6Z�Ƨ�0ґt�i%<�A�C�"��C�\1�6ό�k�D3�DO[,jN�w���!{;�|��Q��O,r"����~a�"�0��V��Ԭ�ƿ�O�7�oUל!�l_��G�_`��tňv�Q�5R�(��Ǣ$��U���]�k.k��!�ll��L�����	j�`�3>�۟���<����-[��6h�6v���b�'���~� \Iu��.X&�ÖD��^|
��Z#ݯ�`x_�K-��=�$ƹ�)�S��nbş>Jdp�V��X�b���I���I;#Q�'敽z��0'�����]�����a^YŃ~b_���r�LJ�x�ػ��s��+vb��r��:_�����6��:���q��68���6��j�>_��G�;�[=���F�g.~��[@Q>n�#����:�C<�{T֧�U?���%T�ħ�[|S'v;�~�Xٴi��6&��:f��9�SeS����GUY�%�@���]�q@��Ӡ�4���BX�6�g�PN�Z�r����+�[�ʳ�&�ٍI�� v����J��Q*�o]�}w����Wg0�rȫ�F��Rr��,;sb�N����w�%vl^Y���~������辷�$�m�����l�ضm�h�46��Vc�qc[�ɯ������̞�׺�f��(���N��m����YJj
����mCn�a��R� �8�*��k�\}n��/�L@�n�2+��kC�~�e�vW ��1�e2]��$7lqʻ��z����|f���ϱ�k6�/�
Ӹ3zƭ��v����K�C_�����'��F�E���p�ι�+A��[i;�P��v%���Oծ=N(��]o'c�<��w�M]���.(�k��E��`�^��/�\�QNm����4��R-�źH��}�������Y�fm�ש�K �t�Gi7���0��)��$��3�����N���9Y�|���!��t?j�w`�˱��?𫳃�74���$��`W7�@o�����M�����s���n�	��OF9uu�?H�-r���Ї]>EG7#�?�l��<��+�o�t��=�<r�:�|h���a?Bk��A.�TS�)���d��D�WK?�8k=&�������y�8FP<̝캉R�8�f�D1���
i����܀��#���:��XU�Q1pn:g8�I���_}ȩ@��"��Y���e�������b���pt��e{�\P�)G��I���Z��K{U޳�Vz����-�9�Q'q���ē��$�5�_��?��b�V�'�;eۚ���)���̳��%��._���N'��޽�&4�=9n�g�,���G�?�W���$�m�p�o,��Y�u���S�]��:�3�A�V>a�!:�F����XzrZfKO�r��m^�D%�e����`��{�
"�+S�B	�y�wrO�y(7�_` ����>d�b���&-�[�OD`�>��K�h�W_?4��Q�,��N�En���C�ВI���IU���w������Sw.�X��[5r%�j6��7��D�秃�LҎ�>�?(�3y"/��
PS��#��͵1��7�"���`%���{�y��������On��l;�[�4 ��I�d�\��������d=�Rt��s��5��T2a��D���t�5����@Aң�ܚ,t+pbd�ܢ9ht���;�H���fN�5��EΝ�:���f-����؊��{����)����.�U΍vZJ�pO\gp�+�w�/h��ۣϖs�<�^���Z�=OЏg���X���߀���׵�Hڀ#�_QY�5�p\���&&�᱓����L�s�F��o�JE��p�M��L�"�����J�Y�jA�3w�������^�����9��;be̱�?�D�x����_.m��V̡>�?�/��XHc�4�����)m/�3�S��V����2��j���(ԫTL���8<�!�Ʃpl�s������Г��׳����eG�f�g/n^ �>t���1�h�I�P�{�zG0}y��nqUCs6���v�?�o	Я�Q(�p��&)�\]e����NW��t\C"%���r�:�u�A�s��ǞK��b=��\\ ��r�q�!{�Ý��s�; T��&��Ԥ^�GH�܇��z�@�Ja��A�ð��g��ƶr�Apq��o�HY�D�J(�in�f2�|'K��k	��R�<�� )�Fk�����nu?h6�iq���wqUTN��yk�xǯ}?�[I��pt���H=�~3w�:t��:@�P܈���Ϟ	`i��y��
���IB 3`��o\�	��1��E����F�����H�|Kt̀d_�N��=Xj��l�[�1sQ���������"��bp
��=j���;O�v�J��p�o�-�y*�s'`��R�Ӷ�fՅ�֎*)0g�w3�u���'
��_��{�m��ՠM=��Ȫ5��œ%����{>�lQ���]BŌ�@�E�lغ|��q�Pm������J�8�n��΂N3��V'�~��{��9�x��C�� ��5����[(�S�������`�u�ر��˴���x�>��N�W���hM��ܞ�F�q���0Vb�n.`�G�2���%6Xڅ���|N�	n�l���������<�Mv�V��nCf|�΍;��^��5�Ɏ%|��v�~I�g�u��q�g�����m�D���I��܍vԑ��(]_+�X��&Su�n-n<��h:�Ԑ��3�L�n_Z�P������m�倬ֲzU�!]��x� �[�L��v� �L��-ą&�
��Y9^��Z���<�z9���!��RoɁd%!�z	�����@[f�uFw�\��`�����̕���n;�׫� D�H�9w�t�]�h�%N!���g?�i0"$��K���I�����Q�ś#��W�*�n�6�]��u|9=��y#�S/�l���iFWM�þ���'z�$ɚ�9����B� W���	���߸��暇�B_}�<Ӄ�+a�e��U���j�hyw�6�8^CѯMNw�g6��A��>W�T�`���m�Ec ���nq�3û兪Tӻtg��������R\�i�^֩��ve�2E�y&��
���D�7U����I1��_tl�M��%��)N��N>�{�|=?#3��#��4j�_O��q�!9̓�+H����э�5�V���k7��5�J�k^�k˵^��H�Ǥ֔�O��ng�ѻ��s��O���	��PA���@��~� �������oܛ/��xC��G7����^�Q!N>Nrڸs4!���9$?��=�4uh���bMj��v�p����l�{����Lzt�\�cۘ3y�,�m< )A��<y�x��&��X���?i�2i;+b�r<�@A\�v���ִSN�������r%[�dh�izc)��\���C���XA|�BX��O�Bh�D�����|��6i���D��߾���.S��_%g�r�,C(�t����X�Jf���w��>���7!1�>�?����X����:��	+F��ƙ���G�H;+Wy��7m� 1�%��< ���y����U�:�C�k��uS/�a3�7�ľq/�i�|XN2Üa^�[��0փ8ε�ћ�h���;�\-l�o�Ĳ0*]X�p.]>�w�]n�{87��s�R~��^Rmd��ݾ*�������
����*P �}κU�b�n&O+4y>�����J����C�b���b9�V���Los-j?ttz��ѭz�/���g�aV�{����za���gO"�qڹ��6C��tB��Ni|kߪ��c�^�zC�4S���V��j��Vw�Ԁ��tw%_�@ɾw���c�J6ͭ���$�s�Rc;�^�}�e�
T�6��Ǎ�媷9��)�^(6I0dm\R���Ĥ[{���'ǎ�[����vH�Aivf8���4�J��e�Ei�&,"�(V�<J�r�Ɇ����$�����;a0ʭ���_Q���N ����%k5�#�đ ̏�z�6��	�5u��5 �TFc��=�ZE���� �vsN�^Emx��P�ΗϜ��Dwߡ����3b��/���\��p�6褑`�ANj�#�^�NA�M�ǝ�����;��5-�0������"M�{���Ȓ�ס&gN��{i�$�J<99��lG�Z�]��K��RhȢ졆��`�u��i�ߑ��=~�{5�e�l�&�Ϫ[���6V�j�#Os#���v�ۓ5��[��@F�������X��Z�n��K���~��s�?�zP�d�/S��k�r
�{���T�����'�0|i��	^90��a�[���Y`G�����q	w���-q.�Y6�����ު�#�8z�n��׎�Od�<iC��`�/�ݴ�I��u[̸��g��N%j`Z>���$�X�v�-��8��Zhbp ��`��5��Z�Ƥ�Xo�֫�!ñ��);�9[d�y!���̌x���pm7����'�NQ{��2�q0��Ĺ���_�ح$r?�5?���C���;�(�#~�/@�ܶ:P��W��6��NH����Ȍ��o�3/9_�i���䳏�O��1��,|`4|��p������l�+�]��d��hߵ}�@,�5���)K^���\���u@r%���l--�Z9�?]ǯE�Q��=<Q3]6��ԓ����fy%�]T�k��*<)4_����u�DY��`  �s�]dD��U�mŵ�&eN��e��"W0�v��� "i�}�~Z�1���f��4y�ΒojG�l��=V�U�Z�%�;v�m����<���9
����� _v8e?��:,T��9u6eәR�l�g
�%��3-K�X<�L?���N58�~?�>US��V�Q�~?���8�`�*��;������5K�V�P�"g�ȡ�� �iy�����L���-��FX��-V��_}�;�����!\�!�xC ����|�>w����$�:��;t�f
�[�t����q�t�3�Ou)b�n��/ �����󎦈�m�����WXz�@U���j���}���LEiY�#��W��H��)��/���-F�Zˮjo�y�ߙ�Z�w�q� ��|Q[��������9(�e���]��b�q�*�}<Q����4�b��Z�k���Ο���؟gP��YF�� �b�udѤ�0㍫ϓ�XJ�֩t�lEF��f�Kp�ϛ{��V=c���Q;ۉO��]��ר����V�q��}ĦS��n'�I3}Heś˪�֡tY�y'�n&v���U�P�۾����ŤG��	}�Ncvk�X����<sp5���Ug�(��M�m6��x�]6�V�vU�?�7"#YB�/�Rz��|w������
R*�4g��Z5{~��/
9������LF����93�R�M�8_�%8��C$�D��׮�ާ����K��5�$���c>�i�|#�/�'��csIU'�Ţ΀Vo���^�vm䊢���y�3�-��-�r��FS�nV]���uP�:h{+b>ݏlq�Q����UK��4�����!	���;/�A	Q]y�_���;�� `#�g�Bǜ�sw�i������v�����:��9�Q���\��o��p�,����p9~�o~�O����H?��W�z;�F��7�:��t�\IQ��>��~U�y`#5$�T�=�b�lM��~'�K�)4�(��g��:����p�)6H��O��.��a��Ekba���D��|��B���I�N�)�C�ӬO�?�F7&i4�S&��y�%�a�������ƵgO�F�l�*�/N���^M�-���S�U�)%��Bs�ڻx����e]|�aȟ�=Q�����T�}ZU��}���w��m� �%͂
YM�ލ�@T������ǐ��7= H���{.��Sy;����x�o$�b2���N���k����e��r&,�#�b����&Uy�������5,�Z	5�4��X	�`y�x.���6�b-v��O.��?A<'�>��օ�zs�w�^B��a(�;�MO�Ի��1�m�\�W�ɕ������g��\4V�-|AfkH��Q�����Tpio���K����$U�m���і1�#���L��)BI�o�'6;�i_ <�>��SԄ�
T%��]Տ��X��~�����r'c�8�n��V��l�$U�=�6�i���<�gҺ�w9ߑ+�L^c@b�a�	�����i��A�X�d���)�eJ�/ŕ�qt0��l��<M��;����=5������{ .��̎z����$w�{K�`O5|�"�j}MfR�ҟ(]�@���F��ūu��� �v6[PeB�U��tY.��;�V�����V���$.��5]M�KPa��9]dXbw���R�ǔ2Ӈ�Ճ��6mYJe?ܗP�y���E�T��gl��J6s���֤X
t)�@�FW�k���A�$��5s����C�5j�<<��^�-����.�~�r�z�&�Aȕ��;���Y���S�/��
����h	��b^�X3�2g�t���.�g��LS�y�`������x�6/ujnF^���$�\vê8�'ǅ�ɢJ^�1��7��P�v�́#���l��.z��ן�!�AD����>�>�,�@{��D'���ڙ\	���c>��dt��@��p�66I\������q�*�`{w2@TdD�R�أ3uf��ƚ0��i���7ڹ8gZ����tt�O�YyO�ω�*E@�9�WL�������i,�|��6��h��dsD��7�Ɵ�L/�e�#ʝ�!^:i�A�.�d'5��X���BQ�R��2�L-��\��g�z�XR��)�ŧ�=�D�����ù4 m�P����cy�ٺf���|J�� ~jhRl����S����,��uL��?'�VO����kw� ���t����,�xR���M�@�[/~4[�!�X��K��c�6�X6"]�!ˏ�\OH��={��"���w����` 0j7v������*G�������xD�,��`'}���`�Q˭m�{���}�JN�3lֲ�3����8��C�1Q8�6�;�&���.���5���8%�ٟ?��m�A���5��E�����?b5�e��S7��("�� �5v�?�&�j/�2�K{N2����3�PN3���Z,d��8����>���qFBo���RÀ|�`t2�$يT�E�Vҥ��/N�}K�A��'L�
\�I��5�Y9��gttK#�[ҨW5SqL��Jwz[��<+��ژ�����$K`�>ڙYӖ�?*]�5�w�
i��G�$��[��1����9���[uxr,�65`���yPy���'�����!,�Š�v0�Pv��Ĩ����i㲢���<*[��1�r���[�ׄ�/R��¦�b����)�?�zI;��e�Q����Mr��^��DRdW�j�&�h�����l��� uC�����wj���[ �^5� �.���1m�SR�K�;����A��rS�$�'�.]���ؙ_�'lVG�Z���^�� J3c#�B����t��H�Y�c&�,_sx¹�a�x�K�ey>^��y�x/x��"���I�����|q��7�U�5��3EK/':�~���Z�1�U�u��Wڳeo�o��� zxz��e>R����w���Y-�zC�Lipv��S(lL�:���8%l�ebQ�q�W薪EF[�=&5g�qU���<��eP���']�r-i�	�<�8���ܿ�@_��A��@#��xMo'�5�9�Ƀ䝖��b�V[�[�h��9ѻ��c�V����1p\��o�U��(;�W�1��ml�}G1�kA�'��$��.���'�p?�����	N&�`R�s�:J5��0�k^#� �3?�����t���6�n�w�_9_��ۂ�>�:���a@�+����{�
qݒ������2�E�F�'[�	MGx��p#[����̙�}n߃�.�ʒ�@m/ǎ��v���A�2Q�P�?P�W�ݱ�?-�\Q�>�s�a_ڥ�6���B�a�7�:�l~��g��0�f�g������n��{qU����ގ��GY��:��ۧ#*��%C��Z�t�=|�4d|������c�1$��f�ΝW�Ai�^CS�4�-�;��g���^��68� ��3f-�����
.G�E��?ɜ�^�~��j:wy�Q	��z%�_}�X�C�1�w}`ge�lj<��,`a�e�9D���:9mick�	E��tH�CWת�ʵ�+�����Sbe���|�k_��eL���$�p�|��v���Ej�>�d"�Ș���M���7�����3��!��X\���/��t�����M���w'���Xu٭���(n�����~�6>97�|MN>o�5�%�{,A͖�̘ ,�&���r�ꕾx���bl�<���9;�]h(|�=)��\Sx���R�i�m"��uQ�  ��?�낹��v��>lc�/� BD�V��u�ۀLC;��1�`Y����:N$y�2i�V�2Ĥ4��oY{�ڟ�@�F���ў�Z������W�XZɜ����2%��'@w�0䌷=��pe�1���4��"�G/\<��c3S�A��!�'��zl/M��^>��P�����S�T�В�ׇ�yYl���l���b(*�snW<٧Gtq��[��b)/�jW�~N�:�����~�o�N�l.�m�x���s���\�f�+���"��M,s�S��՞�{h$��@�͚;ۡ�؎	�Z����pc�ݭ'4�&A�$����P"��r��T����/�x�3����Հ�H��Ǜ�d�B�u����z�O��S��L�:3��#�֦1(�k
��5����4����G!�~��	��j��m7�DtG�x��q���VE^ԩيU�N)�o��ݞ�/���d�q�i bԩe���$��D���@Pr�E��fU^w߹�c�\M���-����X2�����e'��T�-�ױ�*� �l5��5왷�3r���OK�HR_,��R��L��e�k��J�mӳ�b�*k$PDY��B�(QJ� Ag��+�x0�﬚@�������z0S��M��i����'�ґ'����������E�$^!���Y��fd�+�!W�����S��pkJ$��ZZ@*0�h�в��ܲa3w�a�B�-)6(^��<�i�C-`;4{}�<0���������a�nȠ��'��??+��be9�P7�;,��~��{r��N+c_��?����:h���h�9�Ғ�$oX������ւ/gj��r�6��:������v�E��O׻1����ߛ�ɢӖ�:5c=%�0^9�y�i�u5�Y�k��(���Q8�Uu��w�-�N�2W�%,�
�a9"�N��p�}=�`>�U�(��4��B�yE�1DV��07ߙ ��hY��-�����P�U��R�����n��TO���[�?H୐���U�OC�?�l�;�}�=p���j���嶄������o��_�-���G�s�� N8���sǋk(���x�S���2��A1�1~�~��]ː��>����1��	W�=~h�@��ǻ�X�mV,�F��ZG�䤜�lO|�W ���0Hz����+���p��w��7��g!��0���3��6�S�ANpɽ�%�^�&�H2��0&�kL�� ���w|u��p�(�"*�sW��D���l*C��mRM�i�uڈg���s���&���л��
Z\]�,���(�&U�X�L�i�l�Ō�7�<�[�'������KŲ�A��]��F�J�]��F��}0h�@���rמ��Z��x����,e���|�|#]��
N/��I<2��۲X��r޽�7��`��HrLeièߗ���&ֈ==�dxN���2�X'A�/���z���x�5�D깙�9_O�;5[�H�Ɛ	㿚o���W'�iWn�V���2�Y�Vp�.�܃��	BPa>=o!�h-S�@���c����������t�8ѳ�Z�	��߽#��o�<��$�F`��������"sg���3�
2SK�o�|}LL+d�I�꯷�b9��ct�M	��1�0��}y�o���4_�<|4#���>��$8���U>�]I���P�1��5�_EwJ��������G��=/�ɶ�K&�����,�,ו��x���9�Q7�{=��ӳ�s"=�!����)\���*��*˖�I��ul��z߰���(�9��[Z�GlW��w���3:`-vBj�G9��+�5��O-r��S�Ob�O� �SV�x����i�{'50�! 	��,#t�-��޵���Y"�2�B��x����a�X]/�ȭWW��+g
�g�EdWE����D���kMu�8��B�	��F+-7n����$�+��O+���I:b�.�6��hWF�,���?���X�j��}��P�'E���Q�L���u�;��f@vgD�͸L����W,�V����(�M�H--h\,���q��BJk�[��]���ػ�S>�ٓ1�c��h9�� �����&[�Ljqf���	ͯkr���{bk)��~�. ���j.pg{>�yȥ�^݀�*m1~$��v�v�&Y��g'2l?���G�~�=�Aŗ,�E��,p�
�o��1��������c�F���j>��
�w�mk^)�v������7m/�ܾ�����O	1'y#� �����ȴB&[�g��n��kW��ҵ�N��@� ��:�b�*� ��7���݊�*��x��	.:��gq�֌���&jį���+�2/�;-�	ͪ�ypa��1'����y��P���Ŧ�=��8�/�M�Tq���%�AZ��N�-H�?� r&�
+����>N*�V��x���0�סl a!�|�b�Dҡ��>���h%�/����ʑA	9�l�o!~ �FM��&,���z���l��Y�"H��oб��M����a��|�����̽:��F���\���I�q��H����A�4�{^u.X�4�u?��?�sC0a�H�X�FĚ�ZW��V=�+�[�]�&�.���Db����>��gİ�)#�y��ڪ�:o8o��j�LdzI�i\V�RPC�gآ�j�����@X�-��9�f�k��K�H:�n#2�?�}�QoT�����	k�Z��l��o}t���DM>n�.3�ʪ��&�0���3B���' �F��=�oEJ��߅��p���vB_s���H��u�����>9�4d��ՙ�%���5� �v��'�K����XcfcI��^��I�-�i�S�&���:�ӢkCXԀ�/ۚ��<��;q������y_����7�W+�;3`�#�tx�)��@!H�ܜ�k�`�[����`nZ!�*�a�.(:��7���V�4�4*�!�gTU����;����)vR���~�,�<��o�N��Sc�.���7�8��IP�9��28.J�Z���
,��Jl��ɍ%���##�F��E?��7bŗ��_�+��מ�R<��;��Y�u�U�唷@���OtΠ;��z �G��u?��Z�r58H���x�"�� �xz�hw�aZ�̓�F�R���%k.O�W�W�F7��	��O����O�����:hF���+��MyHT}��q4��.��yP���4�I�3dZ�+m9��?�T�}4[�|��2�dG�7E��`����S-��L���bg�	�߭��� ��oW�U�Ϲ�)e)�a%U��<�XkC�u�f�[����a��I<s-"z��7�oTq�!m<��ך�o ��r���x�T��;K��	�kQg�!w�A,�6\}�� #��4� \dXD�8���
��U��WN6çkX�\��WVXIAf�͏FYL1�^����8�������2�J`@� �
ny�/�%i�-Qu��S�}�K[!������
����cB�!�p����M^�B�E�0�ޯ�C"ݶ��^+���S�_��cx���oj5���ZFA٢6{\.�h]��]�#��7��S����р�]F0}֒5f��[����6��>������%�(r:�[���鴕_=�o{��h~�Xh4��U��H��5�Φ�3uV$j�5��V�ez֟t���Vٗ��3������^����] �������q~��+�t��좵�R��y��.1����6�ZC(>��:�V4t,����n-����#F~��80
3��o.�L͠�@��ۼ�9gj�l�����@�G.p�ݫ Kl�O���Y�a�#ng{P�v�	������Z��Pwy�D�� �SeT�:����B5˩G:�ܫ�`�w%�lF =�^R���ά
�Pw��i(?�Q11	�n�����Dq���?�h����s��I���߃H�d�Lp����0ϯ�x�[K5=��i�RC=�(�t�m�Z����~�`��)m�?]
<��Qǝ��Op���!'�͵6}6�Q�z�i�i�:�(�-+�*6���>��M�V�TA���4���P�7��d(f�����'�#��mud4�vLn���T}�0��D�D�m����<�i�+��,�:!�|�Y,p0�ޓ��%�Ӄi��x=o��/z��)^=�YZ�`�p���;d?�4/g�ܼzY����w�8870.�Z���r��,c^x)D�����i�^�TDI(z1�H�k�@]�$�In��d�F�@=:	�Ap�����&�%.h"�jt|5��N�rpan��������E�c#Qw��HF�U[���a��`zH�����d�qnG�dzW�m�Y*7I�(��[� F�������y=s�	�wK��I�Wg駨 t(.}�p��"J��<�30e���c�G��˟ާ�VH+9�y�����8}�w��;�h+i��H:���ZZ�v��*����(���e]�{B\�B����RZO*|e#V�Oc3�!P��Sf^��c�g��a�\%�Yna����*����!I.t��I���r,R^�\S�6������͝����`�WKg�Zrml�ȦO����(���y���5���/6dh��4��c�J>ǖ��.W��޾o4PI��!��7P��+�lh"���b��,�S���P�6�gn��'A��&�"v��&~̄>Xi�=����SJ�7�9�ե�7���r7��X�$R#��5T����x�dN��#2����>9>W�5~�k�l���G��k���P�g0�[ɸv#��IYw7�w���˭� �Ȭf�I���U��5yJ�$�_>%^�=e�r<a�P6x�U��8w�������c��(k<�. u����xYf����O��[��+��e�&/m7q�����U�~fu��6�X 3�R����P�)o�>ţ��,a��*&��˝	F�G���F�}��ln��!�+�V����hgٗ��N*�B�X��H��Y��'����8��z�o9Vd68���%l��v<$D/,�[8��2��h���t0�$�GY4GXuD�sY�lȝ�;���7rQ�u1tpp�u��b��s�B����4�ץ)����Ӊ�q(4yߡVE�v�sk؟�O�<
�.�Oܷ��]�*EF$�Uk�^{�|:T��EZ�:�!���^��2���X|fZ��i������2M0K]�H�!���}�bC��iδ�´B���S��ι��<��(��5z�}������w�Ak���3��B�y,ѵ��Y��<�F��9i� %�P��W�PE+��&.)�m�_���E:��g��G`B�����>�A}��F�j������[_\����V�A7��@@)�WR���3X��i4�t��d��7�t�N�K�|�'Θ����_z1g
�J%�����{ޭn��1�y��7.���������8�7u�}Qd":��<3�Q^�a>B�����S@�Sc��Eb'��u��I���X
�W[���é�}�6#�#柼�Z�e'��[@�׸7�)	Gw�\TS��:_����¢+�bPؽ�δ�C���UL�/�C��7n-�hg�xb���n3���K1�s{ߏ��2EjJ`�x��p1�66��8��c��~\k��-���]ov��_J������c�$��G��z&�Yt�$F���^��D��a
��yV��3K06JW�B� ����A�[�5��o����)k���/���^$���J ��S��oW���ղ,(�gx|YH��^o�F�M��$c��#���9�^̳>�;��9�@ ��ӵ�F��)F����.��h��t|��YZ�2��IEo!d�� W!�L8��Ѧ2�T!�!4O�T��`	H�PN���Ƣ�r	��`�`��`�`86(����}o�;��~����kq�; ��}S��������A]��`�m����C�[�!��a��S��6mq�l1ώHa�H�������u@z��[�~�n���Ib�Fzn��V.�	ǒ�
����y+����wg-��-���%�V��)��2o�Δ������6ۘ{����7�\9e��U��jg�4{{�ډ�� _��A&��a����~��f��������7��L����h�j���]-��M+��Ȑy�O3,֯�~������ܟJt�2�^-���O�K�L�������OO,e�=n�z��nU�ޫ��U�!��97��l�]a�ٝ5���Ċ�vk���:�ОW��fs��Zst��hqm�I�
�y~Y�m�"��Z��s��̘�C�=���x�6�u�9�~~���i��X�\����"�|sw]�M`tK���Ru
������=���\C� ��oL�h&dCA�`i�e�]�/雸hp����K�<H���Q���|�ρsh�(�Ե��2E�;O,u�/}c��I��Ѹ�aG�;w��b
���z�T���CT2��)�a��MЉo�I�-e߮��E�#��;�n��xЄ����T����g�+z'���.WZ��V��n;"�#B��%hC$�@��W0��ʉ��<���"uB��#� �$����m237P�+2��KRH���s�j$�ܧ$��I��|���mCE�(�d���7;���'��t ]֔()����|4�W��Z��:���?����E�o�0�9���@b��'�jz��Rg�QTȟ�d���0��3!M�Dz_W/u�9ܦ;"�k>�55<t��9�{�f�5�8���=:��I�~C�'ͩ��[�lY]r,����%�pD�H�����C	��}�+=mRS2ܛ�Kn��H�L�%!q�ӱ�Pu'�G3���D`�l�K����c��є�v&��G��ۭ~<dK�#ɺw�sW�Jc�Щp����`
~��Ϭ�������e�[P=ciN$|������� �x2${�͑$��8���� ۓk�_Ʒ�x	�oe4��|�Ng�F��>Ԧ+,.���{�a?�9*���Ӛj�Ǆ�Y�y:A{�����L,�~a�v���]_l͵2᭝z����ݣ��ڦBm�hY�1�\��B�Ǣ�o��;"VJFOL�g���JG�\y�Љ�Z���''���@�^i�<Z��}��%2�n�T��G
YZ;d�XM5��<k�5����C?���{o���F��˹���!'�p>���q����S�PK�_����� �7�TyR��V_P��ƴ�P凧�g��KT�zu���`ߥZƸ�|�Љ$s�P/w7�HU
ሞ�_�S�?��ql[kC�uW|�4�ҰލbG��1��Hm� �7�gح��T��٠Z��}  ?���b]<��k�h�Ჳ?0�B��b�FCs�	g�jen��7�����cO�bi����z����0�M�M��N�3��Sw�j��#\[k�L�N^a}N��(�;a���9C�<d2����(6y����-�>�y�t��W��3~�k���V4J[aӃ��߀�H2�v4l���u��gˊġz��K��ۜE�D!�\ptP޶��VG��U���l�ڵ�'q1,��nL�ۢ隇�fo�A|��G'A�bg�T{���O-���K�aě�C<��qm�c ���1@�-�F���᫪|�?=��C\����e(�Ĵ(�H�{9|r��lU�>	#^�FYzer��M6w�z��H����e%rAz�Ǩ�|���=�n����mb��&��&xl:���/ޤa�fП����Bv�;�Ï<�%SР��*:>��XEF�Na��gE����v��6Ob��)G�W<GR+�_�dA:M��g��Ȼu*�s�`�J��^8���W1%`�nws��*�GCͪ���,���)ǜ���r��6e���d(��}��)�0����,+�$� >(�.\�&CH*�~�X�U��K��])�]_��j�L�\>���<Cð�[�*g�/�H4A�j���(nƠ��������ҩ����R��Y(J��~�zZ�M���q��W��-1QV'v3�lਸ਼M6Y~�a��Ζ��Զ�N�x�=J��hm�oY$����^_7�����9��/��X��TB[F��5��eZ��nb���ML��"*��p�L�'�SC���z�E�!��ʪ�&O�N0�"�)��@3�3�rٯ��
�np
���<�z�E[G;�5��BQ���a�-AA<;Z�����#�
�p��b\���Ol&k�� ���#�	#7~�3a���O$ũ�'�di���q(Z~�'z�ue&��`�p!nU,o��K�z�D _G0jw'��4���¬�G;�t�ߛN;K�؊�*�)�����q]�&q�{�J8�o>�T~k�X���SYˑ�?�X©�/��P��L�p6$2��p��U��"^R��v����c���-A�0��(�#�d�n.c�M���:�%���"��)8���L���.��!��b����V����w~j�O$���#��.��K���&|���qg�q�D��w�F'�1�ai�(�^^�"�D;������g1��GL��,{Z~�����Y�� ۪�O1�lT7KY�w��3�.cy���tV{�֫Ś������5}��Q�Q�Y?�?� ����EG�M�]�d
W*�1������2p����}
��k#�<u���GJ�h������qOM(R�N�Yi���5�vㆃ���}F��l�(�J�
 �?c`��������J<��~��_����{��T`�6�����HW��*~��^�3���{�+Z,y��މ�Y1��#y�g ��̸��%���P<}"�6�G�=��/��3L`L�&o_ȅ��Y_WtIB\�;��]ܝ���]w'���Cp���Ỽ[_�nm�j��>}��aFuG==�5��:Zm�ĢJC�bޘ�7�	�?i�r����LS����J��BR=D6҉�W|P���K��e����PRޟ�

p��m
M#6�|�am���i{Ɍ$�,�
_�Ow�uH��"��KywT�2�}��ou�����k��)HPh��^�g��:=�j���m�bI$᳿��G��	���[�ǅ�I<�1�g8�>�������(���#�ԛ�i� j�~����c�yO>��D֭�P����r���c8
=�t��R�������`[��0FSV���xq�0�L���PlV).%�������Y�s�W�������,��'M^>3�Nyn��UY�Q�4̯�EH)�Mo��vu���?�#}�x�vm}�P�|I�Be�)�7W��p���ϻhxz�Io�H]TL,��Ͷs0sg�N�q
�6r�3�TH�K���dd�5>�P��t�]���(^��_%�̸"����ÔSn�Uz��e�{	W��:���L�ùz�0�
��?����z�mR͗*-��/��C�E30�0��z��]t}D�̟n�O��5]��0��&s3j��L�G�)NAQ1vfHAI�]���}��ƣ�{c�Ʀ�	}T������"��ׇ� �e��d��r�Ԇ�G{v�E�O`f`+��E�B(2�� ����C�j5��C)/�8���b�ߛ��A��*6��[�{沈��z&���d1+C���bf��'��39�W������A�ĻM�Q��-1��~Y3a�bǝNV�(K_0,�L��1U6�F���1�dP�E�AM����8i����x<������I���N4<t��������3 �J����v:{��⟺nJ��9����]4b�4����ug�R��TB�a���B,�̾��a!c�[0��/�;�w�X~lL���!�-&I�+-ʦ�m{�c��a�k	�U�r0����,l���L �������Ƒ11d���.a%!�n�.O���C���i���??�E�����7vo� �i��u7O/���p$��P�z2�YEP ����^�{qEtd=�%�ℊF���B�(�2�ʄ���7J�(��"��x�Ԑ�s�6~��E6���HA�ќ�Ƌ�4���^��ػ}��u>����[�\%����)����������%���<x$�uR1Г��?tbJA��>�
�QQ���O�o/�V�םeL��3�[�2'�]�I�7��!�_�9�P�����_���؟�T�����e��\[3r''��5G��_O�� j�[,�t�(i�9����X=hp[�ӓgiiirq����𠤴ԓS�������U����]G�V���w�{*�;Ϯ�l8����waLXJV�z��΂nqD?(�Vbd`H�jF�Ӫ��e�P�r��P�����"FXr�#��s=Ξ��#O����'�+��6;�fm�&�ǉ���8�v<+N�cUb��Ԗ�JN��9j�|��u�0��t���9V���Xx���a�����פr�ry���M��:-]Pq��m&h�s�m������nڝs%��a�Y\<Y�������&�,P��u��ctc��w��wvT�aN��>�Ey��E�U���H_����w;�1�1�g*O�ߍ�&.�ҙb�Wƴi��������6��08a�
�5ļ��&�H�Q�p�P�៤���>�Wܐ1A��Uia,����H��f�J�ʍ�#yf��ūX[CŮ��	{�a�
?-)�7Z$�j���+R9���`���֢��fG4ȫ9_g����� �n�Ļ���;b�n�*�Ď]���ؤ����3Ӯ�|�ҳͫ��m��֋')�3�f��υp2H�~�se���|,%��������*�������x���$�0���������xw��$E���i_�.ɓ�G-��ͧd4�%W�D5k!f˛u���NC��?x���/����y�|Olg�n�m9*�$��'�Oo�T���j��R~�U1o���s���j�xU��h:�u���/�J�V��-����o��(�D܅�1&?���B�s-c�ֈ��.�4��+*���S�����/
Y���Mo,����8��D�����M����\�������lz��0ň���X���>#�IA��d��~Z6��<�|���#qZ:�k�V����c�\
{����E��E1$v�Tc�\x�U$fW"�*��F������fs�^��f$��fPj*�Zy�L �U��*I�b	/��41N�`<���>��n�8m)�]�[�p �j�s�˜����1����bj9T�s]oBq�6(!o�ɯ�⯕	ʩ2�[����.�������=|��N�d3��cc�G2lQ��ْ'K.�s��d�d+����?f0w��q\
� ������p�v�>[:_L��U$�,f�FIUQ������I$!��I��B":B�l�G��qib5	1I��2sH��R~��ߏ�����lVM�B���/��*x-U ��M2ӛ��ߖ�ݴW&4��V�����D;S�@��k����DɹK���mG֗�i�����-I���珞 1X$�ӆ����ͩ���"�
S9*H��9Y�م�s��N�jS�m]1�I�Y
h]�g��Sߤ�L�)�ە�jY9|1x�5xM̑��\��\���B_�ffgɸ?U���<����O��/BU_�,����M ��7��^�JV���Dtrv&B�%J�6-�֋F9��G����Jf}��t� �R��Y<�J��|�.#�(���Sd-��AJ *��W0�)��������Q��)6"�f�"c�{�hh��F�|���,*�4?;+�0��㪡L۾�-�? ���@�_��o��7�]×"�SX _�|G��CC�v��{=.�l2tS<�;;e2o�V �V�=�MWZYZ������?�e�<{��=@<���D�F��-Z-D��a9��H"]��	C)PX�$KL�"�w�[����+����\�>c���G)���<X<�Ņ<�j��_�t� ���ٙ�#qWk5�y�T'׭<�4.Jl�3��3��,q��>�r6�h�-���� g���9Hf��#�U��N���E�	2�{��i��j-Kʵ=�P$!6�G�Y*0j����.,a�B62FW(N'�:y� i�
������e���bh���Ͼ���_��9H��U��~XDld���lEp����e`��b�ˊ���jfn�?̆
��[��TF��^<���q6}�C�S��qB�e���H:�����M�Y!��շ��t(2"�M ��c����`���!G�>Ey=Jd��o���x&|.���)��E�	�|�Q�E�G{�&9�����a�kK�C�4�Y�I���WQ�(,,늷	ԸE(1P����f����|�]b�	�0<�Z�d�/rI`~���-[����a��3��	&��M0� �� �Bƀ�#R��$]Lx����d��H���ޘ0z,�jn�D�`�B"h�x����O�|��ۇ��'������H\?@���CF5�RY*�y9sr/ح��~�"���Z��g��J9�?�}_���"���"�ZpTsx%j��NI�b���L����@�_�U����-��PMڝ-f`�.3p�oc�m���Gut�O�w��T߯��U���Ǌ"F�ui�E���3�h�q�Ɵ��QfL8���.$����m���+P�K�)�^����.}G�v%&�"^�z�����OWW�Y�N(y���������2YJE^�h�&}I��9]⦆0����Y������{�&"���+c�`8����E7��o�h%�â��0f�S�z2N�I���!�M�cr�	����b�u0Sk~\��\#����i��u�1���S��������5�2	Pyh��"�
l\����������	�,}qmP�]���!��)Z�l;,{��Ʉ!<���q�L)�V����Yo\�7�Y%P^�����b��[����1���T41���.K����SI����!�%b7�f�T퍃M6�H���g�dت�Qi��w=�k�e-��l�x��ǃ7q7/|d���9Q
Ʀ��r�[���:~�Q5���U�>���}<kڸ�/s�;\�1ℏ��L}�y�	���T������W�G�]w���e��ȭ�K�]�qE� �aZT�/�rx԰v���3�E��x�iS��G֧��)�&J�l���Җ�NX¦[�[ �ܝV��ZWc�g6CO��� b SIv����sO�H��;5�@Rg#h��%�Z���C$��(t|�|Fס�)�JGk��;���Θ�.1͛������I�z�˲ܿ��*�"N��6f0����Eƣ�ƍ�'^N�ư�I���-�ց0�}q�`�]� �t�l���X�P �/��j���.�'jv��HW��z�$9�؝���Nh��J���5Rq�?r =��SN ����S�!m���`r�i�]������U��aZ�)#� M����⯢�Ә5E��(���,��h��Qզ�|O;#{mX��8�(��w;sq���`�����bqK�TSz��a���5�*���{1B�����/�̪+P(�T���jz����s��7.'&�,!�Pۗ/�Z�\�|g��f\�	`�%�Y�F��Y\2��{��X�nN=��z0{��Q�7�($鿂���dH�'���T�K7��C�ߏ�s���Ct��=��OD�~�	����_��j��������=|d��#�	G�)��E��x�c�Sb�v:ٻ� �<��V�e.��I1�D)�s��0��_���쑐\p94�"҃{wH��f@�|||9��s"�Mv��&^�=��U+��ʨ�'��� j�N�쑉Y��Hd��Uy/1����Н��nF��@�*!�6ҝ�o,s�%��h�9G�(�-q^��ɑQÉMT�:8�4�,9'�Q<����`�35���s0�B쪲��6��&o�'��6��k��I����%�����oUk�#������S$�t;_��0�Tp���AO�+\Z &dV���[a����s�:� �8a�2^�j�ZD��'��3�;Rf�S��#j�>}���&��Z$M�X��a`�\=��/uWZ��Vԧ\O�d����C;�1f�����P�^���~[���˰hF�`ԭLv��X:�{UBl�L�CT����("�/�Z��5]Q>�򹐯��#��ea0��-c!�F��	0Dᗅ��a���Y#|��f0�$�ԍ0�^>����N�S[�r����y���s�:�2�/V`��ս՗�=�@%)�]`n{�ܛU)�co9�R�y�_ 04oޏA��7�k��W5��u$a�����\+�"����7��@��3i��6NcD\R���t�F�m-UU��!5]���7��]�%|�!�cD��.�����1C9$�w�/�!e@Ƨ�Ţ�Y���������fK������9S�HWF	9�hx�x,��=@�����y���j���_���*����@��dF�@M���ءYD&G�2���Ԟ���s���jN/e�E�F��i�Ȓ�����Q^3z�`;���G�a�.T�w]T��<�}�i�j�7m���+�KG<Ycvj�~'\F݌�.'�P�������`��~�=�H�sB����wj�ێ����=��P�^�p�*O�Cm*�G�*�ѿ𹼮��i��>�񯛧�� ]�9}���@����H��.�l������dt��ìn�:&��4�#�F=��ߣ��aM��������zC8')�B���Y�x�?�ȸ�`�����kxr�����a 4ʱ�Ī�K���-����R8���\)"���G�p�L�Znրx'�8y��Qn3!�
���J譃xS-��eZh����wP�t��R�9S,�K��5:�B�۠�j��b{b�V�(�jy��:�lfgw|4 �-���Z�
*��|��|�{�|�>�=1X�Ѭ�B�����y*
gk J s�|R_3&c����?�������J)�	K�Z5��Fq^�y��:����o�
��y���E�,��;�x��uB/`���A_�\(�B�u�zk,��D3�*��rSJk�NȠV�_SJ�?/��-�A�00��h�Yn����i�J���RB��8���H�Mw���A�v�{�8�z�_��!N8Ѽ������9�E����UE�4������(,�J���@]��+���\����e���D���r�fW��t��:�uҺǛ!��Cyx\����uN�	��q���0��H�o���=�nIS��>4��R�>n�����/v���W�Yl/x:փ�|C,m�ѣ�)U �ȃZ"ρ���ٯ��o_�8�oIeWO�����*8���b���	y(�S���/\��0��L'	e�*�v����cA���=��6 z�2��#�πszrl��G���a��GX�%d0����� �&!�h��X������"m��;<�I#� ������Մ��XG��겳U�<�������*�C�#��]�{a���)3�qq�rU*������1��t����d�~ޘR�a���� XR��[t:V����"�!�%ҋ�0>[��4������n���\b1�;t�]OMřҏ��1�s;L*��[���G��JM,qgZz��B�j���pK���I;�g���^^i_�|�t���w6¨5��� ��o~_PEH�i��/կG��^�\�L֕���Ү<�a ����K����]���c������B�/Ƚ��z��^r�r�
��G: �5�{=qvvfLq�,��Q`m1ӫ�l��򲩻X~����&[���̟\[����0Kes{�I�6�&�[���?����WQ����#�	��&Ć�?�;3�㴹&��&ԕ��'���#O���lbS8rN*y�~<�m�IE��� ��[���b%~�A�
��j{�QH�=���	�m�t�Fu�Ӑ�ɬ���4����G"	��/]�vg''"�B`�,Q蓿��j��|E�pM�ϋG]}=Q����/}Ro�K�C%)a��w�P9AAj��(����"2�]��9����˜�ɏ['�h飻L��F��[a0��+j��p���>�w���G�)��!�o�Y�1I�Z"R��ґ�D,B���H獥��U)�i�u��NXtDn̘���Z2��|@Rorp2������UT�T`��n��bЫ�Py4W������hN0:��;�����?���k~�M�2�7�?���BP#��ri��O�4�`�O�
���s�7���;�5:2m�w/�2:DƊᐹ��Y���3�΀�hb��۰�_�!t�U�_�3r �er6]ڰ�3�Wm����+�ե��Q8���X�?�t&��r�!�����*3����<�O�L����p��5���������~F�@Eȭ�����G������f@��Wo~��#8�{�l�u� &	�d̻7*;eح�]�ԭ�d��ޭ�e�&���3R`M�9Xλ����Τ"�}#�w��j�h-��9QB�GỜAO��$qL�7'��zfhe����2�n<��o��Y�Q�mf�ڟox�wC�]�cV[�R[-T}8`w�K`����%"y}�G
$7��R�;���x)!Х��Wb�B���%��P7�6ˈ�ĥ��
͢�v;^\JXOb�Je8�snf�w$z��{fa�q��p#b���ø"�M�Y�廎-��-��7���mQ��/������J)|���z�>V>dx��1�+��L��^�=7���7_��6P)�t]s��=�wM�()I6�.f���7A���戩���2��0��U8�)�N��)�����(f�,G*���ƀ�����*M�&&�u f��؛���Bpm�N
��ahd���)��頻ž���k0��=���+x2����}��d��54�b�������b���&.�ȯ�#oo>`K�55��$�nF=<<~�H���}M�>_���c�~���Mȥ�����0)����������� ?5�!����7|j� ͆;R�5�~���0����'�<G��чF����o��]�9�D�Q&c����%z����DѲ��
@Ǽ}�1��V���/#^o�{�f��EQ���������<�)����1�tt��Wpt~v�1ԛ¸�V��;���PX�2���
�CkG�?�E�
�"�[Τ{.`|�*+��:�C����x	8߿F%>cڡ)謡����I�S�7D�I���ә������x3`�������wI.ՏqE%aW+g���=�v��u<��a�>�8]���3R/����u��|s�p�х�lBe�L�m�@F1ۋn�}���r�E[L� S;g�A!6rR�o��~j��M�}��KWq��5���	���B��<�(S�X��5h1V�l�).;��Q�htk�(ߢ�|��<ҡye�Z`��n���{f~>��ZaX�r�C����j��C����5�,BM/\qu6VV,�M���F�i"��---��_��
�6tG>;[��Y���Q���i�r��a�0�o.jo}�w�e�J�$��Q.� ���j��0�Q�}T2�,� �ō�8�Lq������!ީ���*s�vC�K#����*
/� �����+����d��OF��X�L�,��V��bOOa��TRb��T 4X&�Z�|E3[����j������$�����_��h�6uT��L�m�R��X�A�];�c{���Y���������h��r��ˎ��Ԉ"o�JK�c�Q<�zWD�#�:�$Ɉ�z�A�F������[r����s!ؖ	:"�*FA�;��y9�zX9�����~��;�}b�Vɴ@/$3��`A���D�3/9}���ĭ�Ƴ�r�o�߫�N=dt�G�,k:o�d1�\��u��]^l��kj.z�1`��<���W�ñ�KX?��/&�n=d��W�j�c3���S���c�/bN,ǻ�1�S�0��y5*׈/�a�.�ޓ��ÄED#f/|?ځ�i]�%�*%�6�;)�tW!l���*��n72�<c��:�����=�`�����������ם_�)q��)�%��n'�a]
���3a`����3���.��gs��:f�X߄���O���q�3,I2��BԞ��@2(���Y�7&�\�W��+�a��Ic���j���d��d��>���O%�������PSZ�����u��f'�g��Z�̡������5ۀ��b��I�k�+��+僲J����~vB��`�e��aEU�A>To���љ�Q�{{�8��_S�� ��8��������Y.w����k��	|5�/�8��Uh�A�*�/�7f��B�)��Y�:(Rm���!��q9�[*/wά~p�zJ�^�/����Λ+3��oKa�JO�|ƹ6u'�>���rri�!��z��UkX_С���0�W��ī��)8�Ѣ`�,a-�O`�>7[�D2&�+N{��o(�s5�Bʁ^a�@JUt��"#yfv-Q��a�������?�g�J )�1f��*���-`K��kmm=�I4bv��-��2����f��r�a�]�MD�����H���~{M�ѫ[צO�Y��`�*�~��r�;.D\�TN�ʢo��Q�_�q��M)w���KD��.��yR�ꍹL�"�W��$t� �N\��~?Eҕ���cv�Q��F��;��_��M!�����1@����8�"6�ZuZ����B4_���RB��'0�+���	^jԿ���<:+u;	��?��\��>��"'���0�=xr�@�<Y5����?��1�C׎CvI�$`\�ݎ�} f��Q�M�dO�o�)q��࿛�d^�a2+�A�a�P���@קL�4llnD��h�2�0�KC�DF��b쒶��p�*�[�����5��u��զY=�Z�g���PB/e_���������}�������S���͏$G���1�gb%��츇GGQ�z;1+����G��*y��}�
�BNXA�k�ˎeAA_�� �\��A'n@ݜ��\��s�o�B��|9�ݤ٫Gs��+JX�N�_/M����z}@��:��R�����H ��l�\F)��e��G�w�Pp��2�ԁq�~��VM�<��_��9�+A�O�(��#־�2�"<��h��f���@jMzs�I.�d�#��ɚ"M�1�zI�!K��{�p�r�����Z���SL���.�'m.[3���|$)��)�M��ߎG1�Ǆ>�D:�7 ����y/�ѣn����x��\��h�X����� v~�=��EƇ""���q}��W~���Hy9���H�O$�w��
��x:d|EM��B
��-\����g����!��\�v��.'t�� 5a���+X�A�C��/)c�д��o�z�]�@^��&��uq?5�),��膠ܧ���eF�lmMǈ9�YD�@T�}�쏾�6����T6�8�-�Ք�~�W__@.��t�q��T�]]\���������3����;s[՜H_�	½�[^R�XE�(r&�<�zO�=�o�P���G0́��l��9���|��-eE��OQi�9}��0@����;�r3}��S��CEҾ� �z�]�d�@7�$�vol��³�]Ivoq�Wk#�&�#�'��nOQK�m;��V��l��k��i��=ⴱ/�Iֈൌ�o�_�=��H�)i�Ÿ]�Y���q.�`���U+�6ա��
��]˚��ڪPNW�=*�xw�UN�ܾJͿ9�q0_f��� @��r%T+QQ��0��b��фӋ>�o�}�����_)��P�����H�ҿ������B�
�|߷M�����_�dP�z�
����{�ȹ/�Q��&����ť����2��v6D��|f�`D�xq���|���F�iň�1��g'v���vs����( wn#�3�Vp���J3� ���-�nl}�syE���� �.�qh\�ӧjA��߭[��!���aSs��d�����������X��LT�9,�Su���r#d�E�uI^[���__n06�~�d~��a�N;Ne�%����Hp��e�s��Q�*�H���s.��BfH&��q���z����k+L��TD:we��#����Iw�L���cp�R)�3 2_��lW�	�`�=J��>��N�ؽfPj D�W�=8q�d�saՋ��~<�@��l�u`�W@�o�IF�Ku����69=17a�;�5!����G7}K�QC颷�J�n��!D4Wr�Z������V2�kn��F[Kf���tU|Eb$s��\�5�W<r%�c����R�e}rm�r�\P ����Q2�'g�ܑ�m#j�^ST�va��5n2� ![�Z�{��c��2��(·/1<�2�gvγ-��/h�?�����E�#Rk�y,-o��ߴ��{'��ATA
˚�6��xǬa� ���m��k�"}!�RO�#��8��**d���Q��)��CE*��b �\��'x����4����0|�>��@O�I �=�1�4B=�V1���f�����S��S���o����W�ﭳ��
6R'�2pp��w�3�cy3��]u4PˡBW�l�p�oj�"6Ak��yx�D����0�َ�]����N���)�ՑK6��,Y�s�x�9*�*"��dv0L��WGv��p3F\I��!�00�bo�S̨�H�Ys,��'*��n��ⶺ_l}iU���S��T�ѳ��U5�/��f)p�K�nz�̊��|�݇�A/�w|�k�>'lu�|0�ޮz�J��⦭��;�F�<t�V홈d0�W֨�cC/�h�MBc�8vV F4xs�;G�Y]��C�|��]v<d+�z��&�U���4��k�ğFR,ˑ�Y۟��R��l����J���tU�����֊p��g��ZWD��9�}�U ZV���}�o�X��K䭼[�ۤ�U�"�q{ڶ�$�g����<^�a%��acc��l����_ss����4|#��q��f6?<Q*�����\�P���uj#v�u����F�
 ���p���M��Nx�fQ���֢}Iێ�[l!-�yRM�^I�1��6~�÷�����:r|1g���#�@�����S.l��oKd?���o���\����'�s�UӨG���\f��z�C���y0�-�7�	g3��L�#���D`�����O�=��6�sp���ѰM�;��и3b��*�� �e���Y;K�s�@��5���>�xr�\�t��@���3��YT�vC�+���ycN�~艷~7�b���{h:4}���!#�о�+)5׶F����I��E�>�d�����f�?|�]%.�����Do�8� l!����bk~�b�����"������W%��٦e۴0��0����?��,ȉ{F�<,����4ep�7�v�#���_�־�Aw��%�����Ӈ�a����S���k�yE>������PV�z���~b�J�9"�0՛�3���A"
:��&ᆧ�'t�1�l�]$\?���r������A����t-{}CR����R��I�>���wi@�3A㢤�V��{r风�WC���`\魍��t�����DF�ǒ�-������W��B��G+�S����h�c-�Z1���_U����
��C�ۤ�Y���=T� ցy���|f�Ғ�2k>�Z�|��i�c��Y3��g]��r=;׾�[u9�����.N`�z�G�Zk�S��� lw��i*RU��qA��G��:�O~/n����%�^���ƞ��ڡ%9���l��6�o�2�L�Ѱ Y(��a��Ѵ�7[kͳ9��/!gV�eY�0�ٔ�=�0���}�<�ph�lj�X�ĥV�U��FG��$DC��4��LXD�9���gu �hG�#6X�Y� ��J�XFU�]�ћ	$��W�W�&�f�3�������9bn��X@�Fq!"��~.���]�V�%ok��n�ms����ѯ�,�z=�[4�[Cx*6�]�=�)�6^Kt�r�չ�#���c��ԉ��y|V�o���T&�������v��W�K3EI���1<��' ��z	��-Fa]�|�C�
mJ	v���)/.�r�?���s�  �Y�G�Wg�����M��xo{0��N�|��^Uj��s�g�ֶ���ΥO�����[�	��~��d�ՔCg`ϯ�((+^T�4�����s+��`��l�o��,��D�F�X;�>w�S�n������;:�pS�������w�<r|1�K{/�yB �Im�4�.����&��t�VR��d;��"��-�r�o�5��T�SW�h;���[{�*��f���%ϭJ͂{�y?3���D޻��Q�L9�]��Lj�j���
��D�U���5VR����
�SceMGy���mot�W��k��a�DD�����5v)��ظ��3��Ԅk*7/%���S�b���2�F��;� h(�c�F#g}�vk3T0�5�x�TW���<���~~{�of��IԸ}'�{�Ɖ,]n�K���.�\��`�*�8�-~)�,~î̖�s�%iR홐�d�ֆ�nU*�Bo��s��^^X����-F̂<��d��U��D����5�]N4��k��u��3ckl=�WM��L�{S$i�f���+ɟ~��z=��Ĥ��Hb)��"���Y�|	��Ra.)�;�iXt�MÞϜp��N�#��p�y�l I��9j�7�O*�`i/h]�k��a�p"ᙰ� kh��6�sW�Ъ���v��FΛׅ��l�$~.�P�hIKh���R�E��x�ɞdiy�j�Տӛ ��ezυ�����^nج����g�Nrֵ�&�+Ja�J�9ܿ�#�s�����n`��`��l�+DJ�1P7%�������ZTGȈ�����m�}ƸײB���( ���@+F=]�b}�g���o������ѤI��0���k|����
�O�]���hn�J��3O��Y�^M!Χg=���e�@q3���[�KKKU��M�����_(����&N��g�h.�*�����(Djw��6�1X�Ԅg�dFXi�Y�0u4x
�e
���XV\���u�S��H��'C*�w,��/V����n�Ɲ�ݮ@��Ùt���s�o,�Q��2��鼆��w_lR�2́��3"N�󬽏�|���wpnS�]b;S[}FI�u_l����+¦��qW��Q�A�6�=�����%?���0��Iu7.a���+V��X�ɧ+K�����q�� �F�g I\)�<�u�����a7����X��ij�ځˡ�W�1~����OR������G�O>z�FJ]�S�f�=�q$�:���#�Hm7;H���(��D!0B���.�����E��
��f��v}����x7��v��:��S�gCymB��"	K�T���S�+������5���2�^A~Y����+�v����NdKB�S�K����M�6�V:�tŹ��jM%�4��Bv~��X�
�tn>�Sg�����Z����+Jxsܼ�ȤA?(��(E���(�Z�ZR��0���b��v�|�P���E#����wF\uY>b8^��ę�OT��_ۋ�ςv��.@\h� /��m�W%�\߯J�.LjJ-l�~��Sa�go���g��K�O���<��`�Y�0F��/ۈ,],Y�tõ.jF|�Ӓ��=Mot+�W�����כ�h�1d1U�f��L��,]����	����u�1E�������Ӟ�yq�A�\�;#�p=�fo��r*��ڟ>Bx���)��[�;�7�~.�l���T�5�o=:�V��r���,����A\�Lg�W��r�y��U��e��[�4@[12�fU�s/o���Y����U]��	^�S$\�^`gzL�&�vLO��7�9h���^VFM�{��}!xV/�`�q��}����tg#�Sc��e}>��Ĉ����NU��Ej�K&��W��nb��M����!�A�8����_?�P�;U���;��!|�P���u��,�G�p����(U�e���!��q�/��Ө�YWǈ�
�2Fe���Z���Ԧg�sg������l�����%��h>W�D�~����R�Ek��-CM����_�|Cf������3|�>��l����en/X����k�t����ω�,�&՛��]Wrl��iBsu�jN\��7�@�l7: �1$J��6���F�ȵ �M�l�ډK)L��ik�0����u�NK��aa�\R�M�(��C�id���[}�a������b4�4i-�c٭W�$z���6���}�
Xk������l�Ѭ��a�8W"����;b��c�imB�6�6��g��T�������:�M��Ʊ:�a�PemU4��6�e��
RO���%�kK�����i�/|
�CT�1��[����,�u��z�H�:R�˫�Ƿ�/�(�,g �p�PME3O�n�� ]�?��r�V���3�1������ñ6��K�	/�r�(�*v6=�VI�`��LRo�rņmӶ���8K)QD�����#�
�G4+͌}V�\pr�aBl4�[�X>f���0p��c��T�eM'��:���>N�>&�פA;������q�и�����JCR�q�};��4�CK`�ORF,����s{��Mά_3�
|HpJ�����.�hDx%ª�SN~#8�_9�}=e�ұ��͚�!s�;��U��Ud��ﵑ=����߇�)�jAM�],'B���m깛.57rkط����J�7��S΋��|}#��h��m��������3��BܯG�	M/��t:ɇ��lĢ��AJFh�`��j�׬�حwnf*U��>�Z_g`eo'���k�{��N��0��'�qoWIY�J�3ZLwZd���f$�T��Ĺk���L����rp���{�H�\P<;��uؚ���ʒ~w��=����΋Vd>f�d�"׳�1n�ᬻ������ܘ���<(�U�M������7Z�t�Zl����il��?o�e���Gl؀i=89H+��$�iE���Pi+�D)�+S'pk$����-�e��G�y�I����D�!H~4o%�f�f��'��{(\7}H7���IlNz�B:s�ut��JU6��~�܃�x�E�w-�������C���w�+���N�%V��I��X�wIM�	8"d��;R�9?fy�+,R���l[�-e��<�{�[�'w����w"�d|h-����t�ч�I��F�q�,�NO(��VE5ɦV����5�eW��0t�7&��.~��u(�kA ?�/yƪ�>
���m�Qa����I-A�ь�Tf��㍑��l_-�V�deN�Ѿ�u�S���RD�&A�^�V���V�9��#u�j/iS�~X���*�W�q�j��/����%N|�Q|�$f�5��D���VL~�<�ǜ�t����h��^��]��H�ӈ����jRj�R/ˡ�jSm;�m/���I*O��E=T(�CF(Owg��g�wH�#�ۿ�c��Q��ˤ���WS$X���Ow��E��`���g��u�Qm�A���������)nJqww-Vܭ��;��Kp��P��o��G�
{������O�R�&|7}�2�头'fC�Vp�Ο���?r�E�cI�j:.$���L�u=�R��Y1�2��7"g�o`#�X�.���@�&��ZKL�gp+��u��!q2�j��8f��4���RN:��#��'���w.�^jq��9Sdq�� MD�`C��z%~
�ҕ�	;��]�$(R&v�
%���T!G����f�Ǝ�����t-�"P�����p�]
[Zp˔��M��L�28~�tHE�@�-�L�]�G���f%}�������ԁ[��1�9�����1� .e_y~�z���ړ�
	�c�,èk������:�ǻ�.!�^oO�Ρ����W���*�'�Gd.ѽ�y㠷�Κ`� U��Z%�_V�;}u��	$i���OB2\&�ݬL��}ҝd�}���g=E7i��!��%�JJJ�'(�|[þ���'�����t�'���} �A���H��e�&������i�{O�﷼��'��ُ[��\�D���Y�9T�+Õ�ov�W����.b�|��&�{�G�<Ǟo�n��7#s�:�=�'�)ڳm���X�9�	.�[�������2���1P(�u�,�er;D�%���d!�@�Z7f)@[�����U������oٕ[�I=��P�>�Oq��w�W�2����)�R��lE~���)o�
4!�ȯ̸K������`8s^��n������>|��6���S�B��d�GU��c!l�f[�Y,ZC4�"�z�G�-��W�����q��z�q���v@qy"���1�n��&N`2i�u�ז��������4~�X�zc�?�\ÄoM�k��Y�c�^�os	6-%��V#�Z���.�L/ò.�����l���M�ex��^�^Y��F/�J�m���0�XZ6��>�(��W[�+���o������ݯ`��b�V߽{f���/h(]Cg�����b١�;q�ۮ�����q�S�VW!q�Ь�?nR(5�A+�4g�=��������@�C���[|zn̥�VW���s�e���Yo�$^���x���Y����p�,�T��շ�r�XvCX���p�64�M�ω��߲�vCE���6�9���=�tq�μ��A�a����]�
7���s��Co�a���"/"�����
G�ǥ����t����ߤ"ZJ�)5,u����}��k/<�ߙ\��8q<L�9�X8'�|�e����*�+����iB�3OO�����)�C�\�ާ����,.��O�bJ�;1�A���Eo��5Cڋk���T�an..I��� ۹�����F��ƫ	Z�����#R��)�J��Y�7p��/��r�ܯ�������BGu�, !��s5���!Lo� ���^s����G�5����aQj��?'���"J�����J��.<�I������=����lNp&h_�����z�TִT���D�����	7;��|��cp�F�:�2��г��@�wĀ�y~K�V�zp�w���c�3d��
���C��л=�UH�P%�;��H����u�ƕ�?�}:��:�{5 ��"�`��`��R-��ux����ul�O?����Q��}�� �:��
�T[��i+!��E6VyӦ�L1x��j��V;�����y�
b���v�9���0�uNp�dd �ԛ�uDw7V����m��w�&o�m9�h^����'�2�F�4Wm����dc�ҏ��]r;����.s~Z��&�tM�7� �8�o���_=�O��c����+U5�|��Qe��L�Ŧ����CRx����?��EHUZ�D�$&��㱾��&SC����?�_����{H�0S�/���M��î��t(t�&��-n�$��dG��T��X 8)�Ѕ��u��6�3�	�W�3��'�X#!rh�|�鰜�KaH�'q�yky�w���*�H&���9���y�p����&^��=��EG/�|�1TW?|�\�ɔ����	��7q8}k��+��q7ywT6�����	�Q\t�zܛD�#�|G��T�#F��Z����λg�.�lgB7+�D�o��&ɪ����b��
_�P!���b)P�1)�Q���r`~���z�~V���9�����������˛�sT}"���h}~��C��2��̏�mv8�����)�/b��KQs��ϑv�"��~ޣ/�!��$��3�������
��6ԁe�a�VڅZ׆��i����#+�Fٓ���}����Q�	���_��'I�PTYʪ���r�' T]�?�+���<J�d�?�
R�38I��D�	�q+I}B�ga��S+�bF��6g�*sYK�n��5\��f���\�^�Ψ-��V��GJ^�]�Y'�LM2�5�|�w��[�Xh5���?���!�p�]j���Q�F�^Ls�r�Z���`��,{�h�A<YB���ܭo����%q�K翯��jP��z;|-EZ���2���HH�~+6R��8���Ŭ6k%�M��oq��b쥋j3Av8��Z��F��b���� Sv�[Z܈�eI��!�l�ޗNC�o�[�g�>�h��f�����7 	੃uw�8�	҄�����ߪ�����N��zʼoL[��;v=���c���VȢbOj��;�Sۘ�<{������yo_�+
�b��۞�o�>�&.�,*9q}���f���ª&!"˃О��N׺���N.Ҕ6[@dqu�=ۙ�1	�Ā�
��u����|t�s��}��'����9�� ͟սU�$�ჩ�mր��5?���ڧ_ć�L5?����_�Y�6�dD�́2�� ��X���h酴f�Uf�'��M뇪���ŏ+����,X�|v��K�V/}�q�@!���Hv������L莬ہy�hU���!ف=8R]u�1�W3��N�̈́6�|%��<�M��]U!&�R|��9����}�(�!C�y���w�|�CwOJ�g�˄�R{��<̴��k6{{��A��{y#���Av,�cc��aiDi��@�����64#x��P���ğ �v���3�����O���?z$=~W����p���Y��^V���H'/�T��ڴK���`��`���I�����3���AI�������I2���`���׉�M�i9��K�]���l��%���\��B��h;�:���b��|��M�pͯ�ؘ���m<�[�%=Y���H�T�>����Oּ�҆v3�_Pּ�D��L6���`q�N3`����j��L�}�`�c����"�vK�S���C��ڦ�PY�o^L�*E�ҽ�)����.&�m��6�u�9�N����E��YP	��e#�\�<7{���.X�:�íH��FW﷭*~J�C�����5��^�|�
7�ԛ� �X�"�����f{����O�<���@����H��A�v ����*�m=F�FW��O�E�=�Z�ֹ�v eeO]���?��k`P�7��|+6}�!��D���x��g1DL^v�{S�\�g*�bSV\��
qs)�T��*V�렻�(���cO[����쪌�08XZ�D���x�����c*��@�3]۸�"�7yi�"��A��<̌��[������q��-� ����6�*�O�%slx���A�C��`��(������xE�h ��=�G�2�^�6">6�l��]E?���uO��E����"�ߌw^�1�ߕl�
�\�,�L�#-�'v!5z���pzf�ח�E_/��0��J��,�|�Z?^�t����������ׂ����5�䵕H xj ����th^�d"``�����i���.~�r9�ςpY��B,�ӱo�c������B,hG����*���ׇn����#�鯉̛�щ��u�#U£�ƺ�c\E�e���6'�<�8�[�˄���Gg��-���K�����-�_�d�,���+\> �Ev��=Χ$�dW���i��������M��kӣ�U�/8�.�%��^{����f�|���H��
Ӎ�����nd��87���}�F1���q~C\aKB�5����l?�cf������#N��i}�'�A�|���M�g]/TG���n]�;+�c��c��*��|*���qJ���v�Ղ�������&���:�J��DL5>���&�q6�mc
te��
�$�ێU�WwK�ɣ>�x�r���L�T��K|w5c��$�#!f�]GvyB!P>�l����C����L�l���#��spr1Z�nu;���w�u%�I���J��ޚ��&z1z��c��١i=�ր��~� �����1q��J�b��}����EBeԎ7��(r�k����*���K���Dm��w��c�^�]��N@Ε���7ZJ���RL��.ُ�Ǎ�I�;�H>TWY�'��6�D,0=��;YQ���;w�E0���W�X�:�.u�Qm�Oʙ����w�6~'��[���{\����#	s8܌�d���dj�,=�7J�.?l���=�$Til}2%���PO!G��p�Y���_�*+�V��=�����G���B�]3��3EH�E�h)td�����<�ߌ<{��][�m]��F��
��3�h����
������P����O/(@�2���]�۶�t��J."��Y�~�:ѮnÖ{�z�Y��������Kx:0y�k�?X�-���m;��bɌ��p�nQUU�Ѫ�ꖼ�pD�}L��w�t�~X���vr�A\���dRbzE_V�2�/��i�=�d1��g�cg��h�Gɔ^��#�:&r]_y��#���j�zlN?Vx<����D_�ƴ�0�'���t��w�A�5A`�
�[��x���Y��f�v	��HSN&��sO䊎䐲Y#���jkY�Cť(1l�۾bq����k��NRvK�ʯ�c�M�*n�R���H��[
��=� �ۉ�	b�',c��鋌tU�~����H��������6y����NG���j��A�������]�1-�@�Z�5��@����ZnE$EB�wlK�G���{)θk��t����=��h8�NpAB��q���������Z�w�BSL#"�py�0Oy7��e��nW5ZN����Dӝ�t�Ճ�H����{u�-�'�l��	�t\�V�&�H��t�!� J�5�ًR��M�L|���U3H�E��t�e��GJPt?n�)�a���P�z�9�Ӊz���~X���*����tg�@&�D�h~X���L#��^ݸY�Cb�'rȈj����x�}���͑W��Ƿ�-ST��EPY���5��^����4���P�a�
)˗�(���@tTu��<��@�WE���4��bvJ �l�U/��b|����{N?�<w�������<}�3�hE����N
��L�u�W;;[�<�c`��&)8�l���"�^M�A"���Fv���:=|7=Y�t����~������x��Ֆ��}���m�|ܗ���څX���`1C�����ϔ�w�`}6}�g����W�,�
3����I�x;�T��'��pK��`9�z�RTD���(���6�:�4��\��� y[D�����A�w���m.j{��i�`��`�V9t��Z�L%�H1vrb�#����xh�T~T�v�c놟_�z��p����ׄd�֝x�n���-� �Q�(0�{,�{��&VMd��Qڱ��D�����fcͶX���^J�f�t&dSlLD�c��8sʲ����?6��و�yL�������ȦQ�����>p�cq2j���L�,TK��-z�VM98���\z�W�p�6hr�հ�Mj<���n��Đn6�����ѥ�]��ۯ�2�l�
WjV���SCVe�N�|��!�D����_ �Ds;�Z��*�9�����	� )��c��&�aC��Q����R1L�;-��W�jGǓqt���D�I�L�E���Q�\ˎ��?�|Z[�(�84�^����'��XU!bbb�UqD>��M2Lҫ��Q�ؕ1�-_��*g�̌L�#���|I�o��xa��bb�D D�>����5�1ٛ`��A'�q�~p�͏Ɓr���,řI^�!_��V�P�vl�+�M� $_w7�0�D�~�I��c�^�_�`uQOԄjx�J�ȩ��9Bs�_h�9�7���
�d����[`&�0˨���g�������'��iO�/e�}<��=cb�]`ϯfL[��F���� �6�#����َ3`SAk�Rz���1�1�.�QT���1�ƈ�2T��sT(\pf�^���B��Z���<>�mǿ��/�Xb��p:|w�JAd��!�4e�2�N� ;^�gc�ud�S�_�0/ˉ��&X�_?�R��0xgX�G�<�O�U������P������9�@U�V*>�f��`����3������B�UNl������6ȇS�!3��%�1������ �<��_��FThu�b��ԯ8�3uu3ԃkZ��Q�2�����Q��L{��3��Dm�GW/���f�� ,ʀE(&�!@�	��?��H�:��K]ʺq���%ȪvY?�->1{a�߯]r��T��{�貚�۰anِ��']�yׅK�8�FS�~Q�^��	e����Y3̘��=_�X�>/���@����Ga%���$:ZV�~�WY]�Xdn4�yYj1ܦʌ��"��V��ʾr?����	v.���{��O*ۍ�d�n�UL�|�~�b"�tM+���?/��
�J]��g�l�iVK7w|R���{�Yh��k�B9`ȉ�:6&V��`z%�9N�+"�7J�͒� ��_ԛlj�y��Q�?�6n����,/mFv5׸����'l�����$�E��љ\�ͥk!]FRj�pG/��z�"�}靈_�p�Ә�l�F�q�\���TU���}W�=hv{�%�W|��e�FUc'\��ae��x�e(^e7�����FЦN"���>"��DH?Wxb�`$b��(�4�H�� ����HLy����zV�xϚ�������<�H��IA:�� �z�w��&k0�R�.�x��u�lhm�����qt��&�4%
5�_���|�����VI�-F
�����XE�⤾�{�7	��D�wT��H������?�Zv+N�H�8t�P\9�L��ZʃT�۹>��5N��)��Y�0!қ�J��}�Z'?h�-��W�u�ۿ/*��DF��iM��X�T��%�{��Z'�|�ڽ��]�&xs�:n) �h���U�+�r$�+h9H�L�5QM0�ow|��'l�c;{{dnKL�CCK	���r�P���D�z��6�����?���9����L8�^���h/���	�)�anS�����ݻ�,7��Xz�����3�U4E��������9��4\5;����D�&�ǝ~�7�� .��c�oI!�^������s�V���gb�Ϗ`����P�̚`"�P���kK45����9� ����h�1�8yM�g[���J�A���\��xٜ>DA�Q/�v��I����W9��>G����q��@a�5ab`���W�n�٩�&�
�z)��Al,ʍX�r��&?��?c#ׇ������+���pd�	F؏ӓ�vz=���6�P�o�W�v�?:��5'�ypb:�i؟(�d�>>�nS�����%�z�"�s��V�{Y<hO�'��cY�R���������5���I�@��!��,ft�@��̤�ԯM���g+`^��d���6&�yO�]7	QC����g�F�yQ�J9��yl�T�/ڥ�z��/e���|��=�*$�Jē;Q��Ќ����m43��imEbĖag��XHf���RfX#�WN�~���H�n��t��N���8�bS�Xw-��.��&��+	"sLㆮ*��!0��S���p�)��H,��ד�^�
߯`(�O�+8KTÛ�ŏ���wy�w��_�(c�������M�TPA���K���9|4G
����ஸaHI/S�K���q�ҽر��x�w]�Ңn����2ڞ�RgJ�(�uu�v軈�Y�p�t#��>���Cf����{2΋�nr!�;)!�lh�y�:���0̴��������Y'��v���$p^K�f&Md�����Z.
���o�R��bO�ֵ�λ��l�����wv���H�����`6P;c'����nIҾ��|θDD.�����g%���=��v�n�x��'5����Z�[O�8h����Uʕ�g�l���࢞{�����wo�5�і$~'�fe�j���m�������1u��R�n6�zs�R�i�-��2���k�g7�=;��A����M�&eI ��_dC?�)q>��t�1P;���7��7�4=�����-ѱ2rl����o�ࠋ��X�����چ�F_L3Uo�N�;�p�iT��:�����a�K�߻W��0���(���ΘJ�]�r���&*J�K�p��O�Jg&W̫�j�!�՚��&�"5���c̕�R���]{�E_�z&��M��%T����D��`i��JT8*�G��Ї"n�"J�z�q��\ n&�U�A'4n��&G�;�.Y:��N�GL<yz /��	�}�SV7��o�c�z�H|�d��2Ȣþ}�$���y�u����ϖ��#�ȍ�ƄOj"�#���MSl���fĸpw<FA'=ccV�3X����ǖ����e�u�T��'Q��4��5�pF,�A�5JR�.ͤ!SO0&��!k�!�Ƥ�g�[@��B��h�1Ct����֏�����4�s��Ͽ�b�jN�~����u	�wb@jT-�	��G
�6g��r�SoF��y	����ə
�F��!�Yb4��`���x-cSs��� z��vv+�8>��P5>��� ���l&%,jB�1�I ��A�Y����<�r�G�i����p~�G�4p���������z�$�;�Dwg�(���	ݏ�`�)�/��#f'�!3���&�W���Yx�,�;��&
0�=62k$v1sU�,Պ��1/K����`�2�Eߔ��5����Ř��j>HH+��y�U�6���M�����k]~��ۆ���:�/�r����z�h�0�U�m��I��'�;7	RhY����g�[��I��٬-����Z�q1��c���zN2Q�G$>X��,��n8w��_M�/��%���4�r�	��8���{]�R�]�tD���uT|<ʳ�+wx�ʭ����$l���U�<��x�%����đ}I�,Va}�TlQb%��C�~L�qV��ng��L?�ld�j
�&�3+��1J6�uޙt��^R�Ԭz���(��i�d� �3�BV��9�U�記u7��_���W\��������OJl"�ؓN�>����i	����HĆ��ƣ}�3w�"4���Y&�HcmSx\ڒ��&���������d��q�i�NU�Jy�ݑ%O�L1���q%+G�eoC��(#/�{�ܩ��%ۇ��h):�5B""���6܄{7^�؜B�Y6���2�H=���7�0���q n�`��&a��[P�<�_s^64w�6����H���)�d��5Ĥ���u�F��0m8��T�ihȸ�������Y]�����?���%D���D�;� >)��rp�e
V]}������]��Q����0�?m���f��w��QP)'i�m���,s�Y�j�|q�?n����]4V4-
"}��-W%rfF��x�F��q۟�,_����pX�m"ʤ�%G��y1Z!�Ƈ�3H<�[��'�d>�\�W2��3�bRH,������#[���x}���8�����ȚʷA�LԷ����.���β�"me�ŕ~��`:��a�����o���۫�z�N8�O�־���w��­�O���ݦ����;ci�����T�F*�.���3��Sg_���'r���#o,�6��Y��P�E!����*�_ȩ�⚛���9�,���}�xà�!gaa�e�a�AT�-�b�Ç��w+u��f�;������W��}Y��
���q&��B+&߁��^˃��������4���/3_�WCt��ޛ��9N\�wjSȋP�5A��D�:�Z�o	�O�^ƝFc� M�W�ֺ�⟡\�+��J�Ɉ�~�x)��wdM*m�u@e��|������ÀE����;���DH)�/�noh��~��(ha�<Q���)pD�:d2�X_IhgjJ�"��8Jj�7kU?اO��<��/ʋ���s�ns�-'���=來���Q�w�ia���Q�î&��۝O�eS.ԣ����	��h�B����,;FZ˒
;y�ؖ<"Fy���w���l<(�#*��m6��96���D6�8�t�a��D�np��������{� �C�Ca��kr�?�w���\�t8k�p.{�<̷?'v��N��_^o�b6��(�rm;A�*ǋ)�,X�hz80X�|aN�Ft�0�]��w·�n��5�(Ƣ�o�%���;W�Ƴ5�C͉��_:::>7N�v�eT��� ?T��6;M"�rj�"����E��|u�u�G�Tǁ����V��LC#:��?S�1���6�cF�$��W�˯�{rK������3)�+���C;SؑB�' 
�l�[���Q@��U�w:�5��^K�e���!:������bo,b���
��E^Fm���	�1Ȃ��h�skhW�(�@<УLfF�0n !Y�q�Y��`lvB�5h�J��*>��s{��b��^�9�)�t�<��#!�	�gA}W櫇������}�t�hkt&���\�c�9�ԗ��-��5e\�hv��B³6>�	����e㨯�e��&#�F�edГj�h���,�}L 9O�r�e�m����8vy��m��8�����k����n����)�փ��^W��O���c����n;^����)㒬F�ddd:��\�1����̬�D��(ҏ'+o�e��BdT fɦ7\�{jLs�t�ӊ^eEE(�5;��NM(���k4ƃ�8V����F��D
�lh� H�'�VI��"t2�@۹����u�b0
��Z���a��{E�gI���j\��㽶�h-�\�X�}7�￟���Qe����*��Ŏ��A>�=-b�E�(_���r|OTt��T�wǑܽ�~��9nv�� �]{O�-m�,EU����&��R!j��[U�f��/�7��+ �/��:��x��9`{�DV^�5L�D"�nF�,j���xvj������q����Er�K�1��,wo�֔$�B�m$A<k����s�����b�p���0���)\Ɯ��g
Q8��3��%�9n�<6ի��y="�*�*�4�Uۖ��Y�i/=?,��I'r�EW�*�6���g������S���Cr�K�/�\;��QO��E�SH�`�C���#��vE0Ϲ9=E�^&�~�rSCi�qǃq������}�W�	�=E���`zN?���
�#��X��;�� P.��-�u�M<R���psXN<z�b��]�Nȴ�c?ײ��g3|p�o�gE�,�?K���}k�i��㖅?d�<8u��^��2��kR 8�Y��)�ȹ���e�����h���Ξ����� ����'C�l�.$2G_�� `��)50C~4,��X�7����<v�PV3�D�?�������@� EVn$����l-�f�>Q��BN���$#�g�$�m��k�y�Ff�Ӱ�2�C���>�
�[��v��zz������Z��0lY8����?��d(�%A	�"Ǔ�"C���������ʢRzF�c$�虍 ��Ł�n��=���6:\b���|�2����OJ��@~ LL̂y��*�V��WJ1%
�I�<q��I���]^��4�/%q���d6{�Qs�8C��R=��]�Η �v,����6�v���Y���]�v��;�g�K������Vnb�#~�����t�-6~���Q xF����f�� j��(3��]�8m�.�Vr�"w�r�o�އ�j��D��Ꭼ��BBr ��4�2�fA�z��4u0։K�*�I�b�[{���Y���[�,Э��K���������ya1]p)�7��)0�o���)�Bm&�p>��%��$%+,d璂�.�]�Ο��R�9���� � ��U!q`'���& u6�� �O;=�����fIC�US
�;<?{�����[1&\��xl
�������\x�]̃�R��/n�g��[M��$���M���)�@�Hpm��ߏ�4A��ptq
�ث oӚ��� ����J�'��"lX�3�� �������$/Wo���|�!��x��m��.�����%�b� C��j�gq$����� �UhQ�Q���N`fIk�Oũ �2a��р�9��k���SL��_��v�#�#/,9~F��x��*�;�����v�51�A��ԛ�
�����3���/c{+�
q�{3<I����qh��j�i�����k�����A��h����~���V;�m��ٿH��d%���w�ϿrtT���qR��l#��al��!\���~����B��^� �?;S(�.r_�~�ȭ�%��+�^O#� ������Vv��l��I���M[���ʏ.-F��������'L'�-�|��$D",I2q��L�����ᘲp�X�V���׶A��ūz'�%���YN������r��ݯsx�����&�0vߊ%Z��ύ5��ZTPb���E��FM҅s��v-�k��&1�;��4��v�CZ�H������Iq~C��?�sB�񨃸"!����q 1D��SK���q%���֗��|�G�cR\X�(���������g��vVF����Cz؇[�z�&¥)����닏�e[Շ�J��a	s(~43���g.p��Z����NO�j՜\9�RO-��GO�U�>X�f��ԕ7&ГNMDy�t���"#���H��.��q�u�S��B�+o�>v�W(�!ffI�b16;d�ӱ��:1~3z�p�|gQ��u9��,c��Df���dI(�4r9����w�Nkj�cE3So#�~��a����z�{)��߉�KR�Pￃ㽪N;���0�?�f �e(���q�D�j��v��v�/��^:����av��*�Bf�JN�v�D�d��z27�����LGI�i�ԏ2����\|T(T˱�H����tg�tɖ'+;{5�C05�J(�~c�)W��S}��h�!*����g��|溜b���v�8�cgf��^�w��v�~n9����/�����DQU����� -����F�Z���b�Vf�Z)d>�>�������Ƙ]C!�45V�mQ�/�"��hQ��s2V�d��X4F��λ��Εl7�,��D�4�(MTٰ��9�_Ö��{&	sɭ,Y��D[ܾB�o�Ø���*�C*dB$h�{q&�ha1�I�ß��,W��\�uϗo���
��'sPa��?X����+�-�)��T�!�gȾ6������Qe3_M�_�$�s-�Qw�a������z}�X]�G �d/�x��%�5l���uWE���#��oB���#x��)\��Ά���[��*��m�p!��+L��0�#Kɣ�_��۔exn�5-VD�y[�L�ѹq���x��K,��T ������v�b�]$&�U+^[��Si�o�]���څ�������1~�����6 ?�u3mѧ,�2P1E�6���'_����̈́R���hek�z�a���M�-�Mn�aK�L��R�V�"CH�!#����$�4����ͮ��C����ZS���ォ�����bn6+����n!Jt���8�XH�3c>�G;�N�R�g�+���:�.l�u��ZH?�->h@�3zNh.)���\VQ�j��88��?��0�o�5	d.9&�Z��ςw$�g��&�*i��FO-A@�Ů
EI��3�A]<�ì��>&D�P����V%'�����NE
��9>G�2)��D����3��ŮZ�T9�$��,!��G�o_t6~d��v���N�`!3L�w����Ɠک�f>K���ZL<�ܬ}�M�IL�1p�����}fO��j�/����<�.�����6�aS�۟�L�ݺ"$��0���Bh�nB�}��{���1�h�D��z�Ŵ��ܡ`�����N�����قL|�J6�h�]8�AO1�2�_+�?�촮W�����/�_�������pL+4d�ԯ,��S�װ��/v�퍶t[7�����j�KI��4}:�Y�7�Wz��O�C$L�f��&���7�j�rrc�PUI���g��`a��7���w˱zyȖn�[����þ�_��i�x��F7 C	���,����鄑dX�t�ۋ���A�D����)�����2J�Z��P�f�8M5���M\��"���6!ͫR};ϰ�/���Fv���9�rR�ʘ�N=��"�k�"V�_�qIµ��0��|}>9h��ۦN�K�r�L�~|I	�\ia�k�~��=�'�SWW�Y�"��K�s�@�]cyTIjL���H�E�����[�����"󼎗�e�6��(���y�y8F�%	UY�~ٶ����(�9��jo'��N������)�n2\!�����{�2V�p��}x����Dx�Ë�t��d3�͎Fl_F�8��?ɦ[�_^r���*�H���K�������d	%hhh�F���z�A@�����������?��m�;�᎓s	����)�K�XX�� ���V��r'\iE0�P@���k��$Q%������NR����V/�%�d-��*���Gt��C�� ��95���֏��zpG�9����{ߍ����j��iZ��@����C&
��Q���y��g� ֘+�~��3��\���ޚ=�1l�љK�N�b�a��n��2 �@�[����R���V�Q�bH��I���1_�&x�����<C�}��Z	ǑewU�d��U��t�-c���[�d;:������Nɮ��ʆ?��S&��#�;�~���hBɟ���#.mȓ��#�b��?�\�%�=��D9=�Vq7A9�s�U0~�H��C3�)?S7�������`M'zo�/��9��N��P	>��R�Q�Y�c�v�	��"*6�U��ؐɷ6Qo~ݽ9O�b��\�g�]�݌ ��q�=��֗���^兡%����@?iy�얾Y|��f�6��o?����x�V�t�܋�r_�>St���G�>�����%��M��r�6��!_?�KB��8#~tY����Ta�4'������.�Z��Б=��8�K�o�Et�Ϛ9q�s���+>���[c�wcYs��W2i_���Gl�>�7n��n�/:[��E�x�_�;ɲ��b�$zMer�ۛ��\��\H膿qe,L���4�OW��c��?�-�M2mԈ	�V̾�s��p�����:VU�8.`{F?�'��zbb�冪��F$Jzt�D���(+�:FP׮-���_?�x/�b�I��'Z*�r�ҽ=��E/"&�{~��Bj�/%��=�u+GR;��<�^o�������?�B]u�Hظ5���B��a��s��St>��&	���{��f�qW D��0��p�0��F|���7&�<��Lv��P����.Y��ݷ8t�#��X��86e3�1��`� ��L��As�K ��Q���fe�
N�ȴHQ���_�)ibp�7]�1�_0E�|�/��{OI�5�+[K3���xSߛ��K����=e��>M>|�6omt���#O�˯�20����`���1D���
2�tB7іq���
osaBMOfN~�f�o��6����P�+*���Q��߶�w��Ff#ύ��U)4X��̏���\�P�������eM�{�A
Fx/�U3���7m��hLbv���ģ��Y巂�ɂ$���5 �I�n���� �"��Tubn���$�G����ui�Բn��f�%i={�t��d��fP"&�f��+�-�߉�TUh=kTH���͜��0����a�`�#�<Z%�}��l�����/��%ձ999���-��m2�3"�NLا�<�w��˯7����책�x/ő|33�W�ţ��-�����6���j��GVAxl)/R*�����&BN裢�Xa[�������([�:]�����B�wsU��K���ү�����j&�z�Jʿ����jX�"y��/�G�Z�bDUC�|O�:u<�~�EC1	���x�1���$.���߹��X���/"���*[�yh;ӈ���T�z�p�޸<�lI �8�샣f��C����v��R�ڹ
F��(��Ů���^�l�C>C�5v nmM4c=u������y�N�Lέ`�j�ϡތu�}[knB�v��#�d�pE�6O���h�
�:�0	�=�Cpw���.!�݂{�?�!������C���忻�WEQ<vf��5&Z��.c"V"%ůт��%��PJ�$(^��~�D9�0��,>�I�@��D�^���G%fo{�f��1��#�Ol����ؿ�P���;ko#��ZҶ؜���� �t�f�>����#�ܝ���h�I�e��ҡ��ZP�<��sp�J>�0�X�_6j��gE�@��q���� _ґ����Y�L)�گ�>rtd���m.G4�SJB�ɷ����J���y��'ZWY'�|��/Դ�q𮮮���xiE�j%�Nvk:qaBL�UwfP�M�b�]�p��M�M�M�HB���!��ʅ��ד�̤��QK�i����Qk��~0�ITe�nGS���k�]>��`}��F������6�� J���a��]���d>��&Ts�H
���h��R�"U��%��t�Q�1�R�ˮ!6c�c'����"o�N2`.�wƞ���
Q�u���ǀ�Fq t+� ����bXl� ��ܬ��iG�<�d$@ӝ��C/�=\�I�SN}}��f� 	�T�6MzG��7}&��(Ff���ܴ)���8���"j���8�B�Χ�nʞҗ�uOq����JΜ�&m�-��$���ʱ z� �$�&�1�<���׹94�19xO?�]7`#.Kf�5��$�r
$�ͨ͝?��>�':k�|(�:hI_�ғI��'2-�*�e�ѱRc����!�8�gXo\��g�w�>{��l��S��L��#V�'�73�2.kń�2�ʶ���}\7\],�ݪ?���A�����f����-�ۿ�*9Lf��\c�����9/ܬ0[���n��V>	j�$&�V�w��Jg��쐘-�,YX���Z�55q��x���q�ٓnx���~�Rw����?6HD�Ƽ�3]~s�����@B��+*���x:ĺ��Ӈl)M����g3��bhR4���R3�Mʁ6���#�􀯕NE��ȅ�5����`�AMW��� ip��{�n͓z��$v���R#�0����x�B@7���>����x��Z/�ga�Q_�9��E���E�?�}0͞gz��|Y��ʻ�A�<���o�'���'IC�c�<��^���=J��؉�JooݷL�J�1���Ҥ<=�|��{������(#�\�$) �U�~��UV�-Mھ�E�b�܌ih�J9r�P����죄��@8��ޠ�$�ɨ�H�q��o�Jn��r0M����#�9�Fv��1B�+sSv�a���PV��Mm���_^���z�u@��g��l܈��H#E.B�m�ϗ���Ͳ��/�t���P\N)��l�x���zhi��!�_;�!3>歲G��y8�)&A��ji:�y*Ј^H���X&/����U:�{;`���(��z��U��GY��8�����S�o� ��*eZV��5%�ھ&쿶ܜm������b�.
�����𰜺}Ղ���s��rs�ww��Ԓ���ڵLb�9S�*P��(5��ol�ݚ�7C��>hiK���k{'��!�眊�&UЎ���[B�l&^�Hg������FN ����\������4Z�9���C���`y�]U�g��zi�3��6n����`8��(���X�����^V����BjS�z%�k��F!���|PM-藉��CĔ����ԃގX ��2�
��������.�1TF��Z3�<u���{����`Er���Qi��5]��[F��j\���V�\�)�ƭEYM۝3i���u�u�85���',� ��ӫ�>�8SbAc���%l__�'7]�э��4�M�!�C���L���_\ @�{�4g�P���(ؿ��RJM�5R3>�DV:��]���y({%��Xo�j���R�s��N0�'
S��Px�8�d˜(��JQk7�~,J_O�$?hR����d�]׊�T�/U�<��'Q���@^LY��2���"3B����:u��F$^�Q�\���C��^1����ra�/���\���
�ə"��V��Q���W�������b�xGN�wn�duX��JW\����ӖC�s|킌�	
^�ȊP6�	��^�}�����欹�1Φyw*0PV��6�d?N��B�<a�������4]�~M&z��E���A{����y��WS� O�+��o93��1��PFN�����3�����{�Nd�XژXN*L�,Ǚ��W�|4׆G���b���Mv��T<�qЎB=W�����/��w���",�1s��8�غ�T��̅�Q�d�,{ғ��l:����}vB�&�$2y�вW�0��05�t���mzҷ��������j�e���;9���m������R?���7N)�r���SҞ�[(�:���SSǋv��kRn,��f(*
���qըv�S��2�^���ǈl�%ٖ����͎�y�M�^"m^����Lu�G�D�f8O��,�jP��׍��SZ��v�/d�^��S�>�����*�b�W�+|��Ұ~��:iT��3=��
����z�F��z����:�{��)��`�����?]>��yVvD��7���y?�n���)��Z���j��_�fY?��ⷥ�oƍ����J!m�G�	8��mh��3�c��k��p�)��Ъ����iT���&_I:������wUW7�M*x0��^B�~���4�]��M�b�#�f���V��hUi���Ib��3�p����H(���Ŧ9���)�4.Η��_���#��L�|I1݊�:�H�=�f�D��Hr�@$�9ϟm�!�я��r^$h�3�Yo��A� ��Q�:s�XFv�O�@���R�l(6�9�����r�<�D��+R�LRhI�s���!R�/�\���[3��/XWb��P���[������7�FtG'�@|X�#Xլ�DԐ5��l�w.������W�k,���bD�#X-�?IF�Z���>�,��>Tl.��n]݌�����u`���!�~G[g�s6`󦤦���.Y8hQ�|������֤���	�O�l�R�&�@-���z�ff5�|��mu0�_M-0%8�V,��h�sD=�.t,qYp����	a�2�t:
a�O��u��6O7p/}��k?q,���0̘��$���.1����/��չ��D��~��xx�Ύ��ͦ)6��K�0�� �i؎�.�5�0�B%��ݣO+�{�C}g���q��S�����=��q��=�c}Cdf��a^�t����f�wlcjĨ�Ũ\?�n���ȹ*(v@��%�����)���ٸ�U75�$�~E�U_���(% ݗ9�7��}�ʧ��1c�xI�>�xYm����i�	F&?��$�8�����>F���%�?�H��=�<��7і#jԿ��"�� �8���~����}kO��W�օ�]I~�X}��]!�����(qy�L�����W"�����.0c�����ߦJ�r'�H�R���i�d�d��OL��P4�v���,=�Ug1��g�w� �ٮ�M��a��ؤoZ��� C��SU��w�Yf_0� ]��
�
!�=��=����,l���v�8�������h`�a��R*����{}���Hq�م���oo'�I�Q?�>~�Җ��%C��T� ��A#���J�,׿�hf���_�5�Y�Zl>�W���DԸM8��wi	TU�f�j���3���ގ���Q��$E���#<7����s�T���$̻-޹�2e-��zs0�A+QY���u�	u�{�`���
��]��Ien�d=%Je�[B�HUz-Ŋ��A��Q�[e�G^]�TZ��T��������1�k6r4c	�0����tK��.�����w�F���@��pn|f�|�akj�ȣ��7�����k:�K�C:�UC�GnmC�X�ڦ����85��8�E7>6�`����F|s����.x�C�>�y|��<�!�e�n��$�@�H�m�[����Ue�5���c���5����|܀�z��=dk:�Qx����c[�옍~�E�$�V��e��P�
5	}𦶩כ"�V�y�s��z*����5���Ҵ168�K�{=�,a��0	 Ř�=�>��k�E=5�_>l�>�SBwS}��93t�?���@C��t������ڬ����خ,�4v�H���b����R|���aZp�lE�x~O��O�c�a�/�f�+�-/���Z�ibD31n����/|
ȅ�X�^3
r���E��͹�f��U�_���Y��"���wF��)�\����>
	�V���O�{�nm8��3���K�j�LCH{���0�T>n�{��P��2�"��r��gn��c��e4�R�( >��}���{��E��_�]�^��M0�}�#!���Hxl1 c�ϸ��Ĝ��7)F7ʓSЉ4�9�f����fl�B�u��<C�L����쬓:m-\����Y� f���
�b2-��+X�3�V�́���3/�4��
>�L�}��?���u��d�Fo������R�x��T�{51��V0�8����5v*�?C->�c�y�2���ׂv���I��˄m�# "��ǃ���%b�kd"n����h0J歕��P`� �y��ԇ�Y��j�C�c}j*(�����y�G>'t���c 2x]��~n���}g��th��K��B�z��7K-S�b/�5a,_�(��Şc�M����H�nڪ��?L\K-�(oO���n2��U8�x1��oIݪ�(���)#��_��j*�(���h����s鯁�i�m�@�C@���H��2�a�J���*�#/њ��=Rm>]�FFg�·m*C�O���㠋����[99c�:� ڕ��)���@h�vQ�:��&_=?�n��D$ (i�{��t��Y�F��V�t�#�$H�{]5�T.6e�^���-ɭ�fR��{�����7Z��� oR�Y�޽��a�ێ�C˨�X$�F �Q��|���n	cj]���r�[V�p�	�&���]i��+�y3Д��	���}�O���õ������F�����{������1�7�B�*��&�Hu� �b(HI/�ݻ�(h�_�ߛ���o:��-9	�LOD܏����P��1%�<���oW�k��x�8���0�9='��S���d�����rؽ��/�q<�rH\�|��	v��Sn��*9ۍ�wRc�Äw.]�*�߬��[��4��@���@��#�{K�_�d���j'�t�����8xV�TD�ٞ�|�!Y �ԅԋ�V�֙.7Zh�y[�p�p��P�s-�"�}���Z?j�%:õ$�*����nӜ1(b�����Ӝ(G��˨���@?��*���@Q����e||�'�k�R&�(��tH���������<�}�n���W��zq���eĂ�ҵt������y�i����W�ɰ$Μ�{�'��-�%h�k�%�	��a#�"��U���vnD�׾��e�uA{�1Y�\���ig�*a��
�%/�.AOԜ�X�<%$v�48�D:m�ۯ�ȨiH��d�����R��}�M+����7���3�B0\J�md��	ӕ�d#��bjJ��v�[���c��aʒS�l^����>p���� �_�S������j����Uk�?\MqB�������{�D]�d$yni���]�)�E/B��-����\�5.��r��"��2��� _��=fF�]�<?�{}����
�<�p�S�a}۴"����X�|R�i��s��~n�����SS�+x���˳�k�=�����J&X�Ѕ��J}S�:E��҅�.^����Z�r��Z��c@����j�4wD��H��^��u=����jSTIհ��P��@�K�?����1�q2�m4K���2�M�9���f��"�8o!��W�%��F���-�~J�=3��,(+HM��K�MM�C�}L�����K�,�{Z��8ON_|٦{'8�TV�	fj��3����K�PC������s(���/��2�R]5����埞��V�`��X:�i���e�R$��3Qc�;m�f�L��D�R'��ֲgjv��L�z���CN���d>bb���~kE�w/�:�XK1%��x�J>W�fb'Z����U���C��o0Q���'m�~�|��q����8a�	j�������� ��"��f0H9�B�����x��N� h��	Q��4�d[���	��: � �����Rj�E���su©J�g�3h���m%�5Ш��˫����~-~t�V3NOs.4��su�*Ӗ�5�rʩNA�D�+�X��jX�Fs?<v-��r�2�����x< |U[n��9u+;L�3lxQ9��|%՚��ӯS���=!��جS	�g��ET�n0�f��
� ����R{���*���S
��?�FgһA��hGC3����{�,��@�I	f�ɑ
v�f�c�[ &�b�3`�xW,��f�j�%���z��,e>(m�u��%��[c������<�.b�P������{sn�g0=�&�$��N�_�fw{�`���_�۟Pj�W!�lF	�톯��'\ĸQ�A�(���OP�5������(4���q��{0s�{x5�j4m��<1��W����m�&�Ì�8��}��k"�e���@��$��mb�}��t���
�b�z�{\7�4*��ώ�S��4][�~[~#FU58r�u�<b|����*�ra���X��*,*
'�����f+�Ӱ�e�'r�}����H�љ&�:n����C�l�����XM�+��Գ�-�bB,��SHⲴ���ǜ�䥉�=S;���Lr���K\\��T8�`��?�?���(T\��|*�k)���𪬮`��Y)��vӹhe?m��t�ŗH:����X٬��s�ݻ�,	��0(4�V=<��������u�����o!W,!�3��Քt>|z������oŴ��]���[6��m��v�_�����C������z��z��JMo�V7D�7	:���⦖�'~�y����ou�ߊlv{2-G��*��1��#�36Ql������S��$C����I�aး���g%|Uuƚ�Qڕ=�#�#�'*���@��p��3�*�q�I���?��҃_ض�g>q�`���ę��DV��KG�D�@��:����ъ����gEy�gۡ�1��!�vZ�Y[��	u��"{̑"��jOW��R\Wc@��(��p�>�^l��]�5hd/��yA��f�M����Q�`��8 �����C����+�����]1��|�c� ��{m]=�(Ǌ3'�1'<���k�����V�~	����^`�@�I�EZ��9���������w�OM�Kb���|8n�P$��	c��{�*���5�/Z�,[���@���}� |�SǍ}�n��0OG]Ϧ�͡���Y/�rO��s^��pܐY|ǑSm�椓�O�����1����G�𒗠�H�T��w_O�a�+�9_+���O�/ �S���������/P@���L������QIU��!�E+I���~��L��0����:�W�7��U�����Ϩ�jm��]�Q>�M?�>>�-j�H�l��}���m�К�jm}��?�E��PRR"#//.&v��H�m#�����#�������Ӟ��~`����p�C�������º��<�����&���7ݐ�(�����kt��G��wV7W��e������$\��z���kk�#bf�����H̭>�����e*-���hS�6$@��=;+�ٶ!(�jo��D1|�A
�'x?g_f~���tttl���D�tYK�!(�Ӟ���0��g	k��H�Y\�m�ĲU�����[���&_�W7ԶR�!K,�o���oe��j����y����Q��	���n 髦�0���dI��(�����	l�5:55�>Tq�M���l&+G/cO��v�h����
^�g����c@��]^���ΫF��IR~�k�`�S���t���w�uh�J>:R�h�Aab-��*ƪ���i�={^ ^Z�/�ϛOpUh#l�����M)D�K�=�7���� ��kp	����A25fX�8��G���c���ە'D�3B�Z��ᛂ0���@��^��k��r����J�A���M��Kdh�G�@��� n��_y���nA��(��}r"���B�����޿~�i( ��_qz��ⵐ��h�ȇ�����PF�
+].a��!4�<��R�`�(�-|������z.�i����	�`qa�I���S�^L3�=_�R;��v�5��� l�*�p��y���܏��֖�۹h��C�pl�ڙ��E�d7?%��G�Z/WF�Z�`��\����@��=��/�ܞ�ó�3���4��Bi���B�p���gus�p4�6���+��]u&o@Q�/isʹB�j�D��C���b�������I..?O=�0y;~[+�� �i*�F�B��#��k
F���gM���Oy��K#i�Y���#���w{��a+�XS������g�`S���v�
V"�7w \8���TC0�Mw�� ��#t��}��ˎ=��U3��h�yty]-q�	g���[��+2#�J$��Swj*�0J��Ը�bW`��f�S�O�E�O�E?������Oʶ�Y�F�賺�q�3�=�>��!�p��}�gNKt
lR�^��j�^���M���^�=1�ʈHU���օX4Qʽ˳NG.��'�$L�Q�H��.����5�@�BC�9W�*#@�ы�v�9Mebb2
c��.i�m����N7��ƈ'�t���a����Icc
퇬)����r�hs�~T��gBln���\��[P`�`����)�̥\UW������qǖT��mkP���8��r�>j���zggw$�௸��긾�k��J��3�������'�a�bĖ�;!؞:*s?��D�|�['�Ž�m�6#C���������B$f?�v��z��J7-�h�����M��S��A�3��o� �y�PК`�n>b�(��)J��],K[��������~b{J�5Y�hC�wFA[䂀@���uU�W�J���r5_mS�Rm��б�0ɣ;�D���ui��1-/�� �D�>�:�74p{���!e�(����v�.��Qy�E�Lẘ]�(V���e���+���;�d�H`�зT��!�w�����D!U��FYA<9�3�g�QZ�cɶ7�qɭ:!��h�aj�7�L�Z?wS{<8�c��T`�a�GC�������m��b��T���l�X�a`&X�x�YPL���h����6!lF�q2��u�~�U��"�в�zc�ļ�q��U�ȇ�HC7�O�q�~{�f%��
Q"����Ԇ-��G6� +����V�2n���^���K���K�A��̭��}�Ǆ�V��
i�%�ꬾ����Jr�h5�]�ח|r0��Vk*�k�K��a���P�5Z10�� w�%���Q��Դ��R�xG9f�}Z�p�!R �n�D?��(����-$=�N�jX��YY��&�m��#�]�Od)��E]?)�X]=ͣ�{lU@��s�/K�SQ�ޫ5uě�V���U�S�� �X��{_�+���(A��Qfu��0��4���>�C�u��9��~}ImtK�K�fv+��3x���.U^��W����j�PcƝޏ*�J�-?���^�΍�`�n{���Beg5���N��kI�Ⱦa��O���jAoݒh*&�ARE
����6L��! ���Q%���-���o��.>��W$��7;YBn҃���%:~6�����q�����zVCv��=+�rz��� �ROj���\͛�����C
U=�-�y��݂�n��zn��O��I	љ=�vG�d���S�Pl,�ć�aJ7<�k� �z���Ѱ{�Z�^!��_&G��T�W<�ĳ����=�c��W�����>q�}�����/���_�aN�(xq��C�B!���5-�<+�⑨���\Lf_Q����Fɰ�d4͘����
,$׽�p���"��H5�H����C<6��AѤPٛ1!�4�i�*VN93����p@�T�ɛ%��̗�J��|p��B�����9=�[��%sӁ�OL�.d��^�=���(�(@D��z;r�Ȍ��������ل�H�yn��X: W8�4��)�E�{��Ĝ���Yf?� �@��!y�Ϣi80"�,�j�R��G9��?�"�4E�K�x�BF��|y��\L	@[�ON��сQ�U�GI"T[�����J��5�;y��A{C���(�L�4����n�̝�Ǐ�Z�a�-XJ�bK�E���$����h�2CT��&W?h�#x�1^�T���#t�����1�[λ�T�������8��P23U{
�>C����FA7�S|�:Fz�*&:�b�z��j���jիRa,�d�h��9�L���	�H/���"�RQ�����*�K��#1y�ͷ�U��6����j����i� �w�b>�Y����*N�M��C���u�pLY�˜?��6Ձ˿���csW�����F�7�y^� �;V��ĥ�r:���9�:J��2�����[����c���Zy�B��S��B���M�������K-Fڣ�;�婻���G��_`G���&ϣ8t}��� |zrbNcV��!5�>�W�C� �'7@Ck���t�G��뉘2�Z�ct|ٵs۽�W��"��Of:L��!8]�Ӆ���?^ʒ�-w>�����.�%
��rr�KF7�ň�h���YK!
Xt�%x�����H-8HT��.�XK��<�Ȭ�+1g�|�z\�	i�f�c�2r���D��Un�7x�"n� s\�/p['�r�a� z�t�\^ ��i�$�
A�XZ�l�����}��/�[�b����j?��F�I�;X[R�����
M���}���L�KAȔe���������r��4M�5���p'Ֆ�R1��^Z���2�� @7\LR���H����&J��ΐq������ѯ��gxóm%�Z��Rfz|�o����Ԛ������T�V�\�����Ӻ�G�2ɺ]���TK�E=-zBZ�  b�5GO*�/������X�f.�ӊ�w�̼�e���ac㪣��_&v�\=!����{��
,3�t�eM�-�K��}�_M�RUl��(Y��2	��r�E�!�W�q�}�f�����s���H$,��a���1���
��0�z4Ex��z�U8�J:�*%SǷF���3�mmf��'�pU7���`�������b^��ƨ|���[�cW�G����¥��vQ�Vs95�tn2�t��?�j�s�c�n�I{���u�8m}*�>�]��|g	`��Ф>�U��k,j�I���<"5�5k�J��9�eq��c(�K�Em�/����Yyr:�ӗ@�Z��M~�	�˧ i��j���v�)�$l��X�7��n �0��+���}f�Rc�.�0�.EuH5��ݚ�ث�mC$0:ܘ�H��ꩀ>A��VG�݃�A�ᖂu|䢣]�K��&��S�/	2_�f��~� ��K��Lڏ�(�+������	r������F-�0V��V��Q���Wj}
�G+eD=�:��g���7r��!ϓTO�\��.���A�,h�r|�
�TB����
����N1�89�]�K�<@a���$��R�~�|^���bF��u&�����j��*�c�n������*<�ʈ���X\�����V�X�ܓͳPh���D���u�Q3�n��k�$VEi���#5p��plW�A !�*2g?H�NMv���;��J^9��>Fu�b���.	�"��\*?#����@$��D��ú���{X�."��^>k�B��_�Z	,$ՙh'a~�}� #�zO���M����t̽&gQ{�Z� Ut�H)��90���RzF�O�Ԝ��B����t�h�$̔6��陖O;�x�sK�h����l�&��Ʋ;���TM-ųF4<8_Qs�1��1I����;׏����,���J�\�14��k�ӁoX�[���":b���_��*]��J��h��p$��/U:@!��Z��ӊ���� ���H#�,�,�Q�9ᛜ*;�#�w�X�U0z��δ)�;�s8Q&��@T��Էb�����OS]]�0�!!��g Q����&����+�D�TZ�K*Z3^?[���,G�����`�RQPm�����/��c��*(�J�.�����u	�d}������c�j"3.$�D2�����Zr������C�����z�
�������#f�^<P:z\<B�ˣ�Taq���+Wa�
�s�&U/a[����j�Iu��'����t-����;�G��D 9�>H2�,��b�bh����_Ck��C�����mq�>~���7b-◷�����d�9��s�|�� ~i,�Sp��++I�Q�QgҫG.VP�Ü�� �Ou���zD8u��4:�d��+V�o�ً�B>֣�޲TL�h>kXCa�J�фv=���5[K�����p�.�j�����pM���զ��� T𝬊�f΄5�7ޣ�O�d����)9��?H`��?��J�����;�!x���ׅ狐�EM�d]�;.6�ט;�FV����}�3�Z�=��w�`7�w�`�0�hˑ�`*Ӳ#ʔ�c*���rd)�s�����h5��U%K_m8�C���Tc(l�h"2pV#;�#f^�yw����Y_�v�@z��e�$��%� 'y�� ӿp�@ �z�Se��5r�R��$���
����t���VZӸ��ꗤ���R\g���6���?�E���˖���/�:�@�����le&	�p�G1f��u$�:�?���L�]#�Lơ�Xة�4ݔV{�y�?�H'JvP�� �WD�5��}��;�]�]���/Y[�4}b[�6���p��������EU)R����� �+C���^�b7�qN�R��`���b7jg�(�/.�1s�8s�g)�oL�_���+3��
��x��5%K��<���������{;CX4Z�O�'�/t���_��{��q��!��Ƴx	HIJ�t���J�Ã7;9�~3��naJ՗aX��^���	��.�2g߉� ��ÁD591�YE#NT��,@�$J|0��3c����j���/iB�b�d�1O����C��PªL�pψc~h�����<�Y��ڣf5Ycap�}{eBl�B�r����X������	5�@��&�Y�a�q����[�0��iЧ�4U��8�Cd��ә�7J)(�\Q����*�������%�D��a���/�8{���{����I�L��؉w`�H0w=�▞���)��@�y��82^\`$�e�Kec��2$A�2�7ˡz�c`�k���+Q���t������AF�N�}6�w����\x�t,p�
���pPh�D��y�����f#�l��
��+�a�?^/Fu�6*��S�s�e-K��H���'������a�9��w��k`8��eG8��_$��L�
���<��DǏO�/°�]E�V]��h׳Ei�īU:����c���U�[��(m���y��!�F����f�w�K�H�F��b�S���,�a���s��sZf�9Iڀ�)�9����:��x��+{�����`:�_�]~;d���G(�[��d�t��'ͫ�� ��̎��c�0}�k'�͜�������~p�u?j��%�[f�6�%/��X9*VK�X9�|C_1�7�d���F|��K����C�[���{��W^FzD�fR�&7-��7^��w �]}�8�o)�ĿB�G�[�X�X�n�s�	�����2����[ȴ 6fl�a xnհ����H�RV| ]cCwL�C�ågBܹ�{=6���N���͒����]�(o$���I1��І��k�6�4G���gi�Mn�g��^UW(��B��.�E����3C�hܴukjg¡n�}�C��p���{�<�4+|x0��X�z����L	3Zn	�ks����-�U�ֈ�ZZ�^X߁��Y��!���=~�g�_L��)��n��B����u��¹_Hg��A��h/��a�3n�=�:�z��:�o}��t�kE��x��%:9.H��O�"��#C
0x^*��'N�"�xz|���84�ϣ=��B乼@ue��Av�"��3ۗ�:wp�Sr���(�{�+����׫�A�4�A���E����6��D�b��94fgE��V�+����%�Y�H���F�5�$�k�����XIXo1�J���%��<v���n\�����K�i����1+|^O�4���Hk����{.��a��t���!�\5�x��x�}�D )����`� ��|Q/w��Y�L�un��),%��O͘��f�<l&�Z�bp��OӰ�>k��Fk��X���� ��0����X(�p H�VS��i���P�(�{���������s+S�[�����m�E$��DD����F2=�i�� ����p�F�������w8L���h�aw�|���Uy���"";��Y�wO��a���qۃ�25;bSQ�8Z7� �ǁ�B.D[k.�ΐ<�Ѹ'3z� e��E0���o���nZ�o��HJ���'(-AV��M�&!��"He�ʮ䫉�q���Jh8���ش#3�uD�����^��J��ꇳaާ���Z*Fg�w؉�h�)N�����ُqy&�FD �����mu���G����d���h�vbh�z#�>��@��z2&"�*;��CǮ4�F�$s1��z�����_���"k�Q��}3��j���P�nX˰#E��i;�4���|�׍��
��{ZA/{�Y�S��h��B
H��*�a��Ř�����6��'���̸L[�tLw����Q���sԖ*YʮY�(��!�Q		p_��K�9![����~�q�g�aU�
�V;w7�Ix�o�˼)̑>ׯxl�����=﬿ ��,[�"q{�Sy`�]��αy�@�'��&Hsӯ�'r1q��b�]���n�5�gB�����XJ���b�e���!���w@�.:���(��3��O�r�.3���Q�)� =�f������A�ѱf+zy����r&e��B��6o従�x�{�Vu���%V{�r�����4��8�]�Ȑ��Z����:��M�~5V������>(Ց�^�����W�v����;Q�(9�����&���j�DA7Un,vt�FR1rȿё��ވ1r��x�W�Q\+�xO_�xo_�h#j���s����������>إ�_����"[����P�m�HWj�Z	�E�1�\O�2�m��>�nEd|Ʊ�{j?��}��Ƌ/A9�[�ban���K5�7�����?�d��pYo�������>�v��>��m��$#���>n���`����f4ٛ�\[+�?hA��z������qk����bO���o�V�P�I����Vø@������	�������g5���vw;.�Qw>ag�h0��Z�M�:LY/�Orݪ���d6VJz��^)('e�῔�d�ȌJ�EF\~bf���B����kH(��B����\�O0���L�I�ᇽZ��`��z�p��5P9C�Y]P�A������j�Ǹ�ֈ�~��ƫ��Tl��zw����M�m��+8�bCC^�Q�a����S����H��	^A6�)��ԃ���Q�W���1p�R�թM�c))���G�vnM��y�l��m�jj}lv�"�j�bB��*� �D��M��Ba9C  w���`��f���s�;��,��V%�a����_x�R�xcs�c���7�;ZxL��I�}(�P������k<�.����P���(��gӪ�W]���k���P�*�(Ou�8[8�f� t>�5G/�X-Nb���߫;��,���blQt#~�l���%�O�%�&�@`3�N��-6�Vs>����x�	�z�p��.<^�4�%MQ%�gn�	>�f|���[V*��_��Y@x{|o̪>�W��
����Գ���B�V�;v�h�9����ego�A�j��K���grq�z�������J�/6�2�w+ƻ����M�	j��!h'�\���Q�&~G0G�H�fl9^#'`Խp�"&+����e2����Ϻ?�Jv���D�p�8>��.�wrA�nm���p�b��ǃ�P�:/Su�4��g|U���V�g�FJ�;�K�[�&]��zy"#�@�<��������%<��E}�P�N-����:�5&��_xϢ]��t��,/?�"ۣS��ޮ�t.�#0����ӽ�;�݃�L�O�8�� m�1�(�2x��8Ww�մ�hx�-e¬��I�(	,k�&�3~(���KV�zɛ�O9�Ej2�3=5�,u���ǽ^�*�|S��W������n3Ǌ�*���/r��g-Ɣ�AB�勧��o��C�U���59���0cæ����c����6���������2����|��s���W�s��x(��7�=SDI�U�Ӗ���Øf9û'��騢#�����]OR���yK��n7�^�B���M61�)�	��6j�Ev�N/�+��0��HvVz�$�=7%V.$�9K��	:QtN�g��m ��V���@���C�����"�vw[���{�����+0��Zl��y+ϝMO5^y�N�F�m#�ꪐ��[�S�ᬘ��=QM���PL
�K?\Gw�=]ͪ�<�q�-e+�W2��)-n/H`���qxY:��<7�&�a���_t��͊������4`,�25�UO�*7���x�[����N�{�<��1�o'������'�a��Y���J�qK�Z���v��x0Fn0Н��k=z�;�R���
��j$��~Qw�3�Y�gP��B�w|
�ѓ�k���f��`�_Ԃ���`�	���T�Z@{i��A��G��w=M�'�/C8�ȅŶ�ӆ�=���D���+ �a�#e]S�ƻ�I[�b?i��+5���{���w���葟9�g�����}�$��Lr��f��9Iǧ��9���HM��SǷ^W�Q�T�^#��w����v�a~�(����?ɂ�����F��2	�M���׃D^���������>gS򿳈�j:14��vm#&��<ż�W}��1��wbڱ�j�r����A rm*��P��+jt}�)L��:�!9�?AE븬n4�%7g��m�d��_db�����������?�����r*kЂ��b��L��g�L�^���=N�`��N�	�2���ތ��"Uu"��,t�v��&5ь�^a0�i���$���n�Gs}�MCI���7�FȠE��듽�0r��ο�k�k���w{��P,4����d�]�2���}����W7{c�Z[h�C
��+oh��3�RRQ�������5Yn���E"�$�^���n�ۚ����n�,&�:̕5�H�4�>��1��ayѮ>��)t��Z�sdZ�m#�sgس�l��R�����I<����0�^~�FBs�%�K��C�M70$b�����Uu�U�EO	�V}�C%�, �]�������� �?���7 6	�l�еU"�S�:٪s�̴(�oÈ�����Biat�2?����Y��Wlj7['��Xl�sš����s�j��t�*S�}?�� ����n��F��@�_ 4v��&��Vڸ��o֢[�C�?�"5��ڊ �UaT�ׯh���ʍO���wMb� ��Y�=��H����Nu���IҮ���8�O;���rf� _o��ϨiN2̻�qTVB
�稥���(x�M�q��PD��Kc$��҈$�������s�:�{A�w1q+Z��Q�qx�u4#���?�OgR��pO�2���~��*s`�H�{�b<-���pp�"�"�I���ǲ~^?`xރj9�K�z�mVW��w��>;f� ��Rn����&���o��<��N�����&�AhLo_@NE��@.H�G]�q�|ƙ�N���폎:AA.t�Sϛ���TKGu1j�����I����� �J�P���d0�F�=8o��P���7I�U���v���BgR�6G�%��}^� �x)��7\?���K�����=�7[V���ז��\��;+�����;�I���B}�aYӨ��1�qk\㹮7�\	!^1������yd�d�/��B���N���=_'9�ֿ��z��z��)�w�3,%��������^�8��@Mg���~"݇5-��@p���ħQ�E�)���/@Ec0��]��1�>�d�r���OԢ=��p�E{*`u����cRa8v2��	CL�~cT�Y�p���dY�# ����׆��V7p� ��;`���y��Po���n�tş=���-Ն�k�p䋎��o��urkMPk�����Ț/���s����y~�.�N�QA*81r@r_�^�me��i�I���o/��k�^�����%!�p�BY�׉FP�_eF�����@_�w�z�EwHH 6�#�ќ� kF_-=y@�4N�O�|
C4�L�4>�Ҟ����6��n�C���]�be��� �BM_�7�.���;����ó������+�l��[���?Rh���)�"�q3�x���Y�ۗ��pof��:9�������">��e������BZ���c��\��Y+y~�_�6����XV�gյ�VI��Yy(y��M<��(;�'!�Z�޴��kw��f�ߞ���7=��D�6]�qO���Nϰ���M �v���A�'��t��_�	ѓ�"ɖ:G'�9P�/�b���C�|6�`�O=GkѽG�	}؏�G��Kf��W��0[�xid^��iF
�� (�6�u~�}�^��f��|�`���"���C�7Pb�m�9�9��!>�����|}� $LP�����a�r)�R��g���l:���5?i��-tD"��2n���Ά)�	.	T�Q��8Cb���<��!�?��[�'����l��u"Y��{"��(kvK4�4�dC���_!��mǘi����Br%�¦�	�Vuѫ�+�m'��?>����yPV��؉D ��r�qw^U���z����B_AV���������,�-� �Ś���+uI�;RHP�����I	\��s-��`����k����� 3,�;r��c�׃;���Fb���,�������9�0]P��i<��<��{f�V�_�"�h���_���v[48�ɒļ�/,��k� �6N�Q���r����wy�4^�2��U��fTXh�ݝ���@�6U���q��а1��/-�,&�����Е�Y ��qoN��sh72���3�4��{�}HX�JP(�a/XR=E��[q�-ٚ	�#��Y:f¨|N�����Mo/9zoZ'$�#6��>��c�;N��Bd�܈�ӷ/�ZՕ��pܨH^|����x�:I�qϼ3ٺvn�DܭR����>�
�X��x������P�B�4Ara�|e�$�2����E�ʮ�Y$��'&��~��ѪB�������=Ͳ�$i�s����U�y�ͅ'Ә�t�# #|�$��#C��4,�5��.�
%��ޫni��M���:[����/	��D��\_�`w������+�/@�V��f�4��O�ANކ3$e�e�j=(`���tM��~{u��/�����6�a�+��#51P�K��z��g�r�~<"�(j�w�u[��g��pCy��ogi�{��Ndl^�����?�v��i�����{�7�c��_���)�ɓ�NLO��'�l�e�挰�-��zvux�S-��[��ۢ�06jV��V��	Q�E1;���i�$r|��gN��3]u��2Ҧ��[ܥ�M����K O{�5�����Ş�m�JO�w��(�u9Qa��u���&�� �k�<��׬����s�y���.��M��$���%F 趣��`u;b��^�3�� k��U�x>@~�yѴ���p��(����@%�"��kdDyoa��&K�K�n냰���h.��i0Ï��$����]���v,ط̓���O��Һ�z�Mc}p�8�luyP+��$ƍ�v@ho2a:�,}����o}�yq���H ����i�^ x&��u�/�O��twvvC�'��"�LF�w�H�d�Y�x|��@���*T|���I� *y2x��Z�������R��o?�1�����%���z�|p"��N ��M�,F���F1p�>C(�EPk��eM�z뫭^�����/���~w���ز� �X�L<�>��МMܼ�LQ=�9
�z�e�k�����aΚۘ�]xub6.䓚|r���4ۗ.7%�nO�u��U/�md��a�T�d	m����"�t��I3H��{�R�s�淌��=o-_����zj7�G�gAq�V�&qmE@���0���׾EHZ�Zl�|�c���`�s��xh9L�wv�\�qX��f�a��~U.��QTB����Q�;T~?���&����O;
����r��U5�\�7}�hU0l7�R����)c � ��� bV:m�#C�~٘i�#��w&_{d�T� _�^v�'�n�?��!C��V�	m6l��Av��_����.�-c�9�f����� &�l�JP�/I���+AF�+7��t�f����:$��P4�g������Y��y4�۟j7��0~13`������'Cq��~����>$�����T����Q�t�ţ�U;��Ǧ�W�O���", C�u�qi73��c�}m�uw���I�;���d�e��%	@������&UJKע��}:�t.�U����x}[��~v�?�)U2R������E��j���I���#ؖ&��?C�!�3K_����D�c8?�.� �P #t i;;I�l�B��'�2Җ�P��M�l����X�e�����#���Y���G�҇��o�0g��T���?����=�4���	�[1L;7�/��.��9U���}|��'�/6�'�4�2��/��&'��Ӹ�1m�U�*�Q�r��bC���������6U��C��f���>���4������;����k�2�끮���hi�&֩�c��'7P�k��s�P��s������+ԛь�xP��m$�	T��/v�*zHhc��9@���(������O���=���4��=ƣ��[�|O�N"�>���dцע�qP!58t��	�NVB�Bofo�����Y���}ٔb{�$`�.W�A�i)]�����w���PqC�L �y�y\�_83��f$!'6��"��K����F؟��7-��ߛ4�[]Θ����7~���q��j��.*�"	M*��辙R��k0�K�rڰ�������<����֬��i`&�՗�Pa�ғ�C���8{������%�WƟ@s������ڤ|x{���r��z��I�t4W�h�ꓘ�P=&�'�_?��bǜ(�\7��J�.6�˞���`�_:�fL�X�Qe��c{r�����m�̫����$ݴ����3��y9�����y#�Z�vfA�m�_E��^�A3��xC������k�s�(�S	�+�Kn�Z��D�_i �f3��~�!G�T�
�ڻ�4s���,(�AP0�e�Sj����4�K��U2	���4��A/�JB�O�>	(�$�����z\:'�j��7��ݗ9�T
�XP�E�K��� ������v�,�ϲ�G��ϋ��1�P�/��Ǒ�*�'�q��%��^���!V��M׻l�=�0���4��l�Q$�^Y{վES�vP�}j�S������z}vj���+t��L�z(�3���,|�Gy|��65x3@�ΓIA9	U��ߑG�V�bܕ��7#�R̭nZ�>[����fYaʚ$�&��,����,�$�����&||_��N��������cZ1��x;�x����Y12�:E~갻F[HX塀	���pHx?C��ș����S[`�)2�}�ݟ��aW���g�zG,�XZ��1�?6���lz��9���p��.W���*OI7x�IoZ�hЗ�e�>���i��Y�J��?`��]����$�LB
_��!�'��fE{���{����B���F����?�c![�E�5[���/~�0��!#�#|�l������f��q޵)c���o6��?���l�a;I��گ�H��l�Rn������j�Lx�y��<:21�{�]����C�:�E���p�	q�탚"\�V̼�����@��� P��9�
��)C8{��
� 4@{�@PS8W���n_�(��訹�fN+���55��|b)�����3D�|�AE��@g_}�v֭ܬ��+Z(ZW�8C��J/b�m׳\[�����l�}q�hJc0M痡���H2�,��\}��3�Jh�a������$�������)""�!|!��C�G��Z}(��M���1$x�zi�oA&����)Eo�	��{��{E\�Ѯ��LR��3���n�z�w=d$z��!7����i����^�j!��h'��E'�'�{��8��b������d�Npסm�H�s->�3WW���A���Q3m=��f]k�oK���P&}�
�N��^�ra`��؉"=�K
R�_���󴃛Q`m$jLI�a�e�f���ݘueN���K�_����m`��g$F���8(�q�l�~���s���M�V�ߖ��(7G:�+��|�pf� �)I�)i��#'�\��0�Z��q��v�kb��M�n���=��*��!�uu�q�.�f,i�g���2��ps��ͫ�.��O�z����]�w�5"/o��p��k?x��R�gX��ǵ4�G=��S���������0�������LJ ��ɭ]Uݯc�fp�EkOe�ې.�������]����M˷��Y7=�P��`�KR�9�׊�8�όw.8���+�&�𵲂|��҄�U�L�����n"N(#��S�����b��/9��O�����I�e�����5��<eqNy�p4�p!�#]�����K/��[��.�=��.��㫷X�6�\Y�)��xB�u��߅��v�x~�����>�[0Do7c|k�Wi�a�f�4���p̛��_����p��4I ��Iƶ����Y��UԨN�0F0�纟���aTWǧkzWD���2!��nB8n�S�6$Ek�z���[t&c!+>�K�-z�XC�4�sr$���k	�:�n��� JDmv�N�Lլ�[�kSO
'�։���Q7��bs���/_tU��=W*�������2_S66�HZ��o�m�iW<l�������*�b���*;}��Lk�r�K�lv��|ܚF�zL�+��J���\h��$O1<�S���F�s'���z}+	.ޥq����`��* j hcm������p��%h+/g=Cwմᕵ�>�Dv�w��b��D�,�����v������Hi�����ob����L�&z�G��EPr����l���̽XF�nZ^�׌z�oI��2JT�3*�n��2�i�G	w�thb������t7�R�R*����F�4i�A��;Χ�tN���q�p���K%���@]���uG�A.g��3O��k��30��5gC�׿�_��Z�\�8�$Q�+��(_Ҹs���M���^�}
hc"'G[�8���7�'$�[u��s�%�%�_��!�ó�ɻwQn����ߒ��2�7�e�lU��w(q_r~�n��p�tL`#!3a��_��<]��b��\��-ؾ���g�T�c�̶�X ��jYf��C����Q���\kA�����uv�H"�f^J�g���t�Ѻ�9��eQ%jj���G�2h��>&/[_="�
f�"dZ��r�磓X9}���D1���f�uXX���U�($ќh��ˢ��,��8��\�k�/����ts�mOy���H���_��P��"h��MǙB�B���ϙ[-R#ڬ�W�Ҍ_/-�U�b�ΞSiJcvX#�\�uj��vmQ��1���t�Բ�����q�(�<3���P/��fK�-Ne�iqsb�K�|ȫ�?�Ӕ:$��\��g��
�;8�X��j#+�%z��/�T-p����(�ZT�j�T�Y��`���@p����9B�HacЖ��1�����$��E�z��9���X��Q*�S�;���<���|�~��Hms�H�%y�,�C_�!�n���Xq�Y�ux�lL@M=������D)M�i������	�#B���m[����"G1gn�h>-���(�����M�oe9��l�n\��h����ti��5i�.C�̹��Ybq�N'��ӗ�N߻mx�r7?j^�5�I��lYMJ��<��B���y��u,`͈`O3�Ļ�	��H��E��Ia�
��k�(�# /�����#��^���j���y�Gu���VڬE��?�xu�ґ�s���c&�c`R^4���p�ԼW܁����?Q#�@���Z���0�&�z�5��G�'�/��8륭��(�e�#:g�U�0�+ز��\����LGE#/(C&���Al�'�0E��_W�ߵ����>lqj|x�`Y���K����lDX����l��2e�nm-�����o��*���g}��o�z����Yp�jo^���哦<N_���|�9�MIY�%�_D���6f"���H�c�%�����.<a�=��~����L�kD�gI=�۱a�#0n�zU�ddT{�t洐���~`�!X?J`.N	���T,?6R���H�𦼟qp�&�U�le5��lTu�b֦ȭ׮�0��i�2����}~[����V�������my�a�V��Xwe���#�\��m��F��Ԉ�4�i֙��K��[��H�|°M%�p8�֣�cc���ۢ`s�.���Mv4�P�Z�|�,�W>/n�x;x���*hUi�]���Ӝ�.!K�&�v$���ۊs$�-/C��PbqUR2�6�0�qf���dpmP[�j73�/'��2~ˎ&?z_ŰA�tr� ��b��.o�����/8�<uy��t��j8�x���(^�g�y�����/�$=L���X�ltWT��*ԸJ4�^����7���:T"�I�M��`q����z����V�B�ҕE��գ��8�Tdcaq㺨wY�?�t��g�)�/�,�{�(% �'��P�'��~v��bS�����2m|��1d`���8�]#
�V���c$i�D�y��c����/Տ�?�!f�<��Ɵ�ur�h������N]�I�5V���e/��bm�5{�E~�:Q q�{K�c�~�չo��`c3�lv�L����[j�����g�N�8[NX��H�����-�7{�,5� 1�8k�4Z�UiP-�*��A��=.��v�� ��	����U>����y?�6G��A1<�0���'�]����8�������ɜ���pxM|���ϣz���kQ�;Ņ�	�̄�3���I�p�3��b��i�ݱߝ4���n��=����ό�v�u��DK�ʪ�L�K�YsP�q� �������9����<�c:���o
�Qjf��X��}b�����X@�M���N��Ĩ�O����:-���
{S�ڻvV�<��k�ি[�T�y��2����X���8i��7�S)*�S	:��Qݵb�k H���3���ag�}P<����3���|�U��I���%����e�L�����:�����_�>خE?�O;�:{$^ꅆ���N�����I,��l�<� Z�?�B�
yV��(��U�ڊ��p�F�L��]�i�-?Z3�MwC����.6 ٲ�P�0�eZK%�S�V
�|f�=�7ۚ�9*{a0_�v��[h���z���R.Bx��U��>o�Dh��	G22s~K(W�L��R�k��f3�B���ԍE"{#����A0*�ɜj�n�+�kǕҏ��zs{"�XJ쌧�??ANTV�'l�f��>��HJG��1xQmv����#���j�iߣ �8m�@���r)O�`:�q� �T��
:{*������0Xr�%1˥
�j�~9�'36^M�;���]�EM\$BU J[��@�;Z��#��S�R�dG�R�k��Vs�Jwؤ����ı�:�;�4cF����)*�"L"�7n ��e�9��R�+��"� 1�И��-g��V���ɯ�K����p���y:������<o�<��(X��NS�O�S�h��·�.,��?}�m�Ay֜Î�ad+uܢ!�����I�d�ʎ�N�*�Y����ݷ��``�q�[߰��a�<���}�~.���X.���#=0ۈ�31W��E��2ИH�� l���^qn����]I���[���_�3@%��R����f���ѕ��%���LU��.�&�۫�і>`��?�����s:Y��X��
�ܫ�\��6y�����J�5g,�҈�ƴ%	��10���ֶ*������y��4#,F�5�KUP��/cU�p��H�Vu:ԁ�/��Lf�W�VʙDd�̗��;���=se�C��+�[3�s���3�8����3Q'�bY�/{&����G�R�R��ӽ���ׯ�Y.b=zf����_��
��,]n��0��9H���h�р�FE:=��ٛ����,ܱw�\Ѓ��n8`����E�L�#�g�j�~.������l>{���ͥ7$�Z�JqϻfS̹����0m�.�L����$��I����3<��π�M �R4i���<C �
e�l�BW	æ��,�!�{c3������7ѧ�5�� X2��tը	��=HDN��]NM������.�ܲP�=�4w���նљQz�Q{uߞ�ED@�o\�+�J�}UC���&���i��[oP9;����������� ��>Z:+�U����@��M�ۈ4���f���Q`,�q÷��m�Y���p��Y���ҥ��f��ڰ�'g���R���D����DK��y�]9�XULz�o��!�$�?.�0$���}�Qaԡ�v�T�������!��Z��P�{kzP@�ƴ�d�:���õ�W��P%��d�<uG�5�TXM�Z�4JR���f���D~e?ahK1������]��\t:cO��l���>c�| 7���G5XG��l|`�5�?W��e�ZP=��ō�&��*���꧉Fb@\wR�r\�[r�k��Լ(�5��o��S�l)}��d��j�z����,q�zv��tW�T+�M�SﭳT,�g��R�Q�O��<����]K��n}*:�о:�y	�#��_�+�Q):���m��<�3��;cԍCB_*�]�աdJ??_t �	�̽[[+�	{�3X��%*:�r��� ��N�	�@���n-�h�e/VA�ކ?O�
S��r���~�§Bwn{�fd7��^����֎(!]o>��Cw����pw���	���+���TO����Y@���K�|��gl��Z��'?^J��gV�K�3T��v��-f�c1O�|���:d���C�9��e�}��cu\�C�<����T
h��I�� o-R]��jFY�S�F��p�F��Y�9$~��/��se;�#|��v�8�մ_�
�LS�HZ�]:t���5��L�2	@�����S�3�#��vt��4�[q�A#���;2�w�XV�쒴��V5�rkY����Q��E��I9fO�t"�.��J�N�qY�Q�����;zV���7�y�ʓ�_�7;��Q<6�q���K7T�8�(��\RT�U���{��6Y��=pl�I���%>Z�澅Cz�ۂ�F��;WԤ���=���g��.ri?(�/κ���.����?�y;w(nZ��y&����x��r�}VJ�𗳿����=��÷Z�Π�}�ǅ�z���Wڵ�ӿ�q�1M�tIX�F���������"��/�ˈ�c.��ḯ��U�yp�݊��Ҡ8���t!/�t�	fP�Q���G�]�����Т2�r1�>��`ҧo�|��3W�uז9ş�dI�?�ҿKH�ѾV����u8�~��]����K��(uU��&�'�������TБE�K]��W���Y���{BW�'��"fD�����5Q֭qt��y��Q�qlэ3IN����r�����㠨�ܲ�d�w��qJ��R�?��"�������ݗ��p��k��x��>Ӄ��yY�����DN�n���ڜP_n��֧�o�����7y�X�"oO(nR�kTt�Z��'��Kw0��:�,��*�p�鮕��x��*��e*ƽ#ӿ^�Vw�S�Y��#�:V �����3Y�d�$v)3�{W�zЕ~�8p��S6��I��Ā�gEO��>s�ϓ��DK���׋ʘ�L�G�Y8M(�9��i3���V>^�٩N�H;ZGs��t��k鶯H9^F���4�����)����7y�fW�̵i�\d~���O�݁JD{�d�N�j4.�P�tA����E����4,�Ǳ	ٸ���I5�v���@-x���Uo�5�h��ݟ7�_��@C4����� `�����1�ՋU���<H���n��҂��
���ҹ�)֎���J�Hɒn�f�t|_���Ƃ�#�>�<�"l��t)�CDW�q�u���ΈY�c͢nd^Lގ���ȃ��*�O��νj���㫬��l>�f����	m ߔ�(Q*~�W��7?ɑ���k8���C�`��K�!�۟<=a�V��w���SO�R/v�;�)��N��;���Qf9	^i��Kw���t��YUW"�Y�~u�3�F��FG�k&4_�ҾM�Y[N�Ⱦ)�ɶZ�폐��9b�P�U�_���c�WSr���.����� �3��(�'��r��ëw�r�����{��6Չ`-	(��ˇ���� �2|����"1B�z��������ƻ�7��N�����1t���7�f��������b�f���x�OY��\�E�6�������w�D���;�l�u���� ��R����(!��t��"�l{��t�,r���%)��m�~Dg�V��]m���i#�h�#���-��� 3�5J��m�֯�Ԝ�%-&/����^g���K�y���>��Q "�Y֜�2��%,5�9����NJȅ���of�\N�
�����Y&�Ǿ���Dۘ�Szq���T?�cZ����ƹ꼴Qaor�M_+] l%F��cA��.Q���.k��:����>A_�x������n�k:t��<q�l��&���(�X�*|Bj>ٹ��lqW5��	�c��%=��%��W��I?�2�7Q�/5�9:-�i�Wf+��'��Ό�S;�.�� ��WiݺT�Q�Ju���yO)�{�>��������,%�uQW��nf\(��v�R��d����"�.r���	bR!�y���]���4�Ѓ�or�Oh��F8r��+[��kT�cd6Q�k���<�Z���༵O����3�	?$�4��)̨�%C��%�)�J4��x� ��b	�u�	ji�Y�$L�ոP�z�Zj	q�7��F��,�F's��(��M�_[�'�b/X,�z+�V
�6�{��Dli�I��QqF�M�U���)��]1�d��ÈߪY9D���+^T��|O����Qn�SP�Q��@_�u[}�����*�S�Nq��>ƽ��ն �Sp#((
�|,��`��?{"�x@2�%g�[�%��ປ�l�V^b̋��1��ӷ?}y�����<�	@����|�tI ��Y�	�C����w7���s�5B;��	7? �5SW�)k�|������VN�A:g��r�	��7������wK�'W7a�7����e��O�qM?���[
��Y��ے��ם ѻ�Hy����e&#:�׻ge 4��j��L#cV�DX�8������7)<O�z���e��t�?� �˷���A �����uB�e�_S��{I����tn4�7�������a�el6?���N�ۋ��a�VvWT��%��"��so�K�U��5�߮�i�_��>�YV$nԠ�{�^�����`;߮y'�Y���2])�c�D�S��.�MV�K����^-��]i�>X����P�t��0^���ԣ������֖���/ys��)�w�����e.�γ5L��g�X����Yf�ކ;¾%�QNs6�6C��OR�ߒ��c�Δc�z���$�~ՈY���}fӃ�_x���ߊc��q/�`��Q0��S�\�~���4Ɉ�k̟���l��C�n���ң�NRz���	�����}+.��x(���顶�Y�獐HaK�������-\:�G�O�C|n�?�/,m���0�c���v,��1￝	��>�:{�r��/�zL�u���4���SѱOt����L��' l#1�,�m�;!��'�r�,x�$�5����j��Ō/'��]�<�w'屽8m9�q{��xx����ݶNa�"�ޮ����)f�6r0tb�.��"S�4�@����	��r��=�#��C���sݟ�=o�kؒ&��@{/���������-��ʏ��L����Up��G�� �*�A8��E�F��=�C�	�a��8�>��S�W���rܸ<�l\�f��L�E�q�~6\�Mi�GcxX�ᴿ�at����~]��;���:g�m1F���VM�1I-�6_�l����S���t΃�V6���.��&R�j_Tg�'��̦��Ӧ�=o`�A�$.�^<\�@e�����8����2��~r�h�ᝩ�VZږ7��m�m�w��?Wd� �z�Ԗ>s~��Q��q�T9��ږ�~�3��B�f������@���%�T�O9���b����L-?�,hT/��FQ1F<��:xF���>��q/�O��r�y�sLOM�T�fWVL:*�7�Y�/����T
�FǗإQ�箢=�:ޖ�N��KB7�K��M �<eoIxh�MH��
/�$�h@����-��Z���9�����流��ʶ�����0�%�Տ����%���gsA����� 32��CvO�Z��y�y�j*u^F�D��s+;�t���$��ò�Jk��ބ$uQ�d"��)�4B����sn�qk>��^Q��� ��!��|��cJA��<��4���H���U쩇I��su�X�'˴���������f	̝B��y���x2F��^�VUi�t�Fu9������/�5��Tʯ-�;�u�^����L5ܺ#*�/���(i�ũTW��GN�B��� ���_MN�Db�<�(��^�u9�W�FF�ˢ�YQ�{މ��;�]W�U'�!|�پ�q*-�����(���˲��V�r����n��DV�"���"g�2Q��t�*{V�Ψ�t �{\�F��������Q9<렟��XF㮿�) <�  lV�V��Z5��U��M���f߲�^D�Qt,�>���b�qx�Rb�#
����Q���I�`�y�|jk�wn��l��u��%��RY)���
�%D�|�Z�H�����D�5��ګ���U�04���01KlΉj�V/!8������t���
c�|�6��f��ۼ���'�^�(���LL�ݏ�Xo��rf���23ln�㛏ʪb
Z�(�y�	&%���#��.2sRK�G[-�۵U��h��t�>��w�1N�?�Kl� yg��=V㬀�CN��5D���U�9RR���e`mp�~�]��&h������L�
�RMQt�.�gg���A����W ���0'�YT=�Q�L��{K��aE-s<q���!��7�ܫm�d��4���:[��d�8���D33F]���җ��Md�V7_����H��T=��σ2+$i�����[J�Z����u^H���p�����)���J�_�q1�urjOu�!���I�t��݀�6��1�ׯw��g�<4�̌�������$P0#,.B� 4�t)>��=�����8�0���L+��YO�y���3�j�f}r}.`2�o
�
7rV8����g�?����ۄ*�yr[���Q��>�Yu��e��+�.I��|���`#~��?0�)�ź���� �\��CH!��`5� ��\@�+��%��>ΰ��le+�N�����>�V��a�����TY���-�f��8�ʀ=�K������WE��UN�_�����7w?:�U�N5��&s�;��_&)��"C*�6nq��b���MC�u$�c\���h��(I �?�	ܚ�%��;�������L�»7@T�� �"q\A๒�� 2���n��>u1���Ї('\M�ڬ)j|��3Q���6��o0�"������V�ԉ�k�X� �@���Q�/9Y�'�.�Y͟��또��3����~?�KI�y8*q[�o�Z! l�_�Mf�?rA�uE-�TZ>�4H+ue�t�4u��P�ẉIN�����W^��1�ޏ!l�h�.���P�=?n�:��^�9����VNį0薕�����p�ϻ�4�*$�o��Rƽ6���T�-��|�QU$p��T[w�%�D�5���s����Rt}H�tSk2]������1H5�i�����"Zrb;p�U�K42*ˋ�/�<w����a��Ŵn����C�b���A�ɜ� ���c���!vSc��A�ÊJ������oaደƔZ�|$�h`"u�_@���� ��2Hlh\�R[|�:��mLd3�~��|�\RppH+$��7QF�'kk���0�C�(��S>�{�7ܘp�뫒l���I��C�qTW�S�P����!)R�Bq�*��|��׬��͋;(`x�lϹWκ�NJ���MM���ll��Ff<!6��!���|�.�k�"[7-6bȔ�V-���w��k��_���@h��}��k� J�
��thγ��M�Vؔ���RGI�����a�,��a2� �~жEb��*���Ҍ��Q�g�RV�'�!�X�6 �}�>|��>��N���/xh�ϛ[-�d�@Fd*3�[��+�24r�f �<��D%��MD���;��74�sջ8�c�"L�z�ɑ*=خ��2�4VU�0wtq|BY��S��VP񭾣���V�f��r2��/ts�+�pX�'�7�a��N;ApOyGԻds'uxU��i�L���1t�Ω.�q��r�Z��"$ /Lȗ!�p�BW<����k@�-+�}h�/T�X�~�9Gl���Fq�%�����j*��E��tl�H�.]�	H�@�'�"(Uzｆ 4E@@:��*�%������|��{��;.c0�!{�5�\�|�Z��yEH��!UL_'g�q*�W+���&�����i�rl����M,(��_�ݔU����.df�O����2 ��5�����x�Z��%�|����Υ�sk��Zο��CNz;m�tj�5�K�s��+Ⱥ��X`<n� L�鄯)�M�V��-V�}�f���볁�|�=��j)��9����/�Z��jh(UG�8�?ƣbQ��'Yr��!N�2��|�
�_��s�JW�U�rhXK$��ɡ3��cE��ᦱp����%M��N�J��N�$��?���9����К$h���
�W<K�;���q��d�b�ȕ�u/j�|��@��T�i]l�%{c��2(����Ku�L]�^TI�M,�p�$&�w�x��$�s��p|�O��gG�f���m�˳��a�手	\�hhE�rT��R�C�d�1r�dvdzkDĊGu
�-+m��u;�������<�m��57�P�ed���x��fM���F�z&��̫L��&�6��3��\9����	��Cb�-'����q�F�2��=�A ���2�=>|p{^>�L�µ�%��q��v�./�zZ׎�Fmh�;�Y�Ѻo`b���H��s�N!��y��W���a"���+�PY]�oE�ZU��_�m�`�G���Ōޠs<�E���P��i��;jD�� |! X]�Iu��6+�Ju��i�E�#y�t���}V?�{%-�C��p�n�:J��g2�IQ	�d+X�,���/���CQ]�o��roSu�E#P�*���_�8���၆��ǫ+� Zt�2b�T^'[��vo�!��8H���X���Q *�2W�/�V)���.����L�2'��>�?8-�a�z}f��;�&G��ᓺv�aGɶP�XvZ���G'��)�\���ƞ<�Bf�Y����>����p�a۞�r�`��h�E̪;Kz]_�`�<�����10���@��t�"2�Ƹ{6~'��_�B\�)�����*��4�q����j���f������T��2��8�?�Pe���I�����(3������9�'D?�q�c�[,f�?�`c6�&�&���W�3��s��̑�`�<�����7��Jq�vs�؝w?7�A$}LG��"_�I �z�N3�<}Iz��Bq?V���~V���N�?o;���������n^� h�!<\��qy9b��ڱݘp�J6Xyd	�X9=�tb�E�׆Ĝ���{"\����]*�~ˏ��u�B,�D�>9��k�9�@k��w�/����Qao>%�/�g�JoY��@���|z�� PS��0$���]���	6��^�\7���;<��kCr��ڟ�~�g����upt�3�w�8q���m�E�޳��WMc����AX�p���'{��c�k=%���[.��{qL^�y�ʴ�#���m�,�֪=8���0�!��ĥB��~�����˛clȍ����j+7}�B���U<�;4��W.n��'D�?�z�J�V�Ċ7�vƟ%��,�X:�����@��/���7��> ��6ZwOs�L[��d�H��vm4|
H�w��B���`@�NT;���>iB{����������7�,������0��ۿ86j������B���m�~D\/z�K�_�!r����y�׹�3�;2������Z�[G�0����[��?=��t�L�]_D֜,��[��-v�1X]�_��'w~��_�XR[���:��c�O�J(j�(����/׭foXo�R�ihѳ��=��b���b�e���K��e
%�]�O�E���͵[@�|�آ�/�B�-��/�`�7&���'7֪��ї��5X��gswρh΍�+#�jaY%;6Rd��5�)��+���&��Wt���BZ�t4���I)\lO>�o؏m\�Q�G�i����R
!cIq��3�&��Z�ᒀ(�`�Hc�pQ	:�n�E�T�׫{5!g���W��2����P�=��Lhҋ}j o�p��H�So�˺3̷����r�LI��1G�i�|@�ud��c-�5�����K�k1py�Am�-w�cd���h4,)%�`��C��>��HWqr\�XG����k݆s��E �VB�L�u�wr����ʡ,|�&Ľ�� ?��]����(c�����m�-7
 k�נ,B�-��6���RK���L
��B;G�N��A8-���9�LϪj	��ﳨ���N�=��#DHP͢qN����1��Ƚ�H�i���Jd�S�Q��~��c��e��UJ:QH#:���	>��S4��iq��vw��}	q�Ax�<S0��==�z9��!�C(�=w�k%��{���r0����\S�j}� ��LJG��Sf�G<�!SD�	}�����%ũ�׏�����e��e�3~9#h{�{��;
��SY��q����/�鴕���K�Lc+��7�+� a#0�T��5�}��J���B�i��\ɶ���2
��s�f���۵�U,cbkNv'��(}�R����fʯ�/�`d�kX2�X����XR�Vl��k~VG�>6 �sJ	��<K��+ՏE]�b��k������(���$9z=���Ja� �s�=*E�|�	���d�� ~���unDԂ�"�ؤ8'��CK��=���vc@�nb��U䘉_���0�Ʒ���9�=��q�
ǘ�T����/���A�<y�A7�%<��/�/z���j�-�oG�(��ƛ���<Ƒ��	�2���͂R�oIjJ	u D��L�� YW/j�&�*�8<j��E��<�R�'��|�_���:k����Y� �II��7�Z�?K�l�WBи����*�Xl��s"�o���M,X���y����5��$��4(p��\�Qхk��,�hb9&�m�pŋ����(ߞ�����uEx8�>��6h�+��Wʌ�c�)'��r@^Q�|����&��;�_��k(�cH����#�M��w�2����ɨ9��)��`�_.67�쏜ѧ��8 �J΄*�g���e	��E�hk�'҅	������X&!��J��=<F�adiD¦��b�[e�Ç8�x5��5����)��rܑ+@�/�T��~�6�X�٤wf��f�>�l���� �#D/;߁/ܘ_��p�m8߮! IO�<6�>T�v����Z #��k����ɺɋ�U��p!��2��q��Q�r�R�"$) #���ڬG1�%�1;^z�m��ϣlH�:�ä�"���g9���[�GէׇWO�|�8��"�h�i���]P��˟�h�n"ӫN����Ҳモۗ�ٝ���l��wYׅ�M���p������(X&����>1��[t��g�dU��o0^�ɋ17����dB!>Y������N��6Te	������ 2,�p~ge���-������Y������G�q��G�JOy_j%-Qkcf�nz4��@;��l\�ZX2�+ڇ쁽��W�+_�mu��:�1���t�N^�o^��W���s}���k�#����|���]���x�x���]1����\"������/���L�j�㼕We�{����������L��d{��O���i�@2/�y�#���AD����ٹ�a��`��(���ܮ���zBx��.�u��}%�p\~E
\������.�I�|�j��?hʽR26X�L=v�*�S]��U�� B �Ӱ���F��j"�t������5 c��O访� �,�t�>���A�~��#��)j�)2����WW�Q/����R�I�Z��ȅ�U(G]������`�ST�z2f��'(��]����80����YC�� S.L.�sJ Q��5}w�)i�,{"�K���Nhn5����A�5��/Y�۬�����ЕQ.��W��1�{�W1K�H��	�¶,R�΂G(���!�X���'���&~|
p�F�;O�d����O<��vW�(Z�Q���m��\��gz3��	�蔗�`89����7�-V��/\��_�mYBߤI�,���YK�r8���&P�	�;�((���!����uVmo@������pGd:��4�+k$FDJNZ���@ci�� ۊeN�����+���� �JP{�⠃Ѡ�Ap:� �9����]W>\���LlR1FA���'�vq�]ˊ}G��Q���b�f?u��q^Ho��Z-3�=`H������7�ܲ����9�t(��?�o嗅�����s�X1���冗߭����;��Q���XB~�}�C�� ���T��k�J*�J�o+1�Kr��##%�]��|�R�<m�͂�[m(��\�~\Y�Kղ�
�c�ۆ�^$�)�Z� a/(���s\�3؁j?~�iD#?bea�6-�@:�۵��0E�w�u\���<|6��n�tÇQZJ����~�J�%a5�H��攏��"�\��W�k�W#Ѫ�SB�U��	��##3�)
K:⠷2�ʵ�cﾊ(���)�8�w�XG��G����'ʴX,�'!E�+�~���lX�.J/�>�W�Ft�����]����4�ͼ?�_ ��|?�[x3����t�F��#5�A���z� 5m7�70p"�t�C,����bN���}<����l���Z�5����,i�G��l���A�t}F���>�M�����T��.�Rɸ[e�ƌI�϶ }���Y
�4}F�uV5ʜ
�5n�?!6)Ӊ�U�k��Ű9��=��T�`Z�r>r�bꔲ6z�~r �9o+`_����ۀ�ٓf)/�H��R(�Sv}�TO�>/B�!uawɬQ��N^��U`���&��_��V���=Ŧ�~Ϣ�����
i���e������ES�^�t��ba����3�+�|n��at+zЮ��I���5�Qݽ�'��-�|�p%0D�qǏ>���I��?t����U\�I�xL:=�d����)"h�L(2�c6�ف�)���Ƌ�}�K����+f����Ͱ1kp�����;!�����Ԭ��xI�O�:�~C�zW\�xo�)s!�8��H��e�3�;7韹)�����ʤ���zL����1wF��^X1����;�AD>��?������Ϋ�2قE�� ?���~�.�����?�C���4YI���C^E��=%���2����. �-���t��5��Δ9��:�x�ר@��&�f�"�?�)�z��#6T��u���m��"}O@���_E�;�yH�N��6ޢ����/&=�Z �C��֌��p��K����o)ݿ�����?T���y]9hl��/	�_+�牉5X,<q\�TN�v]�`W�y�/k3�yLD��8�}i����u�����Gc% ⑶����c0ʄ��7;32n����dM*7HI��*'����?l����^V�f��f�"%�4	1h��y��f�	 �Re� i�0��K_����6��r�
�7�T�*�ۯ�U����^��!�1�� �?��ތ���w��.���<f
��ݶЗ�L�;Ыy>Y>�T�.K���^V���"!��r����yr���Ʀ���N�Ţ��O:-���h0��b�z�s/8�w.(���2���y�_��ǘ��2����c^��1�G��r��_[� ���� ��ʎG�j!Y�s���!��!s����A�9�U��'��u�Սop\Z�]��-Ds��]R����M����桀f�d6����|�������*�։_ո-�yYw�K�xr��Up>��Z� ��:ǥ���~f�����p,���%�"�.����>,1���,=�_���94�W�W�˯��V9�K<�x��;J��{��ɨf�<ir������(��{�Mj� .�����(��W���np�,�_�G(�)�����!�SUp*����0ۺ��<�� ��z�nFk�����A��g_PYX�Zl�!���ڀ;�S��������Uե}$��U�1A������IL^�b�F��:~���Ҳ�qg�vw��x�S!�M�U+�J�a0�ݮoLU��	�����mÊ��ޕ��eQ��S�q˫փդ��kՈ;R��qb{א17�U���
�#ȱڳ��Ip���z�j�CD��Q��h��l�5�y1��m(�j��ݣ"B��K��q���Jy;Z���N�Uջnn��f0��N�)5�6�~�����z�˒�OY��8R� �������Xd�cS�zc��:4��%l^y+r`�����P�PlI�*��q�E�z�|$�<�N����Ƥ=len��kZX�`�
|��oI�R��v}�Ӂc?y5/��5��n���8��P>���cU��_������7YZ]_���cK4�ֺ>Գʦ��(�}T��2;D����Ԙ��t��n�Ն+�A��qH�	!���1�/Ҷ�KU���^]��X�{�n��uZ�~
��%lme꘭D�r�J5����(\:�iT��|�-�2O�}����͑��IM>�����(��]X|=��${�5\~$
ڰ�������-Ʈ�i�N)��\$�\5��=Ѳ}�&?�l;���HE�$��	`�f�G���UGmW	.q%��a�[��T����j��
��6;���f��雖\+��a-��\f��5d ��M,N{?(��w+\���Q\E�����'f���p��G����v���.7l�.�Veh;AZW�9CG�ߵ-n��-�����k�����:KD${-�X�W9{���K�,�[���
2����\�5k�e Q�j7Ӫ�r��Z�ui��t���\z��l  �:n<c��J��A34d�������q���AQB��tEu�D�Y������G;^˅�l޽��y���QuPA�N���<��b�/b�<�w/���'ea���-�>�t��������"���w2q�K�Қ���l�R$U�I!xv�W�O���?k��ylf5��zƤ{Y�����ʖ��7���=���[8!9�jbwa�n�c��
���n� ���f��'L+�j�Ӥ����~�XTN�R?��x��V�=!��C���k�J6���(��(�;e9Vp�
�(�DNB�~�X<��7M��äY�� �٥�:_��jcu{ӟ�4z�z-�wcD9�		V;���|�PX<X�%C�k��D��d�j�_TZ`vW;��i[#�N.�}�~��w)��
��m��-����D���7��W��q��0�m����*�Q����wJ�?��~��^�./���b�]>�{[�X���!,k�+�wӲ�зش���rG��}�C�"J�=�E0-�J2Ò�o$�ǒ玁�N>��n�&�j0.`�*;з�ٍSF�����L�$�3�6=Ӛ�9�)��9[�k�:�o/�|%���W���7���
�׆�أa�)?$��� /���b�]��:z���t�>��|���ؽ���#|��.���Dt��lS�3l�Ȍɼ�YT7��4�����iDd��!�O��O��sٟ�]e� e�|Ҙn�雰�}W�ŧ�m"��m:�R�V
�:�j�W=��銪�G-���Q[��҂z�8%�
oSw�$���f<��?C�>�E8O篱'��˒�}?S����БMc�����ԇa�UK<U�@`�:~-�F��3�\�o�+]���,����fVd���R4=���;���W���mI�n��ж�a��0y��X�Pe��
��.������HV����v�MBI�0���)f�����cr:���a��|g��Fl�PEz���ъ{o��[N鹶2I�E�g�>wBt3sS��p�X�֨8�U����4wn���ag�_�c���^�Yb^�J��h9�R.�InO(b}�jm��2��6�D����L��*�����h��a��U��у���0O�X/�c�Ҍ��"�J\������^�q�)�s͟��Za�.�ӡ������oK��g{�6G�ڝ�a<οF?�9=�q�nc��z LmD���`��;�t�╇FH1C)�j0���/�L92�����i����tMx�f[��so�Ȍi��c�S.�
q�i�{N#*2�*V2��9���gP;�PK�G����{�<��� ���zd �ᙴ0�Y>Ϋ�7R��{�u{pݽ�pe>�_6wﮈӲ�u^Y |",���~����V{=��n]O`/!!NN�tl�:��������A���@ֹwN��5"3���e�sK�M�z�S~�ݓ�Rx�2x���a��{�"(zJ���O�6���rV5ࣴ��G��h�����_�ia

�V�뛺��u��[Ӳ�a��Y��&�D�T���M�%�C��[���]T1*~=��צXe��G9�8r%��b��t���R��_)4q)�3��i��Q��� �&�x�� d² �Azn�)�LTՆ�i�p@&m/�����9�Kt�ZCli�^�Vt��"p�^"�M�b��`�� ��GAN����4��p�?T��n< ��\L|�zS0u��x{��>.�>�ΐ���$�����b�3�ߟi�B�3�6�|Cap���k�:�nIڏ�s���t��]�/�{�R��/ҳyx�2�]��VDL\l�IG�y���݁z�������\��0�J���~,�J7�p���8���l����^���5����������k�Zz/�28�۩����=��%,�)��C�����7u]�K�O�S���i��%/|yM��n�QE�}���@^e8�]��<��1M���P'ݪ٭�2%Q�����Rv�t��ҙ;��!�:c9k�cl3��U2,\�������j�����~�W�0�ގ�'�	r?��T��:���>�:��q͸���`��:'�_lݼ���#玑��m�\\�6?qQj"+`����8��߸�b5��ޮ#C(<C�[�-S��nmׁV��]�i��u���Wiuv�|��TFK^��[��7��qxy���Ǚ�H3CV�������oq����I�x�jV��>Xԋ�zI���j�ON�֫8#�e��)��Ɯ�ZFQ�k�z���^�#�|��UA(-�sm�� �4�� ���õ��a!:�v	 O�J�#�ׇˏs�mMvV��EO���*��H�ߖ�MF{;�������ͪ�dCkg���"c�7�#Þ?���M��w�a%%lǉ= =���v>�N- 2���I����`�Zp�ͻ���"{��S����j*��a��߾*��-������dk�tޥ�B�
���)v>=��� ����S�yZ�x�>"(q��AD7�{s_n�-�D��*�c�qE���wt��w�3`�*��;�=��$�p0��,�����RlF;9YȽ1�\S��01���a3��������T��ۣ�.�� ]����AK��RlSK�Ze4��}�7JF��Y����?Hy��jk�	��&>���=>^�j��ȴ%L�;5��!1>$�f	]������ݖlw�7�\d�3� h��VwG� EF�\ݫ��.��~"Q�9��/M�k+��F\��˧crz=5\�?=ԙk`Dxf��}��
�B��^�������+�w=Q�a�nEr�
	Ͳt�֤� �n�?���ܧJ��q�8�r�60`�H�(��7L�	�-;F"�"�(�ζ�s�ؗN�ؠ>���+l�<u�l���{�̻c��R{}^�8�{w�=����zJ �����w�O�L��a�M9�3q������\�߬���Y&U9nm�rq���7;�>��ο2)LW<�7f��{֛K�]����R�*>PI��p��v�6VV���=2��� % ,˙��WЪ��)��B�Ցn�.�u"S�C���])�_�](R�f����
w�����-�$�5�5�`Y	 �w�GMN�'��,]}oq�0�u�o��\���Yh#8dh.9$}���4ډلE@�����ˣq�cӈ8ے8�=�^f�����e��t����}�l_?>�9�y��^��[���v���ŗ3����VW:*h��^�v�OQ��m�������M&��ueߓF\����y���4�A1�о]�j]�X���W��	MP>u3�ПV�(5	���}��^q.�n�M���X2yn^/W���(�OL�`=�*)��MkOP���m <�/9�.�^;o}��~����ФM��C��Y�'�rd�]hՌ���잞�q*���@ӹ��������A��%��*�\��hm{�rD����f�qKE�
&jV:��k7|4�O�_�١�N�g�t��>��$f=^���)���dj7w����k${���5�lyN�5t:[��4q��%_n ��j��_��y(�\$���:C?|�F�RL3j�3ɋ 3�y�� ~F�A"
@��n�Dk�|������m�:�0�FG7ax˘�fJK����^vd�^��.����>��3}�1�y0-�����XAB`�S�:��T[�/�A!�C3����zr,����Ӈ�|C���0� ��%R��O�}]:g	f����Uۛjb7�5;Dg�q���d�����*rg�x��z�	_���{%�$1qe��i=��k��&�{9��<~1���#S�{�z�J���k;+�����/��1Z�]: ��S���zm��V�(w{���~wo���M5S�Z	!�NŁ����.��B����5Ý�|��?�iaj�Ay�%78�C���=_�H���ϱ�5�5�}��	����E��I򽿴���$�������S��P�^c�|?�C�Oz}4e��0�U�?����LUd�	�xJH1é��I����X���%�g��2]��1q������0���Y��`���M�׼�D��O��4����.QF¾v��GR�:���3�s����z0�g���k_ � lq�G��s%I&�:��Gm��c�DX��ua�m�7�a�=<����y���9��Ɏe��sx���|Z:���St���G��=�W���� B:�Ӿ���23��A��߈�@p��=g����x����R�)��{!�Փ&~�I�*4B� dl����0I�}���1'��"�Y-�c$I/�����7˔D̝²��ˋ�=jET>k&*eԱLS�A����l���w9ٸy9��h�Wzĭo��p0�2�R��������*�����9H/���z�~�^�}7��h-���L12�y2� �r��D���5�� �2�4��/�U�k�����b#KS��V�s�
����N�R��{/'+�f �y{פ;@z�Ze{d�{�&6{������\Xw�=ݑ]����_��z�͆+>ͷ���q�ə�p�� oM�+k�yl��K��2]��2��R��P��.�aK�e�L��h�i�<��y]��p|�4[̈ajR���a���ŅKd���zG7P.5��Ê��+=�u#K��+�)d&i�NP�P!�;:�&vj�nGE,�Gǫ=�0�n{��@�(��/��&x7?5�?�O�ִ�-]���|bZ��+�ھ�;�#�fF��0�2���!��)�zm���w��M���
);�=���Oc���b�fn?|^l�9�au���5z��P&��W�4q�Q|�>�NF ��>�v�5
�2_�b����7�_L�n`�O�VGk?C�b�/Wa�lޘ�W��!���Y�y��:�����,��E�j7�M!�^��Sg�X�rA��Ώ��>�ܩ.�U�:�Ȭ9(@�ϑ�99�����ޑW�bb\��/ʷ�6�/�ILڀ�*�����]+}|f�VK�+�ɲ�jd��Jم�j�#v�L�+�ae'�G�nu�2%��d�&j��:�2O�v�R�u lϸj�zH��DN�z����y�c���q�* _�(��SS�sG�R��!�P/E�W�\-҃��_)W��fpM����4:u��ma ��_'�ҁ����7Zh���@��Ƨ�7q�av�3܎�����P�._P��.]'l0"b�z�R�PŖ0'>�m�[�i�b����(x�6p�U:��ɠ:��s>��� �L_-���u=)���`[�ك=݃��O6���/�f�۲����(��x_j����Ō���C�X�ꀲ�^�`���.P�����2���'�`�!���� ����4%l��e%��f���6��u�	M�w>ݯ�-g�=j�Ds�%3��=�u���m}O�T�[��-V�꧶'|y x.�~E��]J�s��PMD��߲p��ſ=c
tA6\@�dnG����fzlǼ�	�.�Y�\?1E���N=�w�Ԥ�?ь�m��S^*W�T�-�t5Jed���FKBg~�]���E�#�)�jO����E�b��%r�z6�M�	�"m��g�n+\/Q:Xz�4�N����K&�Ȥ��(	���PS���E��k����I��ŔJq�C�h�&C�d����L�1p���,��������.Q�N�M�u6��;Su�~�� �O �Κg�~���`����A��v2�S�R��ks�0wp���n��c �J�a+KU/_)\#8a�b�a��}���������p��;�1qh��dgvx�v�����3�� }_r�k�p(�D7�(N�� t$�������_"�̵�Vk�Àܜdx�Q������p��Z�C� ������-���%�H��`�	�SL���N/���o���f�"ǩ�Zv�R�@��~׫H�עjvT\��ē"�'�@��3i�_+�W�C���^,`�|9C����n��d�kŽ����-.Qx��cK�!��Q*�:�Ս����������Ύ]���K��C�g����7��ˋ��K��n8�� ��n,ɯ��˫�{'���܆�m����nqu���h݂��M�̢;1e��g���e���c�O�ѻK�S���E����d"��+Uݾ(8[���Z�J"sf5��t8|$Α�P��Q�M/Sn�.���F��h��zG'�8��'	;��\+���ȡ�˛��`��]]�sA���0S�?%!�u�����/�����!E�۵�n��5�1�5�T��07���XB�xMS��󳢈����!4_o��j�#&�Xt���q���Z��3|�=³�=���K��n5e����K�Ϝ�̎�T�l.)B���`�f�]��F�կ\B[oģ�h ����ٜ�X&� ��%7��YF���:ٮ��Y����N��k�Ƚ�t�{L���.i�e��1X�^��Zb{�����G���p�	E�z���-'�	ɻ�s��+��,P��rW}��9=Y��R��HX�!�#
�o(�Їnб�)�(�ٷ��[�ݘtT	wi�U9�qŭO�� ����^�B� DY���5g�c>�=z����'�qD�̶��Y�ĸc���#��.u@B�QL��1P	w�����,��R͍<����2�Z�P!Ł7(bә^���7ho�����9�Ⱦ	)��``Z&���'bU���U�?`ߘĶcٯ�� U��+��dz�v@g7<�"�k@�p���	�ot�M����VOes b��Ҷ�l75����.�2��ruQ9�1�^�A�g�9�[��R�pumB����ˬ:�x�+�"�豥�W�r3O/&�lZ�a(	\7+bT�j�܈�^�����ax�l`�PV_,/��*���M���
dkWV���M;^?[\��ԫ���͚��57ˁ�$��6qC]�K � H�v��9Y@PW�����/�����{���*��8\ֆ���J9],Mt,�VK��2)��qƴ����CV]]g�r�k�v'�HSok����y�jH�"�>U���s&L��n �֡�$+��rBŕcz�ᴴ�N6�Ӗ3���HjrI\|n�1|�$nq�Mkh�\�����^>M�JS���$Uli�9M��s;���I�tM"z��Uv��1)#�T!Pa���P�i�{D=�/<b���F �y��dB��C 9�x��v��'҈n����g��ن���gXc���_��@�i��3��f�V��t����}�d� ?���[�a������|��%Ү�1�Z�1-��m+��	)w���ѹ�c��Y��)�ӱ�.�k��w�[��zѠ���*X�4b���Z� �;9�h�C�v����Q�pE:l�𢦍�]��=�/-v�O�����{Z�f-ma�g�xg�8��c���keژp��d�f�h��{6~�`��P1S|V�n����
։�Z��"�g��P���;�^��t�dԈm���vU��y7�%�ޮm�6�[�>^z>���]�S'O�υ��g��/o�4�s���\�Q�mYP��`}-���G^ZOO!z>`n����)"���]Z�$�y�%e�P,ܻ^]�rݮF.�ʈs����I�+��^U	YK��g�� }=��7t!/�L�;nD�|I�ȓ �Ý�خsLv9�9]?" ����]���A�@���C[�;�D��?���,�����Қ���7�HQ(�2�v��x�6.���-�2��t�Sq29����T
�I����g��00v�|w��oO��ys#��'���aGg�8h�+( ���ލ�{'{K��U��:4�x���n{�AWp��_�Ѯ��)��� 
�p�љnd���eѴÎ��1�grx��a�95ĭ�r�Y�*Τ+Y��u�G���|	��0�/W�t�(>�ڟ���9�a6�U��`��"w':�S٦s���/sQ�������)�jV_v� �^ *�u�!�a�Wb�HNC�O �p�=�Lð�S��~���{G��Zdk�U���a�����ח�h�$ⷞW56���
�i�fuȥi��N���}fe���v (��������)GX�d�s���yQ� lIA��Md���r�!����#;��乆�!n��.c+n�m�Uŏپ��t��\��׌С���N�7�%u"t��@eD��
M���] �����i��.�9@�-�Z��T�f �U�����&(L�Lu۾��������jy�
Z=�Y,��D�.���Y֊���2�?���6i��E��-G��Z���e+߻L��la�Җ{2�%�2.z�gB�X�b��ou)�'��R�m^���aoJ�4�a���27�ǅ{ǳ.7g9Yèt�F�)�6��sڦje.��24!j��w��z<QF�t?�HY�3$%�xqVwY��eA���r�q�:�yn�4�֘(>�� �Ȧ�9�=�#R�z*��(�l#�������Y�W���s��0�۫�nب`�e	f��m`���f ��p���ߏ���(P�jr��|�>���0xt���m�age�{�>�#7"vG��a�#K� ��sr����2�$��6���z���1 �:��@�xn�]�7}��/>��w{h�-�:n=�IBs�8u��[�9����]M7W�5�����)�Sq4)=�S!��b�'�5�����r��+=�|r#R�実���z���U*�ճ\�*�--����b���^��)��e�SnO�:�ŔQb D�33�Q�]W�)G���Ms��
�b��\���#����5�'b�I�Ӊ=�V���/���%�,��|��_@��*S�H�oi��n�!:8:�~����6�b0Ń��>s§?����#�-��hu[���/*�v趡�Gg9a��"|�|�ZI����,0��s�
�L]��G���M���gىW���!�&��~�"��Ͽs��4u�r���qt�ɕ��bRT�#n���	5��D��݄��;Lݥ�M���E_%��.����V��m�\a�o���sw��J�>N���X�/Qj\0CQ�_/zևo�8z��Wa�~EЫ�ݝ���R4~������3��x��s3K̮�y��irD>�bә	ir�!�M����
{��/E6.S"y]h��V�W`�|��~o0�a�/���jK�6b9z��&�v��B]<Ƀ�}�Kd\փǈk?��֥��[Ș�I�"�<��ˊ�'u+H%�4$-l��ֺo��3-�ንy.B��&0������Ԥ�Ll����]����_r�Y�|B�HS�?�Y�����iR�D�_x�Ű����K�7�R�%�bp[~֚��I'i�.�] ƽ-�t�Ha����%�Vdzt,�]C��՝J*��2p�>��\P{���^���v�~Lsc����۫�2W�-n=r�z��0�+�=���D@�\�`;���0��"�u��,���A�/$� � �mh���d�c�Q��e��O�p��f����2�_Qh��t��H@��-���nSy�E�Uί�-��ڐ̶�n~j���ސ�;��"�k&xͪ@�!!wC�Ȳ��[' �d�?lb�޵֩>=`8� h:��J���H����~j��7�T�l~5T!8`G?UY@�\0OQ���˻�{r��2=(��D�
Ba��[j�	�uKO�mSDW�8i{�M�q�I�j�
��B�Vk����������H��[4�\8jE%V@Ɔ!V���ٖWD�<ʵ��Y�zr��to1���dw�9y���j�E<�_��sFEy�O:�^L�h����	M��ír�:C�P���a��.�`O3��ϴ�E����,B��ۼ�}����,_��|mc��zL�v��F����5�)k�G$g���E����#����L,J��#����eO4������"��G������4m��;�[h[8�D_�4�d�鑱������;Ǟ�a��=��/��u����V��mI�E'dt��V�+����}��T��_���C�V�Ԃ&��m��#$���GGל�_%���˺T��ڽ�vnz�/~�:�n=��(���5�0���
���͝1u�xY�0��k?�侉U�u�Ι��r�F�׼����>V��m2H1V�8����x]���g�J�͊F ���d�y��.d(��·�l��;���i�=��]�to�^�/����%����,�s�m�.�ن�{��:˒-~V�>07#t{ｧ��A�}�Z�p����ص���X�I�G!�M����@LZ��*�&���r������;���	|�#��O�@O�ǒ�_L}T[�7�tw�4HJ7������tw#%%�t7<tJwwwI�7��}�߬�r1>̜���_�bT1��J@j���8c��hxC�]7���-צyx�r��ZD�L/?Xܼ|�3^�M�^͌�����,�b�a����)���Z	<_�g�\3�go�����@+��2 "���0�l����\@�#��fa��MJ��ӳG$]�L��ZKc�֮��?��#i��8��T����/��˷i~L�]9����?,�H$���V��˺
�׿P[H�7���Q��Ǟ����̯N�zA7�r@;Ae%�����_�kߟA�Ϯ���� ��V�v��0���X
� �Zމ��[�j)���zJ�:
�t��P
�b�RP��V}9Y���·��cT�|�,���늂�K���������X��ءx� �>�k�<��)aCW�iT���l�����ŎY�}����O2D��(���v]�Z�hY��p�Hm�ah�S�$"dR?��;�˛֡	�㦔�S)�}y�_)���ʤ�뜲~��k��L���z�7F4��D��D�?�	rU�PNoU���㦂B�A|٩.��A;Yd"���*�U}?��'"ȓ��LuX���9�X!8НH�~�4�ֳO��,l3��ÑC�j���HI�y��)�Qƺ"J�z/���Q��8ee��v4S�=o���:�ˣ����e��y�6ۇչү�ö�]�B��K%���?�[��T�	<���W��h�7��+~�����)oV3RZT��y�u���/�ʮ�S0�v��f���=�SEʼ���9b�u�
[���aJ���(�ǗM��hn���3�9�:k�\�m����%��Yj�;A��4�X0C~�h�7�S�������R0����N��C<�E~3�Gy������g�P"�zlU�����_;�KhW�`��L���#t|Eo�l=���]]��|�TX~������g��*��6/c_3����To�R�9���Ȓ��se�w��y�\�C�ݯ�N�-�w��ߧ�c���@)hJ����?m'�[����R�y�����;�n��������r�fI���V<X1��Ŵ�{���-�����(��<y���iJ�l!�Ѳl:��W������s@^��Ji8�xQJOX��!���v��(��wCK$`�j,�.Wsˠ����B��<�/'�+���I��tm��H��ן+��Y��\��������u�8���s��grT� �:b$/1����|v�������Mu\��D&nx��}�M�>iZJ+i4_O����@�5�եph"��bg�!2��ΰ����P��d:
�*�X8���n��B�C3h?���oq�X6�i�Ti\�wÃ61wM�;�y����Z�{�F�tu`�wN]�P��O��_��K�Q܂���"UUE��JR�I��Ι>a!�����<$	�ו�p����?�a�@v3��e�v��Q��&s�!��:����ǌ����ۋ�@�t\���p��|h;t��7\��3��?�����3�t�?%V�P. ���������Ae2M#�8\E*a1W30vQWL�oC5*�p���!w��'���4cV��[Kr�>��˦�a�C]fM���6C�*Fnph�Q�,`iX������s��⧧���/r��9 i̺#q�8	��c�J������˙��THrvU`�����u]G.tG��o/ؙ�tQW�w�$��E�������};K�;h�r�0�Kp[���$|E��`�Ԭ��D������n���m�r	,f�
-��9ۦ7���C�Z����#ID��o@v������w���_�s�b��Q��rF�˦_����=1���+k�u�.<�<�b��{�Z�N>q`Im�1�������w�N�������c�)�0GgO�M������ANRLc>N�7�dK�U�w^ u����#7ҝ�	l��'�c���6p<�������o6%�ͨOA�������T�8��6Tv*�\�����r�'�=�]�C'������fj�4eQ��������� �'i��y�������Ҿ@�K9ݔ�K��c��R��_Z=D����$�f�~��&Q�����C�#FH���b�#�5�\��u"vF�+[�?ar�Q�Ճ߭�0�8{^֩���^W���L&�E3v�͇�;1����Dm��ܗ���n��%�m���7�����lA��Ҩ-�6g7D&���4��$��&V �a^�P-&�8������$$��]�����j9����r��RV���@�� �aJe�᩽G����J ���^�/�E����s�Y��;��@����3�3xD�c��j�����4�4�����4���)ُ[Xt,�^c�������=�4���1e#K�U�ߥ���)Ȳ)�UU��:?�������"���f�:�Xeq�Ryۯ��s��{gJGĸE`?ᴭ�@,�����������7�>U6�<M�7o�<��
=����������@(���7t�=߄���ڡػw�;h��O�&th��-̨����c����aGQX�#"��SF�N<�+��b���yp��P!�<~Y�L�`Ng�;�Z�o&��$�9p^���f]54\WR��q�>}��qUi�@o7�0��O��N:�d���x�l��X�j����5}�.����S<�7^�&}��P�=�a�F^=�����T�a��m��o�l����/�F$g �=�z�� ����*�_�ߎ��9��F�dQ����afa�,�F1��ȍ��v"~|V.�&�_��a�&8(����9t^��g�G�f��e��pd�c��r-�'dӝ��^{1#�,�y)�W�o�4To/����C��	����u7~���ۉ!�N��+��s��s5!�4S��`���ǯ~a�T�"��_��3�ĝX�I@��s�R7����#��`�L'�xb����x�bfS�E��cF0�������9��9�S��&��>��xs@C�"��d���Y�V�����]:�wd�6�X��g�w���)q�{��^u7Ja��E���{:�lr��1�}�wF�q �>��=y8�,j{��t�oo�g[��$_Rԟ4z5��(��T��6�Hd?��!�W/��qf	R��mQ�?�Ͽ�	���x��x;�q�g�r��䣓���֮ܒ	�Ue���:I	�1�SX��h�+�M"���9�F"��[D`��%�%$N�e��[�n+�w3���ug���w��!�ͣ����/eCƗ��S�iM��N)�³O�h5��48��Q>G��C=6�Е�0�����t������9�Z��ݝ_���h$�A�R%F4�^&�ǻz�I��kc��+�'��$i��c]ܳy#���TW(U{��f�� V��-��5�b�̘k[}ä�]a�ry��RP�Hy��ﳩ���:D����-�оr�΢6�$BC��DȊ�aG�x�����`������	��I��D>Ƿ
��^م�M�VQc��i�|��B#w2�d��xX#+�)?�ݖ˩N�A�[ȑ	x;�N}�m��{����|�hss�1+=��Ń��Ju0�����#[�%���+�Ϟ�}��Dϵ�)Z���DQ0�\�M���"F[,x;���ԓB�q��z��}�� o:��Ԡ�s���~q��U��R𞝣�>�������&!Rf\y5� \�+UX���|]q�*��E[�LH��4�\H�n�ꡏ�]�T0�W:������䟇�<mڇԽQ{��+ _�(Q�W�G���>%E8`�]Ȃ���<��LJۉ@���q�BQ;V:�O�%���S�^��m�z=Z�W(z�)���c.�gՁ��jȁі���Y"E!��S� <Ꮜ����ó��$Y�!�(vⲉrV���4���(���0@��=y"�sY���j*��-'��ԃߓ`�w����Gn�]����{¼�W	$JcW�O0����jaeN����e��յ��[�����[6�[!�'$h�
���;���X������4(�\N�`1�v��E�����Qp^Y#їm�[�\�Q��h��V��&V*�=��[�~	D_^-WhK̵͜�X�d��\���Ջ�{��;>ߏ�MX��K��uCg}~.���o��)��ZnO�}>��<�Ǚ��:�^���P��+{k����x��sQVh5�S$Z�a�� FtJC����tN�ǧ��̍<��
d�{���A8E����M�Q�uh�B:&�MN��DE^���M�=����s����괭���q�o$΅{	L�;	��e��!��F�r�ϝ��kn�&4g}پ���Mh2���P����@5�$���9i���� *�;%|�A���Dե�C=پˎ�۝s��.&��^1��%�Yp��S��ͯ��Ci���%(� Ʌ(�?H�W��D��I��������G��;C��D�1qJL����f'�Uk�&��=�tu��W���P'+Y��w��zF�D�KH�C'n� "�$�!�|dX! r�FQ�MN'��c)��Ʈٖ�y��K*�������:�j�l�I��xT���˄�N �#,�=���E�j�z_}x�9ٖ�n��!5���j��D�s������V�@(]"�{�~:-*�030q�}v��Ts��_�D�U�4��=e8�`YPP�Ȅ���'�ߝ��u=�>�"S;�g�4[�t������}�ӝ}�y���#��ۮ���A�m$�oʟT�ZPG�O]-��"f(]p�Q��[�u�������j��!w�g�<$7�:F��ܬc�jqi�L�˓ ԕS���U@M��'��2n�i;�r6�6����)�񹞍��-�T����{�����:zzT¼o�,�l}��
i�O��z�ڀ�#�N>�ɟ��T���sH�ʦ�C>>٪=�եKZQ}�܌5j�q�_�	����ׯ�y��Q]"uV{ϔ��|��=��b��=v���YKSb���F��O��.����d�U׏Q��B�x"�z^�OC��������K�c�n�x�Xĺ�3�P��h��'��4,��â�NK4�eVc��<��.#�L���H����[�[�Q&��L]k�d�x&�����}�~6�sv1"xF��
}��u�#���aE��q�6��'y 9�	r�X�	�9���~Cn�
����(��(����;�k �ʈL�V��9~����h	f$�r;�2��Q���mg3�-�nP��Uß_l5;�:��HP�K�H�Bq�R�	��
z����1*��FwS ��n�N_Q����w�~�mmYsP�濛��p��t�
�WFb�>��.:@8`�ױ����|�Tmc7?�|n�qT�xį�</�p�>�bF�x+������"����.�[x��¬��⿉F�����&-��%ҝmu� R��A,C����ɪ�4B8�0��V.���sT��]�����(�T���Z	SŽΟ��18�jy�dooҋ�^�R�"��t�̪��,ߞ�Ia�rb:e��Z�8M��\x��g�o�p���^�"�����Gx�/���`1h���^č2i�Лً�!�aG���;��\���ɞȞk��s�R��#�9,���!$���S-�w��3(Gl�w�����F��jX�r��zF$�nI�.�uD�hZt,:��K�[��d�Ǽ��9���ی�;Ô�=$܌=7�E�_��̂Wv���D������=�^-��$�;�*d�,b��m�'V�s�X�ƿ�n���0~]�ד�é�}��{�Ni�c��
r��6��4��Tk�nA6�
J����9��M�gQ����Wo���s�6��a�	�[3�Fo������#7N�{�x$zx����#�z�Q	&zm

v�O<7��)d��T��G��M���ӆ�$�n�T\$}�E$���7P�hZ�5��_f2�|�y�(�Ȥ��fG��/�#/��������:�H��Y^�t��ہ���Y�l���#��<e���G����½aREH����V^���\��R}�����ZH��ŕ�d��8�Ǌ'��tSjiv��ͯ+�+I�7�jk�0Ԕ�րJo�M#�����Ȼ��7T V�ض����n��+�j6+K���v���toL�t$�#����:	�ayy�̩���v�����S����VXԩ�n�A�ZV|�ጆ�|��%���7jG�Q��-�����Z�]�7��#x�D�ǈ�z����+�gS�l��m\x��63w���n����Ɔ��% ����I	��5
�;�1��1N�(P�j'n��[��&�؜�0�9~�P+˓���g��ӡ(XoW��'
$9��'WZy���.�$�O�"ë����bf��_^���(_�mu5�}߃���#R�@0ǂ.��S����;u;{�yA�Ē�v���Y�b�^q�n�:V��w�������&�#/'�2[g�򢳗�V�/��� N �|.!+�l2��C8�
~w_��E���V!b��B�������g���J���+v
L@D��!�O6��'#�g֚�@�gQx�w{$����?8���
��c��\�rƵRG�֋����;�������~(��>@��T�!Q-��A/\]����]���ѥXL����-�&�pPE�Vahh��a�x���eZD��a_�夺{rq�D��&9/
Mq*V8_A���3�'�?��FV���ͅP�d�7�:�D# ����E���Y��J�#Y���c':<~��Zu��oiU�"��B8��I_Eʺ��t�y6��p�W���O��KL[���~P�  )~+�˫�'����S||��1)!!ެ�5��-�.J3ݟ�-(ѫ8���P?����y��k<�����:�����x<��%�;G�Щ!��Z�0�R�-�q��Ky ���qa��5�DU�9���:�yg$b�`k�/�#�	^%-X�v��X��2�s��?���a-~�<���5�Y�u�c�P��Is�J��8I�h�|��03�����N���E���:�F�D��������CܐD�$�]4�|b���"7���f怖@�S���$L��壒���.�:� A��Nnt�y�(�s�j�c��~?�U^������xSH금��DC�-)� vܼ� �4��Q��*�x� _�BV:�?=�	��]9�����;f�x[�(����\�[�$�.e5����aַ�;����@�ij�۩�K^G� �˪�3ֿ}4���dG�G�j��R���Xh�&�oG�i�3DO2օ#�0�m1N ��x������ǓTbs��QN|���5�m��ѹ���##3�)$���V�_����x�s]5��w���w;s�p��s�U��k+��tSB��fHִ3|��-c��t���wC���nKÅ�{8
��گ�4��� S�k����@�P�i)�uF�53�]���v��CM]�j,����.����� |4����_��M�)>���-��N2%�!�x'�?�ct:,�/�'�����'���2/���b^�rx���J���#���WJ�0~�y:��?6/�|��*M����j�FD�s��o2)YP��& iA~�/�o޺�� ?���Z3�1KAJ5����Qδ�TJ [ROP���*L|��Co�E��r�������I�8��M�O�j�_/�� '���N�խ݆�η���8T.������\eGd�,�Z��g��^=��|�=�E�7}�Lo �%r���Btu��Է�s����������%κl�zo��!�,��V��xZ�ͻ�w��T��>=
��z�i�5�nr:�nfv淚F8l`��84-�g��mx�?Q��i���_�edao��1��=Eq����g�Y޼&��<m�Z@���y�I����V��D�i[�΃�H�û���ۉ��턬�����'!��x�R����葔���>��=*�l���|��6�!{�V��?J��Z��h/�wD#:tk�l��W���hx��Y5'<�����zܮ��g��-��@�� �ʳ��ɺrzֵn?P�|r�+�5���牺qr�w�'x��lO/�I��"g��N=*|n �SH��A�CG\G_tl4�r=���]NX�Ј\�N >1����.���j�J|����.=�b��;�ڱ޼>��=�/�M��l�\pl��1�����U��dj��q��>����X�B��S��)� ����[��=�'!�W�V���FN�K�G;�IJ����f��R̢�������>%9J�H-g���k���޺��ɲ��7(�,D�,��spK|1��uL�^�~�ɝ��韽<�gi�zA�[u�׷�����f�Q�AN����j��a&F���y�������v}s�Ǌ�g�㢟���bj�X�J�0<��7$(�HW�8L�Z���N�gr!B��_|�N�3!j� � ��|Ao��8�0�]��eڏO��Ũ��RM�8!V=���b�u��4_]Ц��L��o��W:I};_(-�j�y說}��{Td�t������� �~�v��_���d�f	��C >%5����g�9߉*�&�F��7��C�<��ۨ��+�M��I W�ߖ%�r͑�0��)���sI�&�YG����uld���K���	8�pk��Y���@��}݃�N��R�dã�2�ZP���n��x�7�<4��x��;~����-�ZWf�~�l��;^l�.�q㇣M� �.�(E��; 9�S��٬SYg��~��K͘Q�H�ͳ���c�!�z|�]��Ov�1v51��o�e�"�:#޴9�vL�Ӊ�h6+����ǥYTy��B�?�+j�5��EX�éْт��Z�/�&ϯ��}�ܚ���,���]a���N�{�t(D�Z�����6y`p�-���7��Ϭ/��в�HT���y'�X��4Z��6v+�޳?�-0C�������g���J|�[����i|*�Lb�7�'lb�"{q���3�����g ;�H�4}V
Y��=�:7�[�B}f���>s�(*�ڞ�t�l��M�;��ݏe�����)�2L����?u��{N��?�En���`/�㟸���n�{E7��cE�t��+���B�A
`M}?��$�[���gݧ��~5�.gUvsGY%<K����w���J�;�?�0��p�[���oν�)RG���u}�nKO�b�"��9JL#��,����`�{���G���P��e������4)X��l����keL˵��N�o�����Xj�83�L+bE7��3#�����L��Ӱ�����I�dG��/����`IO^�~%Nj�7Nf�D7��/�w�8P[:?!���
��Y�g��X��\ ��RI ���Ӯ�;'R��s�_4���Eۙ$���$�b�C��T���,x��'�u r��W��S˒öE�(�t��Ӌ���ww�'�!�X���y-�@�X�O�����=_UAL%F�O�]-w���Qy�$��c�'��)�|�[���OP��ǂ����`���4�mM���f��۪ܷ>ni�#uS�C����أ^i�L85��Ҥ)9�ͮD'��o^K���R�#��ym�y�n���р���L��)��Y�!]�h�'�w�=}̶�Z,1\�͠]�4��T�@��4n�尼�+�.��O�:3�c��{�ch��gk��W3����&"]�Ȱ�<����T�ȟ>�{�z=�m�.����eH ��\G\��s����Z���w���%0TʟN��Zra%�7�6�蟰L:|���P�D&��NxF�|%>Y
�n�@s3*�:0V'����g�(X���T_�ɣsc�#����?�[n5f8��
�2�f(?��0^��M;��Y��I��S���m7Ϫ�`��}|'Fx�b,2����O���KFc������f����3Ń{1�'C�=k�덒�T;�Gi�� r��rݘ���B�+�=j 0pw��j��l���y�Fw>U�Os��^��[FD �T�s� ��h/�V���F"���������a�
 L0�6��!��x鰮�P}��\6�Wy[LO���ݶ����<?��f�;��N��s�G����R�� �������@�_}>�aqg��j�*��tw�V"������1�\B:��^m��2��G�s;1�1W=�((Ay�9�8] �^,������}uzؕL��p�Ý�v��{	�4Ć�	��Gx��B��RB�p����~ù�����۫ϗ]��� I�b.ݨ�B}E��l/a$�̱8�� ��7��E���U�e".=�IfN����t�`�L�u�Tcͤɴ/
fW]ؕT���!��� 6/��p+˺2
�LTH9�������sE񖑷g�z9�
��w-m9�2��-U���`� 5c-&.t6^������%���L�',x���B��PJq��qz��=��b�2�q-��٬�����7��CO,��x^沒7Iao�����kHg�&GiJ_�b�&��.�q�rLaT���U������+8nRT{֝���x]��[D-J��	�A'����pq��EL�7�t�����?΀��+Mn,JN�J���&��������F�+�l:�>��Gt��� uQ�h�n�U�@h��B��c%�>�Te��p3����)�z�� Mُ��Ee�`<�\�?��P��������݈����ݮL�+X8�+��1�� �+(Ά�p��࡮� It6�H���hD%^��b��!!�zh��n���3�g�M� <P`u�Z����'�G��O�ƅA�ȂF�ip�^��|SB���}���{�˓+^Q>p�8�ĉ�h��l�nJ/B�. l$�>���+�ռރ�^�����T\]Dy�}�u���
������#6$}A�r�ó+f���A~l(:	A@#Ə3 ��D�/�f�(?�׼W�'��n/x��g�g%)��ͣ�(L$����3Fmg�tdu�ئ�xA&NNFt�I�r���eWK���e��	\���F�Z�)(�=@�d�p�����A?'� �3�}-ҒG�o[ټW�4p~����� 	{!����-mUӰ���^�-���CX�Yk�B+|�H��p��X�?4��+(�e��O^s���ATVwSB�C�*"�%u�U$;Y9P�{���?���z��G6kA�Q%�*��)�L[�-`�$4�B���d�^�d0�����Ա�k�`-tK[�;Z��m}��J�QF�ow}��A�ؖ�j�=c���=|�T��)�( -�͟�M��0��OX��;�;�ɢ����-{���5��ρJ��\�kT�A��h�-2�w�_���k�=&�W���nvm.h�������)�P�C��Y˓���*D��������������d�4yoǍ��!�R�Xy��/?��7���'OXT8#��*�S�;2��;��Sq�k�����B�8�]����Y��o��\���57}�[�̺��@�/j�]�qǨ@mJ�2��	��Y�|7�������,'�?��������T=��]c�AG��V���e_E�s1uJ�����B���!��)	���y�7ѽ��O	���vm�S���A��ٖ�i<���Mhx�Э�2�����Q�)���N]������� ��X�U��5� H�b�*�ǄG�]Ƿ�57�2�O�nN����+���(�Y_qy4���s.l���p��u���8hf�������v=��@�W��G���-F���7�}�pݧ�y>1��񺣆��"�>�>�_#��׃��I@3\(��;~O&�O�-����W���G�.�P��<����u�{�5!g�͇�ڭ#[��0�YYNO��s�l��ͺ셍X�:] �V��^�<usM���O�3�Xzc�?t6�P�|���G����dȝ�
������j�-��ț�m��G ,nVQ>(L�z� ֵ�JX��>~=��L��Izu{-���B�+��HM�����U��!��N��惂ެ�d��goFo����NL,��������kQ������K��	t�?@Q]!��?�VT��2�����hG�ʹ��6i��� �M�O�Y��Em��p't��:jE���Q{qN�p%�ڝꟿ�j��}$��%�n���y�Y?Iש�p*�����E9�'�I�mv�ƞ�E����f+�ʗ���4�\QG�ڀ�{����Ϭ���*T:ե\(^��d�})fyq���V�tg�p�y�P�Kw��mK{���Λ�2{�v�q��NSk� E��{�r_7۬��c"-Wh0�.c�� R��7���9��a{�����%~l�ğ��{�j%�qDӼc1��mTb�O.��٭�c��\v	�	�/f]9��wc�q���K�� ���
���t����]�q�+��G��ϐ�w�D ��t>|�gEI�˕R��#���X���:�-~�_W<I�\�?�r��2�M1�����[��9��q�%4������U4�e�4D����NM��b.[�W���U�oI��MR9��0;w	MÛ�W1jA���5zV���qp�x�E��!��	2y��/���udB@�L��^�F~ݰ�a� �]JT�֛���:�}�RQ~wT���t����1����ۼQ�sk�����a^{��.~�V��-d��!CȖz,��C.&�Kl��n�li�J�M�| Xp�jS�p��=$��������򱏞]��KИ�/B�0o9����?��O������ǛZ����)�y{	}�罶E�R���+� :��?3&�����T�A�?~��Z����'&y��fr����l��"Sy�Πv�>Hv�@��bp�i^%���H�����Ե���/z�H��f�C����-�����en����HqN.�e����%Z<�_�c�@�H�S2�N��W�X��.�[�ovI�8h�N��RI�`3��|OS��wk�~��#e^��s]��73�n5�
����*���B{I��BIz���[����֒�f�	���.X'd1�-zV��U:5]�&��
��j�t��,v*9�g,���?�m�.�R�k\{�sh�z�wR�AtB���R�;����֗2������M_p��q:tԩ��c�99.-�z4X�������kV�HK�4�(���� (���x�Zzc-oK�o5�,��E��]����h�PgE֛�9&Xc��8���[��l? ��^K��Hs��,�A���?z�EZwG$��1�T����7��x����D�r�G�!َ�Y �{��N�%J�AWS��N�fB�H�}�����<6�%��� �Mmu���H��n��!��t��}L�����z틨?˭;���6t��؞b�e�՚SG���d���0�C�g�E�|�vl�./m'����|��Ů�s�
�u=ݢ��	3T=k��2 vM/��$b_�b`(]��a��y5���h �++>r�Υ*u�@Xי���+�|��T}�s$lك�Ŭ���sv��ZO�)(�g!�[I]P��/���7W��WY ŧ���W��0�,w��iD�ȷ���`$���-,L�������ɜ�ї9!��N
���+��?S8�Y�GLK��ٚ�\��^�uۑ����-����
��^��Դ��n�z'Aa1sP�77��|�C��(e��nnO���vA��J�D5d���3v+��߅/?l zW<)���>���Z5zC�Mp�L����턝��[��ͥ����������p�?Ԁ�F��+��X,��%W��/����JێSF�{W
"��-*�3��{	��3�֩+/�q!��7����=�M>U�ë"��pJ,\�ioՊ��iY�V��6��'�s��h�;�k������Z�4t�//wyd`_��^�(/hoI|a�����'N��#I 2���ޠ�l�&�c}��r�����96 T�$n�CxN��'�j�Ζ8ԓpb�'g�T��g���3��ۇ+K�[�R��oI}>������<�p���N��{�iK���k��3b��D;
	s�vy�Zkrd�I�Y.�*�׬�׺�ֲwd�7���g|�{)�ߦ���Q�[,xf�ݟ�����囻Z4�f؉wN�D�P�8�U��<�F���A��V*^�59�ѯ;j��CL+n<���[�mS��[�>���Sk��9�x�ݫ����'�������L&:V�b˿_{ /�C�'�	���Pȕ�2�t�O����Сy���M�	_�p����.zfċ�#p�#���g>C�mm�\�*Tn8[F�YdZP?v?}���8$o樗!�ad�� W~�Jr�È�!ς}����	�{����h��,O��L�0��mݦ�O�b�h��|.���U����"FG�fTW(b&��s|N`Q\�S�x�����\vF��T_=���Cw��7^)�e��J~{���b�
ycY��c�hh�V��"L=�?����&[2-�wM|]kL�������/�<���l��$U�L,ᆔ3m�l�w��s}�-�$�_�Z�!.w3�P�7s�ٍɂg�h��� �L$r��+���NR��k|V�i���S�VƦ�*�V�����W$6~�ۜ�	?��?�iQt����$����b<䦤�A?d	u@��Q�nŃ���l��؍�$�O�ĳ�y"�_ 6�8^9�ZODR"�`$�q�݁+�Oj��c�R���JԽa���>�T(�k��W��;����l��j�v�g�!����$b�w�w���+D�C"�n�=�nC7[�~��Q[���f�OYz�M�n&Xp�Xo~ur㑫ÃvN��Ζ��mJu��,7	�Xr���P!l�����":9������^�!�24:�v[LA+��>����5o(�����j��i�w�ң�	�d��C_���?ݔ1�.Tu����cl�PN�i\"��={�i+�ҌQ ?�g�ܬ�!ڹD�7�U�56XP�Q
)�� ӄ��Z�j�H�q�T�k�{��y�v=�.am�q&�	�)4n}2e��D-���u/L�l�r�f`�T�;�y��S�]r�����0�ٮc����+�*']�M7��W����d$�G�ҷ��B���B'k���u&1>��#��(*�9�Wht
b���eg/jMB���)�������&ƀ�8D�=*�J�Z�w�!v_��.����Љ�e��~�p>��(YN�^p��e�W:�v�b`�G��iFhlù�K�����j�3�ƴ%�$,��^�f�uaT'��準�ɐ-��=�X�����W�#TIG���{��j�՘��mOO��		�C��ٹ����S����W}���q4F�G��%��,xg�ސ�ν)e�]Po�s��p��A2r���+1zUK�]1�߄��p��j�����M�.�����d���2�V�Q2�,��B�̸g\��^��q���^<��.�dy�+I�pp&���.y�6�A���4��N�bj-'���ۥڙ6��r��_/���k��t�I����RP��}�=�W��G?C>�%�k��V]��;9<��+�TfQ���G�G2R�>�@�����o����s9M?��`��� ,�3L��21��	U_�eL��1�4��A���ɗ>�L��k{sʔ���!<4;�r�z� �!�7�1霸���M�|�� /#�Ѻ�5`aCDTS��.o������*NR���|���;�%լ�h�.FNG�ܭwcN�����C�������.�����c�ma�Yɜ���68��#�g����ٕ�H���~���$I}�',6�φ����%̜Z*���о��X��~6.��8t߫�Ⱦ~��耔�*�Y��O\��0�������d�y���d:��V�5�؆&���U9��������ۨG�7k��k7a��7�cZ�ڹ�v&bbzL����E�x��7�����}0"~������=@��Gؠpq�G�K!��y�a�I�F}��Ig.	I����m�����`"���p�=`��Z. �t){v����Ӂ��ۺ�mW�k��	���Y��j�)+���oP��ή�օ�f�H�0y)�- F"$�phhRu�h�b���oÈ���������3ϱZˌ(�.���S���?5�#+o�_;�~r�����S��T�P�C�b�"]�H�'�����g-]j��]��l�)v����%9��&4C ���:��-���%ғ������=R��$p<F���G�xK㥓f�*������ָ_b�۲���Ń��M���W���1��گ�Y�u��6��t�������
��[[g9F]�����ʦewgÉ�9*a޶m�zFW�x��."9?��^�u�ez�̻��n��m�4�����)��Dϲ�Ur2K ���,�ɴb��	����aʸ3&)�<�S��\�%5��nyዘL������'�9��q{�r���֣�V�K��2yi&Y�Ӌ��z_&�U�f6a�mQqi��u���v��_�n5��*�}��F�F"�>�xz�[<�o��Ii��V�#Fn���y�]D�,/F��֓d�~����7S�4��^>�I�3Pz(��������$i�L�q{�!vH��b�o����~`���/~�,�]c�}�D��w�d�����3�)Z���&�Ϲq��p��ἧ+��`���� ��U�|_w���yqB\���机��L[v2f��"U��Z�i���B]4�,����� �H�㕶���>+'��zd�R�')�o�u�R�.6�RJ������`z�Y{uBD3%����؊~�|�;�'������G�[�5w�Ø��RQ�VQP��!��1�iF���H�����F���=|���޿_�Kw]�uo��s>�s�}UD�;p��oK���*�;�S>���[�����n�����^�
_>�+���޹ #%�tm.9��`6�l��mu���g2;��t(��1sT8;@9ߨA�Lo���8�泆u'D���[�nW�#zY�wL����Ees�ev��o�wj���q6�3)��0�ʶo�d&�[(��͋��ᥛ����le��_2^�����_�UC�G��b̆������6|+MB�S��s��A�ss�R�L⨛@ b� �l��f3���W%�v)Tvc?�R�蝖����G��v�2�G9�E^�d�6;�Mיr+ K[��%�9@w��r����kc���L���q�F��$��D���S��%�,S|���K�#dj�\�~<�-�,<ۺ&�9O�3"�b�P��E7xJl��?`�fΤ��)]�)��מ�*"c��\�D5�!6q�~�;G�����6���i���~�YC��s�U�}u��d�
K!���M�re�yue��"c�j�ω(qE�M'ͨ�r�_� q	���>���-��ɚ������_+F��gl��؏ZcS�����Y8bz�����m��r�=�2�w:t�[UQ�ـ�u����w�2�f�lwS>	�=��8�`�e6��=���qj�.����F���W��χ�o��������GQ����_�g�
KP��q�_/l����g'�l}/`?�{�T���>������o�ɋ����i]���}�b��3� D���ø=�>��a����|��������#K������)C���|�i�-'r.8�B�݁�<�ΤS@��aצ�::i��4�4yotH�\�6Ȫ��a����\s\L��p)N���#-Hr�\��iZR����iP��ٹOw	��_��,�k傠�|�R��G]x*8Щ��ڣ]��U�֕�i��@��QD��D���|��mg{�j���}�!5���b�@znKI@-+��j�I)����+o����5�5�α�s��@[\i���f2�tK��`�T���9M�n���ӤW���G٭��v�-�"o�#��/v*�f�#��U��������d�D��{i
|���
C3y�m���Lw8d4dvEi��]��S����K���9ĔͶ���������+G�A�G�72o�ߒ��1X0�ix2��W�.:=H�y�yp�.ԗl�^��>E��[���
�B������zAW �6Ķ�PsYF��/���Kx!n¹%��Z�r�q ����;0¶�=?���`e�������a�uKۑ#������w{���]�yN-Ƞ� �4����T㐼!-��{�B�#�"����U�)t/&��g@�
�4�-�+K�\��LNcܜ�%�o=��R�&�B��E�75��
�Vs�j?�7�&^�����YLC��3`��N�F�.g�Ǘ��kn�{R����2����Q�AlJP���Ա`%���-seűJ�L��;(o���� ��G��~���~d"�Ե���Ǻ� ,�d�o"�qZt��G�S���J����E�O뭷| K2�¦�X�ZB�hT��0��X���Cȇ����^V�%t#�?����,�P�۩�#�.��Rn�/	�>��l�����O�@	i�]u1V�OA�,�o�������	�����i�=����Wt�g�E��m�Ll�}}Q^>&"?��"��F`��Bn]��^�yĥ�=*�����HX9Hxk)~��qBr8��"�w�$�KN�U���9���߀���͹�o��O��8�v�X�[@���}���ˆ�b���<�66�.���;�ϼ����m_���V2��x����P[F5L)�q\zA�nμ��S�3B�x��F�Lނr�_��@�m��k��X=����Ԃ��q�lG�_�U%�ݥ���Ҿ�J���[Q�~b��иz��X?�ک^+J��JAy��U�R#į�>�J�
��`���j.���ˣ�un8枑���ٗ2s�@-(?E���<�KBމ(���?��=�LZ^������œ��)���D	Po5�1�/z`g�ln���zn��9��w������^ߒ�,f����P�MSOղ|��p��`��7�R�6��R1��l��1j����"o���!��=��p� ��
���	Uݡ����<�¯�7R_���/>z	`�Kۚ�U  �Ô���l�?�� ���5�����AX���f2rUY�ֺ	J;�\y9�j���R�b�/p�s���%e�j#�%�����B���_����:���jF� �<��a���iW;1=W+<�Ŷd�
�YU c��8�7��B����������|�I����zU�?e�����a�;�Gz��7//~���\Nl�W|�@9�K�n�5��;X���_�Ɉ���"�w����n�ae�OR�nO՗��7~e�P�4>��������h�k�����v��r�Ѥ�������TU���˩��[�&�ȍ"6�W3��|��ҟ��`TJ��ȟ3`���U�:{�� �m_sm��:�9ߘ�;�]���TQ
	�6Q�q�*Sek��XƇ T��w��b��3��%7�޵���,%�չ ��Ot��� 1~(�q���9*�eK,��~�4�K/�w��j�~��.�U���v��?g��>I5�G����m<�M�Q�&�o j��|7l�j�e��}�/��a��3���HML��w��{|�X��b&pa�M?���l]�ן�A��9NM�U�J́��M���Jw�;�{��Ã�d��k8��')6[$3�J�|����b��|�5U 3IyT��1_Fz�OH�Y
����9�� �9�6�o�立Kg� �<�P�����-���&�����ߞ	߿8D7#JFb��3Z#��t��&���	3���	u����_s <��� )ۇ�ď��#v�[�o+�ҭ�Uv$�(�KX��v��B]RLs�����,�
�4nՄZ�O��a6Qv�'׫(2���h�<I�!e)��YJE��!�[v���B��u�i,�i�q�Aln+�V�@�o#�lþ��7����_;�z�7n�J�I��oI<�le��<9���nt]�0���%�س�����
sb��I����Z6#���ǨI�#J`%�)\"/u���4|f߶�дoC��鈅��1S���m0�dVY�M(������:���>�6��]�^�)ZG����ƴ��	YX��MQ�`�v�G��j�$n�Ug�TIv:K62�5�3s�}Hk�����|h����z������;�t-����{]Nt�3i#(s
?���I��wY#/�X�5�1XHt�h�K=�U�=���ym��?O��l����ςH ��Os�Gǖ�y()GϋҞ&7~__i��-`��^9�����(fv��W�ve7�k&��m�a�-�_^����e��Ռ6�ʖ��lL�`GסW���9��aC[�fDS���D?�k�=�]m�=�y(�pW����zN���H=b���lf!#�g��*@�zIx6��y�+OV��`������W�lҒct!V���{U�����w�(|�$�m`{V�x:�㣚�2��/n�?uF܌Tzꎸ�*.T��7�$�/��M���v,95��|�a�����:���O:��S�L�hFF�y�vR��HMg
��.F��$p�S�8
ݧ�T�>����Ñn�Y��,qm[�k{[v.M�L���Ś1��~�����w�d�"�ZB�7�ק,M��
�,�P�1稐Io��K"�5.~��E����l��YZ IZ"I�	�����ʽ�Ç�C�Ib2>��u�ï�,{Z��?F�	
o%�v�Ӊ.����`IN�p����_��s�������U�]3b�/�����\��k��ׇ�Ci/^W�=���o����Q4`��@BY:�-0�U��{l>�YM�BKŝ��A�ɣ5����`^؄�وW[��%(�䒅r��<a��|�{nMM"%�$�p�vH(�0PN�dUtgRӚ��8ܵ9�L����i�}�ϭ!�%i)k/��l�e��.t8����w����0�5zJ��8�&�w8����x�PPbu2VL�x�e���T�l�&m=�
�e���/8�/�ϰ�|!tk�"��6��I���n�����V
�.k%z��3�Mcn+���!�(�=�x�7�׆c����HB�������(�(w�6�sp�4��#�Y�xX4B�+k��Z,�� ��;��b����$(�ߣ���gRP��㚃�t�9�]9�Q���o�Ä�}f�^K8�O�m	��x�sd�DȎ�������'Mx�,��*���a������|c�Hs�-��V��W_��f��c Bxў�Abʛ��C�_�k������kuWö�E��{�]�D��v󖪍$>����F�f+�'��8����-g�k�7e^wu��l��Stp(��V�bs,�s4�rV=�1=�F.���\��+�O���qߍ�S�S��;�$R�%r��fdܧ ��X�bٟL��(t�:����)=����7:Z���=u�4w�Y������X��Xئ�g���\@N:xzf��j�l1��CB7S �ls��@R��I��v���GNڃO&���k����K��NY3J6�X�E��ʖ%�U�����BOL�*���i��G��T�}�b$s�z.
�ˑ�y]�a[��`�������"8D I~�?;��'	���eSS�˖����|1��_��a��;�k�p�?�����;�� �{'y�@�Ȥ�~�+.ⷁ=V�<;�Cx����%uu��F
I��b��!���+-6��}-�w!f�cX����ބm��;��K�k:?�^Y�2�JOŏ�,�s���tf{���9�h]Wά��1�笓���/!\��c;�r�ɽa�!d���D��!k��e<7�o-�^���\���'Ώ�_�
oO���:$|qg��Y���ӛ9U���p|?�v���ݰ�:�i�HkÔ��]�F����ᡃ�ޤ\O����T���tQ��!P�&������f̃B�ٚ���#�@O��0��uQ�x���=ƐK�u�4)��q�7�z9��������趚X��x5����c��*bW�B�+ AtI}�m����%�<,�[{�&��3&�8�B���z���7�䷵P��2��35�Ңu��$��l�/uN�Vh�o���y?���� �<��߁�{on6#k�L�����V �?Z��X7y�3�	�g6���}�3��J�d�]d���>����U����Ԁ<��k���҆��D֫� ��&��1fjz�Vg˅n��K���GXך<�K }�S;�g�vM�f�o�g�\B��p��2�c�+�v�&��l2+�ĝo_����$���y1 ��2"g��z��j�l��dE��>.�:�p4�
�1�Y �`$�ĢqM�1;�%�i�{��W/�Y�/��Z 1wa��?]�Pe��G�����E�m��y�Q`�S����7Ӟ�аduC��vV��=mM���f�ދ�uw�~��k�/��_��|y�@eZ��:��S��*��|}Ϝd�W���1�C�s������<o�h`yy%�"v.y�ѡ���/�0�˱G�����B��2��7�N�۰�����\�9�Y���Ϧ?�v�P�n%qtQ
�@�6�q+�|-���׆�a��Kz�r蕗�b=Q�n7n��%AN~ 狗�OuI̢����;�g8�A�~��Zxg��T��6 d��yt���\�<#�ed3��VhD����F��#'�y�}�'��Ue����h���I�=�
���/�$*�\��� &=�Y��{����v���$��[�0b���+r#O%H:fV�1�#b�|� @��v��������V膓y��E������f���)�{���)Ek�x�����vS�����T*;���SV���u3����7.����� �զP��}����IB���`�_+�u��5��*��jz���� Ó
y��,�(SSE.�)�'���`�֏9Q�]~�-������Ը�dX����k�ȿ$]�*(��&�.�;��H��h�~Ƨ��?ƅ��{�VH��;��x2n_����,��/u�읮q�@c!�B� ��!��l�_k9{�oh�ඪ�i'\�Fh"��6���%b�6V$6s�"�4 �S��g�R']�d�u�O�{���O�y3���]��	st�Q+4�ʚ��������(�wV���U)$Q�M� �e�;Þ���S4���A���X�=��=S]��9I�c��,̯[wl �\���Y-.M�_ ?=�6R3��`���~���5���&���7������YH7����6��T�mOn���k����{#��6.C���VM�M�UV�]1����vZC�>����͂0��)N��J���C^#�=��;Ń�wYDlXw��e�>U���*|�������=��W�F���i��6��Rm���o���se�&�]��p�%a�e����kC\�kٹ��k��������$ ���y����7�"[���C�n-��(����x�Q&-�墶�ۜ��a�ȣ��q�y�-��E,3��;r��p����]�^��8��t�y�U�� �~s�x��I��p�o�odD=���;�0�e�F?#�h�����0@|�O�Yqu�m?^�����H�#E�1���@V�|c�|� �Og���(l�\m�,��R�?�m��9�b�7�F���$�`�O��[ݯ�|����Y+m�X+�SZ��~�?v���+4�������u��N�k���3  z�5��ɿqbY�
3ݻ�㍊"j���Vn���"^�h$Ա�K�Q�O�@�?��g��YL+w^��vA[�e�,"�>�s?����O�y����x>;v3��d9.TE�b�����-_��r�Yѥt��>�iv8:+(:}�ѿ��t��Xo暂����0x}��b�U�u�ֵ�H�������ͮ}�Q�:�6�\�}hR�n������=L'53����d(
v<&����gH�C��ZIh@�	8���I^�cN�,�J��q}0_����=,�� ��)7�Ҥ�8`�RdTVc
��(Dj̚pg�:)�O:Cؼ$;4={�x�C1�@����:$��v̳���U; w`��qk:�#�w�~�sTy��T����t��i��#�>�ѓ�$q�g���_;�m�����cai�|,[���!�?5%my����Z�����V�d�J��C��,ʅKv����/g��:s��Y~�`~���	�A*|�RS0�����w����v��9x���.t*(��<��a+찰�6�nC5���5���#����k��4��1q������J:�e�-�M�Ex觫+��3����1L�K.����oN4\1��I����J����q�\;���Z��w&l��d�\�G0QC�|^mf���|wtْ���X�!��G�wj\G�xDq�1��f����|�v?���{,]����6�f���ۓ @a� ?u�U�o���i�8�/��-����ȁ,��&�0"T k���ۦ�Yy������6P�v~�3�pK��H��Mli���'��=p�����СW� ��#��\{��B��'�0B���(!o� ��ZC�;C�C�%>9�r��qg̩�A�A�v�g���	Q���e�1����g�Q�J��x-"W��{ݟ<LqY�'��a����b
��W��~�6��f|_} �}̕#�[%��X*�CQ�꤯�ē�i�S����)�w��:|NNC�B�b�7��,Xu�Ĳ����-"��>dK��ߵ��)qw-�r�fn�ZNv�(LN:|�'	Wm`8�콠B>�Ԓ��K��A���Q�~I20@T�M�t�|���cE��y�����;.r��A��pZR��0���J���օ�;o8��P�OO9w�|��]�a���a��f������Ɲ�m����Ӌ�v삶jy6�J�-����xmRm�K��Fj��t���z�Q�2��%
J~Vq��	��Kcq�_K��E�ug�[���s��;k�M�� �)2_$�3N�)9Hhj���&
�,>��u.�M�l}�����!i~au���{f[<����~{��(j�����W�o#�t}4�u3����֘)��:����(}�*T"��a���ڼ���ǟ��+}`wi`W�f�[�5�i��2���礃�+v�ߖV�0u�[a^(���9�zd�!ݦ�10��1���͐n�������lN�"B;!���|l��0��(�s4�s��##H��zZ�B�5acu�l��)�7�,Oڇ�z���t����&J�ļ�"tZ�J��\�l��l篖�p�q)w�Ij��3iƥ���Q�M�]ZFZE �0H|��Ə)���-i�yBy`��鞥����Y�o�CJ�6*����,춡��%U�N34m��֐����|��I�x�@y7�_~d�5vv��j�k�������S*P��_��R���L#�$�� �T��M�ͤ��[|��ϧ5#-��g4���a�u(��h�j���̶����*�'N�X6�N�~E�l��q���B�F|<�%??��6�d��8��ظC%��,�hwE�������C��6#(�F�q���:�~��m;猰
��8���{o���_����N1���Ϯ�uw�|��v-��>��5�1r��B�SS�Ib|�@��@:�,��2}m2�C�H2SY��"�k��UFLpO-kW�|����xX5�k����O����#��*����8�.cs��݋�ƪ�f����J�h�;+;��E�>,!�up�ˋ.���h$�|�#�U�Wޢ�>nѱ.2]�	hb/�Pk�������<E&[�߅�5�\Q���k���@/��J�t�	���%���[EƢ�V��!]����U����o'&ʕ7�l���+��\�mq�X�������ޥ�9��6~�L*���c��K���ז����`��W�63�������>N�@�Ί��vW�ׁ�r¬�#�j;��H�G�2c�h7��x��mp���c^���G�e�5�_�z�r�韡��Fg��;�]^���Í�톩϶6Oa7���x�z�1������<u��eY�a���+vQ���
U�����3X^���� �T�`ej�.���]��;
}Cd���7�b�b�����o+r��S�6p��Na����i�;"��8��� �v� ��#��0��Cj����AAW���x৛C~+b��2��>%-�����S:�͹��YƓzܩ�G<���76�u!']�º�?d���P8�2Z�6T��������{ƓZ�FE�^G򽶁�G	��G�
N[4J��s2�B�W�4�����;7g�eag�޹ѫy%aY�Z�@���ϭC�������)½�7+�&]��Q.#Ϯ�u5�fN��vmc����1���l���7��?9� &Ż�c#�o��j���VPtd����)��>T�垁�3�5&�2EeV�)�7�f���ٟ��zc���%��lt�x}*&��'�v��-�o}f:�s5/f�j7(���2�c�h0�gz��6x��n��~�.��L�d��A�ڡ$��'H1��]lޓ���������EE���A�[�)�˚+��?�?�
Ci[�}i�*nIˢ#E�����(��y+���I}}�
�Y�+�����%_"&�R���PR᥾%N�I�u4�:��-3��Σ3o>cu|IQ����*Z�û~gK9B�¾_�/�y{�h�����˛²W�S7G�\wr�"h
�S0��� �,	,4�X?�.��:�My���f��5��wJ`��E;�g�TΫ��]Q\�oCX�@��@���b�/ڇ{<�wm/�?�����?
!t��W��.��k��K~�Xm��k|�`�1���>'���[Kˣ�$��俕%*^���:I�����������R�����.�<�������̠A���sW ��G�0r�s���0�{w�3Q�HQM�ZD[��pJԶ���� h?.��K��>}$Y��5��f$i�u<%�%#d2�0ir�jr��S|1��Sj�?Flm��ݬ�/�˸L�O���N�2;���U���Q�X�eHc�e��fz�T
#C����۹w�S{u �sh�X��3��
9M��������⾚�Am���Z��dl��3
*��O���f�l�q�b�`��ߠ�DV.�祮a_�R�~�>�_�V�M�����ߟ��J��sW�E����5���$�X�[�Xa�J���
 ���$%4���"�I������Ak�0�^������.]��;��.���Z	����7�\!6�üvP �tmդ���KI��E�爦���ɸ�t����scf�&�4b¬3�g|�~�D�B�7(B럑���1Ճ&���`�}�9f�-t�M�\������L�qtc��֚/�me�ޖ����,$1M�3\h1�;�?>�pi���U`�, 7_�>�>gJŷk���Q��X+1��9�u�l��S'1�� .VZrF
����"֋��j��I��\��e�>�NP�n�</�P�|�?M�I�;�fov�v�xj��\t��@4���8����B4/wJ�EdN!�!Dc�K{�kΓf��؈���l�%B�eae��S��߹k��Q���q��%���f(F�ځ󡄪�<7�\\��{q �7*�MY���ta�B"���&�E+V����
�9��F��F�DI�z$�>n��h�ϳL'
M*Fj���0i�r"M�5�Q��ٺO��!�^�2�]�X['��\.�{����͠�㖣l����k,��0����1m��qL�b_�^җ�R����G�eK�>
}�v�r�F,9qB����*���ˆ�SZ����፻�h/����l�Fw�,bi)�Yj9x3�ĿT�����ݽC�	��t,�%�|�ӯF׹����m��^�(@�&~>�Z>D �wQ���sJZ\�l\�^�E�>��&���g2�(ϥq[�z�~�'G"O��p�&i?�%�ͱZH�(ram�/���eԆ�85��|������-v�\�a���Y;?��٥-��9������$�8�jv!���_HzMN':'	���Tf[j�5���U��p7+}K�kj�L�����6X��>�u�7��i^1����ÎX
梘� Hμk�y�7/��Uu�wR�\�S�ˇ{,~\����2�t�������n�ɏ��_��x�ۈ�M�������Ia��,�
����ya�?��~��2�w�C�o���R���?�6ٮ��5��·�0�V��]?�}Y����Z��l׉�WL9 �w�u��e�ji�a81�=�b�K�'^zl��Nzl���TE�M�D�v���a���]�mO�A޽���s������[��}��CLDY�͓C�vb�u�]�uڛ�'O��9@�&�?=��+~�`s+o���r�#A�$��W��2�+�n���E�#y��uҜ/�
��&�@b�A�B�����-�����mi�B�L�d�՛��Pm���<��õ�o�t�P�m�0����s�u�o����"Y���h7ƕ���ಌ�gQT���
ǧag�+*�2�ݨ��?�q�!��u�7��%5��bo�	`u~g�'���;�/�������\�*-f����<���QD�ݫL^�ߢ40�4�5w����7^Ѳ���:���m+^�q�y忞X���[1}B���"�� �O,<����r�*`yH7�Af;��Sn��m�;���fo�z7i�+-1[W{
`t1��Ty��`b�|�D��_�\ �Z��A�� ����26��o����Ӕ��m��~��R���r��a׭e�mo1�(U[.w%s�<���_���~���@�������\���4��~�k1��;9�ɾ��ϩP��{`��M���(�ܒ=�>Q[ �<ω�yE�~"+�=�{�WӦ���fT.��8n�K��Z�c��t�e�[j���o�0�����d5�ٶ���N:'6+����Ҫ�����#��=(�B��KV+ đ:�	�އTA; ���X��M���)�ꮦ�f�ɄZj�o�.M�bK��Q� Y��Y'9�%��n?6���h��%�n���X�U�$�!7W~?����Y;im��7Mz�)%Vc7!P��7[㨑�u���y��u���1{P��S' I�y�6�����e�m�˩�LT֯G<��S
�@�8��*�l���g{v�k&�ҧE�dv���*�#"�Eby�F���gvz�[��f3��W�(��2�����o���jپ�����0�VĻ�&fݡ%����šK̊�rφ%�Xn��	��\ذ�]w2�
�����7<zX�h{�鋟t�S^�T�=s*e��5r'�p��L���f�0��]%���|�^�}��D�υ��BL�㪊C�ÉB������lD��Kr{~�6�:B�p����d6Nj �W%��������P��{��jUNy"Uq}{�[c �u����Ñ �5W�����^�A}�<IϞ�ؖ�rcŦ��Hb�����S�ڣ�v$� \�=-*��Q��(����1:���ε�$a�W�wd�T�����zf_��V���V�f��tגqSR!��x��>$ݰ�<���oo˞ ��|#xR��ymI�p�^�ѷ"��!��i�V�q��������M5(c��7��H�v
W�_o��岐	�l�=�K���%��a$
H���&*�ť�t�o�zA$�M^�"hl;bW�8��Zx���6�w���;�PG�YU��H��xf�~�b��
�2s�"�ͷ�(��a�`k˩��j��d��Kӎr�d_�"�NQ�_@�����{NS���;�N�(�1�d��Q��%��B���1��'����}�2:ݯ��B硧UV��8��[�U	�F=��`���z��c�i��I�þ�z�擲�	���+^���6�S��w��? I���AߋM�%��u�7m����o�{m>���Ƒ1e��z

���չSء�CCZ��da�J褽H���ǥ J�sp~�)�}Sg���Z��@0-lF��YM�Pl�O��2�Y0�
F�r�����6�	����Zv�Â�3�#<�1�/�!��o?U�r�L�ț��e|���L8��Ծi ���Nc����k_�v� ��[�|��m�v�{" >J��pv��n������Z����ĕ�b�~��,�����WeU�ȥ�� �l��]�c�_�ibL&�凲�����~Y�
�X d���S�V���S��S!x����yQ��U��~e�4��ȃ�YN��a�o������qstwʮ'"i��tt1oI'U���z��(9��(q�Kܡ�S�a�C$O������E��tF�Wg��$v5�܌M�xĖ�'�����ͺk�ٟ7�QWu Í+�TDO}e�p�Jz�W�6���8v��Ѐ����!���5�CI�W��6Oܡ���qP���y洛�BCuo��W�V-�P�0����A|�uJ|���F�wp>o�V4%��ad��j?l���Z��$��(7�5r��]� �Q��o� ,��"�<1���cZ~�}��E�3Ю�������&����E�e��h���j��֘]s��+��]���}Nh���c�Rp��Z(�2��a�> �;>:m2�:@%d��N��T�z(?��9鈧�a���
�23Il�0�y2C�H�X*��df���=~��Ni��	4m�����o�q��0$8�9$_�{Hm�fG�4�ؘA���oH��6����z��Y�a����={L(י,�N��K&F	��b)7(�n�Å,���n�B�I�_y��]�~����ڠ�e�&�)���A7}���#6�P7d&�Y�sO6aZ�%be��ZJ��`w�+l�����8�gtCp��*+snL�u�����rWFț�C�瞁�h�p2ƀ�/x���cf��I�~�uU�1@��.��w����=���5ɞFZ��|�l�&�hϨ��Ю�TA�mP0Վ�j}߃(�#)H�>��&F4��,�5/���ڡ O���X���t�u�s$!�.���C�@`���̣��@,�Ϩ`
2'ȅ\�G��yk��;�8�~ӈ<�^MW�F������Թ�+�O���1L2�."��uD�׿��ZN�_?�)]e�o��I��[<��Tlci%��E�+��ȍ�"����&Z�O�PvZo^�#W.��[�80P��
%N�y�����<pl�P���p�-�kQ9xk�WJ��5���G����n ��-;,�fZ�$@a3���"|�7��`�+U�۹&�m(����q�r�s��1�nɯz��[�;�d]�ͩ�Dv����U���E��ܺ�N��}���3���eb?�Q��P�ۋX�>}��Z���>�7�W�e�\L��=,��[�Ƒϕ��%�3�+A�:is�����tK�I�.�ʚf:<%L�q�G���'	���m�	�g�6`������"3~'�S����T)_i�F�<]�yڎ�P��4A��)%Uu5˶�H�� ���8��*s�O�䐥}w��f�w��7yi�{�O6*N:�#��B�J�ISj�~ɉ%���O�"E�k�PX��@%? �t�J�l�I}-�����3�ג��4�3�.�w��
d�#'d���L�NM{9��]���XW��89P�!\[5RbK���� r:kV~���U�|3�91��
h�Gð���W��Tk����LO�ߌ�懶R�u���@ߟ��b��Ƨ�!�ٞ��k��F��2Ś!��	pp����I���`��g�w�h��;�˥
rݾC�B�zfd�'*�����_�|�����`�B��D!�qwrކX�(�:?�����\X���j��>�A�n���tNֶpׯ�����[q0}8|-��a����[�_c�,�O�F[���tp�u~��?�^Vͻ'��p>fe��p���O�%-��W9ឩ���k�|� �����9^���3��Α���<*���s�h���E��FVʎop$E-1+�ÂN$��;ٚ�<E*��z��� /!��P΢���]}*Ep,w̄���p^N�HA��\ѷ��s,R��2��<VDu@��Prg�f�����]|J���{8l)����]t�z~,������f䉗PO�_�d��z����M4������#6�N��?C���n׾V!��� /ȷ䟳X�a��eB�0��!��x;�V��U{@�L'��>u�	cIV�eE��8���{r5"���[khm�^b���r>��3���<1o�����B��)'#K�?���� 
��ve��y��{H&2��r�B6Z����ה1�ڵH%��,�s��imVw�X~��w��a�AG�U~+_�����*6��ׂq�@�eg������A��P$����B��i)3���M@cO�*��p�yP��P<��w=�k��{06��� �!%�ġ��gk��F,@xwi��3y	1*��W�SZ�0�6�I�ITvX^�
��DL�(�Xe������]����!� �O�̜���+��njG�=o �ڜ�u;��h�~�2��IYM��ʯ�30�%�"o�1��	9�}��{��Vpjx���t��o���ӱ���M8����sb�׹�~��EH8��y��z6��q���+�D�!���a� �i�s�̴�8 1+L�s�( �L�M	]��Ì͈Jf��N8�&BƑc�6�s�s��~��JK�%�LY#��)�baS���IA3|z߾���Q�]#j?���U��n�:"/�y�>�X�Z�:�^��P���W~?�}1i���t��kKJ�����^m�H���wb���o������qq�Ym�(�E�,���Os�������_b7���MA��K`�
\����[���6:s�c�K�W�+P���ώ�~W�ff�偝����a��4|���gP�w25-;gZ�P-���k鎶�ޜ�����^��_��Q����=�*
���ɼ}��Lnh�b��ȲBD���!��q�@.��7M��b�R� �3����'��f�K��YUX�o�;jr	V���
�V;�a�@L�/B��Z�m*)�9�#��;_����j��(�}��bl��I�`�c%���Z����
���܍�� ��*#�De�x}NW�8�[c%�ފ�������NA���ّH�Ak����6��.>�	)Tf��v䨄Ag@.������3N��˛��9��#)/����gk��nV���s;���>Km���WIl.�ä�N���X;.} �:o�7y��&q7�/�I���ݩ"��5Ao�����S���9�C������8�M�?�@ ��9̈=��K_�Y���2��wR�?e~^�}�Ϧ6 B�;Ğ�9=7t�mh�(�����S3Z7�3�jqI�!.�K}������3ί�7�,�-�t�1]�� � �ď�/]� /,.�L^�#R�<�X땥�<!Ȏsk�f���=�~���?���BzC�:ϥ�b3�#�J�sg���o_Z�|��R�<߿�q�������U��,�E�7�S�g�=-2���0�1|��y�|�H�����0#چ����HK��m�B�u�mԞP|���L��c�e�7p�yq|C�������#�$ +>���CA��r���k�"��]�w���c0����.ɿ�T�!0����K�5�y8�q}M(��Z��D�Zo�;�xB�8"쎶��y�&����-��f�a\�E���� �'(?�e�jQ�X���|R�Ը#�AܭϜ�_�T���F��q1d�_�)xD\W����뻑�s,O�� ܌�?'���9�0X��6mܓ���:����Ӿ����x��)�N`)�C�BYn�/_6׿���-�D*Z���\���ם�$��9h�=�cc�p] ���9O��oK,��`PW��c�JV�'l!�=L������+� !�H��\�[pи'�wwNpw��Bpm���en����}֚��XP�V�9��ٻN���?�[��4�#�L4���H��l���gj�_�N�KJћ�x�=�Wry��.�e)�l��(_�R���߈��O:z�Ա���*}q�D��2w�<̹YJ�i���(��O�4�C�4_^��_�ς�����KC$)����0n��'�wF��S�<��[���uڰs_��I3�����d��>��������0���P�g��y�Ƨ���'!���j���t/6,�=5��0����^MCq�����>���Ra��jχ�N]/V�ܩ��7�|�Mŀ?�r�L�_&��\��E-=��$�s���+�׿ӵih�<���`��5��������L���վ�'0ҿ������ {�Gq^�a-e�\��g�]A�^ F9����&KHW���tC��lk���Y/&�
,�'�aV��?��,�s��iR�W����Õ2��5�������,L6
Wm���:b`�(����4��Cj���?n8�dp�K'��>����W�?NH}4�N�f��c�/i�T��-��T��	X����p��C����ߚ��i�����W��\�Tx6��v;a��V�s���'�`�[�%嫼(�}�K��=G5�����<`��'����ɹ��Gh���p6�]��a;J�Qb����ZS�)خ��s�|��ڠ������|�瘸�ۆ��������*�Z��y��{���l��m�ep�n�3��?|�����p*T��2#f��9�7ȅ���4a��~�o�ik�D�_֔��c+�xC��􍼃�v-f/����@.�����]���TeQRW+`����A�!{J�~���WB��Wż���#ΦY1����[/�����?�;�V�h��4$�`�1Gb��A����b[\[Z++=ϣ�	cW�,ܼ�<�)��vު�%��]��}m����M'�Ob���V�н,��QO�������0��IF�~>�m�dfVR�<-���Ӏ���sT� ��b�K������\����W��V�b�@��d��1}lx�9|֗�����S�!�� ������������w`A����}����v|�>�� ���4G�cr��}�����:T�Y�aJ����K��%���V���E���:�rŧ �<�mņ_�D�^��H2�o����2��q2`����нT��a��q>e@�c��G�z�K��n��X��jC�RU*)q�<�ܰK�c3=ET���@I@�&��g�ج� �rHWyũ8����LW�q�裿����#���֎Ȩ��y�&�����9�����{�Ϸ��e%z5.���J��5Q�j���	���j[c(��D�K,���b,RfX� �k�Q�&]���⪄m$G�U:8��!��ƧA��a%%]ȞV���}��\�D�������x Zx7�|�u.��='�#�LhL�p�ep��0��g����/�՝�<&4�]�kpsz�0T+F�>qTw�5�p�ݡ���\q���K��*�T�l2�HC����8v��j5bZH�D�Y]�.?���G5�D�����&�8"Q�V���``hS��R5�^�85u��{����\�EFyM3�������2���G�s�	�T a��E�����u6��]��#�����W�B�΀�c(�s�+�H;g9��/?��hd�PS����7L���Bu���qx�v$$^�ٙZؖU�a\�ٹ��M��B�k�I `�ΧZ��2`��>-[柼���,BW}/�t��@`k��8��6�Q��{�8��y��󾜃�#��[5�Τ�nB�N{/a����k���z��Ŀ;�8Un��LD;��M���u�n5����x򠭼Yㄐa��+^]���-ꔺ�dX�_���^��b��l��s��Xd�zq�B��gV����~�L|V��|�z�n��V>uw�#+��˼�?+�A��%�h$���+жE�YIf���4sVv"]닟lB��ARY�cl��~呗W�-��m3�V��P��1aE	؅ö-����hF�c���{��9Ea�a[� ���`��BΛv�,�����x��ç�4.'}�G��/�F��!��Mm �Z�K4ö���̊��%�S��<��
�ۻ���vCK=��V)�GH�K�O������J�~�b�O>�tr+S\��$�n��mj6�F�3����N��8[�g
sf9���y�	y)���!��R��,������ �n�j���W��7xd;.�����:���#�7�~�\5��R��!����w޾~��X%M�;9��q3tt7�e@�1)�IG�j�T�9t���~,��=�����\��6���,���M3�[\�?�.�H�yM�F��?��;鷽nd!L(�ȍNv�&��
��#j��8�N4��Y<���
�mA�yZI�
�B�`�eR���dk�훃v�5��2]9Y3����>����n�z>�
��l;�5܇�F�e�"��e�����t�>�q,|�����a/�v��6�H!D]wN^��O�g��G�OLyM��'��e��iN���c�fN���B���}�,�����Q8�7�|wv���d?�������Dn	��e�j�a��)��9�X"Λ���3���4��9}{��G�z¹�(I�6���i�I��[�gJ��(/�n0�../0�^_.*D%�|�F?�����ߖ� ��~�a>`3&���ן�aw�2�KϿ��6akS��%,_T2��¼�d��KuS�
�$��Z6����|��>ߙ�<�ڋ��VϿ��k�J���@����{�H�䃗	�ؕF�F�����b�D/�)9�du�H�5s�	���9Aq`�l� �Z�A<�
v��T�v�YDw��L;�[����o�G��#~����7vwr����/Eɲ�?��4���A��U ��h�B����{<��� �"�q�<� L2����������j,��q��?��}������Hd��yG���D�?�k\_��Q�ąN�����;N4�\q�8�P�����L8�,��5��S���uFI�2f�(/����ɕ��x��ǌ�r��$$����}����>�%!"�V]�}ԷW�{�w�˫�x������'�U�X����:�s����5-E����ۂ[�M�~fLxȲ0��a�GZ��pLq(�mJ��1֑�ɨ���G�����ȕ�T��J��"!J�����@���{���tm�����i��>/Q�f\+��㥔)��둜��~b�sL
��s��O׊uD��c%	��Fly�I͢d.wy���P?ɇ�(2	�9-�� $M����}D�%
�NݳE
E��^�j�P����˨�LxYd#����}:8�n�����2��������rw�.��3ls[+�W�!��)��d�6^J����C��?�=�������3+f�B
%/kiv~`C�|�r��ʅ#�)䚼�Xd�����C��~�/����A6!s��?�*�2wRz]�[ƈ�̋X��)��6��?�<��z��a�lG���]vݮ�g)��22`��~7�6�I�XN���*D3�dcێ`�h�٠u��17�ӌ^E<u_M��)��r6"���.^����B6s�,ge��u�m���{T��6*�Bt���q��o��t�6���lj��[
��	��#��o�c�/blCDA�(���;�ͩ�S��Z��V���ב>%/��5۠A�^����X�Iч��Lr�Ҵ�/�~����\�ܴ[� :g2Gv��{�p�gv#��W]���:���~�}���T�yv�6�7����/�̓�[{���[��'�z�O/����#�\F&��͎��q����&P�O��=�i��ݢ:�;�c�
�����J���\W/�ںP��O/仨.!���ƫ���﫝�'_`�VM�<�̯��� �����hs>�'�y�H���#���7�\.��ztX��k�v�u�`���¯��G�����ehu��;�M��a2���$v�oM��)���cA�{���}**�9MK�,��_�����_ �p�� ���y���a���c[�0�����-�� ��V3:���!�r��J:�	E�����
�K�T����|��\�\�
�
�j*m��\6��z�/�4�)����"����x���e��:�&��pͿnU#�/�+��P�NFv�����&3����hY���Q�I���rs���@N9�������&9�R��9$����U�B�z��*�Ҽj��Ͷڔ��M'׾��-�1�A"�f�l��s
9�y��]���{�i�G�!zmk����"���3�Ƹ�"D>4�N���i:h�ǅ<[�J�8�,d�Y��o	��92���F^,㭞�?��Q�N{�����	h`'��Q0}�Z��߳ zX�MJg��Nl*�1taz�5ڲ�r��_i����:�cڶ���|cC'��w�%��EF�WCĂ�y� p�w���*^���ZÖmmY~����dDv}�WWv�S!>�:JO�҆p��(���jۥ�%�w��7���)�t����mB��XG�ή�HV�)���y���!�\~ϢO���m:�x��O�]�=g�h��*�_��V`*��M�zq�9kmk���n��m3$��ij���q��G��l\���p֙A:�Wy��c��y�6u���P���R��f8���,������� R�~��4f22�| 0N�x��<��t�P�E&���b�:��v�[�۪��׵�����~�.h���P����L��ni�o�����V��:���̷�z����M����}��Q�/,|G�$q�2��5P�`��Eg���Z����hS��p�n&ƶHc���N��xuHt�F���'*=q�|��01'c!=��Ɨ�:t�g��f��N�L�hh��xr�q�z�>r��#�/m2�׀�9�~���q��r�]�z>�$�#�j�e�8�MB}k�¦�<�չ8��s�HK`>���}��e���~�'d����{U.3�r���M�9f��!G�Kl��<s�ETR%��7�qe�Ç���u?�']X(�)n��/8��V6�#�����d�VBڪ-^��/=w��ō�YV]�/����z�����I�~���(s�O=��^���t��?zG�Į��4�[r�ػK�`Qy�s��(�[��t���M�X��yɰa[�
_#�4f���:}l�{%;W�����f�2b9����^��c\ 0vSӰA�fЙnri�4��g��J�ҝ:���,)�Z���)�q95T�JCGp3��AΝ[g���N�1��_�=��(ol�R�j�m	{�?��]c�8r�,�7ۮ�!jl��&����8�7!����e;���YY�P��R5�!av/��\V_O�e��܀�����mO�����~Q߸��>���qK������b�F`Ȳ`P��Z�WgBj��t� p� �k͓[��F��<-���4�F���r���<ٱ�pЙ���V&w:�,��T����e>�Jn��s�K�퟈��^#��G�5��N�4�Ș�u�^������L��,�9��O1��E�n$0�T��?�cA��0�=�P:j-5�D�h�����ȼ�J��b��lc�G?"�i�:+��ɼFG$/Y��l�+f��>f�h1�~U�3!�{z�%�G��ָ�..lV ?_�c�P�$����\��4���Q��G���-g��8���]�F��6�vfQ���M�Us����am���N�zp���W�lh��)�p�mK�C��b�G�I.�v�l_��G����%'�K.��ι��w����*21x�#�R��j?��+���g��ƊҾ��~nƿ��V`�t�DD�~9��ڠ���z����~�>k:��g����O`|VH��t�Yc�AC�<�_jK"�H�������F�z/��y��"1gd�Yb�iy2{����U�Ύ�m��� ��~�B(`F�%>��)�˸<t�}�;[({A�Ͼ�)�W*#����X����R����Jۯ��R{ �\�5��f���~����ANLyIn��J�0�Z>�����@2g<ƅ�ٍV{�/#t���~���;lV��2!�0�G�m�4��׹T�b%�{���}�C��-C�� ��t����Y����ٕ�~Ccj�%��El����ä�u�h#�RVֻE���:ݐ�S�����L��i��N�R�!u���ڱ�J@���3��V=�"��x�6�)��0Y���]��Nn_4���~SI�e�u�&Ia��R��G��qj�T�U�k��c�	2�W-����_X	��^��VnfU7�f�5����谏���A��,Q������,Ki�W�h�&{�+݄���}�VI����-��`|����V٦��L @���軼����i(���Z������+�Jn��
�L�K[��O�f5��eI�⓾�@T��i;_�,��b*=T�)C�i��10�S���5B��z�E�E�[�[#�~���O���31�q�����xg�d���f����T^8�P��,�zC�N�FF��ݠ��of��E6g��5�p���A��]�h�� Ce��b�[qےk�@(۠�k����s�͌��y<�]�d�n��e֍����)C�ޗ=W���#hiܔܯ�4�8L�N��f�.�����	��+�u�����R
ID����򀰥g1ل=����,2g�����wn�|[�0�q���T�Lz�>�"�2�-pt�GKXsȄ^���:İ_�h2p�ȁ��s�j�()b'����4�˩2�9���	���
�OвY~}��ft�$$Y�4���QK��p_vvt��Я��P���8����E��F	����ۧ	~\��!!�ڦ��h����d��cW�Y�ynh�z�an�\2���/{�_�H��I�W ��G��v����~ͭ��`�^h4��~�'��A�堟m��k1��X-NF��R��aN��I$|6w" ��r��išɫ�n�[� OK�|U���\ѽ�`d�؞H�m��?��V�K�˥V0Ь�	�B�b*���~԰!P��)�h��#�����e�1�"�@1���R�����������Y��-��ti�P�J^S2��P��A:�{�y�����5�1o�����2<�ؖo�p�0I3��4��[2�+p��[��N��}ݺw���ĭ���Ԧ,�g�lwn��s��6�5�X#;��ʄ k:�sh�B_;[x4V��^Ϩ�Ζ�JM^оQ G��ެ�%ŭ�K��̅�őaPْ�W	ѲW�G��@w��`)4;?������,� )\pԃ����.j�6� �A֣)>cCjH}��d�f�5��r�k>���X���i;�S_<r��J���`�p)M{�4�RB��@�
��f�ñ�!��e{]|�%m�|x!pujX��&�C��̾0+�O�D��<v�PH�[��N֝��c�q���q��xJ���c� �Ƅt6��.���R����J��/��Q`pѵ@�C��'3�c�OH�=k�HkM}9OC���G���/���7HID>����4����u����|鮘׷�Zo�h�i}�*��Q+
�	$d�F�u:�x�Lmj9���s��#�fc��r��wb��� �E�����e䫚��e��� #�V��d(^Tb����r�do�R9B+��_;3�%$*���H*�֪y'��z�9���N�?b���l�״�|Y��t�"9%rێ�� �q���J׸r%�4�\�u��/�g��X�"������#�K�~E�������QY�~�󁹨O*S��K��4���L�v�(�rJw�Qh��2�G���>�d��
��� 9�O@W�=233~�k��k�A,W�c�׀���V�ڂ�E�Ru�#%�A����3��/n�v�F��f<�Y����ODn�S+�s���s���\<HE�����'��^_ �Rv������(�~V�x��E�(y;��P1�ܿ��K�I��pWF��>��Y��D����j_����@L�EI��r6��!h+.��y`?{1.S�J&$Xb_s��$4|��z�a�=�+{e8�q��ܬ�f���k����-ǯ�ݚ�{r1*.�C�w��[�]@z�z 7뛐��wJ�ލ�����Nuǘ0��q�@HGK6��ܸB���*M��d�����P����L����j:�pFۦ�׃J�[u:���"����c���z����8'�W������+�����Y~�3\\�4_��Aw9d"H��6[F�����6B�C�PE�)ϼ<`R0���LL�*�L��Y6N�!�mD��q[�d���.e����PSw.@���2�]��"C��Ӓ&�Y��õ���).����o���t�L[��3&��_��!����F��Շ �2�5&-)v;O�O�G�#6��w{��1�lB���U�ާn.�Wn]1��-��,S�C?�W�?b|	�2��8�$�8Fv��(�I�`�j�?^/�B-��t��-(,�ak�p�:���t���R;PU��ͯ՚�KHI?%��WH��d,�w�dKM�z��i}N�� �O��L�0�˕���1�ޭ���W& ��h���y��Ñ�P����o���:�ۼ�Һ���:ML(r�;�nUJ-�:�e�� ���SH�� �ϵN��T9�����4�S0U[=q3�}i��kDZ|�c�H8�-((贚�n��rw&�=�R�޿�K���I��N4u����8]��/Ox�0-������ri�I_�5�6�̍u�H��O����J~�B���$!��p���&�*�R�wy�8�]��T���%��-��,��1#݂m������D���#��7���L��m�]v�:8$����q��o���/���X2��F�|��)c�����~ͭ�\ʁZ�DFq��pX۾��z�_1�ջ6?���>Oi ��W�GS�-��c����vv6�@��������a93Y:�i;��1��``��-�e�^kI��ėcV������Rd���J��o�퍺Q���Tr��[ʬ"C����k��՟�&#����Ŀ�?*#�wj�P�|&����.���25	�d������@ l2]A��
\'��o�m�em֝��j+�]��^/��\�W�t8��G^�tFN⭏5�z����>��&s"U���)A�ĒÒ����5�*׫
N�h�VE�4-y���b��"	���~�KѸ�:gU�f0�TaRfX�iO3)�!?[��+ѱ�LҞ|��l>�a;0o�A�j�(D��0����'�\����B+	�H~R��9����)��+��~�Aד�o�x�j(�'d�#����=��6�w�z\��MXͦc�OE�-f\�Tm�:�W�J����ٙۙ�|M���d�0cӳ�U9
�A�VTֽ=��B�g�F��<���=��ș%�l�M�����|�I���3)� 4N*�6xύx��M�kL�l����H"��  ��Io%�3�+�F��iI����
7�� �N����ni�9�Z��{R�y�T��y�V���e3�L���Ҹ��S���+�����R�+���
��{�~4�Ksy.�{'�U1�����U��Yf���`�-i�tv8�f8;���!��}$%��D����E�)������U�;s?)�<O��D�`��� �:�e$f�\'�Q�lG|�m̆f����E��@Bӂ@vR>�{+B� *�~h_�x@�	Q/lˏ��?1��N�W�\��pc��5��<+�5j�f���k�vO�͗����xV��3B�贈�L�\;�3����Ŷ��,�2�S$�$���S���O��e�61�WcV!�Hp@���:��F^�t�{�>ߩ�{�����#U�����4�(:=��-G	�4�5�mÿ~�"���*��6�\4l�~�O]���y��W6�t�]�<=|��!H�!�z͋/���q�\�d�~�05����WI~���Ԁ��y	�P�F� �VEd6ud�I�$��^��??o��������6_�RQ���������p��ϐ��Z����"W3	wF:i��.�� �����6C �V�=N�떚� ��#@�L�:S���΅UR�=뇅h��t����('ҹ��I)�e�!��h����n8IׅU�SxD�%�4�V�L�ڂ��>���r]�d@�e��}4Q|�DD((P )���#�_m����3X�T�6��ό�X�k_hE���[
��Do9�f�������G�5(:�����=�7d�=�$���p��1	ILcΛ��~|n�i7:�� M�;�_��ET,
��?�w�YX��Zj�!9ֵ����ŝx>���!��i'@��~0C��=��C���Kh~sNհ2�I�) �6�n��˕W�vy���ć� 	��Y1�YO�/:���h��Z��J;�B>Ȕ����Ս��'J���;;�<�k�
�"��c�4�j�&F��9G������-\��b��"������%tneTpRu�=F�]w�B
bEږ�Ǔl�dax�cvcF'��W�`���/�	��ɦ>9��j]ܴ��C�Ju�.C����Nx|~֘PB�3�b�k)�6Q\�+z��_����.��A@�ȝ���%}�� ]6�o�Ǹ�8��u`�n��A�9}G-�a�����������V|�?��������H�d��4�@g�Q��F%n�N#���&�����~{���Nh�¬�oX�w���:%A>\^�);�!�6!�3�m�7��7�I���Ya"�?�v�U!١�
�͌Y瀾Zx�DQ>�� f�!�VE~]k�m؀�+H��S7؂���Fhw�1�8��ɻ�S���d�f�WC���J�t�����͢���_!1�Щ�#Q��\"#nG=���r�`�����'J|b��j�f���>�ǈ�/�F�� ��-�^��4 �ѽBЃ��Z����f~��}����	�樲���1YX�41zXrj���m����y7Nl�B�K�����J��s��r ������E&���	`���=�c��i4ᵖujRC��y���{$켵M1usUi����u�3�IR}�
�rY:������"P;?iQ�1&)%Vۦw�뎕5Ά5��Mk�::`ڦw�uC? n��P�V���l��&ئ=���!~�'2-J�3���|��|Ꝁw�;��a�>�����Y���ϴ¡�m1HtC��s� jH�~�[�����{@{�u�ב�{�E��z�+�f�_�6�Qc�m�ZO�=�EKB*�ͯa'��[%�I��Z\x�"E�%�O��7}(v�������8W��TIZ�N�gk8mtp�4��sy��ՠo�4�r�O
��.����n���n���d�?^G��Щ���DXG��lL�*�U�oe�����p�^{��yS����幢8����A��ǜ٥!}R�R�2�J�^E��jD���ฅ�$�� ΚdK�����1��yT%�j+�B��f��57����OdiU��2�
�@���k���n߼��n�,�^-R$����9v��O{?���8n�oe�1d��?=�X��s��.kq�j2�G��YːCt����q,�^��/�P�4���[}􈺄�<6Blsԑ�$e��%�����?%�C�z�+�Wn���n_�5���D�TR˅��lҠI$T.����D�Ȼ�b��5w��T�Z��l������貞��Y��{QA�V1�".�1�p�	�Ƙ|U|z�$�z"H��L�+���:YY����G'��{��+�alt�C���#����,uh�&�
eܘ����]Ω�g���U-��;��eX��>�]$V��%�qw���z�qw��0�I?�|����)�C3x�6�ֶ�lE�@���R�Fv cY��ah�I�z�P#�-dGV��_#�^�	��Hx�j��0��}�M+����~ƸC ����b�����i���5me@�f뾧A�p�����1NI¦�w���(�͆Ey>��øD��6�� �'�U���7�����FM�&ϒ) )�mH��=���7�J�;)h��0�4�Yಱ�n5�tm*��q>>֓�E�J&	2��)�� ^���U\�?7TgjH���'vZ�Y���
HQ���b�Q\�m�-ޖ\!�'� �^�P��:$rB�E 
P�v5�� �L�W��bIg���:�*k�A �D��~�⋞��i�q���#��D��>E52Z���0�����Gg��a��@]��e�����C��:^2��T�	�v��d���>ʘm��A1�		S�ԧǫ�oUQ��{��%>E!�K��@���y��^ݪ�� ��^�삩0���UK�	������]����`��m�Ȋ�oyw�rZ՗G)�:�4���.�\��؀�zX��ؿ/{Q�b���2� ��������{wʷ����t|� +AQ^��ho�""�o�Z�^��:=��_fy"{��xˡH�������X��ه�M����,
Z�J�_���.�-��|��Γ��/ o����K���⠜r���~S����)�֏86 ��RY�Azc�=	c��|~����7�����Ђ���@d���)Jz�EU{�"XK�`\�t�'�<�,$����n�Cܺ��h�W�>{�M}����+ܛ5U����Y�k��U_�΍yW����_�9d��r���������i�+@����9�3'��X�WA��ݷ�x~�^x�08Vuk���^ݑ�U�ɲ̇"#�x/x�ްAY���p-�MAT�w�{=?V�ɛ�l�dγ�_���j��'�҅2�����޾Br�E�]��A4F�v�����j��H�J��.��x%�N���:ι�O��%�8,�q��P̞�ܟ�a%�%K'Xe�YOe�377��y}Rw?]ñ�Z�_�a`H_��]�)~��M�1�D�lif��I|�^�ۇ�s��u��4O�FXxL�x7�w��:�Իwx��0���1�����Ь{�O�kc<�fo�E�YA��";S�¸E�w�����[��~	�x�5:i�n�<&��?5c1R��+��}`��w�mv0��cЗ���JK���a��|;O��iZ��%w��	�^�d��c��)�C��n2��x����10����a��zPVr,8V3���,t����N.&�������R����F�L����Cy��	�Xh!�y�÷PM�m|�U�1Ea>�Uèt���!m�}>;-��|V��N�s�MK�����^/9�$D�#�&�$�(4�?+踩<aٓ�{n���8�`G�ɩ��H�,b�[���'�H�'J�  !����Qe?M��_���?�!��h>�Ɗ�
c�&P�_�+�z�80 ~�S�C��cI^i��r�D���'6'��M�|丙�'�߶1��(�W���'���t���AA<���P�ŵ��(>�Py��U��!3��~_A{���k8�V�(^�Xӕ�&Q-U� $ˤ;���~<VHl3�Q�daR� �
�,%$�5���ۤ��H�ނb�o�����H�w�&E��Z��8(:l�����ޔ�j�^52�/��*��m�v}�����mÃnt����%D�>>�h��T+�z�GzY���6�r�}��o擵�G:���𾋘��������'l�R��El��t���:��"U�@[�*C-�_b�v���RR��e?]F�G�uv��I������'�~�ї�
	i�<z��]ްC���Q��5�U�V��=U�l|8@��]ggu�DS���4�3�2^��)-�C a{��tWסu�/�vUd�w��M�`����3RWU�� ��UՄ�ު%��ts�0%@p^�p4\�g�z��v���r8�Ks[Gő�)��Ȅ��WO������H�He�������e�&f����ͷ|����F���k�j@WvS2��i*H�.�{�C�7�:�M�g�pꍴ�6��s�*=� hj�i˝�:Z���Q�V�$�Ya�{�\(�H�b��_��c����([���H�<��Ph������ꗾ�����Hg"¾�����(6��d��)@Dy޲�︫�.2��"��n�uӹ~=���#]"�B�\�G���.<�H��=�1O�,�wϋ<�D�Y�4Œ�3,�܊�!�H��}���^���5�6bǿGog��T��z�:C|�	�O�`��V�`�
N�U�U�4��.�s�m�� ���m�ϐ>��,������S�x�턗��=C�h!5/A�>@^6�>����$Rk2u:�q�������6�-��=9�����9=����u;1$~uG�����|a[��|�V_(:h?+G�U�F�]X�g�i9���[t�6��(��C�27Z��k���{}ޟ^q��>��͹g�.�|�w�8+�R���9�<������46v���"���K�r[=MC~9w�~5�^�!S:��d�a�ǣ	�����D���=/&
�\}����8K���iz���'C��Z	�ƿxn����݂'�K�I�//�^ۂ��t�����3�$�we�=o��f�^5t�Z֔�?�N�8�����zX������f��h�gǘ�4�I ��~�Y�Y����6��h����1i�Ƕ"_���U\�m����FK����Yμ��@ҿ�xv4"`�[Y~>k�qw�ez�3\�Ux�������=����)R����`��N��߿�@͵w��KTn� �W�d�[���L7:��I �cX�pr}�f�F
5^f�ZX��8v������U����*l��[.�������6��`U�|�;7'M�:B���w�z��k�I�<��֡�V��M,,�_U~g)_��C\�\�2I�z�R��*�a)�X�:���ݸC|.�$6��{p�~7P�L�Z������Z�{���^��I��>.��{Ȳ � j�lv��;��D���5�k ,:��wҮH���}驀����qg�h/1��K���IzD����&�n��J$�(Y����b�&�ت3�Ƞ��`�s��co<�_'L�/[� ��ʺ�7�|����.]un�a�.��k5��ry�T���;��� xtA���������xQM��f���R�in�LcI I����d~47Vƫ;f~�@qb �����P��b!�+N>�ീM��&��57S_CV��S��!�ꌦ�ؤT��6��Q���|Tb�R�~��ȗ6�pN��l<f�|ph��(^m�����-n�~ֳꀩ����&m�7�[[��އ��Z���
�a�p��E㨞�[���ā�ClN<1҇·��n�i7+M����@��y(ڻ�/�)EJ;�s@rtҝk&,2 �߭�L��n����b@M��ï�>��n�D�R�>��I#�Qr#���cVeW�B�#%�6%�[1���"��D(g$ײ��� ���O9Fw1H�֥�r�ww,�r6E9���kQ/�<o,(�D*5a6��W����6�52pe�K)Nv����C�}�A=[��"N!Ā;T��+�55��=����;�@�`�����o#< ����;��T�%٪����n��[�b��!{��2C�*}���2����~6�d����)�^�w������l�m��?�C��x���-�D#��P��۱�b�Ā��)���z�s����FK>3����h��=W�.�k�^�p�8�:��&0�M8��&��'�J'�{����m���yW�@���L�);K�����T����1�Й����ü���%g�DE�)$L�W��Γ!��x�X����S�ܻw�O��	]�A�/��ah^�G=/�5�}(��qEX 	���M/Hqj���u�*�Xc��h���Lx���Q0 ���t�!U;ض7��iӫru9.��2�0	�|�T�;�'{w�6�'�Wp�	H���}��pp
ј�!W7���]��C%�����^"az(��/�I�z�RKzU�~�S�@�/�w��%�$�Z'	�~gV��~��������0����(��+y	�⟋��w�d������c�ƌ"ͨ,c�~����5�������FKVYr*f���4v���?l)1XV"�rܘ�Q�:��|�R�W.����럭�r�1C���ɠ�����d�y+q7���0�d�E��cP��8�:5���^��D��S�]
?�q^㓝|���
�K�����c\M��0���L_w�~���v��]�������ﺌO�Q���;�F���M�/���Bb�+�����7)�Z�Z�E5��K�!|U��<@x�7��MʌD߫ՎE,�����R*Y�(�>���&A��2R��z���Y��M?\�0�>��:�'ö�aUd�f!�l�_�p	zE	O��,ڏ�Nu�=�ㇵf��A�� \�=#��V%D7d+#�y�y���
�K<J�������,m11&���o<��lＧ�";b�^��~��DvI�i���+t46P�G��SZ>!��K�ݕ���S��Re�Pb��ڟn��V��RDg��,�lA�@��3Z�j�����pq���o�NI���C�.d�H(?�E��f��Ju�D��lA���`o�R�l�J�`�tZ9sI�f�|ɣ_������"s�n6'�`l�I�WT�FFH��,�J,6ᴗ1q��jf���xe;R&9?:e��r��=:�IK��o�!��|�
��9-:�kϾ2��@�a�T��s��7r�oem��įB���l�����P����{�9��~5�1����h)�Ob`����U��[�_�d$�S�d�Y3��J�4�νs�h/�OH�h��<�'�[��M��yr׸V��N?�t��ѯ:ND/�b�Ɍ���Fk����a�ɓm�vM��l7�5�v3��ɶm۶m}o�������9��>��s�;�J�0�O��p�l��WD����۳�TX/�ʕ�À_�^�'m�5����"�*9�ۛMzj++�Ê��h!��#���@&8��X�pV�?K���SK�j"џ/���й�.�(5�Ld-�W�#�Q���zT�	ain��xkd'���޼S�[�!<�LUW��:"-f�k���l�&&�:��jF�&6B������gZ��	1GD'I��+S������J7����|1�x=�qv+]C����1�fm�s���35���2s=����#7p�2
6WI����o��@��PVĕ���D�ћ}�;�:4 a����h:��i~ys���p�|���)ആQw��K�ywީ�-˟=
�Gi���������B�k4=K�J*T�z#C5rcva��w_�+%+-#�T�Jpj�ֽ���y}��Zg�gc���l���Plad�s����I�D��K�����om3�=L<��X��^�p�g���@�rn��W��ߨ[�8_��1�\f�H�^I�;9�|~;��qͥ���A�����]�1���o���������~�� ��D�3��HI_�X&1�3�Ȟ�3�U�8/2T2Ʊz�?e�-;���$yҳ�Oez����-��I��;hɍ��&W��2 �K��Jǆ~�0�c2��H׀�Òƞ�,�@��\뚀>���g�¦��?k��^mD���
t�u��u�D�?����PhW$� ߫�Q���d�F�/�FzKk�֥#�ùoSCxAM~ag�->lby��x�_������Kq}��ݚz�S,+�:,eF�B��u�3d2�J�a+�8�f)�YZ�7�u�_�IIK���֤���?��ͯ ��w>��@��c�)l���EZ�e��q�q�v.��AO�hp!52����良���J{A��'�����]� e��b&��:���>RƓ�0�~Cu���̃���<2���Yԏ�m	V-we�i*T���?v�R�1�ǂT���Uۃ ���x0A��9aM1Tn��I5K������*�P�H�v:#��&��2^��۲7��W_e��#������#?�]���M�[=�ZZ��kd�nk+��/o5�"�m?jݫ��VUÕQ@0D���S�(�&���SдT͸�^ZissO�U_w�R�>�PTePq�_�
����TA)�)�S�Q��B�?��`�&�1���b�Wt�ޚ�k�1���p,%(a�Pi������S�0B�y��{�|����}u�l�d>ɂ\���G�2�P����m������i�4_��B�L�I��5�H�� �I~�ع�0ʹ������ p�o=!4�n_ ���E�|�?��g��Ƞb���3�,�[��7�(\)Q��ص�	�
8F�-jN��O��cyPa���>�9}=.�ڥ)�(~62q�O?���`��EJA�U�i�̥�#��k���<<p�M�r�����@v:�{������6��1��ݾ�8�t�3��[^�	�V�'�0m!deV��H/m�� \楩��U:L�{r�XZ���4���CUk�Wvr���@��~���j ����u��q�
� ���KG�\�?�������Z"�j��k3y�ڕ�`lK� ��#�*��^��.g�ڬW�1�����:?�J }�ڹ��) j$G5ZOfb3�~k��
�@ڃ~���u��a$�H�};��$^����f)qȍ��+���$4\����>���h���S��d��T�oo0�fO����_�w�乆�C����1�,��HgΩ�l��^�A5��,E;�����_s�x��ɛ�T?�$�I�5�A��x������B��ܭYP�<��m~�J�T#� �ֿ���6�yk�A�o�x��w���W���m?��d�b�n�/�*_So�z�7*����tȂ<�/uݙ�P��G|�^�W�Z׮��@O�q���l�&�s��4���M	(�r�J0����@��,��ƹF����������Z���1�Yė��`�V�,L�v�h�Uk�߱ �9� �Yh6���i�yF���Hw�̨e"Ob��ά��;��\:=�wA�v,זvS�I�M=an`�IⰕ���%k$ڊJP�8����������i�xx�uQ�U���x�	ꡠ����6#��N#
���e��C��ً�$ƝOw�f���&Z�2*���r����w3��D��}���(UH�Ꙑ�k����r,�"�gl����{?*�*��^��z� ��y��{��J��Ğ+	dQNՌWw��<M�\apB�����𛊔i�����v][���])�r�����7|e��SPR��� �%�>D�0(�����!�}��.L!����z&�X�WJE*�zfŹߡ.<�_ID�CK<�PF�f5�{>g�r5��k�B�Q�H��εP���"ĬW'w�R��i^�b�F"XC�~^j����X��,�0�`#h˂ �J��W���Z�x���h�%�hy3�H�(pX�D�lJw_�C`�|*���MO�@�èoWЮ��~Q�EKw
��&b�э�G�p���ӢDj���R4�Sp}��v��uR�u�:�ƿ°�K�s�a5D/�b� q�%)uN��8D�-n$ww1�`�D��v֢�hc�r��yP��Ӈ�?�Y�	�	���~��~ZO`��[�w��R��:W����O�ʩ([r��%�bȆ��P����H����\���R>��L����s�e���W�Su�����8��7�#&`9jh	��3�s�79T�<P�����R��X$���``�u�2v`<Ю��H�������ҧn�B;�<t8�E�0pp���U�3�q�&V���ɟ3����[����U<��E:�
�P ����|+p�YMC����	��+�5��C�
��#�p/���[wB@�D�7`��>�Mz3ڑ�J�-��͔D�,�3���\��Į'��pI�|hTI)@u�ZHF���/��g���Z7�fOJ���iҸ4䉾�lK䨷\� "�=��[D1�?,�Ϲ�`IRAM�PPZ��%Q},��� (��|2���6��&��JX�#���%�����'���;�O��EarR��3̔�@p*�41)�������ѯ�E��������-@�\�K>71�y�3^��v���/��u$:*�SV-W G�����O�6{M|[8�+M����L*t
ۯ":�T��?�n`X���a��k�;��(L�-h�N$C�H_w4=�G ���<RkJ+P1N̄�@����Pi6&�|4����\�G���3v�k�OfJ�03�B��Ik�S-g�V58���$�)}�,�|�C�"C�iP��qT�`ac.��R���ù8�����J��;����pm�WB#t����o�� �`P�M���o�t��2K$wF�"�~S�r:� �Y@܈ ��"�|��'ΪV�Ց��4��tn��K������,#y.��M�����F�e� ��/lJ��c{r���(6�O�6��!kOt��L@e ��C� &�*W��貨��W�ƕr7����Ud�j+�������Y���_'�f<33lh�����R�*�(vś�jq��&�F��ji=�[X�/�O���q�a2rz~�~�~���� ���9�x����?zA���9�����~�Dw� �����mZ�S��y�<_'�7I��(�)�ԗ��sD#.�C�Ő/0��������RD�_�S_+s{�٩� {��/��D6z�#ű,`�%��U`� ;�rx�_�eŅ9�[��ȥ|�%۳c.�(#���D�Ne�Q��S��,QG�"���t�o�D��"��rʫ�(�t��Ш�1@��O�W�$�G�!l�7�����{��IΔD��L�-x�v��4��̯JʝJi� ?�6bP1� ~�7-˪�m�E�{��/#vvV�v?�$����rbM��,h���E:��̍��`�KPFX�`z@f�V	�dl��b�iR�}ן/�Sȉ�WC�s��P�(DlY���i���h��N5��U����2�� �1�A��7Dӗ�g���5�/�����7�͢��'��A���]�8��ύ���v�)���,��3�ൖq�,�A�6��~���@�㍫ƍ��!�E�mxc;Ig��y���'���Y�)��s�Н|���pr�0d��.����n>���0�P������ȷ݁�����I�P�Ћ�8֐����;HI�r؞ڭA*�� z8�0��A�����p2Uh�Ά�:��{T�f�]��E��i�&Jv�,�q`D\�?mC��K4t�	l~6�]����������H��+푩��Ϫ,�V(��g��k+�od���XC̕�R)��O���Q��l�j7Cc�ߎ�o���D\�k'Q&V�!��zUQ�U�����A�:���A$�P��D���>&�&H�㐰�L���A��|\P��x㖗��i��uJ,���4�D#�,J$����:AjTEFN�yd��͇&�JMe����lN��a�d����<�3Ձ>�yGw��aIuB�vG���_<u���nʰ�� Kj8Dǈxj��&F!���Օ���tD���C��D�>�	r^�.�Y��WpvF��ΔOg��!b()�k�_��iB�{��(fYL��E��\B��6<�/p�_�tt=xng�$J �К�U�AAQ�%	�t��+��l��}o�J`�kf����~Ɔ�S9
`�yd�r�錓�f�]]Y9�&�$����}���C^F<�8zd�Mg@�Hl�DΟ�zA�2�����f-L�5��l�}8X-|:��=W�J/�����`���$�	-8`�expN9�4X3BCW����o\w�o\�TJ6�毿=�����Qe�9OO+�ܱ�8��F/�`��S��2ߢ��M�F��H+����ۡˡj}8h0^)�.K�<��l���	�6Qr%��q@,��3�w$���"BlxnX/4<�ⶃ���W�L�V�؝#?�X�isuJTL�0�Au�A���f�o�Շ�kRҬ|W����^�:GK�"��Gg����;�P��s� �S���s�ZL����ƪ�o�,/V�����巚��.5�Jx��M����Ɉ��פ2E+d�����i|v�cD���A��}�|�6G�"���".�ڟO��M}5�������ڙh�Z����L��_�`�!29Bh��p���(�Md;���c�+4ޥ����pO��󒾊T�(�f��g_@7��Kg0g�б�b�j�R�*}��#�,i�5>�T���46�ʅ`�x��9: ���=  �&�K��+(9���v�̓���l�u;�-d�e!K�EM(@[��/���w�/ ���	�S�2"��_��y������oLTZ5�j�U7��x
���uq�>iM�@�s��TU,�m�R�q4Y��I��Y
�3v�k?c��0D#t��2�I�����0(h�@@Ҹ!J��V�ɦ���\��4 �_'6�� 5���%�<�"!B�f���G �&vh�z�rāOѯ�v={󦺉��A&�X��7�u���H����4�陷F�L{���WɈ�}��x0���b�v̥�~L
T�T[�R�7��P�"��	��4���F�և�Z��z0hg���Z����$Nj-nU�Aښ��@����ǡ?p|�T�'�t\}����vka�K���;8�p�t��םy2��~Y��� ��B����	j��5o/]��&�Vr�	^��U��VsV����&H<��2�U4L��������/J��8���JW0у>D&5�cp�n ����@�s� ʜ:b�Lc��$Pl`������\�ڡI��R9'�����ϊ5y� �O�ՙ^%��t3��#��`_��n�_XS��@9/D@�!��6'�����*�u;���7�c-�Q����w��$F5 ��h�%6�jt���d��q�G;o��E����I�ڳ�ca�<޺g�ƞ5P ��~$6�N"���n8�X���9�x@�w�1�Z��
s?/`n�FU��T�Ĳ3�L~�Y$�pP�0�W_k�Nj���Ν_1���G�gj��3�)\�O0N�I��0�Pg[c���A��!�P�Hz{ �,d�PQ�-�j�C�oi*�A7�Z���$eD�� �Sx�4�G�9P�P!A~5`N�	Jin~��P��v��
d��WKВ��MWKP����b@��Ej�a%)%�Q�Qe�%O�N��`ҭ��ffl�z|�&�S-���4}�
�3�&,��V�%#g�'�4�e�D���%*���['���p�#Z�30�ޣ C+����\����m���eA�79���j��|�
&�5WUj;�4��2޲�7�Yv�,����y߁s� ���3.�2��oZ��<b����ZVLyI�RRr��ގ"��$�25I%��|�A�x��RV*;Պ��g;x4�ϑ�]�j�+9QQd���>-]�L|e���A�5�18L>k���4vo5��)Y?c�;,{t0�zb�)}v\��u5�$-Y��b�n�۟(�i��x�1��%ZJT 1d�%s��Y2���*��e��i�R�|��˄!�8jC��ha��Ѥ���H%���b{I�Rx�."��M٨-�r��=ܕ�Hq5T�g���]wb�N�$0f�_i9$���g��^������&����Ь�߲�Sq�a���6q{��ƭ�\]��)9��\C�ja<~�T��;�\NUxrI��E,9�.K����Օ���!�q�ŗ;�H��~M��̟�����#����x�&Y�u�=,F��.���"&�d�HR��!E�~۷���W����0���S��[q�t]�.���J��i,E������宫$#w�0�DD(� �f�e���ݔ��3!��B�� ��^;=�gYӞ����R/�.E��`v�-��q��c~Tev>�&��4u! 7�}��n)P��+��Rbm`�?��߫���]��;��w �f0;��b��M�����v��<3�O��?D��!���*�\�S��p]Of��^�Q�����4�3у���N�F:�DI͏�ؒ���*A�֪#��)��v���/��ԇX�V!�V����p�AuL�2Δ�
^{a4���j�&�=��6�'�Oʢ:/{B[�Tp�T�I���ilc��`7O�<��YD���,�yl�I�*��_Z�rܯ*J�Z��:�_{h^RhS��9Tp���4y-����DACpi�=l��|�⸎�~�뭠3~\�����9��1����{��9��l׬c�[2H6�<�:2��ׄ�#7����!d�K:�̉���<�|�RN�V��y�OE�o�e֢�(i�3�8f�}&��K�V1��PX��|�(�3x��"�g �o�P������˫�_kϯ���(:�/��b�E�_"���A�%��!D�w��D�������S&�����
�Dﹲ��<U����SM��

oy��-j�:�{c׃�&L��=�WR;FFE����7��tf
_s��\{mWO�-ߝz����t��O�R1{�7���޳?�a�J
AA���ZY����%�����-�����3Ft�Ig�h�.{�bݴ��*�l���z$��|��߮Y�����[���K��kt�5����&��b��r��b�\0?;�8�Ѿ�E�F��7��.�f���8����LV�L����#e`�{�p�ݢ�<�L���F�]�����}`�����9Ű�֊�+�:%�dO�l�����ٳ@$��<6�&;�����w�h����^���T�����(��S����
4��:+:�Z��,������ʦ���g�|��J_玓j�/�VP
��~͌|ôU���^x��ׯ2�.�Rʺ�����B��s�TCs��>�uD]��e�\%����T�]6���H^�sp��z�<\w�/8���!��q)�e��%�lLh-)so(F���w�6&�:�4���D���bjA:�&�#����Q�m��̩'�/�I�F:"�[c����ĭ���H��j'����]�����L�VT�;��W�B�sG1?~16��>�� ��¦���Q�w;�1�G}y�C�6�_BxE��ȏ{;���,��i4%1=u`43����7�ɕ��s#f�$g�g�ϰ4l�I����L��*�Z�6$������mST������\�v��i��/���|7�h��iҌp��D:�3�%�b)i�%��p�r� K�;�6��e�}X��(�f.��
jis^���rep�c��X�����te���?t/2�"/���4�g�Ǩ�q�-<�'������]�#+!C0]�OM��ǩ	Ƴ7�İ�����<e!��;���9:��x�Io����{~,9��SHx9�a�\
���>�I���v��!�G������Y�|=D��!�{LW+��?3�_7 ��&�s�"������
��������n;÷�wI���GV-ٵ��2�v���.fT������]Z��y�Cj!�w��h1��așiO]V����V��E���R�������� �+�w0'm�1b��4����g�w=\{��h7�hq�*e��if'�K9��V��uC1L~A�R��k�_|�c�
н���9m�+@��:r���6+[����/��}!�X.:��A��
����㛔�f��q�IL�՗�����'���&'��/����Z���U50��b�2?��ͫ)�l��m׆�=�ŝ��0���_���~O�f9~I,&��[��&��#3�U�nb���)_�����vQ���������d�/W�~W$GK`|�j��?u�0�ԗ&ޅ$�H������^�k�Oшq5�靆+�)|�O�>���h��ߧ5��\^!�{}^����@sMFG��׼cR�⭻J����<�,��vK��y:���,���un���$x�}��t����!�`�7h����e~/o�?��H��.�Yk������=&~\�YҀ��E�A�A���}�K4��S�&��� P9�E�%�w��f����G]�{���u�a����B���o��o�Z���Wh�D�����r_"�+~�	Xd��ߔ��@j���/2���r߃ ���<.E�3ߐ�3�2�o��ˇ��G]�)�/$)5�s�ff.�4dgJ_��'	ڹU%5��`�m��+4>X�����mi鹿&�����wغƺۧVu�SH{6�i�	J��F���� ,���NPE:��
u�զK�	.G0�^��!�oC�5���_	���}xt����+��(���ӝkV_�B��9Ԫ�ɐ��(|��";PW����k?n^0��ςZk���o�:��"��:[�~G\�X_�͗�+��J��p�^��*��k�Ǔ��޵y���^.�d�S�)=�Zك��ѵj��P��)6��2n����Vl;(��X�
��q��ه�	�ߵ�꟝�O��Q�v�L��Yj�5��iϖK2�x!�6#膺�ݨ��3W��Y��K�A���+����si
�('�B�֏�  �ܐ
�i;��{��G�:wC�,i�/NA'�H,�?~qD��&�t����..~��;������enÕv���V˙��=�t��V2��(����&���gU||�+�k� ��h��5��(��{杋�y�	}��	.CI8f�|�W?��K����"E�Q,�5T�� N�������֮:y�͔��d�LK'!旸���tT�R��c"��lvV�x{�*���Z9���޿:�l��a��ۦ�
O��Q���������c��c�J!a����bo��d����0�$9��ʞ3{������|��d�OH�ۘn*�!�ET�9�UN�}����sx�t�LzS��M���Â��4O��4�.��a� RpX�W�Zf��o�C5i:��u��-��3G�i	��b�+�Y�-ec�����l��0���v�೺c�{K@�	^vrΗ\��ZP@o�0N��8��cMm�)�UL��~�����暢PJ��4�VT������r���ޥ4�E�����AA|�IJ�ү0�2}ʌ���/��h�gc������_$�vG:�L�&��惡��̃��G�>{��>w�8#8[�&��H��9�3L���\d;���1|=OQ�A$bg_���t!O������W�}�Z\�.���\�
��,����� ����H�����6�Kz�a#1�ωǚ�/�^��\���\�MS�኿��A���<{����+�����Y�ﺮ��{�xa9��f�_JtG�
==��08�"mh�D����"dNKà�x�(�Y��&j��[�1�{X��X�/��������o��;)ԤX�	�x(�"z)k����LC��%[��|�2�x����o�"\�s@gӒ,�;4��<*�L�1\k�a�E}���<�3\��u+�;��SGz�V�����jaZ�;ȟ{������Q�r��@��F��"��#$wVjd��No�G����j�G��+>��/��k�7��gQ<6Ǉ����ى{�������x �@���nXx�O�T��Tg8\�P��kpxL�T�<�%0��.�����`rs���4������*.k<w7�q��v/��g�<����M�2&o#�_�1�d�u�A��ZD�K8�y�h?��L�2l�wL����ϗ��|쏸ފ���bA�"�㹜����<�<���Ȥ;Q���zW�U>��s̀���պ����ȭi�+�g��a@�Eo�m�-C�5�sC&� �l��=r�w�nwd�ũ�7�㷕��_|<f@�j��xvĒ�*������UH�S��g����Ǜ�c�8�6���h$Z��li�N�+�h�ɫ����A۫�j��UYA����&�h��x1��H��v�|�^"��K���0/��`j�FM
��Y��k)e�{�)wj�}�~;/�N@���ҫ�~�;�_+M����_p�F����+�J��<�8G�����z| O�9@����D�Zwh��oR��O:���Za9RfZ����{F���MT�l��� b��9�8X_IΤ�>��|��'&��_P[�%}��~Vz	��f^���xi=�s`���\˂/�H��1�6�A��/�tP=�	����TO��
G�ʼԏ��{q0&�cJ�����jگ��\����{�6_߾�B{�Q:&�0�gWP�^� �`Bx�OR	��Ao5�8��h��z��/��C�����CG��7��w��6b�Rn��Nб��<+j������CsTS�#�
�xA�_�)Xu��3�5�y^�$k�n�=�Ӎ��)�y�)���T#)-?�i�|R�JZw$Y�&[�����@5�a'�j�T5�2�
K���Yz��Zv�S��DY	E�X�t��U�$�G�:��B̬ܻ۴�<F;QT�A�����A�Z�^��M-��z%���"�>��,�Z���M�Bj����O���5�0RMX[�j�VZ�'5P7���^�8.����>���V�����b}��
���.��۲秘x�� y�	��9���p���0�� �a;��KaN��F���󅞠֮�urfs	�RF�މ=�&��DYW��t�Ѷ7�O��>0Z`�9^�� )���ע�tL��ǜ�onE�1*�����6���HY��Ϋ$��"\ڙ�d����7�l�6A��(�-�Ym�����m�y�}d��u�Fg�J0~�̉��J�V��1���-�C%�i�5=�a����Xb<�yln!��1��������h3��7�~��l�&��ӵX8a�\�gc�Hm8�Z:�>���Hz^Q���_�V�mF�� }����Sh�B��U�09|�,��kkm���#�y9�O�q;�]�@"x��}�Tr0{s1�;���_�0�vL���|uz�O~�tKG-ݯk*߉�ͤ��֞��~z�!�e+!8���>i3���j�:9�����6�y:���G�}�
:��qw'%}*�~�W��NUh�Z��0�=������2���pZ5�ݜ�' �q<;����si&S���4ToI]�U�z�(=o� 8�^�b���iHL}ɑ5�[�^ae�Q�8.2�Ъ�dwD�����DOy+��������c0��ƚ}ri9{�I�k�����,`�f��5�9�<��.C��<zc��o�z��(�h����<����g����C�\)͢S`6����>���U��d�@�%vs-�F౾�I�ZD�0A+��?�2�`�}���^�	V�3Vl&���펄ǐ�x�� �k tTD�G�Pd�����T��S=)�\�gq�2��B^6����������]��i|ҧ�nq���z�3����G��{#߬�
�o�	�p4��n�m3qؘ��N�W�\k2��.5�(G��X���R#~�2N+*��nqp��(�7h6Ì9��W���
�ޣ����+FV3���I��v0��
��N��`�3�	N��雅��p��G�BI��`���wȔ�t
2Ԃ����?�.3��5Wa������v��<���L,-o�ʔOo�@�eՊ��D�%�{��S�ٙП������/l���fq�c�8XiA[�:D��l��v�y|��E���ܖ��FT<�C���o����A-��η��Sll�����q�������L����:6�#>���6��<c�)5b�őxݕ)bΗ�Y��n>�	V�36����5]^��u�Z�&�߁�Qw�r�h��_�������lbq�Y�R��J5Kr����}	�&kE#3�"v������x�<�q�\b6rf�D vq��˵�*|7�-��������z6���$@�#�mh�h�����΂��'x��Ix�����?<���Sq�R�}����mʉ����M[�:�]MEP�.��Tq�K3����	��5����#+4YvF��^�~��Wyy z����&,+�,�`yc�dA�v���Q0�-�[�2�����N&;d0�����q�-E E��Jb��P0�q4�����S9�Jŵ!"	�DP6{�?
�\�k��`��~��y������;�"��`�PWHHE�1���Z�����Lt>��C SI�:��!~���� ���kK�/��h[~sw5�֎\�T��C����c+��0���7��. ���:�9�mЎ��>�ײ�����h�s����;~�� :��	�M�5�����yE��3A�4&[�sTmx2��9M������AP�t�[H�����ј#�/,����)����%��7��v�#�,�I�;���۲>G3 21#�!N�a8���0R��v�i(A�#��#�ǫ�>��8ݑ@�?�Ͳ�����G����+��>�Pb�������yN3P�R�S�o*����28I���reMϽ�4��0���H(M�^K*�  ��b���cM�/j�8�{p�s�T�6������k5���}l]���BLf���6��I��r|O�ļ-),>⡷-�߇����5N�#/��@~��Й��ڱ���$';��>��Z���Z�RT��@�4�_����&�<Qf�C�>��28��o��Y�7�E��_����$��|��+�^�X����{G��֫�����p=����#F��{,����g�/�6HlϬ��敐[��m�}��]%=����k�/�4\��91�����d��ԴT2/����%ɫ������]��&Lb����q|��C����O�o�>��%�y���y8����a�0t��++g�6s�k ȯ�n���p��I%�/
�q� I���J�.<<[V^I.��c}��,D���IG��|f�*kͽ@E0?���=�1b79��?c�P��<��.�5����<�=��R!�Nɵ;���n�(6�'Y�T�;�r�	�
�pS<+_G��HᣝH���L7u�d3��j�����y��Mh����s���.��Ј��Yȝ �nACӧ��]15i����U�n<!���,�s�+@]�҂���Q���G�SƴŁ'��̮�6q-bj��qUp���&WB��P��	��� �Q�3�X�٧.��D��F[���x��U f�_��m)d
�q���.��� ��\�>/�W{�9r��|��k�e��ە7����� �bnBS�#*j�S���i[�������k�}h�{CtǾ�-�z�סͥ�}�󤙇ˉ�C>�H3��
���jO,0½���M�|D?8���F�ƽ�������t��>�B�B�[Y���������g����	�u!��_�DE�H@s�.�z~�N#��dG��fдQq����O0hK���k�>n1��z�p��ٿ՞����ܒ�|f���t����3���0��;�]�`�t=U3ST(/�'F�A��
�K�BY#lS�ZC�Pʖ1���&Q�7b�*b"Ǆ��{Ol���
�8w��F���@�{tGN�f�EyweP��C��#��J���bT�����?W�t�{�o&�#���O+��_C��3�� s�ˍ6���1Έ{˼��J�F9��|R_���ڮ6�_{9T�{���C$����6q�5�i*��%(WX>ɳ>"�ˋ���BQ��4O�A6_qGL-�,��d��,f-4���z�@Ïך(��H%'f�΃�ܒ@	.����\_	v��μ�j���RU����a��w�����B����Y�^�;�X+n&��ࡠ@N�N��Ԩ��
y�57r�.����\�3�j��+U��7^=�=�A?�������!�!����n��K��p�m�4�M�Hb��[���P�e(����{��$ebQl9����S���?_�����w��<�(+3�JQʠkFyx�bl�@W�R��Ⱦ��8�رY~͚	�e�K����$9�;sځl�PM����Y��(f��UHA@@AG�=�Ta��t�]�)�y�%� '(�:�O�f?%������7:cN;��?�\Ŀ{R穴�g����>�-�-`N����ةc/D��@�DUJ$x&Cy�=��WqA\��/�(*wy��/�[���,�7h#�g�l�7|��ڊ�"��V6�r;�"���p��#�����M�%. �_9<v��Þ��~�,""+�@_N�$="����9�
���:|��'��٪ͪ�!i�w�J�������6��%xѼݨ�9���nk��j��)�=G�ӁM&҃}�f�0q��37���`��O��v�Y)�ѴjpG@́�P�۳�<�/r��޳ջm�֠�k�u�i3��Gv9@m�6�)��Xh�L�+�Dsv/4���3���U�� ."&�z�p����xWX�o�O�(���dy�~�"f�I�
Ҋ�u{_�J���������Is�7Ĕ�
}��H�$�x�*�J�����n�qop�$<� �ٔ��3���7�d~vfPG���<�F� Z]�8�ޯ�~�^*܀}�>`�7��^xĲ}P�?��7R��p�+=|�ǔ�%��͂�K6?��%���4ƴ]�#�`���X�L��☏��5�=�.��g�X����}��k������w<~tF\ݗW�F2���W����6q�Ap�&�7�=yJ��*=��,eHs�@��=����c�j�gi$y&#9����;���~���:w3��n��m�=�|�T��HK���ͼ�O+�*����$��5�� ��`��XXG���zp@UY���i��|�u�%x�SeD�����/�Hm�"����O��}'���$��p}aq�>�	 +����]��%N����A.�v��v��P�X� N3�G]�rb�B�{ �K�:�x��?��Q�3Ģ��a3�H�[x���5g��"a�A|f��Xc�Hd�B��k������m���+_��Xe�;)k,�,�T2�7�K%C�mG����ovY%jV�W�-�,���ʄ���X��L�g�w��p�gV���.%�^\�
H�C#U�(�������*��A�2�����?Mκ(`����#0��|�6�P�Q~y��#ث��;l��K?��튂��L�:�Y5Y��=��5� Df/�v_�����}�k�!:7��@�H�JB���a��C���~4��(#-����	��������Z'�9�����)�/�Ct�)�$V���v�/�e��=)خ�׊O �x.����;4�!��X�!�Σ��Z���%��s���5�!ɣ� ��/�5��O�A�rX��t1⦢5��6�c��@���i�R�l%��uM����tSihU��z��2�Hr-�2��x�K`!�:�z�F�^�Z@eO��ia'A�cզ09vr���*T9�y��λ���Ͻ"�twc+p�hA�sBr�׋f$��zq��=�.
Jsq��k}.�lg�@7�R��;/[�fmp�/(�e��G3�B51:�V2��VT�s��;�ɥ`����m ė��=�6�Q��>��P!��3V��4Zs\���~�ek��-���lc�e�^�m�jqY�6�����>}~�ߟ=��s�s��λ��\P�v���!�{"@~jv�m��X�r��K��8�\x�"j�j6�1@U�:No\=j�<��?O]����\E�I7ƺ�!���O��I���٦�`2�+�v����[�)?�T>Ϻ��@W1�&�ᓥ���!]}VF=�������=�E�ZFs�<4��)�&Dm�W]�7%�Y�l3r��O �|w������Ч�	�Q���@"Y�����R�`70�5�O=���dm#��H�:$�anR���R�����2Յ/ʷ%૵�(�B2<q��h�BiO���E��s�Sf���Α�(����
Tɴ
�p~[��e�����}�V�J�K4��A�Yoq�����|Q�ذJ�}�%�ǬWA%�@Y��&��0}ȳl?1C� ehK,{Hw��J��D)�bh�.)̀�O����~��~d3B@c�=lޭ����ő�=�Kߜ��]Rz��r^�)��	��au��L��{x�'�_��Ã?+d�������]i��P=�F3��C4s��#|��Ȃv�A��}����cXяO����[�9�]��HԻi��	=��?�Í4�RΕ��<{�BG��j�1$7_X%4�2�c�|��ҝ\�0j�O��Ӡmu��ev"��� ���Һ:|�XG�騂FLC�'zr<%$,3�ɢ�\���$J�Ab�K����{��y,ܴp�܏��2��yGH��{�,�	��9�ޯ\�a�Xy,O�hj ��q��p��	�-X'Z9r�D	�.�m��-"�!��:Y���ۏ, ?���2z}]�~V�6�D�͗�Ì wmP��6��8	�I�Ds����<]O�*�k��]�3)�(�d�!�Ň3ˢց���d�
2��=�Ek1��:��6JR���7��Cb�O�uc ���j�%!�j�\����_�>�H�90!��T��z�U?���K���D����z/x�;�ڪ%C���LEZ�߻���Y@>�eCW��q��2#{Mԇu�B&bуd	����GЃ�>��x�>�X����麲�?�МO#yYz��`	�dq@����pWM���4T�~�h"
�Ĉ A��l#���P(�_|u���'��1���ԭX,B�J��\d�G��b֬M��LL��t��e=�h���O�_@%�g�dHvJ@?���w~�Zܪ�%=%e���`��Fu$�����̰�w+>q0�]�ZU�{'��uQ�@Ww�d����jA�\}�q])Ж�x�q.ܘ�>��n�=Ϛ�_�a��`�U#�:�AMw�H�C���3C�r���?H� �[}?e�=���Q*��>� �!4zf�Th']���{�GUo��''�%���<h\�4ȱ#�][�%/������JO�H�Pd�Ē��g3�Ϭ�m���] �gI��lt���;!�`#n	����V�ՄJG=ܛ���C�t��3�&��`�(��ͪ�,���0��nHK��|3�5��O���1�c���	���Nb�0/D������K+J%[�Q}��S�?��$�d�l�`6���g��H�pD?ӄi~�c�_�ÉB���V@RV&>�)�s����Z%/�x��
��{1ՙ�:m����M��gt�IR�8P`�odC�(MFk�Nأ�R��l�m�.��	�r�R�bO�-/]R�6=�E�	��p��d�g�RG� 7+�B�zInv�պpO�W�îv��$�W�~����Mb��Cd���d׽�T��	yZ̑����{t� ָ7���X��a�v���Ui-#�52S�v��d��)����䏀K��ʏ\��EC0����Cb�E/���V��8Įub~O!�X�]y��#ĕ�٘�$P��/�h����֚F��X	����׸��6�
�� $��Ѡ�� h[�;;�; ߀�������>-��)�S��ԇPRbu1Qa��5l����R����ʄ��b��Ӄ@��R� �V�n)$�P�|�~ �}I�n�g�34�lG���!�(n`�P�d��01b�c��Nu)I�q�?y(3?3%�� Yޤ$��L�xLOK.�:%Œ�މ�ק̤�C�Gf��������co�Ї�_�M��4�vM�K>6��bR qyEQZ��:L{O�abj�8��Z�9pӖ���?�~���5A�j�lwb̓��z�B�2n�v�g�V�
PѰ�Z������y\g�r0� ��Qi�%��ux/��4U�G��_c�?L_\�{��b�)�L]i/V7݂p�_Sn��AM���?#� y���P?v@፱�3B�*���Lq�h� �x�����ߢH_a�7���s1Ff����-0���5��x	�*�	�.�Kb��?��hl8��+<�$E�F�l�ٴ��3����g�$�{S�����u"����;MCe|��;�a(�[J����hf(����;"��, �����L�bZ)5@�洔�C[���tԝ����e0���Q�����}t~�zw�Z��r�M�U���Ir�߼Eb������j`���C�Q"�ܙ6A� ��Շ����ϝڐ��HH�����T���H��l��|�]���uĀib�~��@�~�136��P?�l�]ߏ(��s? �b�nF���ݒ�I��T��r_x[����z��������Vi��wD�u#|�2��>@0�ӹ�/j������B�d��֧��-���ւ#�w�ձ��z�� *d^�N����&�h�����ɽ;���R���&h)v�Y�>Ŷ�������:�ALVg��0�re���./�e��=�H�x!l�Ƹ��,�-�fh�,�<fй@�bR���������Nr����f7��:�Ҝb�M�����h���,�6w�#�����fG����	v7T�>u/]�m����sI��@�^�&��i���i�J�D�W���4�]������3p�I�=fo3�P�Z���7�Ҹ�T�F<��k�� �B�$�GӚ@ U7s�%{��X���bF���K�N��[��5����rc�S�Q*u��1�}�d5n�r�M�R[���I�u.�b/{�`Axw�D!L|�@�Γ�An�]=1�v������S�t+�N�ب��%�Tq{k7!8SW��><o�ӣJ��h��<��96�MF�p/�av�C�is��)YC�����
Jo �\�d0�� �V1)�u�f&� �D�Ks^&���5������r��is�.��8!�|)��f`h���Z�\4iS����H��rz4�QHdf�5��q�[�����a� �kl@�#���Yfܬ�����$zSƲrN�a	O'1�w���������U:���@�*����v�e�/��)ZB�m�	k��r���W�H���;������/�m(O��1�uy������.+و��1$�k�*#]y�抻$�������s~�0����R�=��r
c��u����/�0�.�y�ʗ��B�̶�m&23������?	��Y��gQo�B�;��F�J�im��������/�g��[ f	3����
(��)`�0R�Th.���5�Ձ�j5��+98�j�0��z��D�w�`����o܇D���AÒv���϶I�t��	�ъ����YlY��"\�6�wZM��zF�����������\�x�:��i�z���a���a|�͓/��.��`AoM�Sz>7��ޒ��EL^@g: Փwv$�3�1�L�+3I�[
{/�}H�=/�����5�0I6�u���\9�荵�})vF=HgH�kN19{�P�������y dz0��ǡ'B�w �B���������慯�/mZ}��a�6�B�8eOԁ��#xU㑎�qng��Q�'M��Gv���f�O�W��#&{�S��&5�_{���Iࣜ���7G]j��M��ozs�N�%a��)dgTr~R(B]]��J�R��|H��&��\�ќ�Q�4��B���d��M����c�e~��A]C�G����a�^��p��l�8cM7�Cvzh�+U��]r��c��D^�bL)K-��E(.ϰA��"��2Q��!iI������2��,���(E�*��vH	��@]\M2N��霻�r���<y�g6D�3��I��%���41�T����ej�����?bV͕�^���1ǔܪ��:���r}�*�rX�i]�Е�o@X>H�z��f����1H��3�4�j?� ?��>�� �s�
<2�`�y6;��f}��Ej�h_LmBL4�MC��;�,v���yK��;�+�R���Al�����1?���^��MVnCm4�`Ј�G��Q�&/�����W���]iM�A~�f�y	]�p)���!�}� �oCCg[��o�S{�h�j���b¢����l��KY��kt�"����/4�|Y>�>n5���O\Z��ԲAR8��C����;�_4�9����Ud���*�p_[dp�r$ExԵ
>�*�L&�	��� ��;�D��wp�8S�6��6�EfM�{yP�)J�zB6>i�s��W����ۛ���xi`}�4��Z�����n�޵�:PC����ƺ��PF�����{��&��.������@\�_=$�Mǭ���`?��
��3}!�8�2��3�e��R����e����a�)(��������z�aoZYq�2��;���N�$��<�.nTbCE��_ �@�| �h���h)��R �	�9	�5��G����⬢���D~*�`��[�Y�K�=�b8 ����\%���#s:F5,oeH�Bi+r|Sb}�Q���=�+$��u̅�v�n�B��ؽ,�ś`��Z�9����uX���>�{p��I5�.ey�9s�Q��ߋQӄ�jG4��|b�������۱�����#����1|���:h���K�T�;�M$��3iw�i����t��1[W3��w\ �Y�c�GE�V�����?^Y�W]339�	%|xl8��� �->One�%��fJ���Ϧ
O��فsZ�%"D��z&[����N>����"�<�kF��G�MP01A	ع@@��y'�;��r�X��I
.u�G^��ɦ1�^��n�2���.+aLyo܁�Oh�o�a`ş���q��4�y�?R���S����B`��@�϶8���n����ǅ���%T�s��/0�F���������H0���)�_��h}�]�9�������"�N�"C-��l�^�/�NA%��(��C!��ϖB� �T/��xYӽt�l"uSk��R����@]��2���Q�c�7����u�cRw}`=�vl��z����2��N����HA�Y���7u�*q�]�����Z������H��z����mt�e�}5j5M���;`9ܭ�nx2��M��wc;��%)���Bf�Z���x�.ߺ��6̬[�;J.xS�����r�ߜ�����X'� A��B]h�hx� <��&���ǜx �:\uԚ�u��mm��@��^���2�r��[���3[0��c0��<�wcD��� hL��|�Ιp�j�{֓Iow;A�\�}?����y�_��hG�O��sT+�](�5XZ*f����b�~@��"<�)Y�|��%è���)Z�@�_*`l!}��@��G_m/G�\��G�ல-��n�A8��UJ2���7M����sL�LgS��u�����Ed�����8��.��Gz��~������lZT�ܶ�������O��#�#����r���5������gj�s��>�#���+�g@������s�u��p��������"��s�
Y�rq�p'Ҡ���+,[ЮQ�w뎨Kz�o)u9A�B����&-i�YR�ޣe�23%��>�a��!᩿U�Q��بx����o�����]~�[B�JzAV盨$��&���l
��2���>U�����B��M*�U>�)�B��S��o��W�S��Z�Zv��M'�\�+j�E�4�E��t�,5�p+_��-Ʋu�z���(����Q�Q(Pɲ�0�'���	�2��S����V�Hzf�{��ԾE�ԁ@��_��clm����A~c�_��b��һ��+��TS���:�'��x�dyQYM|��"U�����
M����"V��@��3�	c��0Cg�"�_�=Нe�]�Hz�ok�?�8�3P�D�o*�Ϟ<�wL��*MO�h3s����dY�$����5Q��w���A���17��#?�����i&����O��/nY��Z�� �f.c@\^:���1�Tu���ߟ����*�GTvf$P���эlqQKLk3�v!���n�=|�#���@�­&T� �?�=��((�rG7Ƴ�@q�X.Γ���2�w,��G>����Ǐ�%t�������'�:�|���,�{Z���Jů�d��Fߟ�o�),���7���f�8�$B��(�*��-�&$<c<������5+cFU�%U�1��9M~�x�漗��+]���%{i�?(1��r,uØ�-~�Қ̕�z�o?X�к����j��|pw{���2�P$��V',���~�fA^�'�Q�*����g�q����V���7e�#��|��@F��9��5�;g����٣��?��c��z^s#�#������h�r�#��hm����*��x��3�Q,���O�T��S�ȇ����<w��D<FWsU�'�>��oIq�ݧ%;�N�����'���*����1�[�#����?��|����;.v@��Z־Y��c�O���s�F�Q�
�[�Y�!'�;���b������i��<�go�#�����o�IrI�MT�O�`I���/,�k)��N ���nn�Xf4�V:��|z$�4)�'<;̀����݇%E$�rѶ�������)�A�"���&��O~������~�H㢐Zbjݞ���p��@����69e'�<�I12��M���`���4�l`�)��,'�����#oFg=�������kw��/�g�Ñ'g������iɵ�ZKna����13�+�����IK���SͶ�$��U�:���GV>J"��Wm\ui�ǁ��/��j�|�,���?�,�0���k�K�b���}\��`��yl�y����8��[��1�
�5MhE��O�6�O�k>o�����`����S.����M&mc�ٰ [����##���D����߾;=���]���)��TPkt��@����T�=��~!�;���faɁ���8�VSċ����,!��K�jX��b���2q�0��X��U�&̪�p��
���W���#�]�F��(�o�'u,���`�f|��� ���*���,*E����}��A�➖6j�[z÷�ԧ
w��ޢ���#��i����v`�ۘ�[ʪ�Y�����
�hs�����]K_���޶�~��Zf�m�kt�����f� w������$�e���T�&�W:_��)�@���-K�(E��[�7�D�)�ּw�`�E�e=g�Q
LV{�'��D�R��*�C�sy���1�]o8�Y��XvdM�|��}�y��(uz�������,�����<����&�����e	�w ��7��O�+[Ѷ�YF��N8�t�m��8L��z`� �0��͉��`J��^+[}_2W4�N[���,t5x���=M��ah�`�Ǿ��˪�x�J	�6_�Ra�U�B%iz��~7?�n�c�^2��S5�����c�W��|u�K��\�珚s�6[k�ds����.�0����p�+i���*8��qۅ���U��k�2�),�@�!�ox?+�aE?z1��8��������k���d��C/k�p9�P��CeuU�5G߫>ׯ��s�"�}w���daȘ����tT���������j��nʌuδ}F�h;m�o\_�l���lU��C*�h$�%��f�U�8(��U@f'J;bbtB�����&�i[�/8\���Wj��&����Q-��_C.9OwM]G]����3W}�-�\��tȈ:�js\E�ؔ�ڀ�������7�ĉ��ڈtmv|���<|�X��5ٍ{;C����zE xfw��p��!��W�{�Ն�$����^E�7���i��u�7e=F�v��>y��&tϚ��j�<�WZ�۲�|��r�2]��x�}��D�k��(��;���2��0Ҍ�W����A\�_u���!���K����#Y���4������;9���er̶��@��D���Bk9jI>5&jX�:�ܑz����y{����jY",��V������c=��խ��ؗ����lK��?z`���J����NU�� �;�>O?V�f��I�S�=�b@c��9ywU��x������V�v�m;A{�e���8G0�M��I�'�:��_�φ��p_��V�e~G���u�r,a�q�z\��|�;l��L�U��n*+��z������DG�����Z��� �ϚJ���&m�����d&g��$����K4����^��|�>���2�͹��|��-uƶW]jy'��ၺ��g��f�Z:y��s��5[������ɻL�@Q[�~ml *Ұ��c̱]��ǎ�\����;������z���s��L�����z[]��N��A�:!����Sb��H�k(�������bT��&w�hSTl�?�;�%�42���7�/����~��zM�%��_ü���i���~�£U�8�J���B.B w]fD��ӸwظX�����x�3Ά��v�c
f_n�K{�W����t�[^Ɡ�� Z�E��C�bi0M��TP}���ڈ�兎N-0������=�-����8��a@#��B�#fFcD�r�|a��RXt`6��3��B��fϞ�f��^�F�� �D��Uk���`�t�!"FbD9f� ��
�M�����-mjeۯW������3^�O�r���,�K�4�Z�Ѧ6ʈ�q���0������)&JG�s	E&m���y�k��\��L)���f��3�����'˱��=�s�S�`P1� b�e�i���*b*F;��Xo>eTN��7��;���q�.<���{�<Lty��d��[���:4f�:U��f[U���XsE0e�hq}�g�}k���yu�z��#�U��u6�xB�J��W\T�8֊���74.��~ե��|���Dl�K�ų'-t�G��}zO����4���wߋHFf���[ZQ��4v�@ ZC�T\�,��7UJ�G>�-�7��̜�6g�L��ģa��J6���I5����Ͽ�P�,=�4q�Q���"�H��x��f���;�D�E-�Ί�%��J�z��ʅw` �!D׺�����=��y����B��'�D��i8d�����o�ͷ�#Y��U�W�z��������\��gxŔ��>�n����L~S��Y����x�QG��)n��5b�q�o�:c`�v��^	m,�l��'�[�hq���Y�������`q�Vi̅5�f8�������cy��3��J��m��l��jy�_�y��8��>")],cp���)�w�g��k�t������$,,-U�K2�F��o�j��Dߊ�����w������_����rR���p�~����b�p�)k`/������u���v<OV��3S���h�T�U��j�H0j%D�U������cX+�w�s*}a�z����ס`Ev;rIK6H������ml�Ζ�gA��^T�G���8vl�-^e�A"�޿��'|]�R�.*�K�t��RS�5��/i}������'����������F��8� /-�<?4V%���k{�P���>���W��H�X<���D)���X��IQ^��U{h���R�j�t(-~�z��eiit���ARm���v�c��F��=�>N�����(f�H�+��iN�5��#uK�)Y�Ӭ�7��mB�)!�}S%��
�O�`t��-��h�4{��z�l�{���x��;��mܳ3d��E7Rt �:��;��ߣ ����w���8xV���2΁J�:� ���v�a���"**v���^���N'Ŭ$'�`N�V�E^���Ϳ0R�Dz0,�p>�2��
Fm(�
�&)&��̱^�� ������s���g���F}&��y�Q����H���eA
�K%4�;��r�dm��gA�/�)�_�Gl<�<��n��2���~��.�/�%=�laED�+&-�P��K߹d�k쨈�ӮW#��_]����#��.ϱ]7�3�f#�$IN8��Q0�$�������Gf����e~�U ᆵc	�"�5FLѳ�c]���"^����ݶ�Oxb�[8:�ʿNVO�׮�(\�2�&o7��0U��<���b��&��n)�:�-�b��3y���gdjim��X�Ex�-�_g��\f�w3�����,b�V��
[�����/e������4�(J��n)7ި�b窊_�|U<a}1��07m�v,�};>�7R�-�ذ����^�\b{P.��Fv����O$JU�M� ����Y�[��>A]�XqGi}��Z��|7�f|�[(%�R#,�;<0+�U���K���@h�m����mN9[����<�����2q�w����_��jIXq��5�w�>�@��E��>��"�"��� �Oa���ʴ�x�A���q� ����~c��hj��5�U^�"��n�� ��Bft�m�M�ծc�AX(�����j�'���p����)믓o���k:��|R�p?.��W( Mc����Ta�ড��j�����<�3�w� e�v'���N��ѣ\�(	4y����T^�hwG(j�|A�!���vw#5�f�@��3�]�U�-�~�������/ژ'��t�?g4Ś�����p���D'�ᖱ ��8f�Q�#=�Vm��C�W��|�%�F���3�x��f��ZL�\�S{�N�%��[ק�D��C�c�⑗��]�k��&���6�e��Q��7FAԗ3Si���N%+3�z9><$kv��Ƒ�ZTy.kZ;�#/YH����'3j����j8�;-��F��FJe���ߋ��LeHf��6��՚�z3?b��:.8yֻ2�n��~4m����HSkd��7l&67��9���o�ғ��d����"$ oy*=���ߵ�.f�%R��./����靮��m��L�\|���~��#3�·��;�a�f��\��7A�y���^i�̽�)�n�0c���0Â�Q�'�rY<ށ��n��Ԧ�=��h��I��^�-$<
O��簥V�7p�V`����1u���-��FnO���q�����7A���w��}��5������L��N�|=��F��#}��WYo�����H�jl�7�p����C��jA��N����Q��O�1OR�����3�cɼb+װ�S�+cY>3�j|�^0�:w����󾋛��NL�)R����q���lR�$H�\�P��tp=�g,<��H����;k���<P�9�A
Ў�g�[����d�j�e���d���'���������ki�ߝ��>�����<�&�����-S���L��_q��&�S����,�L6�0��?�^k��d����H\�n�c����Mg�-½��������r�V�ŷ��0��j���-��ۿx~_ŗ��z�# ���bnۍ�@�\[��{�_�|M��m,���P�4��������oM�|��*��������gg�U�� ^B�����tDi��QO?g�օȧ�	Q��3
M���5���=o>*��A���4[��d,G|7�Rz��D!��b�Z��V��Cc/���Ο�8B�=dyi�W���_��^Wb�͗7�fú �[#��9�"�2����ن�Y��hW�����e����[��?�C�1ש�oq�u�y�KH�u�CN�ע?��-�]�*�|{������&���e7�5;V��RC���?��l�q�����ұ������121��/!��-X��5�n�*.$�G���$A�A��$3C��ɟk7��;v[v��7�B�O�����7�i-][�Hg'�u���9���:��p�мŃ	�ߙ��v��1���<�ٚ�j|��<����P���߉�I�	:8�x��:ٱ������^k�k�O��������J�Z�����v5)����D����.�|�L��r������M��e5g�a�0��%WM��<&�� ���F�����62�t���WM��/������i���e�V�������b�.�q>Y�����h��][�5�K�A�E�IwVp�~�V~�_9<�p���7Q�Nڃ�c���?_h,n�Ʌ��OQ����Io,�i�H�~|2�W$_(�U���2��&fL �@�CK�p"� �T�ËJ棟5K+�u[H�)ۏl��q��ے��
Ul�?��)Q1i&Wh�@�`�g�P%���Z+_]�o�P��LŊ�U���fw<h��!�S�Jbf��`��������4(��d��hS���n|g>��

�d����)�Ι�6(.�F��n�R�R��2��=:8"CXky�Ch��Eq�;�kh�����拃�diui�����}��k�$����z���"t����@�d�U��C\fa��TLfC����ܫ�srL�	f�|
;�qcb��f��T����`H%B_C#��\��g$Sl@S�z�)�POt$Q(�[9H"�_nԎe�a�"&��^ �RZ*�nF�2�k�4iy��@� ?:l�/ �瑠$��وq��N�R�;�Y8�x��6Ȓ�셵�������p���0ig��X`e��Eq�j�|y��5�Y��#����c�p�j(���J��AlN)e���#/���2M�?�����Q��e������0f�$�ȕ���!��E��Qp��2,��C��.�B��v>�s3Y��l�.E��J���Ĭ��#Ƹ�v1��l�y��� ���I�?������ډ��k_�i�L�%!d���h��a����<,�PU��K�lȦ� ��WR�D�Uߟ�҉�ϏuʓG�D������uB"g��{�s�n�e�`���(�V`r��%��r;^�9(D�?�4��4)�_�p�?��L�������79lΉ�.��p��2�����}�����wK��a�G�z�(3��lYSaP��X0ydP"wR�n�iE�وo�%�-$	~�s�Y!%/?����P�iy�~!�1N;�y��E߸(2�H��F�?�
�h�8D�r�<W��!���|JrU4�A#�CM=ViN+�Ɯ{�̳̀QI��[N�n1�tN��⟒1�F�VcC8�?io}@�%g�l�)����c��9�K�i�������+,4���~�w�	�3_�.�9�=ç��V��֐��hƥ��k��wTJN�bb��څ�~��5�ϧ��i�TK�}�b��US-?���	�5S��&�7���l��z�:�c�hzۅY�4����sD�L<4_�)�AԊ"�aQ�G��������3Z���_���/K), �,��~��z�s�8�J�F�qd�Xk�e�*�3�����ن��S{L�;���%Ou
����q��iD.k��	����î����[��f����G�����a�Gf�W9�p�h�����/Z�ї��_�8�=T�� �y����Q�X�\��X�l�ɟn�~}i�W����L r�U�`հ?�t��i ���4Q}�>��1��!$��ᇚ>R�!�͞�ɬk�����[ؚ�Mwi$��]�|�(ac� ��#;�z;�¦���S���܋�}��4 qJ�����W YmY(k_��ޯ(r���v�9�8�G�M�KJn���k�|���8k��:�&
��-��|�K���8��9x��]�C��U������t�O?�S��䗤�;)>ИR��f�>e�00���V��,��0|F�m�$�^�Ȁt��3����̕�mߣAf/��_���EQ�P~w?+Hcy��T�<���b��Y��)��E�a�6B��I��Z�;w��췘�ޟ��+��^���ӡ�~E@�h	Z�%=�VX$�֪a}���ٰ�\\�Vio&�SJv	����RHA��qO�{�jL�  B����OlZ����.f�������KX��q����c��w{�6W)0oKغ�ڿ���3L�Ns���G	A>�T$��%���-8������X�� ��.Mlr���|���u�6=�j���;7����ײ�1uq@Mq����6�9!r���<�u��y�}S��,�[Y��^4�H���h�́j���kEǤO�:�M�,��h�ۗ�u��(��l��쵡�Ӌ�=����\h`r�^��i�]~1=tn���^W\�>���%��i�V@�B��ܽ 8�a@�s�7���g��Z�%�b�?F���e��}��鄳�C���J���z
�[�Q�胴��"GN�;]}(�gO1��I�\%B�9'�1��l[�b�w-��6(@v(��_]�Ɯ7�e2�u.�߉���(��|F��ǵpA.��e�H*�GG̝"ZC�kq�	8������)8���d^*A���C3{�a"��/�b�/�2�{IB��
Y���*s���=���� O p%,�P�{�OS,�m�1zY���=���A��ר�C)���IL��[�:L�E���=%�6f!�b<9�$RU�\Q��]���r'K��.�ć3Jw� �%�L��fg�IXC�(��p���߀����o����! �	����{ŀ&��N�ۦDLc�7f���g�/��K����j����N�99�Z�b`��&$���7P'�k�5:ݟ{=�0����ӕAa�tV���|��'6R��]$�r"�z�+���6%�A&$�c^��X����ƥ6DDQ�� c������?�/�qk�������<f�Y��y��_����{�gd�Uv(��6�lh����F��`���@s:�l_��7&V1�͑��=�D���աM��i\#�Ifj�y�04��E]:�Qm��F3Zm�����2>5�aQB�}"3�&�68�Ƿ�٦ڕ e����f����)/?F2��1k��y���&��H�?��TU����^�7���-@��4{+���՜ᴶ�:��[+u �z�6�g��*+�e��m���OW��9���5QX��8��P#�t.\E��ws	���
�!�8�������f�i�d�����m��'^cG�R�v�)l�ȅ�$\NT���+����,L;X)�k�hs�ث��iQ!sS(.�(CITٗ�x��,�mw��C4oP�~���z��߀�t��m��[ۺ�E���ߍ�N�r�����1P/�R��S���)��
�>�R�&�����sF5ޒJ���DMʅ ��d��&�����3��a�$�]x@���1�9�) ���8�:��ݥT�I�>�r�0+��� �[f�9����pR,�W�>D�~`
=�D�^͎	�Ẕ�ڼ=����Q�����}�zDEɠ�/�V]
ܾ�������������o+��`~�n�+����+��?���g�u(�ؒ��|��|_͘Rx�0��/4���j��w�Ez���?���oZ�G+?*�d�E3��x� ����:}���l�%>�kS!.�	��w`�^�� <(�g@��c�� ��éO3�=*��}]��h�,�R_D���"�B���v �y���<΍�;X�Կ�uX#س�SclI
Vp�m����S�r`�Q� ?6#:�2�?N���c�Q*�Ԁ�h�>2�2���/��X?���!�'���oe�YX%K:��֪Q0�Q�;�kف~�j�Dj�=�px�� f&����`n��3�r���~q!���G�����
R��ΑB5�}�[u���5L*R~X��E�$���'�]����8%�5�0�ed&΂�	���Wm�R���d��@I�܄?�ݼ�l7��C��ZN��-PV'��t��<p-ΰ.�r��T�[���>��P�~��Ĩ��A <A/BV��:��2c��c�ڢ�&��w�Kz&�z$	��xBP/�n���	vs۶��K/�ƙ[\T�c�#��'̃Ho��z{��f:����/ɔa@CQ3�4�k�#��3uS�3������J���0
[��~��~M���14�^�:�Z��@D��,�V���>eÚq�Uz�z��%�;�CA�[��^�?�����<�,"=@����c��3�_`)�y/�E�;��D˚f^LnX����]qC!�tK)��T����I������!P�^da#_nX�d��������q�uɕ +_�|6k:bI;���2C��]�my���&�,Tĩp��C�,c�O����c �.������s`�:�� a���\�U�Ę�
�aj���s��:�3q��:'�0����*���S�+??z�(A8Q��_
�8��1�Hʆe��ʙMx�X�1�����H�xZs��)_W�4�t�QPpn��P/f����ɠ,�f�ǉ9ٮ�[9E��,��@~���SK�������=?I�᾵���Q�����t�:��{��vc۶;il�I�jl�hc6��ضm5I�w�}����䮕̃�������<��M���! 
ܾ�d�8�|h����T5�����*M*W>k 9%BR^()"���=��[?������}��?����o�E�ry�}�}�^�a��g .��{A;h.KYX0�A�g��nJjkHX`���-G�������6��)��p������M�AH�%#����=$�n�F�!W~�(�x႞��9453۟�R��6~H�����(փ�0s垹�5���D���T����Y�	��9j׎�Z��
]��dg�=�帶��+������<��@d���HK�#� �-+���i�/���"\W����p%��=o�5|-Zfq��Bi�WS�����3���X�<2Б���� ��ĭ�֢b4�1�f�����P�m��>}Mi��W����p���S�rE;h�U6�դ�r���� N+ŕy�怗N�^�q�Y0y��l��|6�"EBA7�1i�bu�R���� ����r��q�x�~��-����_�O�B�� h4nꋸ^ Jk>6�%��o�Olᵄw��z�(��4c�QГ m��('�poV�CkS"s���)��pF�+m�x��IR������\�Ӏ��IW�~j�eS��_��Ѐ�q	�S�z(`� �P^�O9���/�D�rR�^׹anWz0���,e���kT�'AZ7:�G!"��9�����^��DZ�O���-�ܣ��9�	^MU!��$qDK�1�8r�X�������%�^��Z�$hB��r�9�zJ$/x>��CR�ǐ�J�+�.!h�l�of�}z��ц���=�w��{4���|��IUa�:Cٕ�:Cy��k=�̇��7�Lh���Z�����=	�!؋1��Y ���Q�������$�d����݌�m	���r07���y�rXD�>����W=��3��r��`wC$=!E��e�f�5�$-G)������$�yn��^�q�_�HӞhM���u�ӫ�^����`�$ۯ#�Y���H��I�_i~>��l�ʎp2V�kF�F�	ME�w��NB:�m+��a��D.k3�Ν*�L� �DaּIO8�n�u%BM◕� [׉�>"F)�W5s�]�v)9I�Y��s1m������wP�`��N��s��y��㰴_(vtyJi��
()��m�J-x�y��Rp;�� ��zv�&�ŨU@&TMEPʠ_i���sC_�>��p9P�׆�xK ��W�	��$���b5����f��;���b ��d��!��y�7Ƀ�ԅ�����j ���G&�s*������1���?�W{�9�JG�!�9	,���������S���7ˊ]�z���ކ�S�:��l,u��-��y�p�C���Ԙ���s�D�wud��s�̟�(�X�`/�K}Q�� -=��E��{ݝ�ΡA�5p���C�H��-�<���9R���R�n�3\Ҍ\F%�)@�M);���[(�4"p;�Z-��F���/Pv'P
��*�9�-��s��8i��"$c����ɜ�Fy���Mq3g#���ݚ�h��'��tD�SVM�Zw�R�pBn|��eT�X�Pu��r�Ϛ,��(�FQ���QC"�#�Q`yrl�r����8�=���=?�)��Oi���l�a&���E�.x"���+��aU��$AG��Ƶ�糃�<�|�ܞQX��$?µ�)fk;-�i��.q����4�5d�6���~\D%�L0��1fKĳ���9�u'/zz����U)�,i��p��~q�0����0TM�E�k��R˧&�+r���"~��}���Ay��;�D�(��	5*>%�A�D�rT'so�ݘ�-�q� 2�¶��0�v՟�d�j�YC�V�wL�7>(4���������Ꭹc�3 w"P2�L�K�v�2X�k���P1���ԛ��P?���L�e��4�a�7X6���݄��a��4Wcj�
>o.c�Dv��̧�JH�������d�4�:@m�BZzT�Z�G�9[7�y��̌�4
%G)ǣӶ(�-/L3�	���$��dm�9��]/R~��c��4�����E޷
y#l������!y_�[)���J�~65��o�Šd���c"�:���s�^�J���x�j����qR������|��B6ʛ�,0�8�tp���<U��cy��6�!��ؘ���R����{K�Ϻ|��m%I��Z�B�BmzSOK�S��Vn%�t��\Jk��R�n��W5�̦��N'i��6���S��J�
u��o�!G�e��RpM��Vɖ��9���n��ϒX����8�����v4�H�.D9T'�?띨_�4����ۈ޾��}��Á���1;��B�
��� �͚$.x�Ȑ�7�4���Yߟ{u���<9�Oc6��`v %-fj�6�9��RT*�2I��� O&����}Mp�l��8$��I-z����Gv�g�:��4�j��Oi!
8������Z�Zsꏺ� ׂ�#}�����{"(.�����:�ih&��մ�CGVV3��*����ȤT%��F��:�x�MQN�߶����=�qO(�G+�@��^�T��c-.���W2ν]#
�JDɟ^����=M})�E"{���P�H��O����-���ٿ�� �`�+�ѶA	r���^ӈ�|���0U�.��3u�bm*�`G��W�F��o�xJP���6��wi+x��%td�Z爸g�ǻ��` �&�8�!���;����3�Cq���O%�1����y��SWc͑׸��Y�0t\�O��.���*S`������e�}uʬ-mC�烟��!V� ���8����b��K� ?��{�]�O��}��UE�@�����÷4�ԌC�C����,'Ŵ�~�����
�8Oӝ�+�f��晽���~�xoDR�������C]��q(7t3,:;�]�aUY���_�z�J���o05��CA'���MB��N�Q¶��ե<6��"%��S�0J�����>��؊xߚCp�g�)$`l Rq�ijf)�A��QL�Hn(O�$p�bR�� *_Z���^E�����g˛)_�}1\y+�V�c}:x�HdD�cLtrUo�XIK�}>�#���,�N��zI�~RA"���h��~�{Ŏ��Z>����uB/�������������<V�u�3祚���Aߪ΂=����<��d�6Ƿ���[a������*��e<_���{e���}���v�̘�
. H��Rqn���ٕ1c��8"<c-�]0I1��8�?�S�X������E\U&�.�ҧ�2��b;s�iI�O�1 xң��b�*F�4s��p
u��d6;v�Fj��bt
5����,��gJ�!U�2�Bz@�Ԍ�hb�U��gz�!�L�ȵbP䭛�uZ�9� �IBl��0:�:}��S�1��C3,ݩ�U���g�bzd�"���3r��8I��6lkE5����� �d=��Wc$���.f|~B�z���Zg��/Kλ5\}8�� 
K�wr'�~���}r&�d֪l���t&�4ˤ�>u<�1���JP��F~X�0�;�'%�bE?̸e�>S]�S}�\��ƍ�������Ћۀ5q�WR����SƱH�tjY;s�D�P�F,����-��ԡ���U��eקa�R���F%R�L^ np�ݐ��i����˝�zj����K�'����o�"�Ⲡ3_}�z��IQ1?,p�!x��` yP��!(�P�­���-�2�Oj�~qNQ,�}�NR �X���+�NW=�l������>��+�f���{�3;r�g�����L�daK\��IE�ء���z,�-��,oHu�EC���8J������ܷ��7aͻaC'a��V��EsePΨ9���1f<Q��I�h?�Dsf"=%x9qS�)Ȃ"���ª�k��3!��!�\�čb��-��c�,c+��Wy�����t��H���<�y ��Og/�#8��0�$��{/�y�(�=��>8�+�c+߬z�{d��յ�`4?!�w��q筦~��_?M�r��3'��{�$��ٸo	����U}�x�?���|�}�!/�}�|�0�b��ޟ�y���.�S�@K�H��>>w1���.T�:�ڷj�[�X�\���ˈ�ɘIF'�W��(0O��H�̽v��B^7���ټ8?%`)��P@�?�^�5�ޱ��h=ڊ��$8d�8%XEM`��Z����T^�h%:�<,���6����8��$�S%�G��a�[�w��OW����o��`�2�S-���ފ���}y��Ql�d�DD?��D-%Ar��"���-��)E�#���PQa���ѐ��БE0����aQ�̡I?M���E<��i9�'�����H�K"�ch�R����e�(HC�܎̥&~r��@��	u���s��V�Z\|�E�(���b+̋�,"��f}>N<�D�k�4�U9�D %Ϯ������������3}Q�[���ߩ��	�@�+Mw�P�{�q�DF��+.�N�k�!�$ܯ�];kӫ����H���"�����bv�y�"�7[]�(���~!�o���R?������u�K��n����/�A�hQ�&��6Ѵ�!�;	5��w�;�z/y�@�h �?�AE����]��":-�(8��n�8���p��]�2��������wd�iĩ����h<߻h�3���f��F!�0+��� �ʠ i��}zA|���S8���m���Q��-�L��R�ߗ@���4D��	�dP-w�ב�˷�A!�젇�� VE���س�i�?BӶ�����薻����M�����:���|-�Z�J��/����a]a����0LQ4@�d���p�	���x���W�+���6���z:5��Z�/�I$>h�~��[te{L��XtG�B��ӎIVڇ��"�_�G��?:� ����{�/�:-"A�5��DH��Ʊ�M<��X����Hi��/0.|�Z0E�p�3c+�k���O���3o���#m�36C��>��5\�&�V�����j�O�~
�q���'�_E�ukƤ&�)����v�\B��U�����c��s>��w�i�:8ɶ�?������D=��ʭn�eR�ٹ�P�����?@r�6��)�x�~��ϛH�`���R�*��*��Ža�)���)*6�5n��hc^�a] (�B(�/��I�/�$ߒ~e�����~L]�'3��!�þuw8��o�4U�œ������%���6��4F�!@�-2����5�������cJ�0�5��F!��M������>	����R�e��t`n�������I�	��s�C��$\�������2U����?9���-��R3��1�{��_��$~���2[CYe��-�T�7��{�R�
$sA��I�2���:axS��!���6� ��ZL�����M��H�ŉ@�k,m=�8���ퟛ$8�.����)��J��k�Hd�A8�D�o����0v?�.H��/@@!��$�Ǯ������׏p��*�A'^��#5i�����H��|�H�w�t��ir~��
DƟlSe09p�b�w}n�S'�FJu��(�5�~Ğk��? 6]01i��eg�����e��c��fCj/.�6:a���J4�D���9=�=P��;��J*���0�B���%_Vc�5��������L�#�W"	p5��z�,lp1/��wo�"�)#2�j0�C�&�ň�U����I4*��M�����,�焯!dM��h({Uʸ�p#w�||�O��^mU-oK4�}����jY�F�����u��B�3k�!�㭣���Ǥ�΋mn����H��J�NN���OJ��[��g
�
0��u�.Z+<�o��*��r�;�/�,C�X�!f[H�2r%�%�B]�8���l�>)&<�@�kv,��a�F�h�)�\ؾ��pP�pnb&��5�˽�|Y�x�!�j��r�b�j�w!c�vj�j��d"��t@�Փ�jM��R635���g&4���˹̂�A.TD�Ri���ft�mg��5��qyR�K �,Q- ����A��@ �ۗ���9����-��6$�啠�y]�Jː_�#����".#��FS��Vd+�C�sA#!T�2�ߎ�"��(�u�\٠k��Qϵ�dG�>�@;D$کh��.�ת���bdr���� ��/�m'��ўG���:�����e� ����4���m?�u��vk��\�H��������?)����EM/�x��#�0R�|U<����P��r����}����"�d6���C�r�b���>?��k���\%�2�@��`�����]Fѹ���	O��o�n�Z���y����iO�i�{�K�X��Q5�7�xr�[d��ML=�	�O������x���v��1�]:'QiĆ���_ o6y���`�}V�Qk��@�a���%8�U2y�cc����
I���N����W��m�s�d���	M~g_d��'����mBg�p���qj�*�@�� ���"��ot!E<U �
�h쏪�4��s�}n7\�O��@���(��$�Ȍ�mc&����p�8V�v?X8~���6�2��Qt�: �᫇�i���p>J��x)��\�*V��D��^W%�B,��(�,nr⮷�kwk��W�v�/.���`���S�]&���^��C(Y���ͧ?-_��8J��gpaw� 2e%�X���qn�~�_����X��4(j�=���k���ƒAw��8R��G�9��H��	Z)
:��"����@w����$.
�'��52��|�7��F��\(X�_���L˸:ޏ�%^7��p�����75�ӳ�f�kA���jf�;�Ŧ�	��>��<��uѱN�ؒ���1�&`�����j��~���O��=�뫿����_n#>���+4�u~��^�RzX�M�qy=;�M�S��wU�/;��9JDY�����K��@�l�fG�w�EN;U�UJۥ�8D0F�t��׹2��  ���vO)�$���-yA �c�M���7�?��!IB" �������<v��N9��޻�S�]OT+�'��)�r�.=7���L���n��.�i����#n��r�����穳�3�)5 ~���x�MK3�0Jh�)df�w	Ȋ������~/�s�hӿґ�|w?[{�9g�z�� ���|��}��S$J��W%wC�9)@l�_��~������3�{��欦��}u�-�IMJ
��IL�ʋ:i�1�F��+��'��'�#� |���'*I	*I�㯱�G���+�1�ıl�/~�����c��ckm���6��Y3�֛)mQe,�!��,�\����md���h��Q�D4V����2n��GF���㵎�<g6�䱯����)Ư���>R;#��vD�Z��V~M��e�K:��6��mU��b*�7εW�o�����Xk��J-�7!�$���E�­�1;/C~��?�ff��ZFEב!�U�2����z�����a�6p��*��ς^���M�F�nܹ^l#��N"���  �?#�]����k+8��g�<F�5����K���*�kٲ"�����&�RtM�0���(�M�'}�=�`9;)�)8��L��9�x ��2}[%<T�%��5s�(�QT��K>�;	j�Ycw)a�?e���e�a+�I\�6lȮ�W���K*����:T49Cƴ��*�����H|�F���[�� �!����5��i��3�&G�T��`-�5�6<����9A'h��Fnn��4H�0���Eɶeh��8���6��V�����A�@���ri�㸸�O��ɨޛ����I&�H��ʪ(�ۅ�xja�P�*��M+�5���������?�sUc9G����p����l��-C��&,p�b����ݖh�6�,���V���R;�9*&[���n�&[VNdu�޹�w�����Ѹ�Bi��J�4��(l^��M��@,��!�� KЕل����K9L[&n��r::�gz�VQv��8���!���|E�!��H#�0�؍Kb)��V�{|�:M�'=�����-r�|�S�L1�m[jw>�c8f�fWD-�%ȷ��������{�����L��n�][$I��e�t���l�vJ�*���˳R��Ռ��*�=WH?��y��u������ۣX!�Y�cr����4�F
{�<����3���y�x4?�O_l|�}�Ql}<�s��-�� �g�:�yy���*�����L��g͟"��.��������wj\&\��J4��\u���:��Ua�H�K��y��MZ+ܝ"���_��6'�:9JB�E�hW�]|an
e茲��ncD� �";aIQ|�T0���d���?������_���gq#�۾���=�ͻ�R�3K��wWFZ��k<��Eɱ�+i�ЀXW�����i����s��Fx����0;n�9�&��Ґ�s+��4�߿q��K��bA�k�G��\����g��I�~?C�2���.��
W���eT��@�)䜢n�j�= ʙ���%܄��j��j%z\/��m4����2^\������b8�0D��fϧ͙'��m��9I%*3�\���'�𶸏#<��c"����Fz�@���9��6zo��VըE߇^�����v�m#?10aEm=ۦ��\���B9qy��ʍDК��#+F|7�Y}��k����G��}���J��m�=�O*nv]b����a��)3�K�8/����q��5�˚׀bk6�`i��;�&��KKлA���G��:{�{:�3�ۯ*X<woUi�g�ώ��*�.�&�x]��Y�3�!C6AHj���\|
j����b[o���O�yX�w�B�r4����>y�"�e9(��;��$��,��|.B���k^<LU3�)��Î����s�1���#b��8�#@�����,�s���Ŗ���˸B�Od�UT��y�������"��M)�o�/�덙	N]��ܾ�afvD��C�=�_���[j`퟿�J'N,KܒXI=�\u]��Oj��]�1�D���)�ucW�H����M.��9=H���yL0F�i��o��u��$���>�5��Z�9�e̹HMr'�!F�P��w/�ŏ�Κ�D�D��:�~Q�_8zu����q�O(��jb�k���'`_/�_�r �����fU���[������?F��1Ag���?u7ӾZ�Y�?%q��ⅱ����E�����7Q�}e�:]��'�zRf�o�wͻ��=��^z�F�؉��w���D�2I@�����gUO�A���M�l#1��_)����;^�8t:/c��O��5[a&�V�Rc^��0�6{�!,�Д����P6vYg�*�";.?<��W��� �+]��HNEcݭ��"�&������`޹�I�h��]s�r}���nں���k���_�0�n2]H��ve��𢟓&���uC��͒��d����� �w/:���1��"W���Z/�x��޾P\�Xͮ���`zL{,�4Ħ
���~GasR�[R����XX�����熛���UG��:x���7���j�/Ai]���S��(�:��(z��2>G���R} �
�9��e�*��l�oG���%�ܵ<�2-Fgۊ���.����?��N�_���,�kZ/SE`YـR��l<���Ӎ����>e�n!>Ó5p�����?�S�w���x𶑒-�]vl��x�ϒ0+;e~7�i�R��pr��&\�.F���U�Z0N�����(�Q�mmЫ�����GyN��q6z&�.�/��5<<�=�:���
mz�5�
�&o5���-�/��'z�Z����r�`�X��{Oðj!�oմ�_��؃��43�����]��k"�����=��Xو9�0P=�(�����/�gSD�c?�~M=�f�3"�o�'��FC��xv(]�r������lW��wu�ٟ����/ܡ[+G�y�ѡB1�U�4ۘ���[Q��?���@<K�!��H�����n�8̤L�h�p��EFq̪V�7:��z6��j^ 6���j�[�w`���f��nX ��q�����U�T����ܬ��ӓ��1d�(>xS�1���\/�]�|����q�L�5.r�%�s���"Id��_�5��qq��2�ǲq�� �9�~$��|\�
��&򂡫/��J��&.hdiK9M�xC��V9�>a��<�xZl�|٫y�������=8�M�A�h*��F�$�GX-�q_�������k�/�`�{��[�ji	E��DF�
Q'E�1\M*�
�����hy]-� 4��K�����O�y����^�!PZ!���,4v���m*5<�����ek��v��8�ņ�C���aк�Y�n�����m��|A��U�3�_���SA�Y����=�N��UOR��#��N��+C��]���'��E���-�w!s��*�[ি6�Cy6Ѱ��#��.H-��f �9{�Ez�@��fB	���qQ$�Cc�$!��	q�>���T��]������Q�-_�xVwZ��I���t5�pMn�5ntQ��*Yڟ�f�+�S˺�I�Vˠ�cy��W%y�Z^p����.�{�Q�+�8�0>4��]Ǥ�
Ɗ��'Wɷk�Sik��9"�����m�y���U����=��WD�I3#�!�y��?������~;���xG��[m�$!�v8/~�3?TT:��R�WN7*�1���<+�<��\�ݡ�f�����0a��p��^���Շ�٫��bcMo����O ������D;#�ɐ #S*q$���Wy��Q�1�|'ۀ�����(�Tw�%��A�[�E�z�{����ɚ�zs����8�00�,��;��`���c�:��r��8l�lR�K~=��g�gO��%�>XL�q�b��e{����ls��M�����1��a�Jc���ۂig��g;1v�ҥFW��#���e�Q��wN�U�h�.������{��]*�dH�n��*Q-mp�t��܆V����nDD�kqu�jZα/	���ض�GWۀx8��/��^cb���X���B,ֆ��AET[c�ۜ`� y�P�����y��M��K�\�$�eO6�S�k��q�e�82���f�k�ɕ���(��N6E�É�"���Y���ͨ��Ml���0��M�Aj?�]���nԪ4-Q���ԯֹbz(k?��o�/@5��jQ�A< ���}ʅ�+��R"��� 2Oޱ� oE��9��i��ǠX@5�s�L����c�^"n�$�t8{b�)����8�XJô�珙]��˚�2X�*+�#�F꙼i���Ӌᴋo�Nl�\����:�_ɍ��Vu�*QH���'�Q����n�aF����^�Uֆ�LNk���3����� ��O硰��3�e���hk�_Q�('u8h��'D?޻�},�^�Ŗ@P�!D���A�G{�����'���6�!X�ks_=������_�PuSMo*!-'�us��C�����65��ekaWJl�")��1����ok���7����*\�P����R�3Q�T9��ݞ�C����D޷��C[�-�d_���/yo�.�K/�mE�|�ڋ@ɱ�p�B5��1�9���W��=p�#T�^�`�X��NL��}��K�����]��Iә���1+�isG��"�b�=HZ���,livҙJCn��q��X�����g�4%{�[�܅�\`���s�^����o|�����0b�3#���r�b���	�"�S�h\��!��A�?�zr���I�QK�գ��D�+��2l�Y�bf�v#��A�k��=��zș|�#���vDgTx�	�y�z&1���}���(��$8�iWb����t�V(}����]�B�9�}˟w�H�����^��N���p�HS��*��d⍆v��B��}���t�[��W� m�h�p�Ħ��0��	iRi?�@�q%�M�)��7K-�����=pRh�-tUuq�G�u~9�(N�n�s���(�)�1�ƕY�
D��ݟ�B�ji��ݝ��Bj2h�2J� �77o*�1a1� 5eas@K��� kj��.9	a0{�  �Mr�k΁�Oeq`]�ǰ|�����qd>_�ZTK��*3AKE���B��xu�FA&Z������PyW� C�ë�{�["��C|��C}Z���Q�HY������ך��a{?��l�.���M��_?dG�W|��Έ��݉�dY�V�|�Y�rQ��*��m�~����;(!�,T���'��U%!��rs�*��0���?:ǋ֛T}��Ef���,y�(�|NV�I��Z~G9g��?�M[#/���?�e̝�4�1�ښ���<7��aR1n5�3�I,$5���V�ߵ9��c��v�%�skk�:ѢQ�'�[4�:�\W�Z��y�.���U���'�����eC�/���.,���/�<�W��C�Z��~�0���
ƛ���h��I?~�:vc(���[��z`��u�!Z���镝F3}b����XJ�@�r��l!�Sle^T��?�
0�����%����3���c=W�9[M�����]h������82�����9IW��ybZ�����:�u�=J�^	�p�>~w��|A���I<�z����3�r�$�$7��@"m� �U�Bv�G=�՟��)�k!:��F�f"�5�~�\��P�E���^̂]Z��9��uG���d���;=ޣ��b|@�>[�)/D�Qny�m8�k�_�3L=V���9�ZiY|��	�C_�<,��O���`��e�-��;;�Ug��oOg��2a���t��431�Ƙ���)�_[Ma�7��4�uC�ٓM���Sl����d�p�1��4�~Ȝ����x�n��"�ֹc�zоׅњ���FR���Ed��ꌏvRwHեN
?t"�^3�F��yn>:�����SY��An���.�)(bAl�w�-u���ݴi8��J��-��R?�SF�w}�->Tk�@ϳ$:9�}�W/�Q��W?B�A�p��
f�n~��r���U �qSGP����Ѕ�f�,D>�$əؙ�$ 8[�B|��i��CW�U�\�Q>�����,u�x=��&�8W��Y���R�<v�|�uS"���VJ�0еyA�.��[���B��"��<H�tq��h������y���L����F�-ajӸ���]ĞET�`�R�w�c�/BU.�� g����d."�M\j*��j�D�H!�_�HQS��o����=�O��H�P.�=���SI@��U@�F9��f5g��?FH,*�V<Z�⎢_�4�9g���8;ʽ3WD���!��Y*d�)e�'���l���M?s�
�>�T'EK_���:�x���A#����靷��Ἠ_����lR'�ZE"�=lT�S�I���"ܱ��I �'� ]Ĵ�/�B�RT"�E�,�����s�#�ky��V>�_��'c�N�Cjy|N�&�5���A�����އҚ\��sl�9�����Jq T��1�W��b�~�G$=�Zϱ���������?S�����^��8���-�����S���%HW���#��.��iI)�OYH�fݟ[FI�Λ�t���;�c.&d�Vh��:� =��g@����ϔ⎣�������.��V�n���|����=#F ��NJ ���,�\�d%���u���7�����h��'!�'��y��P�U ���w~�����xƁ�v6M�����n����7q����А�x�^�;���Q��R8O��S1չ=�<5H��fBA̹�O+ȵYXƹ^�3ll��FΧ�Ն�ǆr�:�J�'�quė;D::�ǡdj�KE�� R!e��pW��e��y��A8!���[��^�fx�w����b|N�]K����l�H�t1*�.�L�p�G���/����R��`}A���/�~\r�L.�>1�HomȺ�-��9"�9�2?�8�H=�!�w�3Ε$5[�%ML A't���B��\z�B���HI\;���	��Ԭ~�_���fC�؍ԃ��5�)!"�g7��!�?W��f���a�����= �@���h�R�OU3y��ϛ����
.1�j������l��	�����UvȈ"�,x�	�|R�8��4�F��\t:��k��#y�`����2� �Z7#��e��g�)�I��ә"N�c4� %��º2���0�{cґo������TV�C��qّ,��,��Ok�����_$��)�EFp���3�z����� 1d�$�t��m?����zD8S����)� ������q`!��K �ʃ�L�q�o%��oe�I+�]�>��N�Q5g49"�Un��ed��,��_�K�!�����E��oW��Ќ�Ր��N�.�N��G�҆%��oG�9���4�̳Kx�l*u�4�`�E��-pE�����`p%dZ�1R���>��MY��&�r�o�n+�m��Z����̍oa��q��ʠ�g�-���b�+F��<�sz�ȩo���%نm�0K�MB���xm	�.I�9�쾞u��ޘvalp��UY(�#�QmO=uH�*��"�!�\L�ӧU�g��!?.2�ݵ��oV�\��e[A�����1wY�=�s �����Y�-sk���4Q���T���<�%�19��$�4���q��|C�(�>@�^��%�^�AĨQ�CD[���u�Q`e��0��-��+P��I��ȣ�m�N"Hn>g8IC�6G�4u�$Q�m�Dʰ���(�Êo�Vd�+�*�����k��g}���zѤĹ���a�KHH��&B��  �{A��AZ�?��k;�l�-�W�m;'� p`_�Z��tϗ�;j�DV��:��n��u����)�pa~,l���1k�TK/�A��1�C5[xb2z�x�*h������oni>�ޮ��%�������:�sӃHX�ť�(E	Al��]��k�v��e���1X/���3E�R��'K��� �e����1��A�Rb������ !�^p��X��h&/*�Q��U$���'��8����c����- ��Rb>���-`]<���f7�X���ҽs�����������Nd���f��
Qy4����GN��B��u�zx"R��U��I6�U����fX���\��-Oc���ō�z���0�M�������b��7��������>�Ao��=���W�����2?T 1k�#��q���15t��>&K	��\���~eδ�grmx���`��5�@��]��Y�H[�l���]�j�}QY�Cǀ�Tud[h�l�F��+	fnRp��ުD@mF!�]%�1W����IG�;"_#��T�AdO��;�I�te�廒��S���e�1�xɇI����r�ͱ�����+4k��~XK�]�I�c�Syt��-�?�Y�L&	ϺH��E��`��j;Ĉ�`��V�yA[� f�a��EN8����I��J��<��\gj���{���I����ׇtg�m֩�����R���O�v���3ő���.K�Q�F�c����vC_��-q��;]O����s��aa(��q�	G0ͦdt���@q�U�K�A��݄s5Y�vy�?���!�n��^ @+>��#[��x���r��r�I\Ȏ�-V�=��4f��>�hs�d~�|������}�I�2w8�e}�j_+�z@��y9L�Ź����c�*���c��%���T���U�5���gS5�Yq��.����lN�]��o3���Gr��<n�`����uiK��	�M��Qs�@��W�#�
i�6P� ��.`.������)��^w�Hn�)�WN�a�}*{Uk�}먮��Tl5� 5fà��5���#��,�P�̄���T|�n����7��Ӝ"Y��.2��'y��]�'\�f�X�`�>w��Ҷ�����5`A�(�?E��6����ШM��K�b9�A,�M�L�!��U~v�
H����Wms��В�G9�V 7�isS{Gvx�_d0��Ω2{�ǧ�RV/��jW 37ސɁ�,�=n%�Df�'�R,�H<�-��7���� # ESd~,�<�P|���S̭V���8�pջxx登W�>݌b���ÿd��M�r)b����G�yy�ݯ�p�DF��ZP�{��f������	�AA�dT��$�(�|�i=��h��m��q_�B��u��7Z�vY
� �D|��O��mX�a�}\�)�ӯ)O�!`|�V'U5>I��!��)S�|�Zgj��*\j�!/+�1׀Di��O0۵9�|T�͈='�e3��ؖ�u�Dc��n���6�����8Ew;q��B�߻�2�q�?d��� �w:�(S9�;��6s��t�E[�"V8o��M�X��U�G)���:uiV�5W`�_������t['�#��`�pڌwǙ��@j��1���D@����zr�tu2�ɜ�\�")�+'���E"��[�����J������1�19�*�__U�~=��Cw*!=��H���"0  Hw(]R"�")-HݡCH�Щt7��<��z���|��3�����^k�n����R��,��ng-�$��{�K.�hA�~��3|]O�f<MS|(��'�+�Z�<y\b����-_&����V�tq1�Pb�!�=4��S�f��G�+�;�g�l�c�\���	+�ޠ�z�>8�ebu�'�ym�؜�âd��Gϴ���JW�π�p��?4-��-�*�^S̵cz�鴮,�C�z�tA��:z�͙~��X�T���B{�&Nd<����`��'V4�ƻ��|b��j��b��|	}��4�2���,�Q��i͞n��AI;י��n��qE0<��o���$@b���<�8��G�K�X��c�t�XJoȦ��r�b6������J��v��G�)�w�*+w�1!+�=��
q�m"�ni>�]]WJz��Fܶ�����}Y?��gLh�L�r�~ܨ�@M�*Hm�o��֜�[����$��>f���#i�-���()�bA[0���Y�0�p�8c�i$b��Z'[r^�-V�#�2L�ȹ�
I�5>��%X�[�r_͐��k��7��n�S��e|�ߔݢՓ�%z��Ȅ�|o_/ ��6q����Wzo8S�#�t#Rd��*�Es���Q��/Ϟ�z �ރ�c}y1&T�R�ʏnmO��կ���>B@l�h�!_\�}(�`�Z�4����ۼYL'6xA$���!���k,\�^�f���HD�*iD��v��>��Z?����Tu��Ct��i I��E�ڲ�Z�[�K�zyZ�kR�1��^�M�_�|b1�ҿ��!fU���AO��108���=����P�Ϗ²��!"�=P\��]69��%���|,3������ {$,�7��UG���&����)�İ�oz.��o��z�tSh���/���Dd�E�Q����BL���>H?g��t���S,Q:	�l}b��M4�+Zk�E�*�^Ïv���t�.��1p�
�l�s��$��s%z�D|���"�y����o(J��kO�����Ʈ���F�]!,�=�1�"���
�ȟ)E]�z�&9����?��<&\��oQ�yJZ�$�Ab��#ب��h!�S�j��mαõX�&�i�!�C%J�Y?����YM���S9?YjLXAq�*B*����6�@�Q u��G-���b�t���̍+ɥ����[�;t"��X�x����t7!{���i���R�eΗO���ㄍ�D�VW�>>Aag������y��q7��3���rW�ɑ�L��~[��ìo҇7-p�a����.}�B_����y���M��qz8���| ��?��+׭����p�YQRuN$�q�����*����}���/XlMN��0����M�����*<*��iY�)p)�Q��zIÞ�~�{���uָG�X|����_?�#��<��-ߚh�E*!�{�>�s�Ի뽝���H�� ����\�
3�^I乔~>��tQm�g���ka^��씓
��$zUE�`u�}`T�EER�,���p�?u��:�D�֢m$ǟ��f��OD�A���O�g���G���NB݋�f�R��߂�1=����&��z��>JgJ*5c-�M����qP�B�U�)��0I~!�p5�u��Xf�,��{�� ���I�CcB�`�doR<u�aז���Jߨ�ǂ�3�j�^��ޒ��9�>n�9��2�+p�קLF�$�k<=�:���R�m?J/0��6"O>@�	�ݤ{�z�Լ�g������ؔ�U6��5�S�ғ���i%�a����!p�^LH=ȶ����Up�QU�b��NqS3���F�U�T�\�T*Z���j,�;�v��3e��[Q����D��JCN�XI��uT5]��Q��n�W%� Ɩ��n�s�/M)�K6,���˩�v�;~׸��R���+�Y޲H����c~��aOJ� �e�r��4���Fp��g���GH�OA�\URT3��:֢;S��A.����3N)�*1T��lCb,���?��[���)z���8�%��ʣ¾��͉bjPߵ���z',.�/���	#�
�ay��H�T>rU��*Ս)��t+>$����rs'��obݸ�$�O5���/�9�%��5c���b�T��8y%99����$@������dȍ@SP�k�g������&_.$4%���T�s��(���߶�-��lJ�ѓDʎ��ȘU��+m���5�������<C���j��ɷ�xr��"\��J��q�
o���QM�RF�����@@_?�-�� Ҽ&a/�v�FAk7�6�5C�����Z�-�(���]��v�q���K'��ϕ��^Z�ý�li��{�6�"}v��/3|�W\AY���e�{s����B�w�$f�=:�z�	�m�X�Y��GA�$�y�f��ِj��n��x��ˀ��a����;��T|NU����)���3z(�u,~�T�� �v-�%�Vs��ՕOE���*t�ef��e @��i~+�&��ȯ�,	Wk�[�vE�u&�r�u47�i�u�WZ��V���iA�A9��f��>%!���s�z������٩V�Ģ�d�^�%{�5�k�t���0�G��Bl�4:v��m�R���
�Oֿ�6�R�1k��ˊNv��T}��|)x��x]ξa�����K�m���� ��ͨ�+��De}�Jdrt:�q4�x	��wRڏ �<��uc�I��7s��4��o��Mr��~J��6�ZJ5�ɱ�ޗ����P��VJ� -����ڢi���	Y&*�wCu�jt�o�o��Nȇ�Sq� ���{~�<���߾�gC�2Ti����Q��X�4� RM��=|=vX�{J:��KXU�3��S��s�JW���}�U�dq����bs;J�§����4!�USEj��=���~dG4JLA=Y��Z�y����l�8'�eٵ�x�~��o�DK5k;^'lǌ9\�|�����`/�>4�usjq�t�S=x"�G�	�h'�A˝6@�o��]+��%�} ݲ�TYc�SqqS��`����r����Q%�����V�#nhCL�f��F���;S���H��{+��V6���o��>w�p��H�^್�� ��{I���;�_���T�!xn���­̽R��F��#dm�^w�Ӷ���=yE?��KC���a���4�"�Ni�g��$[g��̣��d���@cL����J薊�xn�L�F5	-i��o��xM��,��v������S�!�@��p�3?������,�=*�El���W~mr|Y��^q��p��f�$% "X��~�k&��
k=��5-�`J��^w+}�c�<V*�q���?67��M�,�C.6)t0A;o���~�E��ŏQ�O�#k�` �4�X���;��&���)�<Pϣ�@����-���)��{���I+��@&�ld>��#�|�����T,�ⰳ.V�� o����ٹ�>�W}B��_QLC���.��5�ڏ�Z�G ���c�w#��omo/�9��I3�@��"g��à�6���P���H.�7rW��.��Z�	dwwp�O*zϒ>�����K2E���>�~�p���x�*����E��d�a��&Z?x0���w��6�>#����-�գ��4��L��:E��zX��cY�\0|^o1��&��9P�L&��ý���I�N$�96�33�6Z�E��TH@��y�U�EΚ�L��D�4j 2R�q��7�����U�m'eꡌA��Fl҂g�X����ƮcL\��|�%J��j�j�w��3��Þ`���-��
GZ�^�U��#����~�x����,��y�;�6F'6}dJH���3g��P�8�(����_^��J�ߥ���%�b���Y�oL�c����eS�t(�4�\�e[\R��,؆�/x?�R���8�6F!�;��:���4S���rj��F��������j\�b�GJ�ĥ'�h�8���UҤ1�m�h���8vN=�m�No���0r�r�ls���od�(��/1#�:�����l�D������x���R����+�|��Y��z���|�p8����XƜ�Ն�}l9�E�o�9����MN����1
�ܿ�_�,y�UZ��=;m��H���[Ý�pv��u��\�I�uv��9���Z���WǕ����U����U�d��ɡ�^P4�7O�Wx��}��1�V�'a�ۥ(��;�r9�.\�̚��GPZgX���G]{���ѕ6/��8������f��D�Wj{�+QLh�0����vl����L��6H-5S3��U0�,N[V�c͈�2L�SqW=�6$��6g�	��}�2���˟�H�
04�%�TgU����^�����ti`]���v��.�/�������M�����m�I�c4���j���^������W)q��مK�^�C ���ש���ZT듄�#�����M4�K	�g�7�$A���x-��h��KNzT���\N+P���F#�I�VZM��	B�t.ue؏s��m��2b���:p�;��=�_�'�Z��a��C-�v����3^�&��醂�]v�n�\W�O0k*o�!��(��>��Ǡ�o'��3
84fμ:��}�j��9]���y��I$�Nv4�m�T��y\ �"G���5����ݒȵ�TZkQTa���Y���~��Q��������G���	̩�ܼ���YPP��켎�/X��h�z��]�s#;>@�,�3/��f':kk\y�э:��Ş�X_�L)���	�	��
�ښt���R�����5��
���y�4:$y�m��꽖�kᆇg*XA-�g*c��n�]	�p#����@D0������1a���ހ0݂��'Ck�wMJ�B��?�e�=ˍ6;䆴�� ��t<����/X2�ז�W?�<c���I�j���ft�K�8�5觛����a���pT�a�;7���4��#Rw��t�����'�����I�Iy���!a�3��6�G���t�a��c��y�vy�+�٘�N�Q�{�����8�����?T����
X�U���یiܠ����\����U�Q:x[	��q�H%b�'�E������	4� {$�
߳r��mYY3̱&�jy��]�v�:/g^�J�.;
�Ȳ��ޙ��S��"�9��3�_��Lw � ��G�eoj*4����vԞ���r�i\�BF簠�ǚ:/6F����b7���9�p鎩�H��*��R�$#q��uX�xP\��n�;�����V�M?~Q6��ehܿ��Dx�1QJ���U5�����k��<.����*��l�.�Z����-@C�_��4|��fV��=��Z['�:�]xa61��kӤ�];a[��^�LN�=�D�Y��X�A�hY{��E;���j�6�4�����^4�.z�(d�To�pp��`R<�\_���S<��������!��f��|�5ٟ�9*~�����1���e>t�d���AV�v������Z��������Ԭ�+�'����^J	v]5���b�d�N�J��ֶ���>Øh�oa>���Ey��{߻Jd�A�gN���;��	#bP�j�Ds����k��Դy�s�=]�k����P��O��1���5�b�Ű���8�^\���4x��ߜ�Jj�m���������&�R��q�f��H�x�x4���yD���+"s���c�u����tJ��?����� Yb�����<�Do~�Q �����Q��o�C�]�ڦ���,��uܤ۲=�٥����>������ૼ�հ)��T�����w����/; �ZU�I�5/�������b-{�XIVC�G�Hf#�%��q�Diy�F�
"E@U@y��
���]�y'A���=/�m���w9OR��\�F��(���ʧL��E�f˰�PeZ��yh��W�/`q�5޷�E{���__�ؓ���j+2S�;�a���8s�K�O�_v�ր��!�EbD��~$����Y��R&��<
�ϟ��>�ia�h[k,���b� h�WO���}��n��ĝ,�{�w�cG+EW=l�t�!|NP�ݛ�bOy=�5�U2#=�:��r~o�Df�D��|#��wx/��ٜ<?P6�b��Ւx7�n��֭i�D o�dy����՟{��&���y܅ r�̛��$� ��6X~NM���~�Ԥ��5�w�'Ӷ�=��/�OB�!:=�{�6aEk�ٛ��q�W�%�5���5�w�v?�(C]�����ak:��I�!K�����^U��w�����ҷ5?dC:��%���:C��nW����9п�

j')�l�\n��[�A1V�_��h��ǣ����d�}�h?|˼����&�)�r�;}YA�p��=�8�#�*��%�����5��0aT��ih�q,�����&֊� �>�0�ڻ��E*}`�M�N�L;�)�Э���M"8.��ۆ{l���C��:[�o;%'�M����C6�C�)u�VFz��uXlA��E��[xƍ�Ϙ������-��_���K&���W-NM��ى��,Z��D��e>�8I5�ӇUlJ��ͻ��f��N�sr�^�B�qQ�{�x��y[X�j�|�(������C7Q_&���y� Q[�pښ�#��-]���x��H��$O�	���/v��������}�a)�&���`\w�Cjj�bh�(�0�2�y��\E�(�}��p��C�e�̟,eO��w��&�M'A�&h2b��t=�����>�3�3-�B(��$9���Km5�h뵄��v6����SZqƀ`bU���,���(�[p����#�V�l�s}�n�_�����9��a����<�V�Şa-uc��C���
����+�;V��d���R��ϼ��K1�����N_%Gv֕)˥)���I�G�\D����~��z?9�fF���Ք�5b)\����3F���5K����=�_p�t{��1���]�D�, ?�=n�f����;��f�Z�qb	C�(��_l��� ����Mo�Zz�嵺�x��OE�J���N�]?&Ո;?���7&W���J������;	�a(w��2`�j����S4л	X|o���SL��/!_1�	��m���G��F�q6����}]���U��?�¯�������)>!_��\�н�� I����#71�ޏ̷)����'�iX�*���Y��L���*�O_�wA�X�T[�{��q�0O�O1��3����\_N���������Ӭ�k��TW�
����T�]t�zٖ_�:��p܆�x��ӤU�b ���֖�RL3Z2#�k\,?4ߡ�Y�6߈+�eÝ��O���Rl3�g8�0�J���*�v��z�݉������ݠ�~1ix����>��|֥�̐��=~\TW]L�ٹ��i�kMZ�6�]�(�
}]�Gџ7��!1 h.Z��㺊$%�&H.����ϫ�&����
��4=����$�'Z��^R���ߢ�Ҥå;I�RJ]��n�p��S���/=��w.H[4���5����B �$	F"ԡ1AH�t�?ŧQe0(����.���j��Ob�L���=���3�(x��)Ԓ�w!����hI�xԷ������B+"������?�ٚ!�&����,�K̀KJ�۴���.y��)P�Z<��~�-<=�ñ�z*�:���p��*��Sn�*{'��Y1O�����_�l�nS�l�S@w���X�	���'1V~�I���� �wf�Th��q\������V	�2�{s����ǡm�X�m���L���\c�,�ӑL��kQF�������t��2T�BQP"����w�r=x�К��{׏l2�t74�$;B*���ĺ.x����S�`6�����xTL�k�۳Kf�N�����ݏ�	c�l�Q��l�����$/ϑ��oG'E 5��H����E�4PY-g"=p�=A�ޔ����X��F��"a�M� �5c$�+���C�[�$�5���9RP�懈��J����
��=F`[�6�ݑ�VKY[���fͯHN�H�N��5F�v	L��hx� �����d[���`{s�&zׄC��Ɉ��>nc
a{Q�2���+h���Ys��
�B�7�Q�(�<�6�S0������7�5�����)#wmq�p^ֱq��[%��^Em�6�)|čBp��2Qq�3�6��:�`��~�Ў���7U3LJ�>���ƞ�J����U�ο��S~{w]N �SQ��°aÃ�W���i��c])�;�RJ�
�l���qM�T�e��M�����ԕ���
/C�PK   vOX�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   vOXǐ]zd� K� /   images/972a987d-5ae9-491b-9c1c-35ff468aee03.png<zUT\���n����6xp'�C� �� 	'��4hpw�����ǽ���sN��N����]�j�WW���I�	  p�e4  �������u��Bp��$���< h
2��^&'�h�����*kE�g3"��n2'�5�k���}��z��k��Qr*��zQ�E���P�AU.%}�����	�;ޓ�k�EA�������5��Y����� w�+H�UhQ`�����	�dC��_'$�Hn���o�)B�х���Զ!b�`�[�������߰5��:�r�v��khL �t/�����v��K_-)��i7�8yol&�ө�������;�FF;����d�^#��D�a��|�����i�2���O,i�B�K)����SJ���	�d�`�-ǺU.��I���_�a+^��G�+�X�Ǹ��K/R>2��W8G��R�%�.��*ou�G��/�H�9u��{<i��'�G���'�*KR���k��n3V �6\�;l̊�n��K��x9���r���9�/�J�h�~В,y�t��J����L��H"ˊ��r�k\�}ff�ƟgVH�a�
�q�,T�l_V]z��)���<�#=�B�6f�z!�]&�5��.;ޤ��V�������r�{�n���������)Y�km��~��$�� �gz�����̸YN�#�f��x��~z:ٞs�t4hӨC|rS�ǅ�9?�UFr��?M�?����|�>\�5En�$GF]��O�=�_-;���>|֧=�!�����X�38x߹�s����SǮlћ���ۂW"K��� �r)��pﺐ�9��_��vw���ֶ�NW�Η��G�ZVe��?����Qۅu��|E�켙Qz����̮�+N{�%��U�ݪ͚D��L���Z"k��Ǆ�J��%�k���< �z1�*���Jy��DͶ|Z��1��3��
�ٴ�d7��[�7�s��y�j�sL�kH�\�o���H8��t:�5<�+#��6?̮>`�H��&)ο�P111�WwN��ڧ���*$0&}h���:%��d��d��۱�5���a쳨*����'�A!�+��G3�)�t��]E�0G�4|�@�����]�=�'n
3ާ�����0c�oi�-3g_����Y��8;q�t������Bt1pVc9#⣙�tӷu��p&��������(w6>�T��i�
��i�|4��@k�lHش?m�J���敒9DX�\N�(�
<B��T0�+k�.e���3��	��!���*���l������Fυ���w�o�Yz�]O���)3��P� �������Y�E��a�k���VUq��in(��L1q=�5��s��,'{1��L~ ��d���<m�t��n#���y5��ξȸe�N<�B�x�h���0M�}��]�C����4�|�ʯ�;~�\���<"1F��0���(����cCgK���;cqC�d�����5IZ�ln���_�Q�����Wnr����Y"�ٞ=�%���������g�)~-�����O���%ȈA�����cRdR�}t � bn�����8U����d��>��i�����IN�_?!�}Â)�ӃfN�j��z��{	�E/�vj�-��gBrh���F��FX��AꜾ��h���G��I[�l�Dds��if+�Ṳ�q��>�l^kE/ݧe��>��߀e����·\\�������<�!���GPeG']4��k����F����?TE-ݐ<8'k+s�0��Ш�����x]j��U`C����]�D������/��M�'��⚊�y��26\U���~@
ش�+K�S��CZ[w��`n\���p�A�u��h�x��fcƷ��_�c��N��!/���*~G���Le�Aċ��
2����!"�0m�Oq�ّ��o�v��'���=�r�1Fحt�i��BC���يO��]sB����n��@����1��VМ��K(�}������	�}�(��V���%t�p��UI'�^�P�7-��K}�:>bk������Z�S�W��T��sW9}���}#�>�~�����Q�bР���bBt�rF��Z%~2�c�����������B�!
ؙ��μ��pu�S��Ɏ�PF��Yۅ=�5�[�e�J�$����sC�(�"�tc��2'v����%�A$d�9�z�����w�TmE��꽍#�)LP-��>#��W�.vw6=D���
	~ �l��"�n=w����p���Q��Q,��j��LK�7�vU�6ϔKX����{�����3fݥ�VH�����W�+�s�ȵ_G���fz�+L7�e�8�n.�Ґ5�2���#Λ�N&-�Y�P8�CC�g��|-:_,��{���4�zb�Ð���Qң��P���I xP��� �@��pR�=�� �Pm�3��|��l�Qd��5чV���A0�}�v�{wS�� ��jX �)�s�e��"E�"�����kF��/Oi{ �n�*$�<氿>�O��4Hg_!1�fc�U�8�c��ke�R�9)y�(�6N��T0�tUi�ܜv��]�e5씪�ٓ�f��%��,�b���Ǝ��/CJ����zd�(���!=����*$�G�kq߄;����s�r� �QZ�V��]��zE-s9��8���ɛi��侮��չ'~�A�s3�TU�����#�(�G)�-�K�=�m	�S��S5u����U�ܮ��T�}[n{���H-�Yc���~�ը��{�����=����\�����3B-����RNB��_i�J���8v;*k��g�ܶ[����AU;F�$]���2��.dA`�� s�w��8h���~��x�~?Z@�뚸��\.�pD��O�����h`���@��X�~J��K����|O�_�᩻&i�1d��>[�7�:�1�6]�bW�RC�E|6"4|���l�tn�#]��u��J���o������a5��/����o�{���-i�{nu]W�; �z<	���_��(�֫���F��nM��d0��۵�@ ����ˁ�2�v�t�Oܦ|k)>��+4� ��=��o�/�%��~���[�92��/]/{N�ק��}���ވ�&���jwP
��dm(�AN���z8����%�Q�Aܕ�����@�/�U�s��D���gK��N�����WL�G��un���!���O�U��f6�2�*�?`�
ui����^�q�*_���ٷ� n1M�	O�����Y�|^[��~�R���_1�~��~��|�;��bP���"�g��訬��b3,{tt��� �O^)1aw���rнvZ�q� Jʗ�)�5�+0�n��y�4$�5���Ga`�Y���H
e�5F����~<��Z����s[�a?����̴�P�^{���>�r4�]��f�+�l��1�tߖ��o�W�{q�����0�Eد�?�$E����.��;w5�R,8'T	�?qepF��zf�!�UX.�i]Ͷ��S�/N��{i�����Ǎ�����sEc�7Za	����B�	O͐�Ւ����=<J����fE���s*�U���2�
�'�N0���ߝ���m���A��՝~���~���ߢ~M��ņi��j��LŊ�k��x���f��{�s|s��Κ&�K�-z�$/�g~���T�5~*�+�gr	����>a�܉b�*��M�J=�Ӊ~��^�7)z�f_��$�����5������o)�Fp�MQ��N�B���u/<��ڬ:z���='��?���J&�:��8����U%���� Oc1c]�O�z�h�/��LŶ7�h�\!�~�7)�II����"�����S����y�J�M�`���]�m�MN{�xh���Z�s��ƚ�u�������/�D�r��s�2�`S�s�7c�>�	ճ�'�}S����Ӥ$�����J���WLV�����5��t�����K���x����q�kd8U��4�?��?�O��¦�T��_�L�:�,W�^��l��H`T�3��P7d���3�����(��"����N(^��S�Q���+�K��������⼋�Ѓ%��	�y�9����݉���~�}oܴ�&k�;\$rw�J�`S�����A�ۯ'�u��n�|^ú巏�㧳n�k`�'��S6fV�x�M��� �����v0�ړ���*"�9��
ٸ_��`n���9x~ �e������\o��:���7�%&^���k�?�,܉V/�B~���Ia�3�q�=N ��t���=������-�dU�w�$c%���>~���O����c�)�#�O��4���w^�H�R��I�Jq7�@a�E*o��u"�E�F�L����̬m���M~���;��J���S0HiJ�2���lB���b�����OW�Lfz�g��T�m��ԏ��	������-����;��Ґ�(H�I`�.[�%���(�<Pr��8F�"01��>�/T�PCS�:�b���(x��[?��I�������_��5O�)����� �=�m7��H�y���c!#�Xm�p�P7<`��EPD�����Cm�?!���[1�.��^���l����p�6� px:v�ⱡ'8T�,���r	��X?b�@��@��&:�̛�L�*�׹��4�J�e$=�{�
:~|g����|�!������:N��$a+�9������*Z����j[
Kg�����}Eze�j�lM������B�Ϝ*�I�@=��6�/�N���D�W5m�}0�� {a���W�q=?eHP`9�!�����VQ�?����*rJ9�q`O,��L�H�����������K�ݱER�a��@r�ȴy��P^H��`P_��u�������I�U��bD@?.��^�Mv�wN��n�p���[��a,� ���B]X5���?�qzP����I���m�wcK�lE��5���OYh�,e:+���靏b�HA�^eo���ybW5X�9��YBޑ��T�Sb��{ni��z�p_
R�o�4pc����i�Z,����`v�d
ėbv�W�!�4�wj�N�*���y���3�A���[�/��&���fX�d�oC4�
���+2Z�B��$R���
 YSu��P��G��L�m�*�+���mVp�]V�ix��%`�/�]E�-"�w��M��< V�7�ȣYL��k0�P�g#��ڌ������`~o4�c�0q#Y.�4z�������e��� $4����㪙��f��zǕF�S6E�)�+T"?�Sq�P�ߚ�(��l�j�����{��w_W  ����K�ru���-!fjm��18��="K����ڿ���Q������k�uFDgD���?j�KmTk$J��	α �X�����$5�1,7��~�����d��]k�����)p�\�n��.������F�{�jƎF�d̴���mX�dvg8�����3WHC__!�ԫ�[��[�	B+>E�2��@��3h��5���'��f�}J���zF���6>/M�9�ϝ��^M��b����[�j9��9-��*����Uʥ�+M�J�m�l�U���&��7�䢺����P�b&�.��_�1�N�y�>\�z�9.[	���ǫ�K�<�����Im��:�m��?�+#'?Q���ǟ� �J��OXgv�>���{9��=/q%l��C�f�:n9�*)&]��'�j�LNz!Xkd�&me�<Ԉa�J���O'��O@��4h�wL���ZYխ��xQ�C3�.#QT��R���ٚ\3	\Ԥ���ے(�����_�h�
��}c���U��]�_���Zj~�jr2eec+��d�B�:B���I��^�$I�#� �N��0�fe�q��gOT�U6���� �f��]ۑ���}\���b����:o��ɗ���fb���\�茆�ژ!��Y�x�������P��?8����nch�i"���շP�Άh�'eP{��̻����{8i�wa^�b�qw�vt gls~n�����@�7�JƸգH�_!�����t3�V��Ȏ��T���|������� $ ��r!�8����Y�X��;�7�2W"*���+]�Ի���2������o�P%����C���ҍO���6v��V�)�	����X�$��w�<�l�/�}��h2ǟ����ӛ}�K���	��Ҷ���]�(Wgf������Ѓ�	�zmmu�%T(����F�sY1n�O�+hb$�$Yon�w\2��Y0��r�9������=m��������h$���Ğ+}���ǭk�z�Y��Y�+Ĺ&5P:���H`�%r�|��%�sݛ�t�gw�i㊗��]S�t�B�A�g^M@�'��@T^$�_�l� �x8=�"=M���w�%Z�2�Y/��O۩�'u�:V�2�U8֊���c�v��C[Y���:����0�����Xшo_�������Q��<���Lhܦ$ad�{&���w��E�<��*�!H�u�|�^��M%AH��7gk�8��%{�� �o�̸�)�����	��O�	���	����)���@�����A��A��kD��>�t�m �D��8�A*�m&e�J���<��c��U�I�p'<��]�+�Y.ܤp+����MB��~���=�cN�3�������m\�lkB����W]�ǩ�P`ӼC�gЈVֽ�&���b��p��.�<ߟa�/ۣ�6a� q�L�o�A�L�^t��y~��e���������?B���:��?#;
_NS4{��/)N׫��Sl�f�'M�2�X����<!���ݻ�{�F�W���n�'6՟�����6�̤N��t1h����e�j���^�d�"r`xC=By��K��L|?s�����卟�h�xPuR��r�}��nc�0;Y�m�	!8�A����&���O�ߜ�)x��!2�:������=���7{P-h����bШ�h@41+��	`���}4WF�I��k�!WhS�L���}�9��"v�[��m���Q�6IU�m�gY\CT���ǥ�ĬG�)B�Gs-�D%���єj7������/>a��/�:��uA��
��Y�3`%��Rc_�x�3{��d�Щ�r��p�i�XV,�L�ڨ.�[�n�r0TS���$�'�x�����]�	O��w�\v!�FFDx�^�͂l���|X&N��3���P��^|��؅��:ϑ�\ ������ �Yq���-����q��C�J�z�@�7�+&mk<�e0��~��t!�b.�OY����R�[̘z��p�&}RUm/��ҿh���ߟ��/I��_p3$��#��Z��&'p���ɴz��o�s"�X2�)q��z"O�)�.GP��X)m_+����'G�u*Tŝ�kHҭ��.�mȶ�nX
�gg�P|���,�%:i�.�"����i ���3��qS�W����4�R� �v���esCd�~��w�.��u"�=s��bv�NC�  �s�0e��h��˙g�h�� ���8x*���Ծ	���R׊�5��᭦�{1g�jֿ����_�{�Ǥ'lRc�z�#0-���Q�4�41~��-���)��.��������jFZ}RJuq�L�*`G����Ҫ�Վ���r�J���9�ի�h�������m)b�/u��.�<��6��2�BM��-������s�O���U���~��͙/�dyd-����[�Kq�mXM{Z�/�] 52�"�T��-f�\����J�k�V�k���U ��C88/u�H�Ġ�@��y��n�/��(�Hq�"���ȗY��ea1B�4lOeu�g�kJ����s��͡�8��"�5D�{�����+05�L>M@��Dy�e�l�I
�ȶzw�����A�����a��{o	�=@U'���Sd�^�����ytz_�_����u>̷Iw��mћ��܅
�l9O�sF�����|5�:���	{V豝�A9Z]Pg�{��~�C�Ƴ*������1����3!��(>��S<WcQ+q��c�վ.Cy�qP4.�x��ǈeh^qU��w��Ƀ�a�rN�d\�%�3�D��]��	� �4��fv��E�c��6�^1E��v�	��_�
�@���r��l~��h��{�Ag RP�~'�r��p���1*�W-�/
�(<Ȅ�ʐ~�Bu�켓� ��hx'S��A��6;F�q6�E��>տ�fUZd?z� ���H�E�9,�GE��S��$]/�Wd]z�{��¹��Ju�1�|�9>���U#��E�����?��R!v��%�
ٜ
�hE�"n�漱����5T�-�ٖم�ݮ,)J�ܨ:n��$�A����h������vK��z�GS��+&�J)������z�H�T-�Dج�4��3�LN9�u��`�y�
�>^P<�I&7��/��%:��F#���oɒ#N氎��d�۹Zs>o&�4�#�'A���)�f�*���#<�Ͷ�m�w����?d[���8��ƻ�U�ET��L6�J�D�:go����&��[����(�� �D�E����7�y�P��;�Ks��kn�m�*��r[Q�Q�"dH� ՙ��t�_2*(�:��z�n���B�Qi�N-�;B}�ژ� l0ZVnD)���
ǐ�2����[�;[�E�E�,D�Õr��,�%ܸUx%��&�H��:�e굉������'#�X<�7B2�����R����K�Xoo��&,�T�1(s�<�hM������+W!R�g.:�O���";#o�~ˎ���a<\�{�iP��ś��<3;�:�=��nzg8l�aC8%Z�*�ŠÂ���o�����4�&�·��X�*�㢶B����츉�˧��lo�a:�3 ����T�;�)w��C������R������y���Wg����.�n�&<�u�^���rr���zȕk�8�|S���/�� <�w�L�Y�;ӛZL�)D���k�V�����\������]�I��ӹ0a�t(��\�j!̾��\�x�?�G�i1d�T+(K�<I�,�i��w}���k&G&���P%�D�Z	��5˘�����g4c�<�۔c�;0)S&�K�;�����<���Q��ϻ��ZTt�]j��J���l�}|��\��UC�y�Z[�Kժ!�E�Xhucw4%\2#"Al|��ƀժ�.{���q�L�/E.TC�oI�Z�x�b:UQ�1�!�)�5����DšR�*��_�z��$[�)���M��1n������cbP��4��
h�����V��"ǜ�?}Ǜ���߷ߨb���Ԇ)#���j/�����ٹ.��>�����t����Ƌ���M��V$k։�$[8�#�7YYX�z��q�n��L��Ɵ��.�?��>B���s�8l\ϧX���ZBb�$�]�8T�nLm��'|~?�ʝ�K�����-��������u[�X�6�Y����[��K�m�$)��Ȧ[�'��c��cɬ8f�7A�W^�|��p����?"�WՈ[I�$�2�w3s��a.Xl�u���CPl鍍�[���͂Lf�����Px�Z�������;�4<q(m�o����+��%�w����:T��=�9J�4�[v���@M���Z�<+��#	�Y�\gzj���;��%W�7���v���Z�����gaG
&��o������uo��\�*�Ci�Sd�齅�X�K�x]~�k[Ä�������pa8��'���;����J]`�}pF�$k�aӿ�]�b&j��ZHJ����[�Nj[��{u{����m�s���N�Y��&ݙ��qw���x�2�Ѭ)��W���g1`KzI�-nzX���_N���-�#�?7j`��r�/[�D���\>�u��L�Z�13�o�B�9.���h�4�$i2Y���"�����,C�؉Υ�-"� ����u��p���ꢁ���g@�������۱�`�=I;���&j"����NmJ��am٢�2WP�&gr��#�2�D<j H�(W���B=]��?���Nf����/N;t�"���t�}�tOF`��S�+jRԸ���d��G�����i�H$= %Z�}u{c	M�0];RJzD�<S���u�v�Q~)gʎ`B$��Hf!��+Ֆ^���̠���_=��8ABL���Bq��zb���R�W�rImK��� �WpK �=��c��I$��3��	�Q��_���z5ʥ�4辉@�:,J��'&bY�A`�xr�s��sm�hD�&�+9�O����tk����q����Wr��`~��� X`������֛KS��������������)��ő�x/eV�C+,v� ���*S��yW��<~ �4� ?�$�i�C���V��w��`�����Ub�`������Y�%��}	H6��P����B,"�G6��xW�C����'x�H�T�����e��W�<7T�GN�����'[�caE~Ks�3�JGN��t9���3M�_Ռ�-�y�;o�S�������zC�c"k�%���6� �b�e��x\#�� �q�|��9�s�]��eM�fV�E�/��ą?&s��:U%0Q	e���F'�ڇ��U';�C:+��wބyMy����*Y��|ǫU{L�e�,�9e&�n��«4h�&�4Rݴ��&�K�N.�%�Z2����\،�z4G����lk/V�E��e�s;�
U�����du�`g�sҾ�$�9	\�������beJ�P;ߣ�aml�P�y[�#��������_�a� ��ƶ�s���� ���n�
��	���nҠYD�OY�aM����y���u���>��f<ݽ	N��Y�&�����eq���{���9O����(���&~M�� �Ѓ!��?����*��!Ѷ#��!Q����V�C,H6�7���0]���ϭh�h�c��9���{N����?�����h� �z:57Bb�Dy�D_%�8HB���Ys���ęS[JsY���@A��O�^&�9�+�k���e��(�n߹De!*���-�a��58��:�C�~��p�fiF�1�1�1Cn�������DJ�m!лTWN'�,����8�>���A�
1����c��񥧧��f2����e��I��������"���=��!�� H���=c����rj��,����|6m۰�8!\˱��Zo$�;G9����mmy�cm�^�QgHTxIƕ���N�8	����˭�Uܐ=�N�>le>�|�i�̀�ާtt�x�7�u�<�o�es���"C5>��h�c1"Vo�l|M*��q��wk`Q /-���$�y�w1�@�����Y+��]w/+�� ,��s�׺5)�}5~T�a��i�o��hH����?�b6;���OL��5�|C�i7X�<��Ϩ��<���+?7�kao�`D�)@Խ�ː��l�?׿��G��_֎�A�PAD��Hj�#-��-�xi��3 �'�H�H�Y�-�"b6�y9@��=��zW�A[O����P{f�)���*¯h����3�B٦_)�4/�E2m	?�M2�h�#d♍�L3�����G�7㏕2P~.�3N	E����������ܝ�B�y����yO�TA��z�/&���BP�d���u�;`v_7]|B�I�]8��Xn�2h�87�{݀�%�]#��;�����ʈ�0bA�� ����#i�a���D}?Gћ*ɻ>q4_j��^q!��?n8x;WR�@!o��(��B�Z��hh���_�|��§r�/Y�(\���i|���S#M��5��O#m�@} 
ܠ���E5�������'x��\���'�y��̅y�Ɠ�ѧ��d�>��*���&�Q��tI�_1���3�`;������B(�:Y�P��`�<[�NŘ#Ή(��op��Ѥ�y��M�M%�j�w�Xۘ7֬`����R,���/Uk��0z��?���wD�0�V�~i>�"���/W�S[�?V�DHBzs!��5�(v����\������fDh�PG �������xۙ�����
�WR�+�j ����x�Tt��p/�$���������ĉ��;	j���j �⎸���ƊweI����	��k�X�13�\��ݓ}�
�_w_�����=���HO��m�v-�S�-�U���8I�N�����Ln�
ɭ�s\d�ɸi��`;`�Y[�Gji��ґ5�*��o�!�C��)�������p��a�z�Jز^%ʔ� �� �.��;�X�I�Q`�G
�y*�xf�3B��C��@���%"�<>ܜ���7��MƮ��b]���o�m₌O�<�A�@�g�Z.�u1z�����D�΍�u�S�fo2-���I^�R��t��0��M����8����H��h�ff�8��<�M���"v��Tؠ���f�����z�՘C��Dٟ�xɡ�oe�����paRD��W��1m�����* �k��<�.� �wo��.+03�W���[���bUQ�g��,����T����џ��l�-�+P�	�x�Ar1ЀBc��1���ˏ�wJ�� p�oN9+:@���8��RKbBN7�N+ӿ�crrO��[�=.�w��d(/fj�lV��&X�;�ϱ��ຉ±��@�;�D3Y�bCY�L�)��@Pa��6*�S��[d=#�["���R74�����&�֦$I��1S�d��[7�;t�]t�^��7B ����q��u�N0,KS�\�X�(�8��C�q14�*!�B�^Ϧ�������ę^I�~\,ߦ�Sǀ |,l���[��!��z��[ɲ��JS2��Ԩ���L�x�����6>	;�cYX�S,od�HK�0�i��ᓎ���o�m�Z/�ӻO-f�U�F�c�7m�����	����;YXj�̓(�$���H17���x�ӻG�.��Y_y�vv�	�tww���mrTRFq�+ι��nY�tj�?Ŗ���uY�{砑y�o��6�1��"��5�7#��1Yʴ�	��ϙL�x��+Q��&+��Z���Y�=�3�֖q�K]�*:I�����$!���t�Z(q�oXI�jdB]t�0 "ÛKΊQ߅��	jɐ�>�!Tz���}b�d)�`3�]��m�Łs\��=��=��e��m슧ў�  ��vM��*�Jҧ���'C�y\F��F�*?r9;�uM��I -v��R?Zy�">�IY�s�ʍR�=�-A�<�?ݓ���)�P��vX����{��1x̤j��Z�c&��O��{�j ��c>�4wp����Db�w]~��"�;j4�^��r7W���t:�0@����;y�o�/�xzX«��J�3b�v?�
��Q�^n���8��8  �y作���5H�TT��\U��XNym�3�����k~��ƏwC��J�H�Ny����|�l᪑)�=����'V������ ��^7cI�ǧ#[e��̜�O���!98p� ���欕�`eF��E�Y��z���b7�(�)���1Ż������ԥ�~4�� ��$21{P�[��_=��V_8�������%����#
����b�����3?��.�Ow@�^���H��t�޶��/L
dW���_��I�:��J�.pG�}��`�eQ~3>�/��A���:Y9��a��5q�Lpr��;&U�a�6*����.����a.C	��u�ջ"$3"0�2F Y(.R�^*��;��+�E�h�|��7϶��]-��\y5Iư,O��2F5���"oڶ����P�/����=Ah>�j%��9��
ճ�����T�����C1�31�w����L!�����
l�ɚ&��s��c����R��D�<RS��:�wc������W}�Z�ꊲ�ȁ��>���T���1_�~�w�Db��޹A�v!<TA�,^<E��BF�>ZX5�k�~Cd�Y$�
wÎs
f��&��@v���v��s�� �:�+�Β��,��yw�5�xr��G�a*+.�pZ:�B��/�?"��Ⱥ�F�ۋI�,���xs(�0_J�v��;W�3w�-Y��\����������Opr�Ao����5�čM+�ѯ׵�P�^�i|�puc��VϪ� gd���������-�9��ɗU��0|Co+�b�o�2Avn��ʱ�H�$p���5�w?Ұ�����+�
%3�B�q\i�>�8�@��ꒈ�q��G�N�sYA��5�(�"�Hy��l��Dc������9�b����>b&fT��Ȧ2�C �(��g�	�
%�$�襒��QU��Sد
���K[�a���p(2�gr1 (��z�=�9�Ш��&�H��D1�������-��(�".�ءF�� ˋ�و��S�W�P��������m��N����<u��Wu�x����H��S8D�܏�q�;f6�4�v��հ�uA��%�4%5H"���= y�1���������*����Eo\���uә����I�F4�"�#b�k���,��g�f6?�;U}�j{-�W�� /	�x�P�nĠ�
��n'�+���\J��OQ���q$"��$�S�J�8ƳD���C�. ~�o��$8F#��/r>󞆫�ſ�A��>E�~K�;���&����Q�ꛡ?hq_�~&s$�V��Y�|Q%u�i�B��hM0ۆ��"/Ɛ�O�'=��Եa�I����J�������e��%�ҀH���EM��,/S�?�D���O'�AO��g�h˔4�A�\����Y�b�:'͎����'Lc~�3^�D���G_�����$�v�OC��-�����?���@]"��J��<��A�����q�Ue)s	p�HbԽ��w>Wćf�/�u`�JA[w�o��u�����4�%�#�4�.�RJg�-\/��g�Q��{�|�gTN��[�)�
�MҫA�9	���c�W�zӎڽq'�E;HG01���-���+p{
6$����Wo�:��MF���fv��f�4»Őh!�s�g�A�p�IL���c-u�N�����)X'k�ȖYQ�N����7������7��B���R0z��	�:�8F�o���ԕ�)��keO��ӱ�MV�S>po�/M�J��mJ	(U�ӎi�V�A P�N_i{ �H!A����s�;ć_t<!��ƥJ�3��_.�$����E��:����s>�S��<��+��)�/Ma��{qX�1���e���ڧ��G���.S�>&j"��~[�´L��onYu�n˺SG�0����jG_����+��#����ی��N��t�9����X����k���g�ĳU�we,�ڥ��tM�ӾV�{;+ks`�h�K	?��[�U"u��#| z>6m�}��z�]������)��ltĉ�O��I+t\ac&_W���4��-U/cO�pܜ��U���J��ݸog#=��s�Bh-�(�TyuyS�@��{����BES�l0�9OBPqO�B?���5Kh�n�3��B��Ry���ѴX	�
/���w�VB��"��SY�e���t�8'�UG�I��W
ζ��H������#v%3*�k}n�coO�j�g�*ptTN��"n,�W4_��;bª80������[�D\�$�:��Q0����S w"i�x������]������X�-um �}Ko�P�b7�~�3QY6U���P�z��R����<�U� �)\/K��w�L[}1A��9JM����y����=3������_,�[�#�w�Lm��H�wEiV�8W^	;�2�ն�GN臚f��a�>��(چ	�������'���r��~��I?++����<K>j���O�B}iW&�ڶo)$�|�4�۩�;Š)dc�!�j}�vs����W�U2�=܋$ooL��4��+TΡ,݇eC���|Į�:k�5�I�?���Q��o�� ��ٯi�������g�u�&��՝���cL4���{ն��.n��Z�P�䉨�$�P��vzK�r�D�%��U�f�=�Ps�~0H�?�ԙY�����Ȝ>��#|nh3u)�'u\ד3lr̽��g�n�Z~k� �mrXWtߤg�0�xH�z�w;�7)�+ pIJ��: �e�ypG��޽OI׫�H�\(�'���Ua�S9L����] ��J�o@��
]'��ꊆ��Ǐ�b-D9��~�)
쯝!�D�XM�o�����`o� �b_K�_��=�������NQ/�ڰ��ķ�T*�WS�0�s� |@���Q��T�kTJ�$Tcq�?�����=����S9�Z]�[Ə�����?q�.�%����?�Dwǎ�裏&#�p�F�(_Ck֖R�����9ulv>?��Dh�J*�ї��VBy��>8k��2�N�|���5sf�|���>ӊ�U�.�� >f�u�LW^y9u�O3N��2�F| �"5�a�z��gì7H55u��2������?�T���/���������C�a��.����A��.a�ʕ�F�U����w�Ü�
t�Q���ߓ���./��t�J���~��ʶ�;s?�0d�զA���=���1*�#�1�
�����i(p����������ߗ�)e��c��~�q*-]Cy>����0��Ր�)�z�L�8�y�B���T�R��ǐ��<p5)�*���i��/����P߾}��4z��_��W<�x���P���V]�VZ�t%�0 w�o}M	D3��`fa��ul�[_���<�\�p�$����@�^�CѰJ#��B��Q��������~���|�̥р�}��%ũ���f�z��<��^�֮[Eu5���ϟO�7m���uDF-/�D�FO��/���n]����x�*����Abp|>8v�}�������$(���|p�Y����}��E�6��үi�UL[yL/��w�U�6��y�Q$lq�#p��}z�,Rn����䂿��Rԃ/�U�v��m�/嬟�d-� 6e%b��E�ԱS<�
��x+u�`�r��d�9_�IlH���?�<��xz	�q�i�����oyQ@>T��.@\ȁ	��W]u;s�>7��i�TX؅/YĻ$�#%+��d�jJZ^ڶ��:u)�+����� m޴�����iM��j��ch�"|��5k֌��%%	�*/���ϙ	����M�\{���*]J��EG~F�֮-�Ꚑ]l9@U�:*[W�Lⴶ���4�P�+;Ā���9�1 ��G ���'��'�� �����6��;Z��m��+)T���nZK�C����p�x�h��-4w�����A�!CQ�>�U������j���z���?����W��Fz�����30(���ѣa�E�xS80�z|A2<�o��CǮ�.�3y��(�08�4=L��,�mٲ�����8�^�o�2oPC���1�%�/�0��0 ��\D��y�ƏF�:���ҕ|m���(&-_��j됴.E��A���N��������իv�m]�w N��JQ����W��9�|n޴�^{�E:��)�>Y�a-{ư!(�e�__���	�-���#���C�zı���]���.��
P���JgMǃ���Ac�r�F�֮YF��WR,VE>R�&ȃt��o�<o���~D�5	��۱�0�#0aT4���j�.��K=�#����?�����G���V��+nG��䥗�kdz�s�"�t�T[g�דφU[Q��8�$�[n���)�{��٠[YY�.\��Q�F��(���о�m]t�>˖|I��7?[�N�hU�reo���D�)Z���o;ڴ1D	�K7�p+���y�>���|��t�L?�}l�#p�WΙ9�QW�Ϡ}�G�z�^}�?�����)�{��tđ�r����5�LD�A�QUU-���@���ʫh�I� h�>�(h�6<�r�<��s,y�a��T�38��sU,AL��+3n A^���i$��IR<
�~,~���h���޼�i{e�?����O�K��u�_�=�Ye.@q�Yԛ�C���#x�k��o��ϋ��a;�@:��Q�1��ø��&�
GԾ}7�2�H�D=���6�����2k�!ھ}���;��4v�g�}�����w� u�������|����u�d]s�5�[زq=�{�%<�7u+�H�W,���6;�;*�%h�7�(�C�_������^�3N��y�OӺ5k�8�����r��!�Z?�Pv.��%]L�J����?��:��R�n;U�l�bҜ���i�hݺ
*��Fյ�}ޅ����{���w����d�>x�W^y��}��!0����@rA��u����LI�C��6�	~�@�$D�'�Q�C�(C�> ���K��oSUu��� !=:\���7�J$��������i�?�۴v��'N؟ƌ:H��'b�1�<�����d�Cy��dz�9:���q��H��g猷�z+��C�5ft������4�#���nc��*�B���4�d"BK����D-�UUo�H���>�c	2� ���Bk�ld�m�Y���I��'�y��ѳ�=G���6� ��Fh�$ZG��O��舩G�9g�I5U���I2'�u�z�Ek(/_��HY^
��Q����P^�*9�l�!�4�����p}��]v�et�����T^^��@;�� " ��. �C܋#�2�[층C��WD
zUvB����:� =OЖ���ʸ�����S�~�bfgVt�_�>�Y�q��i��8��<�ݾ��:w�gy�5T1o@����H$T1x�l�k�Oe��y�*� �:�;�<*�ѝz�!��1���#/8}`�=��C.L��O<��:�(���5�T^V��!�����C��C�E/-Y���7�8�|ew�i���胏?�pK��>�x�6��7��ɼQ<�d�w��t�Yg�AÆP,RK�U[��r��8"Q+�d�^Г0�F��H�G�������/���x 9^��	��#!�����R��X���D����M�雯>���j
�}*7�O���─px|D^?8��L���c��/W�w�t_��8`��7�?%���[����U�D�Y!Ês�GdL�rN/x���ٷ� α��T��OU�CN}�ʉ9��g_PM5损~��0�í;|�P'��|0���do���v��`��F�j�����G��W�i�F�rĀM6�~��!�P��9�D����#�������z�x���4���l�>`�lauG�M�<�N;�T�ٳ;��VQ2���3G������CAC8�î۷��	�@�g�[(��u xб#�� T]�u��JE/|�����2�2В�g���i���H�8}-��y��L��iS����T����={��h���>�d�@8)�'ڎ�$H�I�'6��Y�(��2qm��R�Cg$�|�53i�hX�6�PR{�N���R�G���<<�˚�W�ʕ��r]�̰XK��
l�f<�D�Ka�+m�}%�0�2&^)�g��� ��&��NU��ţ!WOD� n��#*�ߏ$��j:��{��, &g�M ��eRׂB:��cXY�=��Gh^)hc�n������!�O;�:u*u�܁�-�џ��L��s���^�U�V����`�׏��Z�1���i᢯�w��[���1��T �G��:��?�A,���S�$vk����*C�eu��WL�,��փ����C��q��m�����x[��o� F�!���oLd�|����|�s޹��c�q�8 �A0 J&����^ �-^�m߾�>s��d\mg�yLQ���@ｿ��a$*A�i���z��co����D{x�n���[��7��&/��A[�L}�	���:�Sg� Ε8e�Ef�.y�)�+I�dao0�C�����p�ް�����"�8O���[{ђ�幄�D�ޭ �,��G�^Y�2�������	��l#3J�F����R; ���<d�a�MR^~'�<�p�/Š(�|\���\1̲8h�w��s�,��j�5���!+�|�|��ǻ�5d�`���0)�>E��	�1�H�_,`�eH�P�����4�7��G��)� �	w�ѣG�ĉӞ8�M�3�H�~�U�Ѕ�ϋ��%D"|=p}��G��(�+��������.��w���3�������z&h��iC�J%��1�DurMP?y�v�F�;�S��Kp��xRe�D\��bٚ�����Y`c����r_�/�#�s�^��8�3W|'Z����8�8Ydd!�׽+�,���@�%ͷ$��;��v�eW�FԂ'�+�"���) �c��[v���󥾄 ��&� iJ�E@[ȿԻ@_�x����kQ�I�O�w�}��_J>3E�D2�>#)�� %y����Qu�h;�б�<� ��GT��~��ڸ��~w�oc+�?��G��]��c��ǜ9s�D��_"��%0����!�"E�eG�>GL�E�@�{,ؒ.�	��
������vR"w�ഖ�6����$��a0 �m�F� gܸ���v���D͐ÿ�b��z+}�����/2^���g��#G�y�����Z��cၫ'4�>"�ҧioJQ�f;��B�(�f?�R���������>��:�*����ۧ��L�j�}t�Z�P�|�  �F.�s�'1r�}��/@+�X��~�i�jc�$x�#�
-����E��sJ2.NyN]C籱�H�~�|J�|�� ��� ���Y}7%�,��]zۤo�|��ޘ빂�|?�To��c���CGR
	�L"V� �RA��ku�\@E�=9
�5}�"N��r���!��&v����O�;�z ����pA�0�y睼c�Dh3�;�v��(�`d�1[�h>X� �ʐ���?\XTpe��i%�������a�hDe~T@Z�dᓉ*�������<0T&����@�2R�"�
�P���q�����s��>���O*߾��"���@����j�"ڼ���*D�f�Fzo�'�d�챐��Ճ���k���K�]c�	}&�4�
`�J&�l�dLu�_^�e�B�H�Ut@����:��6�_�r�����
l��,$2�B�0�E��.� Y�t�^��m���N�Rr�>)D$�+�Q��Y(	}.I���`G����+�0hp�	����G�+���@G�7pu+�G^�H!/��F�n�����;v�	����{��x�ͷ�G�|���#.�����v����(ʉ,��C��O�%d ���� �%��HLͿ�c�\�^�I&\&���ŕ�`�֪��)��,&%2�q����ė��q�G�|��CI�!�i��G�d��8�A2RaZ�v)�Z��k��^Z�v͝�1��*�����5�\ku�d��'ͽ+%� @���g�E ����`ӵ^L^	�G_bl�ѩI�����'=d_
wX�s�w𿠦p}�nF�`<ڀk�}E9�3
 $���e"�c�w�L�_��SG��<�h�����˞���~�/���P�}w����x�V1�Ȅ�X��=���~4��IdQs!Y[�s�X�9p�>���y�F�����@�����[hђ��������@�z!�3(]��t-� n������@d�q�$�t�v?��

��5k��m��9mz��U���f��(���D��\�.����f��Ź�q��`�|�ǵ�L��~�v �>Ĉ�E��^����P���6Њe_S<���@�JK7л�>J�����r�	�plk<��L��"�Z�k�a��h��������ݔ�1������ୁ������v2V� }�<� ��y�E�Ƃ$;H</�{8�%���0�b?��1��)���� &;F�%��*#��L��DD)<��(4rd;O(h3�Aa��]��c��㑘���a�d�v E>�z�J�HE��&��7n�rD���C&<�z�N�(�x�����|ҢD
6b��kp,j���+�p�1��9�}�)]����B�!��E��cA�� :�J�CY�kd�(��nW��1.���"�4�6��5|ݧq��G��k�2x�Q�V_���߲ʋ�&a��	m� �#x?�t��P�����~���?L7�����Q�I(Բn�&zw�'\��4����O��;x��V�G; ~�?�8�O�X���� _{��B�SO=œOvm22Q��Ȯ�>F�$�ɵtZ�Q{�^` Zl��Q�M]�������N���0��er�f'FTD}��w~>����4�u0?�s�[ ��믳���_b��/�g���}�a�~��/~� Bd����K�&��v�(ϔ�=� 8j�6�#����H��b��b�^����P"�����JZ0b�TVM.�J���y~���p+J����g��;{�%R<�.��5�,��GqE����x�]�Г���c�1 S��w��߲����;���`3�ْ��)�.���	��B&���̚� &2���|:_=G�(��|/m�\F>���&����B0ОV�*�y|F�*�컌�?}���&��ښ��<s�L�P�\QO^�LLq)6��	��l��0�Ђ�r����x��y�B mF7,$�uY��#*Z��a�9��LP�"`�äǳ~���gM���y�~�I�&�_D��,���]`����{Pp.�{�M��rr,vx6��xθ&+ v�9�ոq��Ya��������B�+�'��Xu���h��)%�{1���t��jN�fQ2UG�L�'�"�7��OI��ӀA#�������@�s�@6�r?��@�讶>�M<v��s�����D���:N	���j�Yz`ZI�_C�ʋ��>lԁU�vݒ�!��354���y.@9��|�h����w)���D˗~�Y=M�Q���Z���U������k��b1(�8���j�hъ�m}��7�A�`Q���1�-0��Ȑ�K.I�'�Z�,��t(��Ď��������f`��O~����#�0��?b ���3�h x}�_Z!*���\W�S*Z�Î�B�Wp���N`� 9�v�L���n�İ8��x1DPǊh��B9��7�a����]w/��=��=�=�-���P�K�����1���$vK$�h��h"�t�㬷�t��`�R��]8���A���ߟg�tFb7esB�8�9��͝�믲3���z&;  �k�uA0E�[l��ؤ�z�����'m��w�2�]�a�.�������$��t�]u:(� �3�Mhcp	e��j�	Z�b1��[N>�E~o��Q���'��|;���TFY���Ę�4�?s��=�@h��U� S��16���x�@� 8A�������>~�\�VB��K/����cq.���(�@��Y���������_.��_q��)������}�g����TԮh�h@���{���
��BH�,B(����X�d�õ�;Eܐ+�`��n �� �yj�̺�)�@�����Z�\�?���v�x��<i,E�8�c�R�&�׿.gWϣ�:���	�n��~C1�_�{����>����_BpAD��E3�>�3ĉ��XY�Equ��
�~2g��'2��9|�%G�\�	�E��#����%�.=�K��m�����Ȁ6�����	��@�d���b$h��o(T�|��f���]!���\����y�C����O$�5�N %�֚iDO#H�4*�q�k;���KJ� $�;$�B�t�E�@��?!�4=?��#�W>��w��~;����?�1�eq�<�{�w HaW�����ڴi������T���x ��1�(&LH{��>�"�	�h<�	8���L9�98��-�]���s.B.�+D���u`�s�y���E�w4���!�0vM�:�,� ���
�t���	\u���'R4nq�^s����#�3(�?�r��������8�]z]��y���ϐaQ:uW�F4�p�iO�BU�d�}t#��ً6���� ����x��; '~YY~��;�` ��Zj�o�����27    IDAT�(���ƊFԾC7Z_���.+��0"|���߷O۝�u�t�xa ��I18
� @��M��c)�iUF�����uA�����y��ǩg�^�9#�hZ�׿���TPX��x�hh��^�S���c�� ȣ��,V��@����5cG��K ��\�7���6j�Е��5���of�4Y�s�-C�c�wh��E`����i��c��;�B"FmQ��ZN�;~��zVO��f���NЏLJ�$bI�s�.��#�Q )C��<^������b0�/]�2c//ڤ�� �sYGd|:G����~N�aQ��g??��mP�o����P=bm��
t�1�g癑�Y���89'�^U�ro�l����-j�b�0����!�9H��Q�<������˧X"ɉ��O={(͂�����Ř�P
�/솤��h�H�'5@р�����c� ��9@������y�^��c���`���7���� p�\�]Py�߇~�;�@
P�1c�a! �ʽ8��&�馛ҁ� g|�Pa�B�kKIP^Ai�3��#�7d�G���>��)Y$|C6�},hX\�N�+�K���E��}�$^�I�w�﹂��硔!���R��ԑ��d��~��?Ծ]g6�r��]��J��rTSU���s�EC�|�wI:8Ѿ�0"�� �3[�n�'��􀓟�l�d��X(L(�x�`� `�K�-�X�w�q�_�^�8�'&�cnJ�ʕ�i�ܷ�&���~���~;�Y=��mՒϛ��%܏z�(TG��Z/�Ȑ�H�J�ᢿ�cE;�/���>c��!T�ѷX�la=x�Hv�D�\ �C�@Rn�H������q<�����������<�'�P��*<_Q>����Ba1B;�o_\[E�p/����!��RAN�y�� Ա�by�[�v�W_}�89_vI�����F��kz'����sp��D-u��P���k)�qv[D�#�-�z"���ǞH�����s����<~P�w���ڎ�$��9��f��3;�Ocm�!�9�W��u�7I�늑�@��ud�\=ۮ�C��l�d[��~�cF��ɇM��p��l��2�!�xSL	��N��|ݗW�� b��DRɫ�k�Sgٲo��l5�=d%c�1*H�={��\]A�|�5UVE8�F���Ѐ��Ͽ�k����q � ��N:��W=�I4T�%:�b��X4` �5j11ax=�i���L�`��w5vH&���ջ7�
 ��~���.���i��;���ޡEc\Q����y�B������d`�Q]����?��ϋk'vH���(hY���C&���}�;p�0�"�0��XH$L��+�
	@�	H�*�7�<�&����)i�q��.�\V�*e/+�ѣ�҄	�ϓ�?�����~�~k�}ߗtB����� #�ҝaT@@ �E��8��1&�0Bt=���â��d�I��{-�W�V뭻��|���[��Mխ�y[��=�Ou������<���<�͟��T��FƊ6o�b�����X���I2�����=wr"�ց7Y���D,��zW���;�|���^�}_(��yԺ{{�g$Pd(��e�d�+�V�#&)zF<�����k^�j��h��3aae��3�Kֈ��8R鏍��:`���W���F(�`<=�i~29��F��UO�!T�x�N�d�h�\���(|3��Z�r��{�x��6R�K:���z�+(�E���qu���(a��r84�g���\t��y`>_�!��0G6Z�={\�%��G�eB���#�g������B���8�	��^�{�ġ��ݻ����QQ�0i���c��*<'J��SJ
�;4yNA�%��,�Q�<��r���;&B=�p�"dyw| r�J��u���p��5�o �չ��g�^�5�������`==��÷^�͛�{y�L��Ț�綶�V��P�YG�l���W�x��{9���fQ�4{
�~�w��<31/�(>Y��}2���ԟ�w��VB�5�f�:W*�-[�,�xa��T��*���l�����s{)�R���)�q3�f�@,�f������wO��'">���k�m"���m[��*L����X�`�KkU�c�a6/�	�S,�ȨdQ=���D�;^�[�z�N��ju��Y�~��^-Z�����y�sx����6:V�F�bfk׭��+����]ҙM��I�}��#"'\�C?���f2��į����#�F��ɣ�C���@D4��v]�M�0�c����;~��qo�q��C�&@
 ��ً�Z@])E�KX�S�XZ��}Շ�"�uP���(�1��@����n��5{�!͟5��A�4Ԑ�p3���<�G���z���|&a��y۹�^�-�(Y:Y��n��Z��iu�9���q��24Hi�X!����Ü������uA�l,s�k��f�w(a�;�B�e��((���n��;za�cHpO��:���6�4��������mOJ�6��ͥ�^��/���0]3%h�yX�t�z�+��>�D�N�:a<�]ג\���m���U��\�ȑv7á&��DGH��h��Ֆ����p|��Oʢ������n;3�P��\�;��2���}���6:ְF*��TճQ'R�Ǘ�T�̉F�ɘ�zPYߠq�b��`s6������Fи�����/|�A�Z��U>�s�\���ż��������)@���8v�r]���'��7�r�SWh��L����G�#�'a҇
QE�P*�wı�D;()KB�{f�S��¢�^��L�?Z+q�X�X���c�<����>���͋��7_w��_��V�^i54Vr*u�ow�g����~���y���˦)�@?�e��{������b��ɢ��p�ʅ!��S��#���ظ��x�����v�?|�P~��2Q���?�8͙�e�LچG��g����M��K��ƍW��;<�R��U��̳OM�8	:l��z�>�5���w*�_�4k��K읿�v��l�T�a}G{o�J�d�Lڵ���CL[�i�������y\ D� �4
�cҵQ �"I����w���hf����<9筷�;u�ی��H���;`8���q`�[�Ɩ/���|�����7��K^k��y]�	�Xiˊ�bnЖѬ���7�D�G;&��_ו������	�����?����^����-�ͺ����l��:d��r\�[
�h�0��A(.c�x@|�3���'����J
��p��1�x������c	��@���IL�
�M���� ?�O�u�[V��T3���<q�>���5sI%�Z��nW��F/�ݺuvͳ��|�l���dl%��C�8ξ��x~���?��I����eng��f�XC�x�T@ɲc~8�d�ŋ8M{��I{��'m�L��ǜV�g۬X�x�E�����l��%�\����V�Xa�Q�X���i�={�xhh�����dO|��׿��v�O]���~;u�=�k�ϟ�S'�˲�H�ldp���Z笥����c�S�cO��dN���N1�_~4�OZ���:�)�3���#g-�L[&�a==��U��86��&������ݏ-�Ϙ@��1�R��B�㌖̢��������LlEca��b9��7{��; �X�YE-���͋�G��x�?�2�gh�>�`��gº����7���;o������ODٽ�i�7k�����)18�y^����ONe'#9�6 �� �!G�
����B�`)�
�F� ��/��K��M��ۮ�-�iX�D+G�ի7ؚ��Xjxm�l6�a�����yFm���(l�&Nw��F�}"m��G졇�^����J@맪't��uyn�
�U�kTG��w�����J�UR�V-��[�a6^(��c�v����7���$��_��_��u�Ȣf�'.�v�����/6��O|���=�������&����Ä��}���|�b�U��o��/m붫lt����?�ٰ,5AJ劝<~ʆF+6p�lo��o�9@�Z99O�c�������R�?��Y�<f�d�Μ9b�=k��l��Y��?mc�����������㣈*7���`��%rg��s P6'��E3f�J�D��QCu�K��ht<�?�g���#��2��ٖ�[=�h�O�s��#��ޫp�2��١c�����J�'|O��BOhМ�c�	*JH�� @IF���}�"@H�C  ����]@(@��	T��8��|��O*Y��������K�Imݚ�m���,���*�`=_B8�;:]��5�8|Q* ��z�(��o}���X;U�|G()��k��<��J���=k�ʈ5�e�;�g��H,sK2�fǏ��b�aǎ�[��N۾�j��=��<H�G��d�ό�[���������J��{����ۿ�V�n�j�?�h�]���"���b1r �r����<6`��,;|d�6l��)Z%� ڀI��Y3�ACCӜULG��^�÷2^���\�a=={���V#q(�m��� �i�B�2�>�l��e�F�9��h�܌;>8ru�b���,B�(@���d�Q=�lp�)�+ |��;��/��"��=�:B�G����@�a]P3�?4�# �5Ƚ h-B1�.��8�cD9�
e��\�*�rh�q�����p�N���`9p}�'h�XXD�`A�(�(i��fM��B����i��E�D����\�m�Ԯ޵���%��m�u�Zd�_q�Y��J���HeL��'�X�Fl|�>���@1����o���Zd��Ԕ"� _!����c8~h�����l�ڥN=��+ǭ���}
�Z���=쾉ѱ��Z�����wXG�l;yj��z��S��[v�ghx�C�4Қ�+�W?�^/��ݳ���7��y�c�{�4N(5M�mhpغ�{�����c[�&�I�X���h�T=#��DLl68q�ԅ<�ٜ���p���IT=sq�8lgN���[+�[ �筯�k�����sV_ �_�3o��4'8{���Q�)�q%�B�=�*����P. ��������誉
�g� ��C�q�j�ε8O�;�& .JJ�E�9�/�%�&��r�u��T�kI �x�St���C�����uT��5۸����|3��KY�e\�#
�$,a�PO�8��������_*[.�r�/��յҮܴ�2�v��	�C@5��8~|rQ����sv�0A�1��94|�֔2���r�X "ð��������|�6o�`����w����b���B�n�=w�2��v��/7�S�|�
��7R����۩��x����u�݃�C�>��=�6�j����T�f���}��u����^�����6>Vp��d�l���9r�R�Y����bӎ	�gS�� W����H�4�8�S�Ntc�l�yq����D�j'���=�X�FB���Ȓ = ���z���J���X�("�y15-�8z��[�x�d2���_߻�4Τ�,��TV�����k�������Щ�s���y�����M��Rք�		��1���ֈ�wx|�<�YϦ���u�q�[���Tb�����*߅��`_�g:���/Xow�����l��Wx��<�u������k�o���h�r۵�Z��Ky�Wwx{;Ԇ�������D� ������U�ư�H�D��̄�B��88�}��_�(�9sf��C�}L�wTm߾nK����Q+V������jG�#�K�qԺ����En���}�|bhh�7��=&���������w��_����~�N8}�J�b�O��P,ّ��66^���5��ҫܳ���I6�q��MQl/�+���(,���*��'~�^�h��>���O=lgΞ�������:M�H[6�n}GO۷�����,��l���d�ǛX\<�o3� (�T���&i��p	����څ]\"A�^��N�y�ֵqB�-v�K�I�&���h�uX��.V�tr��}	E�85F�v���,l���8��^=ח�YA�r��zg:p��y���m�%�b���'�k���C͈���ވ���uA���n	+Z�Z�(�T��͌U�)�5�~��W[��o�6+�	���x\����#�4�^4���}L�oYc8�J×D>�|'�D�#�����)����b��-����?y̪��[��2/�O&�e�N���K���?d��s���1�����+�_�p��fjI����gQΞ�i�|��l��%�ޖ���_�+�Z�6�_L?�;��Œ�����Ƭ�t����w�㌍I�6&E����LD �S�� ���jT�W+��h�,sm�<qB�9`'Ou��\)xUO�Rx/��}z�>i��,7:�f�r��?tBJR���M���P|����Pb!�zC�V@h;��&�^Cm\�ǉ+�Ix~��f�s��4��u�P#��s����9�/IJ���P�,�����	�PP��-�f�L�j(�4�\;l��K��b��Y�{����3~��8�{����|.e�zɮ�b��ܹ�s`���wȵ�{M���k	[�z�U=�&�}/��I|��>g��/����;��N{�k~ƅyDt1O�����N��O��r�>��}�ha��S	;5pʊ�1�1� �z����q������7~�k](}��G=˻T�|�/��$���w����Ї'���j%�F�[n�����6V�F�h���sV��G!X4s��e��6tn�N��5Kvٛ�����<B�T��E ȓ~Ы�
�:�Y({���I$B�	gQ���*�P��>Lzil�Ν;c�:����Y:8�̒�W��И������k����k�y�8�E�}BS?����� �ٔ5GY��k~*�����E�7�����e�:�����t�/KA>	���-�
QNa$����)ԶC�Z,�@W���JX{du�,�4���JP7[*/U�!�/��kVZ�&�?��7��O9�R�9]Y�;���uG�xT�����Ȗ�x�t�KĹ�X |::���@�D��������O��!��R����������ر�����;2|�
�v�d���7Jʹ��:�y�IK����s{�E�?�V[�d������w����po�
b�^�ɝ�n�����M	���Ă^�|���]�b�ͷbaԆG��#�|����D#2)�eʽ���c��̳k����L2�rl Ջ�!�VzQ�S<p�lZ8B��r�h���6�&����5��g��=K'1�Փ��|QS�0�k��B�H�Y�v�z3��	���"!.�� ���7���4�f�#&ː��<iѡ�>ḇ�G ;-���}�Ly����.��9�C/C�<�eB���Ofq�<�q�Ӹ���BJ(����T�<%��f�n�g�Q�����-�({�Wi|��u5�Q�e"��b�b�sl��^�'s���p$����V-����)��p�b1�Z���C6:%�(#��(!�����[�*6p��>t�N�������6K4�^_��Jf슍[l��U^���@�,�p�M6v�Fc��h�x��TEB\�u�ַ���Fm��.;sf���N�BR�}�Nۺ}�D��K�B���u�?� p|�m���P/��<0�	�ęL($Rǽ�b*��'�}�8���Þ^�j�ly��b��6^�������M ��������{��Es�����oH?4[�=�/� i�D�6-�?3QP:Oc��!@���|�eYH��y�V��]�#��� Y�u��K��*,�&�3�4����v+������m����L����E�H@�X����,YBmh��F��XH�@�.��a����z�T��W�	��I�ܰ�J��[�yKPJ�����w�    IDATa�1�>0p�>��>g�Ҹ+R�Qf�*�K�w%��P���	�ݳ�+�
֖�X__�=���=4���âF�+V���o���̙��B�9��E9tz��gF��n������_�J�WU�Z��Y,�{ӊ��Fn���I;E�0o�Y���p����=���Q�(&���:���P%,TZ�7����T��@�ؖ���5m6ɲ 8@ǿ�~�N��X��=q{:�p���{���=f�c��f�^%��[�bu$$�+�x�>���GH��+c�����;�R���m�N%<D{|��K���t/Γ�PXg���<��s��9�<r�N��J
�yo�y�B���C��g���ZD )�?�~B�*O�
?�'�����][�P��7P��J�D��U��j�T#�?����Ջ�}�e��͖�G�I���w(������1��"�oo���>h�����y�����w� ����16�C�w�hb?��
7V�U��`���J�IgG�G���%'%0%�����xN�9h�o~���v,��%�Qѹ�>3�o�s���{%�D����.�ȭ[7{���~����{z�%HĿ>���.��nB�S-5�&,�E� `A�!J�Ϳ{��y�E�ڏ��T~tޟ�rq@�U���,۾��@�/�z�liZ?&���s��i���R�膜7���K�)�-.nIg9 
9cƀM�u���D?1��Y�*Q�xJ �2��/ R�fb��p"��P�G`c�q<�AT�^c����9��p׆� #ƞg&v���]�~d��X(�D�l5�x�,lz	M6� �g�W�%����[��{�X��D�����pMţ��Y��	���?W���M%
��g,�G�J��%ͼqnX�q$�AIz/]������	O�"ڇz��,А�y^}�&+Ǽ��$v5��'i�5{�]�e�G Q�n^hހ?-�3������w���ٟ?��M���\@��G���}����Ԍ��E����[}	%oԫ�k˻J��7�I%��D}��oG�qw�tTl���,����i��1������+lێ�v�����Ʉ�g�r`ч�t���A�%ٚ$uQ3���L���OD��6��#����[5s����#�m�T��k%��F-���B Q���}}�v���c�굤�]�>���{�.�CI[�j1�� �f �qz!`�v�V$)������a���G13	U�Yuo(�FF%�qŜ�: !ay��l<
�~+͘��l	��������͍�M���4�H ��zTڤ\��}�A�l\(��F.�$�OB��|��'�G�Y�Ō�Z6�.܃�PuX�EX�=nٲş�h
"@�*V$�+�'������Qh��'�źe�B?��Bk�8� Y`<Ϗ��5�j��U�P�0�{'�����&�.��	���Q=���m��N����^�皫7��)ژNd�TnX�m���3w�OC��:��6��j�Q����g����w�����n��V��#ܓcM�?B����߉R�>q�w���Q�Q@j'��")���ɧ��y@�Jd��]��'��L�󟺼CӨi@e�+CVC�c1���dܵxMJ=������I�' P��?�A��{|)S� �0Z�����j���9}�z?g�҈�57sm]v��xTۇ�΀������3/ry�K���j	���Q@���#��	�c��ËEŘQs���%@�	� 4(�����E�y��G�MŘ�`G���G  Ҙ�gxX
�Q����� U�m�|��ا?�ihr4e">���fF � P9���F+$������^]��C  Y�J�`� ̈�WD�.��@E��]��A�I,�Y#�1`iV����r8l��y#f��C�I�����Ġ&e#�;�G�ERm���<�04ɅX-���� ��$�"��*��9����g��zz[6ٰjm̶m��v��̊��FK-a�L���Zn�6l��IZ��Jw�jO�?<;�V�
��}�3 P1o{���C�kpg<QX(�G�&(�ЂcND)�*7�NtR@O�'�1�¨�h��o�u�g���?�#Gd���Z��u՛9_E�4K_-��-@`�g�e��� h��[����W�j�d]�.��������iTk^ҹ��ɉ�nQ3�FT������.3� '�ECcs��Y��� �G?�Q{�k^��-��L�� F�B[D@0/l@�z��Z�	Z�� 	@��Jm ��4rd����c4��kM�b�U���<� �l� �(�v-.B:g>@(����;k�͏@C�N�0@���Z@�G���'
�!T~4��ތ-��&H��d]!����ð`X�|�*���I_c��cҌ	sûBePH��5<7�KDy��"4��v�!�0@h�>܏�X�|Tj�#'���J:������@TϿ��r)�re�vn�ܶo��C����<.���XǬ�6>^�j\ٓ`	�ѕ�j9�ԫ^6����
���}�{<��g�b	a��֩�
�KM	X�5s�5��q�~���w�5�x�}Z,�j���XͿeU�x�B���P (��9�Z1�!'�̿q�����j���aΫQ�%�ܻ�����e��O����Nؓ������rVk�����#66vk��bY�����{�}������VҏLd�l��y�&
�r���D��� � ���1��$�Q�8x�cs"\��;�U?y>,1�h�9�ȓ���Ei�*;V����$n\��h� *-3P�� k �x���������]w�����@�g=�BQ	"@��L�6M�i����]ԑ�5� f���tPj\���E�	���L l�������a�b��bC��@�1N���xƇ���ȉ�����'̎n�W�6О]�$�����L\�?�ߊ����k��+��}�Wk�^j+�\i�:%*���4�N����LD�`&�t�A<V(x�^��GuPذ:��+S�RZ{�#��X(B4��/֏�����G2�5�[v�~Q�\����hIi�k���P�H�7��\
�G��;�1�, ���%��l��ג�M�^AC�ٹ���'�F�>�ԸOؑ�1��MN3��zRҙ���3�p����d��w��0XGP2l*U�d�Uvm ��PѪ��DB�;>|  ;�8�0�k3)���C@��riV�g��M-M�gCp��w�s�� �?��s"��]3��n���~Ο��������D���Y�\��P\��<��E�@��z��"� ��yg���̀���JQG_,,31��5�c�b�7��1�Z���`e�<ļ3�h�X#<��1Y9��J�\ɩ�B���������|�T;�k�F۾�rK����9��z�[��*�6�V�'�A��Z�����#~�<�b���r�|�9ғ���wG�S_|ƞ�fܨ.���|�~��0�K�-�I��!� ��hi����o1N����wF�����#��T!�#�r���Q6���ߘI�\hQ*��h��X
��h���k��7,�6;kǎ����yR�s����3�?�����������F� � ��)9 d��!�D�������C�x @�#xo��c��E�b̠'�ș b +� ;ԉ����� XC�\_�	�q�H�h68���������@��9~�"���t܃ka)��o�[����g�Fk�Fh��:2�� �j��
Nj��x���NW�AG��}�N�O�ϸpm			F���X.�(��@���c2�|x&(N,+Q��������&�d*Z�����q��1���*�^<����F�*6�R[�f�͞���;$29KT�zD�e,��ɦ]������>_�zT���c��T�9U�g�{	נhq�a��K�F0�\Kʢ"�Z�����n���}n�whh�=Sq�tih��Zf��t�Ĥ9M5��|Y ���hB�)'����A��7��ꓨZ�6j��!;s昝8�cV�!�_	�Kz��Ѩ���>4��G������@�KfY; �$�V\04`�JX�M7��9�GÇfPC�8�~E��^6��0�8�c�9�s�����8D���<#߳�)ԇ6�?�v��X�Zͩ�	x�ݰj��p�h�8����K�X��@ A�`=�}�4d=���7�e�@s�R �yg�1��yXT�3�$~���&4 ŸBc��2�9��	�*����!|��4R�C� �emx�z��~48q����2�p✃pVn��k̉O�S���9��Ba7���{���Q+�V����d�ƸY��c�,a��$;q��<���ͷy�;��h�T����;�z�h���P*<4�ֻ��Q�G�:o�@	;�£C�AX���J9l43W�e����{*�,���w�Tܿ��Pp��C�˹����5YD���s4$L~�^���0KT���G�T�eSu��j�&���NB=�����oT�?k��<� ������4PQ5
d18E����� Z'�1c�E�3�aB�) 8R����	x"Դ]4���
d���V���������w<�V�/4�k��b�p=��`m�vۻ��?BI B�{Q����Hy�6c�?�*�8[�l�J��G0����;����F���?A�T���gM3X<�/��cqM���r,ϧh"�Hh�r�ù�0h$�3��
���'��O3��[OOTҹn�y�Z����I��`Z&=�GJ6g�����a)��I���l��g\	#��λ��9ͷS!7:��yY�
"�~������؇�������l���-Xxیl�8�K�ntw�0�q�prB�j�2Y^2��[��8�l<b���h�o�bO?y�x�?qι4�a�nƶ��0���o����ڻl�P����g)�����S	.Z�DHP�Q22��R�o���3����^�"���dI�����cj-M��C�h��+sqmy9�B�D@������~���uq�P*PC�,��D!�y��XD� ����=Ѥ�%ᫌ�Ve�� �;��b�f�xVU��$r=��wFH��ܛkb0g֢��/���a�w#��5˹ⶹ&τ��傠��X��"��S!C���/њ��D�Oe��/Xo�a��?:v֮�z���S�l�0�;�L֪��n�:V�,���WY*M[Ժ��qͭ{�{��G�c��Oi��eh���B!�5�R�C�����R_g�
��֘07��ߕ��
[�y+����U`�s��ܥ}6[�'��,*�k��Z��1���N����A� �w����W-Q/��fuം�,�b%K1��ځ���Ǟ����'}���r����b5s�F�C�$�Yc	8C�����@���Q�ތ!�E�	�7��ax�"M�0И���$ņ|� ж�x�T�.�A̛�6�^f;@Z#<a|j̃���%�Z� �ϵe١y�
�û���������]є��.PK\ޝwCx�[ ��&?m+�֋�5�D�qo�K�1�r@h��:NYuSh��W�.�$j�ga�3P]�{��	�����Ԯ����=�MĚ�y�5� Z�w�*��^�vݼ�&8��+⪞�"9|)��qGj���M�m��+,��z�o�ޒtK���Za�dU/�\�|[�;~=�2���pl�+|��&ٓ<���\�Q�F�	�sQcr��]�5\g���p�$E�_�F�Z���,\����җ��������i��3�,X����Z�)TO&1�b�i*�xX��X��o�y�%幷��l��Bi6�j���h��IFo٪%
WQ�6�`_�elp�`�D�ʕ�,q�˗-�����0�a.tލ�6?!��s -�b��@	`@q��Frt�'����� T�7 e�����+�G<`�#�EH	\4�2�����hL9^��O���1�z�C[���%�U���yމw D�l~�#�����>Pp�D��`�6M�)`������P.��揟 ��Z�̬]�%|%aƅq@�p<�
M�{a����0��<B�s�P�^�R���A�u�_~Q'-@��\<�g�
/�|��D��Mٓ��kE��H��Ymf����)����@�'V�&��HY���\�͊�(@�8>�}F%�P�%ӕ����(2֒
���Pȅ�(�kM��0��f�*��Y����o��o�����ӄzJ"��*�]��f`s�  �]Z�jvȡ�w �4���S�!�P�tp�:F�)a�`���CV),�m�yu�(EͿTI�h�j����3:-_F���.nw9
%д	xW���`C! T�5 ��ln~'�@�)��#��i�r�|4t�08�*<6�~� x.�A~��&����>D�i��W+B-\�7�E�p}�(izh��MJ�뉱A;�U�F�O<�:�j�+34
�B!��/��%�9Z������� 0��DQpO��\0'�cM2����X�#Qb��S~"�p8�ySY
���r�<>#�V Z��h.�d� �~X4��XOO�u�wX�4b�d��U�4<J[��h���g�Ξ��6n�f	�zE���1��eU/��"n�駟}��|ܰڇg�0�����1d����h3�Z�̍���a����1dO�\�l�߳珇�o���+�����ĝ�Q�d^n�^���t%"�́F��l��
ȧ�Ρ���-\2��*ɋ�'��������Z��Z�D լAU�l����g��R#�n�/Yk+�/���HR��q�Ffч�Ei��5#�_��4om
EN��F����Fi�:�ߡ(�#E\pOi[�V�����

-/��d��y|�dѦ���ϵ���s�4QMat����QD��$�Bk��d���T�A��,S���hL�!ϫ,w���3+��Q��9��q_�%��k��Ƶ5��;O�o.�����cL�8�S���s˹�(چu���K�X�:�e��(y��i��;��x�n�V�}��N_�"h�h|3n�}�'#|h4\@Wc+k�C��;�
�C9\�1W=)�%�f�0D`C���A("4�(7~�20�OD{
���Ok���f0����%����:�� *�y4=8LņK L�
56�xa��{�c!���I&jv��S6����esIKԫ��ʣ-:���}灇md���x������5��bT�x்.��ؠŰ��=���yKi�l,�IZNH�79w%�Gi�y���X���ϩ�' �Uǵ��#%ABBڜ�Eq�l��tM"kI� DJ�~���7O���Z���9�g���y<oi��IWֹ�+t�A�r@r��Y'��X1ךC�'Q������ʟZ�Mt��:]�l&a�ڸ��v��tnT"���m�7��-�=�����:w�9��Yq�lt�i�Ko��;~�-���7�4AI���� 1���"k�c�
&V"V��=QG�&(�'(B�>�Kx%`*v�e�o��3	�+76��8��Xf��&4�"M�c�˄�z��8��H��{Q"'ؼd�NI�$��w�#6<|��U4\VQ�p����a����~�
cKg��J8��{��b���N�"�i�r�3C8��j৸T��j�(|�kl�fB�I�� �����p=6����k���mq���G�&��E �@��8_Z��$��>�X��:N�������B@E��}��r_{�IK0!Ƞĸ�4x����(���}=C(�$����$���CKq* �{Pҹ^����aˤ���!�r�z۹�*K6"��)�\�P��l��e�e�.+V�6,��{�&���F�-�?���>h���֬��N�=e������C �J�#c�>Ƿ���^�Z��QLQ4�����/�����>��>�B�>7���v㍯�&<I)�aw>���޼����_h[�l��wy��5�IDy`�� e*����A��c( �*ԓ�t�3v��a;}����/    IDATU�c���(���\~����?e�Σ�Б)�&��K�{}.V��(i���%8F��%zi�i��t!�0�3��K�4���e���I[�!(�u�*�%���s�kB�c�f,����OBCt����9*�gܸ�'�{*��"ǤK��K )�M�U�c��)�� ��Ѹs=	EJ5BY`�B~ 	E�I��&�?/ ������D�oV�M�а7Z&E�fT\.��]�,�d�lպKl���f��&b��'
�������OM�d(�K��d,�ې�Cd��Y��ɾｷ[[[��mY/�|��q{�{߷����o`Ū��;���a�t���Pw�����o�/h�/�����S��K�w���p�l�D�������Ν0h��� �U��⥫�k^i��Q�)�q�L��~E���ӂ���Q{<9�ظ�>��V��&�����f�L�Ϟ�Ç��b��k�C�g+9v���S���;ԓI^5����o^��¢;H��Zn��n|��@Z&?�'p�w�G�d�:�j����- ����F`���l��d�9N���Ӑ��=��7�D\O�o��hQ$�^xvmx	{i�>F��k~�ֈ�AE�	h$T[�~j���� ��.�z&���%�{zڧT�m[/��;6y���r�b�d�.{�.�5w�e3m��ztl�#���z�j5��l�C���Oz�s�LFY�a���5�ߎ+B]�Xw�2BUٕ+�Y�R�Ju�~���l���V��-�H�u��>�.�|�m�~��)A�L�����O#k�g �V��=����F�x	�¼��֭o��
�C66|�N���޽6Vt�ϻ��='�v����+I�;o����q��r�<�f$�[���Ą��O#
ca�
 Ĉ��*�� �Q:e����ؑ笧�+���\&c�|�uw������6�sA& ��F�L�A�����H��}fuF��DE���V�(c#�(cE�	ILQ��W�6E8'@U�i��[�7	ݛ���*��n���s ��Һe��9
r�[�{Y���k&�ώӏ1����y�$넱iV�uC��z���Um�����q�'r���m���M��b�F�/]mk.�ʒ�v+V�^�'�J{/���X�)K�纎2��Iu|�Ɍ;g�KE��z�����{���g���;�����ș�G��{�<�φG�hR��
R���F+���]��M��	+���hѾ�կ{QH��~�VY�/gny��J:k�9O�_�h���i��?��-Y:���<u��e4����ㅪ=�o��������.�p���夝J��-��c��6�8T�>$<v-7w#m�T�����Hة�����,����$g�ݪ��&x~a7�FKs�����'~��S*VX��ЎD��8�\T�����U�� watl������Bg��q�lB2Y	uĤ�C$���$�!JK�ҶC��{`��k���;D�8%�qo���x��Y�8p��O�h�ٯL�� �N�	��O���d.�?Ɓ�2j"ϼ�S�p�a��/O�U�|�R�Nh�����?��zy��;7Z>mV$,�Ҷ᲍�pɥ��tZ�R��D�9���9���s�t2�@Nm'������=���y�X(z	�H��LrY���?�����z�F�O��O���Ҹ;���Kh����6pf�j������b��^����}��H�iB�_�I�t�\�of�aK/�z%��R���'v�+��$M�{�[�i����cG��V����C�e�.O>Bsd�PGF&�f�_��8[4?�<�Wm�B��>��U+	�fR�˖���C���I�T�L۱���f./,��O���0�����O ��fc�H�v-���������C����p�#:I �Xq��0����>e�)����x^�&d]s�� �ʼV�l�"2b���z>6*N8������%�9aA"�W6̝�"	LDl��u��I��Z��#��x���A[�j�+!X'T�Ĺ��#������Ci�G4�L�LK����C3�-�.�]�l�|�zѬZ��K����vX:�?8��Rz��>$|�͒Q ��4��mDh�];=�\�H�#Ɏ5E2�Ah������.��w����_�����C����s>�POc����{�::�ّ��v�ƭ�����^��pw����:u©ח5�Iv�-{��l�X�W<Bf�ʕ�[��[�j��ࡽ��w��j�g�8��&�D=i�#E;q���>=G���;<}���Ԣ�
�(��d����pO��� A{�yal-�z��&��l�'{��@��=s܋Y	Eu�W�OU����1���S�S��r˥���Xp���h9�È�j6象<���pp��.�(�' ��LZ���'��0��"��|
��tE�.��JHK�秢v�`��D5���`�����/x6�9��<6w��-A��P�L��\_���A����~e"�MO$��:�*�#~r�>ƃ���ь�������j�yrc\Փ6�1��s	��kǕv�5��j��UzZ����m��E���T�?�ō[-f#'>%! tJ�D4e5Ŝ��F�&un#󙪬R�Kb�c��.�?5��Wl��ˬ���{�.���3Y2���S,�j��g�-����;u��M�pj���!�
�̥}��d�F�%[�z�}���3�(��O����W_����w�5��d"c�C;v�U*i�>�?Z��o��J��|���J3FC����/�뿣ɲ��rQw��k�^.���3���g���&�!��N�[w�@Tҹ���Z�Z�}�����Lg"39t���+����dI�h�	GlowNt��elr�)�S� L�LS�js��M��B�@��	L������|<;N;@\8s��]Ř�;����u�������Z|8��9�g���|hͷB?�t��Vu=5�x'��8`��6

�$�D� "N���-���pή��*۱s���-���IZ��0Kϲ��V���Kl����9&��F"�0S	s�k4�.ؙk����	س~Y��]��Z�R@�,��s���y���X.��cǎ����HФ�ܡ�G����ђ}��`���V��Mh���
��8c�8NG��,��d�:�������u��/~���~��2;ܽ��Q�=��C�#v��	�V3�w|Զn��5 �^�E#'��@���h������{7'�ςB�g���� ��M�$��lh�%%�g^��z$��������X�Ƒ�nk��ˋ����
� J}�G�$�86�\��X8/��:G�XDu�0�Rܚ���<�� :�%���c<�7?
J�P��&��͇&L������A�����q��=T���/D8V��!U'+�9���ޔ��܇�D$�p9�~Rl�|#����(�-�$�Ph���z��Λ�q�;
��}�9��7�у��
�]�H��
��$jhZڇ�==n��#v��+lێ+�Ny�l5/�l�U�d���]`۶�Z�J�9�T�lg�J���|��]wOXz�e�4��p��)�֨ΊR��l�)|Sp�(}}{��o�/��ʵ.zz��Z�!�����Xɞ}%`����Y���5��5�N��v������T�`����f.�3|�!��-g����ys�X�������֯_i�cC6<�OF�����;f����l�n~ÿuPB�S
�pO@�C��P,V��͌_Gi�L.jD.���E��M�qPKT���'�H�~k�S�d�3}]�E�I�[O7���9�����Y��<_��W-�kw�zʣi�_�-Y��n�G&Q|7��MC���p���h'~2n}��@��]�M!�F�6 ,�	�Bgr�+�J4WsC.�6s#*Fs�d(9�$�(d��z:j���J��C�b�K����8yk���߻��.�8ʹ�����.�}>@��%��`�'�7�}��1��_�mۖKm�+<�'A�;B=3yk��l�P�9�ث^�+)~����~b�� ��wMT��C2( ��)�>�$��K��`�}�"a�(
��=��7��3ms�̲��38m��y���#�ldt��O���ڛ�g^{�7�yv�>/��E,+�e�o�
�U�L��J���M7��n���f��k�#�$h�,K�?[�9WΟ�S�m���������S>�Z`�q�UE8A�
y9���'��aѱ8�j[��U+E�7��P�8bV/Fez)��ى���s�mx��>�锭\�ܖ-_9�����_�� ��r�~�~�ߏŷ|�R���W��Lԯ��"�І� �z~�w~�#��}����&���f�`m�	�6�h� +?Q>h�,|��\���&��1/8e��XlR����1�jnx6Υ.��k hb|$4$,ࢱ��D��I��d��q�a����PH�Ї�}�O�����w�r5xq+%Vx?�k��1�k�߈�Q<7�w�>����V�h�t�๰4�o���PP�;���M�>�a�C�#Ը?����Z
��x�� ʵ'�L�v���lTҙz�����_��.�b�7=�륚�sY+��R���ZmX�FV��Q �RX8��t
�>N�5���N�@7���ظ+����cL3醝���s'm��Y�JH������1��=f#�{ǯ���`����}��}Oa�Lc�-X��/���|�L��9u'�F�J�Zd��Kv���/���6����s��SO��J�FTK"E�� �,�]���;V�dTT���Z�1�p���lf���" �=�7��b8�y�RqI�L1���U\@5j�*{�?B�\%3��,w����96^"d�b��|��X��
�޴���}b�R�ģ~�	���t�Zf��t����h��i�X�� �u����ȣ�� (m@J��!c��� 8����В�3�X���&��y�&>;Pо8_t�TH�iL��9<#�}�K_�,����0f�a9`��� �`��B@vZ.�l��=�Ԧ�	�L	`ʈ`Ma8��J�v��: J�φ�2�D�!�yg������.X���˚�3�Y�Șk��z�|x�3���5��FR��Nh#��yg�@�E��q
�yE��T�a�^��d����d�$�����V�|J2ac�g-�M[��4��z"��(K��-�J�*�/{�$<q��dv��T����xG�Sy:�8S�R�(41�˹0d�iPT��[W{�|�z���(�uKeӖMe�\%���i۸y��[{�c4�_�K�7���Tz��;s�����}ph�]2��xs��HZ%n�<>:�����z{���R������������������a�V��׾�&K��zł����U'���bƹ�4���'N�t�s�� :6��<�q�8M��mu�?q܎�v�?�%��:��L��600l�t���B�
��X��J��:c+�'��;�t$!pQ�����fuL4� \٬$_1ԭ��"d�D��%2�1@�ط�9S(>*��;0�h4"���k<_���ƕ1Ҹ�a��3��x�d��0[��b�)�E�C��*j&`I�c�I`�d/4Hx`@��[h�p�1T�7���������h��8����XB����.�hu�s�?����ܯ",5y8�G��p-|Mh�{� `�����u m�lƁ�&8l� jd4Z�\�5�����>��D�0F��%P憹b-  ����IP������V}��k�9s;�R������V'E��t�=�6o�f�k�v�Xs)��	�60?�G>�)�(�x�b����%HY袁yO�x�޵Ò����{�g�'�ǎۙsg<�c��Ev٥���l��n��Dʾ�������}��E=^�IF`:����|AΛ=+���|s]w�5�������>�4�����uk-QoX�3~�644�?4�o��f��h�y�r�ı���h"^����ب��	��ھ瞴3T�L�,��Y�R�Q���t��C'�������^��s�-[���5#��Bm������,b�n"�`D''�l��e3�b����Ip��Izcs#h ����3O=�&36r��9��	P#�µxv	�x������2��46-V
�E�/Z4��D�V�GQ�G�]�[�/�����y��Ra�� �x���&ƀ����# T�z�k@��X^��>�4��LX_<'�������1h����'?� @#��C�@� �8�Ʉv��������Zg�c�Ag�8?� gm�[�_��`�P��(@�o|��'�SZE�fj����P��>�4���2|�N�@��֟���x��/Xb7��j#i��:���eg|[<t&���½h�B�19�qd3��#ㄦ��\'�(w�wݾu��!��(<pp�����  W�Zg�]�622f�]�큇h��W~�H�L�3��۪�{�0�h"Ж	�$������WU�^6��ѱ1���v���kAl��,Jܒ��F�q|��؀���������`)@�xDJKͿb��>j���d��5~*�B��l��=���=aC�t����YV����ޭ48����Dҙ��>���'lvx�
`ġ���O�k_�:s���׿�5��W^���F������.n���ccqc(�l,
�b�� ���>�FT�]���VZ/�B�)�/�e�h]���Q��SҘ�8t?~z</c�,nE��,<?�����C <�ll| Dƒ{2�h��?����k ё�aJ��̀P�3�!<?���&c�u��6�;� J����F9��`y�����8Xdj􂠅��:P�Xm����{� ?]�L������"�Zh���t_j_U��^����Y&I^J�Ն%3Y�d�FƊ6{�|���<0�.x(:XfШ�?�K��p_�v�ڭ�[@�yG��S�>���������׽��8j���A��j7�(a�"s�\�H��������w��Q$*�MHw�O��(�\🦍#`Ƅ���h���h�L�Wl�-���Ƥ�_D�@E� �*�M���j`�"�p�hЄ=)a���Xm~�v��ΗҎqJڧbGz���'���4�Q�!w�&��p�){��O��%�;�Z��V�p�GV�T�?�@ |�cI{g��n�J���=������G�,Z;|�-������Zԓ�?1�)��q��c P�u@T%m�t�����"���wm8�ņ��A�0�r��@��.aYO�<��q�D�@�BQ>ʁ�'�O�K�s \z�AK���|���s�m���#��oG��G�=���Z�ǃ����f�l�a��5�X�PwX�� �h���g�0( �\���u�څ�йV�� �=��P�Ϛ�jb,v��I�'��xX>Z��͍����f��;��{�r٤U��z�z۱k�%�eW�Ru =m�ɜG�\�y�ժIKeڼZ�C����G���}��_�E��G>2��b|�g,w���*ժ��,T栽c�]q�+�b^�v��x��G�`V�Ç{���r
S��N�
��gl��t�>��,2@�	Ne��F�*e�1Z8v���j�}#��бǩK��Y���9j "�z�$XR��?Q�BB%�[q����lxp�FGO���i�}(E��s�Ġ}�[߷ᡒ�ۢ"j ��UK]�F�i��cݐ�Ef#-���/~8e�Xo_�or4B4M VM�т�� 6���骫� �	�-	m<�m��;(��h�|�8��8��^e���f���]������N�7�6�W%P��`g�a�+GA�E�T\�(#9|�;�׀��g�~�%�)*��b�������}��|:
c	��Ppli<*�O
��u�������r����sq_���ZQ�@�J���zrT+(��eMqM��g�r��8^TG���O��Zͽ~j>� ��)3|[��v�����
۱sS��e\#�?a]]�mΜ%��5�/Yn�z����?�L�ӗ+��>�G���E@~�w����)J C�bY����)6R��1    IDAT�gfnU�;��f�%B�#b�����K/qg��X��A7��SKD��{ǭWy&/:���?s���;��/Ȓ����'���ظ�e�У�^�s/��p
K)Ւ4���b6�������ܤ~�m��T��tf!Q�`J�oDF_[&�)�=m�O1_'���#>n?�d��H[�T�K.Ygk�E叧4�X�{ m���F�n�3.�0��~�X�[Ex�A�Y�߷ϳzh9,l�� F@���G����E�1D}��|������A�I!P,a�Q	�ph> j�N,5Ȁ�����>����.�ڝ|xfq���tM����a�����W�ʩ-��+?s� exVh�2��zr����"����uO�����&|P�z��»�""�k=N����h}��� <�ƃ}��%�����; ��<�s4��/^Ѥ���h���)+m˖vݵ���;!��x�ƆKw��+�^��;��A���{�tųR܍����r�{��`3� (���r�χ��KOF9@h��e�q~'�8B���3I�����"��C��7�֚d�f.��t�Ʋ4�x�ġ�?��g�b�4C���D9hCiSPd�@5@6/+��s�펅%z�Ο�:U��H#JZ:��.^�D���{��g��+Ke�Xo�I{��ld���Od@�l�b��}����X;:�"!��c����B��[�0�<!nJ�
5}Ox�{Ȇ�����������T�V�-����t�{7PÇ�P����59_�V������\�MO�)`h*��s��
 6�j&XQE����_�U6�m��6��::8Xq,����/��}�����d��<q�>��(×���d�9j�� )�IYq�d�/��V��l�R�uJ_e����q�6I�����]�=Y3�j$0���Q9q4�tsnTc���3��?O��1g�k�{p��-{n�����`���y�����y�'6������U(  ������
����� ��V��  	N��h��4�G�U[.e4j:v�:�Uk�3���}���>j#cD-D%�q��\N8be��Sq����.���=����*m�����݉R�g����N��V�2^i���xL N�WtL�M�gCX�D_ hy �)�ĵp�J���j� /Z8<59��f���¢t\_�S?��'���%�-����Z 2
��jG7�waX_3�s���]iU
�ў1�
��ϛ����q�Į�f�%K%jV+���ˮ���7Z�Ay��[���(�V�|�#8{�O�O�uwT�5��=���DAE&)���Y?-�gk#0�YPJG���r|�N���Kj���{�ǳ��<ON硝�x ��O@��������ln�"�Z/덨�U˦y��uz�z�z/�l�͝�ǎ���<�Hk��zfŲ�����2�3n�ieq�}�t ��C/8��Ǌ��Xw�j���CZd�I���55�ԊQ��6���e��qܪ�W�O4x��AX�i�xm��F���vQ/� @j
�ć�Q�ZΓ6�spO��p�S��X�PS�<�P�#P>|G�?�1 b�1;��$!p��_�z�mW����N^���-���s�c�ev�u[�V-X�Q�J�jK���U�l����6^�z���N�d���8%ӨW�?������#���M�ɨ��9�J� �&-�����?�9�?���5��[&�:U&B0���⣨Y�1��)Z�`�B ��p���BH��o� ַ`c#gll쌝�?aC�#�6�JS5Ǝ�L�?U>�5����eQ�H�M��3�ȑXuax6��lt>ߩ&>�X��H�
Xm(ƀ(�ƈ�_Xn��f;P��G2!�d��A�uE����	��P�#A��ɠ%f��!�SA7q圏��kh�xo板au����;B��@Ӈ7��z��Kr�	Łkആ�x1�J?�B����ի�z�o������`==�Q���]��J۹�
�L:a�j�R�v[��޽Q�\M�jn@����I�әk8�H�'��"��d�b��6�<Z&�|�=�|�%��.�{wk�֙��/!p���:�VB<�ł���'��3)� 4�?_�����R? ��؉���@�Ɔ���G%_R�6;�7`߾��Z�����4�˗��ZםJ��Z �@,*%0�|h�Ӂ/K5R�m�iu>����ب	�H�Nw�l��ę�6���G�����P���gW�>�V�6�=t�J���S��r�</s�ld���Y x�Y�sg<%��.�v�۸/V � �Q��t��O"�_ Z����45p��9y��7�|��X#�s�e�u˥V��{�b�����*ik��U=���*��oo��J������׵�����r�7�H)�\���i�_�������6p���!�4���F�hB#�nr�'�جh�a�n����q��4K�-�"Sr��������8j�Ҙe3˥��]�;�w̱#����S�BUh�+����ΪY��C3BP >��je��8N�p I9V�ĮPs
AZ!��C�C�V��i��DA���y���ID*a ���E�*�F��(,������~;��k����s���������_/�!�}Ё!�F�^����?����ʃ�k�`~�����\��������f��A۵�J���͖JT�FD1�n�u��x�f͚g�]�j-�-��p��{�R�'��:�%I����)�p�7��LE�|&���[S>��(��S8|��帝��A�C�h�>��Xlbi~�z�@��V��^{Ķ��mլK�g��Jy������j%��LZ[{��}��~�)�4)V�I�'��B�Oʣ�������y~�a�TdC�Zn�y*�G �	7�+Q�l�i$����xEIp�q�M�Lo�O<t�4q<����&��$_ׄz�2�Г%#�E� �*�;��է`)�@�yF`p}��*Ĕ��0���r��B	��@l���.8|U�'������s4pﵜ[ӣ��o߶��ch�J8��Ixe�f�����M�Z�Y"�v�8U]��'�G=�{/�]ȘJ�z��T�P$T@��iGd����i�}��}�����00��(�	���&�\0	/c�jz�5e9��kG��d�h��h:m��wl�*�#F��$��g�R6{����B��J�l6��˩'ν0�������J�*��c�㈆�����w�C�1/p��7p� z�(+��8���y*#	���&�Fq�Y(Jl��⚊D�#Y��r$��g�A&6�|���0�H���r�9��W9�0�D������h��=�x��(r-j���h�{?�E�,���Y���,�oV+Y�2�Y�:,��rw��/V�\JX���L�ݪ��er9+�"���~~0j����z�S����d�˼`�[����jg4�O�O&_��f����K��f�vv���8<<��ZWW�'Zș'`�����W�� /i��AܫUy?-{��{�"�4j$$%��5��.�'��L�#3e�j�8Y%���w`���ݿO����
��^@4�v���4v� E,)��r%1�/JbGCb���K���`��wfgg��������~��eؙ!�/��s]{�Ιs��y��������4�dh:wx��܇���K��s��P����9�D���}�)��H֬\�bi�RP�UK��̯Y5V���M-�m��,;P�Z,i�x�^ۇ�<�\32���*cS�L���W��/t"4`��ɣ:�.0���
:=��9��������Z���}F��?�����2|�s %-%_{{���'�oނ��h�bkjn�b�`'QX�����>셖��Z��mJ#`�ʙ��D��~�]1�p�Q����G���?������Xv���ɘ�ke��b:�����%;|�۲y4#:=Ǽ�ϼ���/����E�PE�g}�$�h<<H A�?yF�=z���q��#f���>5/�]�	�36y�Xˤ(�V��Y�,f�B��?�.��f�B3���h���O����G��?~ꖺ�&�!�o~�o��@���������&3]rT���j����cC����Δ�o�׎>f�==~��Jf7π�?|.�?yʤ�x�?=t���f.$q�������
d�-[�£+H�bQ�z�=�ڹB*�&�v��qkۿ����7<2m=��"�H�!,��pp�*� �?8OTI�7}�fC^��}ʶkףv�s���ojL8�{נXʒ�&۹����v;q�ߒ�Fw`�@�3;������q��#N'���E��f�Q:�
N�@[I8�
���
�g���
�7=Ŀ�ᛈ�l����v�RkH�;|I��KY�T�ɓf؆�[��D�56��8�b��e�X���S��)E��:F�i��!AHTAx.o)�''>�/k�3?c�L��!������d>�
�B�f��zh�}��o�B`�ވ����G+�f͂������R{�e/{��$9�6V�y�R�d���8���9,�xZ���X��O</U��%�0d�ǆ�4.��i�z���ݹ���>dU��J��V��KZ:�b:���������[��٩�ٳ��O{J	�����U�S��M�ld���#����B��X�N��u��7aȹ�>Gg�4���RD���5�ym3���c�u�e&��S}�y�_d�
��)��i�4y��=4��t`8�u���J,@��<���=���(�¿r��J����`-#jzz�F���������>�;u*�&�yt�����G+�K:"Mq�^��^��ߴ�&
d嬘�z�*Ijjij�~!�7�_o�c�Y�q�;R�i��z7����&Fm_lJ�aB�9��C� 0�}�$�{��>��������:h��)��oHc�P,Y:�jm{=%ɋ����-��>8|�?R�/B���Ĵ��8�t�OC�ۢQ;Q�����}��Ϲa�7��S��$��F��ty���+�T�ui��5�wcV,e��u�57�؊U�,f��Oo(�G�m�稱��~��?��p�(@�ƴ'e����Om��Paޣ���D}g���%���T �����jժ-\�ȦO�i�M�J7xe�}m쓟�����Y�q�uV�>[�m�����Z�
�8aV������������y;�^{��?��J�R�FsC�]�b��^w����$�P7 T�=��s#D�j�rS㇘a�ˡ����|caRu2Z�-/|ڱJѱ���tٱcv�H��v����Z,D, ��=�e��+���T���s��
#�w`c)5D/����y�_�.~_a�}E��2Z��#�����xN��������>/�y�J+��M'�&mN-=�V��d�w�
eknj�dH�:d�!�1V���GA��د��Z��l��	����G��?�yg�r-��|[6��B~����:w����}���㌍�0�^��ټ�����Ŋ��=�ȣv��
�CB��.�?i��t�m�������xOo�ug��B�Rɸ���/�+.����Az觶{ד�L%,�ΈU���ռ�ґ�ݶh�{�^7�%J�I��ۭ�B곐�T�;������g�d|l��r�$��/@����U*v��k߷ݣH�u���{��6�CcOz�r���>Ϥ��(6>�����ƣ�Ȅ	�|N��Tq���F>/:8j	����C���b�97�g��v��\�_m�<`kW�g7���d�j�l��O�j�nt��n2��3C"��D@!��By�������
�l�r[�q��� ��@�6
UpaB&|���|�j�(��jκ�qő���sߙ�6;r䘭]���ѓ���n��K_��=��9�i_^�u���oV	�ل���}�-[z��
v�}w۬����T�:�a�R�q�%�iJ��;U�W��k��/>��� �$qू#� :,�Ph����8�}Ī)K�O5k�N򪞅b�'�466[[�A�����=A��@�ޣ�����o�z��$y1.�K'�W��;�E4u��te��2�yM�bcC�\�9{�e����h��%���=6X�9�ۜ�X��6oZm�*��kV+Vm��%6k�*+V�V.��Z����ӂ�G�� ���G�b�[�ƌku*�� �3�u!���T�_�?e?8�rΎ����`:;;,I+�xh��Y=|����g-�/����fϙg�x���;�5(���>g��m��zz�����[�O�<���G�q���������9z��zp����w[��#�y$kK��R��Z��7�<�4C�P��B��ҡ�����]��<l$6E�p��覧�l�z��b�͚�v�H������}��W,a�;�����S{��X���i��U��x�Ё�+_��]r�e~ppӺ񢋶�&�l���/�9�a��&�.=CY�r����-�0�c�S���+���˸�r.��Z~*�B�V�a-���/�t4F[y
��U����������*�Aa���>����4�Ud-���I�ɀ��i�pMeG�*(�.c>�x����E!ߌ�M~�9�����-ާ�E)K����՞Pb��
���p�O/���f�b۲e�U�}�L&,^1�>k��Y��*��b���:=s= ��Y苡�B�����2&���y[�]�W�������N$��O'?U��_�����'��&Nh�	�Z��=���Y�6Y6W��;;�RK�ɓ��v����rNM�O�3�x�VXt�G��,�}F�PՒE�?w�]�u���>�����]v�k=R���C����fX2��S������i��q�V������R�'�:��fs���OO������'�����r Y�7kH&,��Y�������;݁��4���uڽ�?d�\���Й����z���ꆍJF�a���osС�O6��m��^@G/V�OMz� ��9P��<(<T�) ��-0侀���h"m|���(�34�@ 
K5v�q+��ļh��V�ͅP�ƨ�`	�A�Q�ƭ�b͇~�<J H��Ґ?�s0^�c� ��:�� ��
�1N֌9�s\�N��t�%��4]���ֽ���u��C���D��*�%�,0"�O�흼���7sQ'���%��X��+ϳ͛WY��o���e?a��]��;y�����/��͵r������~��)g��⋼�<?
g�fCP��৒��g����}������ov�sm⤱�c�ϭR����l�v�9`k�����\���B�x�����=%S=j���Y���>���[���v��U��@�}�߰�/�`�X�����p���Y;r�U*��v�5L96:�ޮ�_�MMo>� @�����}׭��8��u UR*��%gt��J�����}����SGͪ��h0��X۳'8|��g.�����!�s�h(��h'����c��<c�={���;<�B~�֕$�ѺR�BQmz(�I��(xHs�ʀ��F#�� �� �!��Um 	"��Lt�+�O���{�nc0	��J{H *������q�"� �p��B�u��2~=�,�cM�^�F[����?�HT�%��c�\SV��������e�N8��p���u����+��P�!��6�X�p����o�8�4i>��x�ɚ�L�ISfz#u2���N�C��g7̅yt������-1�G��G�O�'���g�+�K�X��ڳ�q{��o�ʕ�l��V۽g��$��Rͪ��=���4���'\���
�U�yٮ={�'����G2Z��Po1X�{�����?�^�ɪ��>�����L}���'��[.�#]�A�G��ѡ��,"�J
�PP��8|��l43q�j���<b�o�`:~f�OX�T�LC4�x���i��費�}����&�T 5�3O�����P�\�4s���6���^�!�P9\�k�6����0c#���)o,�|G7�6�4h��@F�q�'j�*�,��QPR䖛�ޗ9lE*�vQ�d���
n����S��PU�b�    IDAT ƳH;}$@�΅��h.���q�
�|J�������o�;���X��yn�8lֆ=�ƪ����T9������2�%$������{�{G�uGC�����z�۴q��q$��|�X"�%�s��G�<�"�z�,I"g-D��kh��]]��=�Wu@��8;�[@YC�!H�f��e��٥p=����<��~������ĉ���m��KE�R��lޏ��w���2������A�����mFֽ��9��w�?�GkK����&O��η�n�S��Nul��D���T�:1`��d��/��^�җ:xP����o���'u����$�:����k�7��m�ڑ��<h����&;S��//��'�#��,�Y*�|$�D�G�9��I^ݧr�L�X�Z���9�3�|��_���_��_ٛ��&[�|���b��Ǒ��9��	~e/+�M�T4ę�( �
�J���h��p@�4K��z��4z(��c�gS�(W/*Jܺ@?��.!%zHt��*����BF 
�3o�>�����{�y�% ��2�����.�2�c�ŵ٫p�\KN%D͝Nn,��O ���Y@Q?E�ϴF<�z\h=�N�g��O�{�f�qo�N��WY<^�r)��=e�c��/k�c&��/~��*���O�;�D�P�+����i*���Y"�A��F�'��g��|,<�����8��}�~t�]6}�8ki�XGg�ˑ�PW(�~�C��ȱS���o/x���+�\j'Or���/|�N��v��|�V�YL�����&�P�xʶn��^|٥��sº�:�����8y�ʕ�%q+{S���c);~�{���&�_��5N�pҹ��ˁ���~���XhWl2{��A�_u���=Z��r6ƦM�BM��7<C$y��8j�	�$k�JIgw8�c�δ؎���;��;g�t�K��S�'1�#w�Ղ�O�UW]��� @���w���C{��"��j���E]��1����-��0�QJCܺ�n6���Ґ��^`!MYZ��q�9�w�;E��q�v���ʚ�`":F<u��$Ǯ��k���`�~Y%|�W�bQ;r���FAC�X��`3$��0c�,9��ή]�|��@�{I(���[ȱ�Ϩ7��G�,YC�LtMt]~
�7/��:�|:"��×f.O�}��_��Ų���CSC�J�|�y��Y������V/�\)ǩ�˜�7n�;~�~����zg�@߲�?�я:��<+����}h��h�����u���u�ú���l�+������	;��k:�X_o�^�����f�2v���; ��*hρ�(�݈v�I3���׿�Z�Ҿ:�ڮ�OZo�)KRʙ�o޹'i�J�j��󗬶+��!��D�s�{�8�}� ő�/��O��/��n��&w&�Y�!g�{��(�U����W�R�Y:�D2f�b�R�F+Wv�D���5wX[,f��p`f>��>h+��7�!lj����r�']�|�;��!��gy@���A�C[=r9(ꔅ	ˋM�5ѐY>��h�(�A���|>�;c D!�!�9�X�+g��|0���5U���" Y'����Su��S*Ғ�{��)J�uHj͹�"���s-�s͘��s4K5|ѳȂ���]�z���&\�R"��s��PEX���H�p]�IT����v(9o͙�>��Ng�)A��D��(E!���8�-K��J`�4E��.�8�O���~)�L��榘�C�D�O���|�i��U��(�@Ѵ�eZ\�O{�>��+���A�_��Я���(+KJ�g���I<���jլ���i���Y6G���G�Bɚ[-�/{��qc'��������;��A��3ٔf6jU�xh�H]Up��ۅm�9�j�����O~�#;��a�b�-�;ޖ/_a��l�Y�X_߀o��[�V�?8|�q�I����?���]w���x<l��f�\(���G�;�k���Y���T�fU��d��h?GtO�,��д"�$V%���U=�|F�d<�&Z?4����N>�ʳ~�S��tTϏ��\2� �Ќ �K@�"��B`��}��ph�'�y8�&�$� ,�.-|$��0�9��LBp��"hq���c�)��cf��G)cz��\�3�G �<��3���Ҁ&���V}���K^����p/��K#`"K.v�ʘ��ʕ+]��pD������sM9b�����d���5t$��{�;�\��9���5`mn|�y�����x������e�l�B���`�����݊�8|�	��˖0�Eђ���b�X�
Ţ+J�Z�&O�i˖��J~?�%�I���Wc#M[ʮ����u@�'�����W5n	tYV�=B��[�E��ﲥK���wn�n��~;~�;�)�BH�̙sl�ʵ^h2F��Z��o_��/��t��s��!0Z=6�Lu~�u��i�F����Bo�́�����k�X�&L�ds��3/�M$~,�& ��X���ȍh�lG�I�r/�o��o�q*�tp�}v=�����I�Y�R�)B��ԩ�=��V��_f��˂�l��V.#��8��WB	�fӽ�5�sڈ��9�����;�0ǯ�إ_��W�Y8�D(���@���>g�|�+�
 ӵk�:� ��CMH�A�O^UNB�+�xrσ%G����kD�5k�g��0gPvX)j�~�m�����6w��hx$��A�%�C�@C� \\��B����"��p=���q}� ��? ��e O(@+ׄ˿���z���گ9@�RB��<@�#��Bp���[n���F�+���A(�,W, ��A,� ��]����g��,��3��E���������}rMX#� ���`��=4[��ૈ�D�)�oO�2|G���[8o�-]�Ъ%:��=I���R�f3gͷ+.�;W�����)錒�X����=uʱ��y�E���u���/�gy�����\�
�8C	y�k_m��u��\(�Ѯ�v�P�𠱡�.\lc�O򂊍MM��?�/�v�ϕ�h�轢��^�4����$+��~P.��W��!�6��M�ߟ�����������?~Jq�lT6?}aqS1�
�\���_�ʠ�)� ��X`��\|z���_�O<hǺ�[KC�J���ͦ�Ix�۾}�=��G<f�B�C�jη���
����C����׿Ձ�g��׾fO<�sOhan���@q��!����t8�� _��v��)�2�4y@Q��p,�\��ܓ���'�=�y�s� ��.�`ܙ�\�w�֭x �	5B��9����T�y��b�/�uh0ƈ?��lXH 4���S L�}XX '�A���l�F�'���	��!8s�<#τpŢ �����ٯP��9����y�#�*G�o��o�}X։�@�s/�k�6�����,����1�&�N�}Ü�̿���ꂛy欈Fb��'�)����f�G��h��v4���Ϫ��m�ƕN��I_��j�wĬ�e��]�Ɋ%B&���|ɝ��7�C�;��n�[��H�?a�$Wz��ST${�3L�?���Žy�W��J�9a�Xߋ�Jy��Q(S��[=���;��g�5g=��h�6W������ji��0O��!�K���D�������^�>��x*�>��'o;w��~��v����2�i�p�ho�xh��o��MZ �D����}?�
��hh�̑���l���Б���Ү%KŃ�_���j���{~�����=�B E����B��ac��‿�s����::� P|ի^b�=�<�����h� 0g^8$r2����a����G ˈ�Vh�h��6 
��ÆF����%�!�   <րC��"Дo�sO�t@��v�o4~�eВ0P0��� P�V��r`�,��5f�h�h̀>ό���	B >�3�@�4N��5��'�)$F� ��AX"�����Cb1�>�����D�p},&����A�#�{"`���9�^��.�'����#9��� b�y&4c��Dp` h�OΎ"�$ ���;|)�P,���5K<cߪy���Z�a'�P�z���u[,�i�r��u'�' ����?�1����,�ٳ�z�7�6���|�c�R�ϣ\$@�yϿ�.ܼ��iTidM�p��v%�$Mŭ�ʺ�w&!pVW��b�����y�p�O��Or>�is�Nu�9cƌ�C���lX���~Sf�Y��ϡ��&����CE���� ���Pa��4��p�n�R�֒9oP�]���x� �}8�2��,^|�M�>���G��PB[�N���k|�2'X��O��2�(���������{ #a��|̫,$@����3�I��������Ƽ1���
���so��f
�:tȅ��ڱ�rJs]@���1���9�p#���c�q�C�kG���P"$������=� �'����~ m��S��Oh�B����F�h�PiD�(D���[).�`yp=��8q�<��ڡ�h�X8�)��E�@��B8 �/��s!�z���j��=Þ�o�`�Z@X#@x&�-
7)oӦΪG��9ڇ�ΔQ�$����R�Z��W5|l)��B��1c'�KVX2�h��R�Wt���op���|��.(YC����}���d�27��!�."���f���`��R����B��X����ΰ�E���Z<a}�Hk�^g5�_~�����j8�?�$�v�"M<�B!;�~����t�oEˤ��TZ��B��_��_��Dy��C��h�����-�q"z-�x����U=���Wky+�؞}O؉c�,ӀI�������j�,�ޤ�+$y-�3��V��h�?�q�$y�I�1 �}�� D��PCc( Q�Y/Om����������I����Y��]�Ce�2��e�?�C�p� �	x�
#�@c:s���4n@P�|O��1&��[�L�#��z ���@`��h��A	N\�ﲏ?ό Ch�>��2V���%��7�G��X�D�H��3
I�E� <PMF@]{T,4�dyvE�)Z�9�|ȷ�ȗ(��'�s�gB�����{�L�nY����O�����5��zl��e�y�*���Z�jD�4�،����ɳ����C����k�t���y�5��S�7��>*���<ɡ�{�_�A� �a>�'='ק�K�ۛ���!D���+,s�9E���r�����2���=|�]񩞞�7�nB����Oo4B:}����K[?8�нG���f�)'���q���9�8���X@1���5�{���G�R�Ǣ����s���ai	�fh��n��v��S������>ف��b�:�/�&R	����11^LN�����(h�������"��?h/4>Q��h��1�����%=��b�a��
	�o
)0E�ֈ��'�(��Xt��U�d�H�(�C�T+�� `|Ou\��>�Z��\GQR$����r=��M֤"�؛\K�+t�g��*���r�!���e�!D���h�|NJ��#d���?`�gEI��<p-��n���:��b%p�}��i����y����}�+�АIX!�m�/�u�.���_�ڤI��${*=�jP<��;�G��@�<ɋ�?
������8�U	���U���B��u���@���38���8��h>���i���@Q��4�)�&_{��f�������I�����fU̓<�0s��җP1����7eZ���wP�OA�
�xk4A8Mi8�������>��G>2�@h���*�v&��"a)KZ���L�b]'xI�b)�<���?l���'^�ڧR�;(�R��p�����p�vc����b>p�AO *  �Qx
��ϡBbJ����7�����[U�l\��aN�	3~Ɔ���@B���u|�4~w��+|
��;��X�@��*?@Bٰ��W������)M�����ݮ��{K8z_龾A_��q�����T��br�	�
G2t����N��!����G�Gs%��s�̫���{�4����SF5SM!Q�Q�$���[��8^`k�,�t�jTM�C���KmּU��W���d2�)-$t��hL{G0��sS��O����� e_�w�5�Y��`-�|� <j�� �J�=���u���zC�
�J���B)���z�s��f��m�>�����3j�5����^���
~BX.FA������]*�tS�8yN�IT�d� Lp�*(Հ���o�;~0U����UճZ���=Cq7�>5J0c2;z�ö?��� ��2����{?[�D�����/tǫk6�vc�\�y�X4�F�I|���s�� � Z<�,��CX��@ �
�s/zB�%��i�:P�'�4DJ�LS~���e�&d�E�1i_|A��4Ƭ���"��rUn�������wyN�/��Z�l��D�B��A�/E���" x�Q8���e �������J���a˜��+!-Ag���|f(x�<����tV��Z�B�������B��p���S$'g�-�իϳT�j�R�
��-\����_c�J�2���C�Fē�z��Ԩr>��W/G(Z=��,Z��!�'�H�#��u��ϧS��T=��s���)�����M'�<�s��030�'b�$n�
�w+�/�ԁ{+�U�6�{��O&��4�W��{�ő&�CqzA��E��u���ٗJƬ�����s�>q�k�P��H���G��w�o�Y��]F�9#��� �5�����s�n��R������C��� �04�Q���H?��<#��sv�P:�kp �� ��f�=_A��m�T���z)dt@��ӜųhW�\h[6�6����)U-�j�9�۬��󗢇�r���p,|����`�̠q�T�,�`�?���*��n��di5fBR�W�> i�I�=�B��C�����ʭ����y�p��B�	� n�bg����!rE�* ;!��<�B�������H&��c6 �?�hrI��a^����:���O�c�d/�J��il����=���
�PŇ����_d�f�䅹;r���ND�?��NJ]*�ϸ���,����m �_ڰ��у�\�g�5��'����/�n~6?�pc{��O�R��{�nظ�jeJ9Sч�кcl�����:ަL�a��YS�8/�\Ĳ��W�lx@������9T`�4{�9�S�Ƈ�#�NTD�<gIB9��"r�T>���Z
V�5����OX�<��?i�|��>;t.��s���?^�`�U}�tTN�`~�<��S�.y%P��K�e�e�G�;�F�Y��l�-( 'Ǐ�P�UG�v�P���u�I��Q�J՚[&؞������C=�	Vb68�PO|u�p$�!$��5�\��Q矿���0�I�����""H�h��Eل����^��p�b=Ȁ;�q�z4ƿ����* I^O�����C3�zd�mӆl�����ސ�X�HDƊ嘍i�`7]h�<�C��*UK%3�h@��$�|��A�od�K(��ɏ�)�Q���N)5�y�B('Ih!h!j$�ǕM|�жi�Џ�7p?K�$��J<���3A�NXA�w��\� ��0�j$�}���$�37�k#̐�I��Åz�����G�\���7�-V/�[�O�l��'��{�%�S�&.�g͘�tV�p�����f�����t�+��ꡉ8��w��ͳ@-��I�l���<�8;�� 9N�{�����ϥy*�?��C �vklHY6�m�V/���ά��(
"� �X��Ŋ�3Ѷ\x���!L
�'I^|	�-�s�\�5��;���9O�����ij�e��+��R*{���	-G4}�ߛ0�&�:�O�2�/����{�i��D�T��o�+�����'/� ~P���N�B�#a!� J�@��G�'`K4�����B�CT$o�    IDAT=��5f8��'Z�����UK���֫Ikk?b?r��z�I�}p�͟;��1�	�EG�F���ybŊP'��@<8B�������AU/�+��{.��sm��טkY�RZ��ϵg��2���O=,r����CU�T�,ޒ-^0Ӗ-_d��P�Y2��`
��?�2��l����b��/& V ���_��C�dE��E�I�Q��a��b�!(T%����G
������������ng�O=���n���:���$/xp�RK�)�Q��G�"qy)|���(� Z@��(���Ђ밍�Y)"M�Q/�ŦË�
��[�Zo�I/�L�(�&V�ZKZS�D��/x�z�@%[�p�͟7+d�B�h�K8y\�<�-�08^�|@�':ģ�Ik
��B�P�gb=���2fEJ�Sʌ�tT���2��8Nk�Q�9���:���Z�2��%S+�<d���P���Lc�%S���<�*U��:�� �zb� /�y��Y⥈,�a���5�.U��AqW����x(9%"���g���K0傥����O�4����G+�P����h�l�F��S�jH���-t�pnii�E�e��,�;�vR�66��uF�5��Q�o�j�x�I]���v's��}m�����>K��?Md���d�}y�1�'��Λ�%��//�k8�G\����o
܉���\����X1��p4ro����}�=���ϊ��"�c~Jy��U3�O�����>��t�Ϥ�V*g��9f-�)�2�+18�A��ĩ�f�z���cA�S�z
0τ�=�aťpVi�Hi��E�D�Jm(d�L��ǒ��CkS��\�ԦN�l���>Ι��<�4�87	���{��4N�R���U���b��v���`��fO�m��_�9�f�E���MJ��kRH������?�I�#�H�����iq��+��n�,�pm�6Q��?b��<i�l�e�^�ө�QJ�'v�c]����gΜn��~�3F�	��|.�WQp�����_q�K9���@��p��B�3�����g����w�OQi���?3�s>���:E�-=��Z���� �C5Oj����9k�]z鋽�o2I&P�p���!ڇr�p�(e仼���p�3�T�q�?����G��	�$'f��6�lkl�0���X�ʢ{���?�'�[���B�D����Io9+9��K:WC&/N�J(�If���+^�r�0n�s}D��S�N��\2�0Ƕo��}l	o��%�dh�
� ~�EI�UGvM�̹t���JV�^��b%۽�!��M�Ȃ��|�7N�f�ut���&%~��U��G (!e$�׭e�~&?E�Q|%J��Z��
@8ʔU���� ��Q2���
�hR
�>�@�E���~r�X�6�(��CNa�<��!�\���F����I�o9�d��}�C�+�\t"�a���C��d9�"HX#Y����"K�<������h�g.f�]�|*��퓴B�7�wX�ܬ��n+W,��X-�h�bŒ���[(a!�����;`�&ݟu���6Dӕ�^���W؟�ٟ�Y�B�zq~ɘ�ҭjT)L�(��m��\��Ək�=��'�0c%8�����;�)���`��fa+4t����Z����ꎢX�3M~�_do|�묥�1X�>|�v<��u>hM�F�=w��w��:e�KUK�3��J-6
�!P�v=un���S%�M�g�?��O�#�xp�>��{��ah_�x�v�z�N�8`�B֒�%c���IKc�x۳��{߃6�������i>2����hN!*~�vv�u�ɆV�3�B��E	I@ոK��(� �����åB����G�5%PD��k1&e�J�]	/�[��響�
�IX*ƛ��B�{�:�k�\OUe��7����s�R��e)Ei���sܛ�Y��ҳ�7����SB����5�	�_O��~�O��P�t*f�B�mް��o\a�b�ҙ8ͳ<ο/�9�Z[�ٺ�<ڇ��yXl,P���Tۇ�Y{���k�[�盽�P�-@(P��o��"�٦t���Y�\�\��k����<��,��#X�����^!V�>�
�P�`}O�'M�r�Y�u�֛�{z�=S���$��y\�)S�7_�*����V-Yϩ���#?�'�|�Nv���f���/�bp�]�l��^��#` �������
�S_���ԽA�!���fΞ�%��4
�C� 7R�'����	�9u�N�<l�~zc�V�X�XC�kk;����Bm�~(��}��3X��Z�lF6;σp �pg�R߈�a�J�^�q�?'�U�+����Ł�����Ɛud>)��f�9c�GF��!sH����q]擒J����z|���N�Q�D �_�� �}d���&L|�^�ʳ�ٽ�AV�E�����B�j��{��� �oX�� sĵm|Iܟ�9撹C9�w�&*/j�L�2�+�j�x�$.�mP�_�Ϟ�<�G�����S�e�r[�a�U����$�����i6a���I�@��垓!䓤O/R*�y�k��G)�����y6�d��A������#�@Nb)3�I���K����{�b��{m����s�c�굶v�&���%�Le�;��fh���BEÿ��ugga��[?���s�3|��aH� ݛ�'o|�l����kk�i?{�^���MQ�b�jI�!�j��_�%KWٺ���9����}����)�P�p��+��~͵oqI ��<hm�G���zmr�U�=�޶ݎ>�!��$2�&ۻ�34sɖ�ݤ�ϬuW����q �ď?��mkmE����u��9�S8(<֍�u@�������=���T����>�`��6�8�i��e� ~��O:�p㾔� �ɑ@s�z����cԴᙼ�s<X`���Yփ}��!�(W�㟱"����������C�s;�^MI���O>Z!�{�Y�ʝ�	z=pO�hQJ��_��"�3.������X�p�wXc�\��&h �%�����5#y��O-�b��3|�}⵼��x�fM-m���6v�T��˚�.�֡�C2c���,}~9��\������;n�Az#�����9�;��B��#���<��`A�R�q�i{�ч��'wG�1�K���z�5���V*�l` g���?��Q3�a�
��{����m���~8�w����Z�Z�7��Ͱj�h�>���������`��KK���w>W���S��_��lŮz�[h �]9�2���� ��y�k�>��O;� ro��M�D�i�=(���?Z��Uc�I&,�(Y���־o��j%�P��\��G���)�?!��_�X-�FJ��� 	��j��@?�Y^��KD��h�<� g�	 ����e��?��?�k|��?�/�@�i:z���ŢMQ�N�� ��V��F��É��`.Y�@G.�=�3`]L�:Ʌ%�)����\��hX.T'eLX>T[���vN�̯��9�K�y���?�k����;4|@��`�ױ�G��P�Mj!!d�/h@ ����{D�QdA�r�
?t"�E��BbL������g�UF�}���)�`���Z��֭_j����9#0n��l����a�Q!��]h��D�F1���:0f�����Vk<eͭ-���WzIg�?���X��a�{�ö�\>�O2Q�#��m�欄<u�{C�|��kv���,�����~�-Xx�o��|ͅ>��|RZ�(�svk���?� �i��ٟ�ɻ��a��}��ٺ˭Z�Z[�.���]��Y���v����f�tۖ���9|�2aY�K_[�G( 	��}�{���ń�۶�,@��06�\ФG�},n�Z�j�y��v�X��k{�
���
�����q����M� -6�G4?ټ<�f6���ƾ�-Fh�@�2ln9����̛@t��j)@{�'?�@e�5Lj5�ȸ/��T��µ��i<���+!r��E�s��d��C��-娱�кyV��5�y��_�6���ͅ@���u~��<��'w� �U����b>���p=,�xz#�Rv���c��+Wz�4�{
���PE�!X<(X!������e/1G졨������ь��?���D�V.[`�6,��J/x�����Y�-o�V��{�s��sJ�y=�9m'=������s~ޒ�}��wT�,`����+�	�|��{��߶���)T�N���o,�Z��}V*Ǭ�x��ʥ/�K.y��3����ӳ�i�r���=��붭���a8��DC�9m��p���J��:q�~��o��e�������ug��R�ӝ����l����6w�b�r��g��jY|�EW�q�U���e 0���"� �5����DȌ�Ex&E���:����y�
�~�E��D������i�_����
�D�'��.~_��&��w�.PD���`i^�3���IVh�h����g�xa#<�3 >��(�CA3Ѷ��];��� ���}����چ��h� ����}$˫\)�8xa�߸?��3X*_�Hx�G�((��K_�VԞ��#�lX(T<廔�� ��Iz%�	j@����}�.όe�����)8�y߳k��=#�g>��\ ���G�T�'�Wq��zU�P�'I!�ꀭ]u��߰�҉�F#��Y���u�H4[�d0�Xܳ� tѢ�&g�g~���>Ŋ͘5ӕ��v�g�Q|��P|�s��_؋�S�'��c?�x�-_��&�c;v�E%�$䥬�7k��t���v�D����`���w{%�#�N:%�s{h�?^��?��������y��m7�`�I۷�q��[_����V.�Yǁ=�M�S����Z��C��ڎ��KVx�T �k�Q���w%�GQ��b��C�븃D����>�P�3 "pJV�����Nkk{Ҋ�^knL{)j�留�}Z_��`i��l��YV�~$�a�W\?T�ҥ��8>����^��Q�]8oh4_�X>80�<��&�"(&N��3�	���C� � f��C �e_s�N��v��2� &����ϐ�?��$3��j�O�<���������G�:S��b]� о�7_��^1����h�?/�A�#��cg~^��K��_��S��茙�&X!(<B Z뭩�ѝ��
A�傰Ta����������B�Y�*���N^T�ݸn�mش�j��OTi��V��9K��������4y5\b�CE�������hwkݣ},a�}�����7��)^�q,a�S�	5��X~"�9�(��{����a�2�8q����J�Q�L�-�-��]m^|��'g=}y����ߚ[�Y.[��|�c�Ѿo���9��O/�r�Gz�{�:��_�7
Y8���Ʒ��g���v�7���������|X�j%i}�y��+���w���e���Fʣ��������B��h� #��Vv����v���@�T��/9w��y��;rp���V��Rλ6���X�ہC��{�L�LC�
Xϛ7'���k����+�ꪩ�%����'������n�Mp�j<�g����;��w�P���] ���,%4o�V�Z"�`'�1 ,C�i�p�{�X�y��o��8��>%�X#iϬ-�`�<�Ȝ�7Y�'�{X>�=����>��<3���������+��F�0G(���w�� �N��Rr��ޔ^{I���B�OE�9R�آԠr:Ȣ B(�i�U	��8�D���c�#fӽ�?�\���(���O���[�fm�ʅ�y�*K'jV,����V($��a���0�����uʜתa�]!����٩>4�P2� ~ᅛ}MX�T�jemI�"�G�����??w�z�~t�7lŊ�6}�T{��G�Z�'/h���,�h��G���d�'n�L�����ܳg��&���ׯC���_����~�<�d��Fx������w��55��Z�ٿ��?�E�-m�W����!y���~��~�ʵ�=^��.�
�L6a]8�?��X�K.��M4/�M��p-]��7����nΣQ@���Wԑ�{T�|�������U�$%��*W�6n�4{��6��COZ_o1����m��6w������r�у��P̊� j��U恟�gW��*��h�\W	[��G��F���j��\ �\��o�D%W)�_��Z����
��}�[���9�џ�R�38e�)7@m�J@SG�~݋uT8��y�3��5ŕG�A֏��T)�?��b�?p�T��	�g!c�9�H$���O�mUP�/�BC׋�c��14���H,,�:y͝��N^�5���Ջm��%��o����:M�ן�1�&��~�R���{��J=�'a1����[�p�Z�I�я~�[�2.|?(������s*kN������g��g����1}�577Z{�^��(��T�1{�g;-�i��ǻmݺ�쥿��Ǝ�d�v����S�N�?���[g/��F�`�1aM��r�6[�v��,���ʀuu:���]����J7ہ���y脝8U�����\�����)�8����H���щ���ܻ��ݩ*f�/��hn�t���Ås�}�N�Q��s�
�>76���L|�����x؎�pb��Ϝ19�i�*pÃ?�*�#�s���f-j`E3�=Z�Rq *��<)��M���P�: #Z/��?@(�s}����=s����氢a�!�=�/�&��X
<#���+ˁ{�ys}�+��s�;�Sy�ų�󀇚�3V�����%$��3�¼���{pO�Y;w˴�V�,��ʭ���7��2��J�����ESro������i�E�:�Z�(���~	����?w�i��U<�w��́���W,؆u���-k���'E���%l�l���j�/Xn�\Ś[�?�Y�����[��Af���!jg�	��Z��BAOr�yvĬ7c���p��+���'-��B1�:�3ꊱ�-�c��?o?��Þ�՛�����S��w�|F����l@��Q�&O��K�����N�b�8�P<ekW���\s�UJ9+���c�#��Ȟ�ŇO��	ո�eK�(���.X������㧲K�����+�� �N��p��׹�@4�����pM����f6���-�g�'��b�ϓ�0)S�9�{o�=�}��lt��l���6s�3JZ�� ��p�0Y�d�8q�/���9p�lv�`����������9<�CB� �t��	��3C����4Y�(������*x2��a�������<BN<�����rc\|�5b�rƁPC�#�/������@ �(�7~|!̓'dM��kϸ���S��d�TB�H�W�>�a~� "�D@/��f�j�0�`��٫Ap�7et�������b��,C	,��>�KSԂ��W�N��ГV++Hc~
��4�o��L��^[�`�-[���P�������y���<j�B��O�����ʁ��k���k�Tj;g��r�-!(�=�S�e��Q��3�l��U�}�־�������',CK�B?��ez��6o���n�fkjn�����˭_�g��%dߟ�Uo�r����+>������8O�f�KUZj�<���T�����~��ֶw�e�h	w�,�`��۰��;���,.�@4HT{��%��F� ��c��M�1݋E�� ��!���>�i؃A5���=�i�|����!b�b�s�X���V,�(ڢ��'���5�>h�42�q��
-��w�r�g(0E���n����K4Q4~g���l�� a�1�e�XHD�`#�=959��4s��7�a0�����D�0��:"��y;D��	��B���p����0v7B�8k��e�#܈���K4 �{�
 �m���5'��H/�V���A� ��׮Q!5��8h��J��u�Þ�E�;�'_�T��@;���ח��U��5foHj�D���	0G�}$��\��=b    IDATG�ߟ1mz��{���������T�p���^��S�*�����z�2��6~�Tki�h�}Yo�B�x�O����H�T��Q�z��#��"�e@ԗ(4YF(6��Z�`Ǐ�����ܹ�:vX:�r��YҦO�iny�-Z��b�����/~�KFU"�Fz���?ra7B�b�@��@s������:�?g�d{h�`'O��G:�6q�T�>m���0�
� �qڢՉ{�@�9d ����w~�@�8��� p�1�f��gpͬ}�>{�G�����U�9�N��Œ�u"g���x��*U"�ʶh��={�����5���c�U��o��Vki��I���p��Y �Z᪀. �Q�A��{r��	r� ��L��;L�� �ѦBݓfP"bEEf1���y��Qr��/͔�� >�q�L|r-7���C# ̱$�=������N4"< |�|��)��%�M��~��pX�V���yf��1��x��rҨ����s�8\W&�0峚	)-eq�Q�_�蜨�XV��Y~}G�CV\0�0	Y.<{��s�����P��7�v<Q���36ab�ūeKg���L�<O�P*ٔi���/���4��>�XҊ����T"��n�5��jj����'c�p�����|D��(�2��o�iӧXKK�u�:aǎ���9y��Ek���lμ��L|���;v�W��ekko�Ʀ��p����+F,�������F�m��������
[�t���9-^E����꤀S��O#Z�*5ʉ���&�Xt�.g`А(���녺�.p y��H��fO>��>��V�D�f2�Gi"���\���{к{�Pn�g�3g�͙=}��	��4���Bp�]]�|��PG�k�dx�MJ�����? bM �p��������NT��ׅ���a�p1.���4l~b����.f6�:V �6��pFx`�Y�ϸ� �p����j��u$�@���s*�-���`a<<'�\�
Q_�����-%�ː=��QA8��9a��o9��KQ�;�ы�����×����t~2�*�w&�"�)?�׿�w��`���'F�[J���p ���,
�u�{3f̪w�:s=��\�ٚU�m�U�<x��$Z��^7a�]��_�^M�c��A��),2�����@_���;�|=�?�>�x�;˺D��x֐u�|�+��+�!(����l��M[[�z�Fj��FX�߼�۱�I����G�p���)��;+�}Fn悃,t��@�ĭ��j�9k�4��.��6n\ocƵ���d/c��'�w�s�k�Q�5�Iy��k��B:|0�OM��W��8sB=���u}��V��;~f'�z;G��	�DXa2����~���!��@ uP��ϡ�H�l^�3P&���}�k_qpE�E��	��xf��d0��M����{�s���3��X U ��2P$� n~"��_���9��\��.L�Do0� >Z5c"��sPX ��'z�g����7�@p���\!w�5�8�@�E�>'���Rh����>� �b`��;�[�M�	��H/�.�0@��v�sF�xi�cBԌ�'��Ⱥ�x�τP�rGi��>e,������ʘk���sO���@��B���I{e(D�?�$�,
B�4iJ��^�?�N��n��ev�5���Z*�L"c�r��u]�w6v��Z��� F!�Y:�`U��jN�p^?����A��NJFdh��V2�{��nͣ,){P��]�K�㖑Q��]I?X1w~�N;x�@(��sX��b���j�Z�2i�gea���8R�#����K�ZM��%�Ny	 b�d?y�7���{,]o����,8��& ���������h��f`S����7Ra7�:�&>}�����FS���������?��T�
�!�J:��q�9G+��a'�u��� �E��3*MV5  ��\xm �a�E����y�&��� ���=�@�= D�����YE�p-�V��=s��m�{@�0���	���,kD�Q2�@�]����@P��C �yc�h�(? !��"���hrMb��h�0i�\��M"�9�惤D%�y< s�P&"�u�>\ۭ�tz����9o��~/�c����S�eNX�B�����J��ҳ�I � Z�5�%��q�?�f.���[�������X������R5�i+T����-8υ���i�BD�"�����7�)��66X���^����U��^�0?��^��b��;��Y�g��:8�<�´������Dw��U�EK%C2�sWü��[�ʒ����C<�)�t}ʋ��J)$	ł��� ��kj�;:,J:�	p���x�l���z�'k�U�������$�z̳�?��R��d����;R� ��4s�8
�s�eL�P���b�n�*iH�N �h��zդgNWϼ�.�Xڧ�4F��84�����gĽ2~Ơh �3�7��6�h�pW��r�	+��9S�-�仌��Sa��}$�枊����O8a,H����9�F)���h?��C�� �&;���yQq!���^e}��e���~��{�}�s/|-�e�K��B`" �h7o?�:%X��	+,�#�	�G`�Z`/Θ>�����!bi(��鞵5+��u�\9Jz�k"��է��isl���ij���B�l�J���S�롞��>p��Y���&R)+�r�V�/��5V������"��(b�>7D#y�!�h�4��M��j}\X�����b�����}����
fR�%;���j{��zCo���A
>��,H����^r�Ձ֏���D��P�#��'�[>4OBBh�7O�<�����{n��y��r�R�c���p��u�k���g�?��q��(ِ��IA���<��m��1f7��|q�q�r^lz�I�աW��(��p99��:5�L9�&����j��:�-�V��Ys>/�Ut
ϫ{i��$%����D"m�46�����N}nDo(�����XO��G�W���}�;4Hi�DXae<���^��1 HZXS�?�+�Nܓy��}�53��דlV ����ʇ`]��_���,�:8ЙX}�M��O�0Ux(�+����^�2�X�X�Z(�i�C�W�����ﭽ��~���v�4ѨkV)V��e�-Y��2c=��.^iώ�z
����	sa���ߛ��S��\�W�d͘/�rg:���9��N���+8X ^&\��H4�Z�{^<h>�P���(�;��=�L�� u͟�^�����Hl0�������F�_�%^��A��g8DD�l��B��Y" ������ 	������w���Y��S�*a��G��͜5���B�؀����w� /LH�=���V4:>�Ӕ�D�h�p�p4H9���B��h)�(� 0��VH"��eP&h�P9�Q�T��{P2h�h�P��JEà���g���c� Uċ(\?��c��l8kq�)����$��1C��S���U/��% �B@�F�Eĥ�S_��9�/�{(�ZV�@_�������#掝�����_[*�v|��I��E/r��ń��9��<?Bp0��r(i��ի9�%��4�	Ʌ�S�5�2��$�h0�/�!�G�k!�
-���Â?�/��Y.{�6mZn7� _��&�*��]a��-�l�l���Rҙ��U"D�Q�Y�����ł��
)4n�+�����S�J~]��{�H[]���[ �
_E�Rb����>�����3k��^v?��CæB�?U�L:���o�����$V]�ߞ���۝�� &�qSۣ��{��1���y
��Ъ�{�d�VJ�`:�����'�!�\
�Ā>�ihy2>��������"�	�c���w�#4X��8�8`|0g 	�K2���g�Q:T�D��!L��Ǣ"j&Q7X]|W���h� �N�(�%�b�B���1_�7@d�h��;�	�?�G\�U�q){��8]��'m�>J$����hd�?���_�h�]����O*�27�?J/�$��o��{q��g�x�R��pt{�{�A��G2�`f.��TL?���Ǉ�~�~.��%N^Ԣ�!/���b.�k(I���6uZ��sZ�W�o��C���/jum��/���J�d�r���/�CQ�������k�p����`�>)/�m��� {�hG�Z(��K�'�Gđ�9$1h�`�����?�_q����t��ax�B�Y��/
8/S�τ$�@w�0(��
�BY4`�)�C�Aw��������А��0�5F���@"̀��y܎�g�r�A�fko��K��J:W-4s��l4�_�9��V}�e��1���o�fO�����I�*��.��E2�J@��U�	`��4����@  ���P�8 �d Ѐ�*��|�*Aa5����c�!��.�
����3s-��  
�@�po��8H8�X/�<'U������/�3�����%? �$�ƺ#���!�g]�2UrӾ������lf�q
������Z.�����!�%��ĺ!�A+A%`�ܱ�]�/���|=��L����^w�y�3��ZN��
�cF0c�!DP0X;	��t����N���ok�.q�'Uݮ*��
��ҍ�_�zMj�s���רµ�C�p�cu��c%Z(�U��:�pܑ�߱�V��7f	�r��C�Qh(Q�N&�5pf�0Bԋ�&O��t�nݶ���==�?#�ӭǝ�1��s���>8xc!
Ӌ`�D�������%�@��()�;� ��h<����9|)���1^���v��n;y�Ò�rp�Vj�H5Y[�Q�羇O�%��?}����f�h�`0�n�r�cf^���ޅ  �s -<?`Kr?q ��7MH�͠�-��`B� ����E�>?4��5 }�w��� �.s!�8�l���z�j   �3r����h�|������R ��x&ƅ3ap	 �e H?����H��b P�)!�b2>r>��u����c8w����A���Љ��n!q}�A�s(�J��Y��,XM>������M����S�3{��W��khl�<ւ����{���G�����SXŬ#g��V��8�6p'�+��Wm�t"n�j�V�Z�߄�-��Y�Hᴄ5��n���Vs���Eע`����{0;��\{�gF���r�d[�l�$?��9�Bs�$�%�	qbSB���P\���$!�⊻-K��fT�h$M߳�>���=�myfd$�����5�=_���y�zֳ���փ���V�T�-TCX���gT�O��H �;FX���k��]r�O-�/"6 ���Q=����ܲ��==ݿ=2�G:��+�y�j���@�x$��[�lSo��2�'+�>�>��8m�U���ΟI0j�7V�C�vX{�~��=f��R*V),�Գ���n���������o�h1��gW��@ �D���-�' �{>t���j�i&�B��` �X�o�� ���%`�#��^2� �=��my6� ��� e (�}��z��K�P  ǳ�;W ���� ذL�2ѯciC}@��?1�U�eL� 	m�c�i�6�jG*.Yi���:�����^oL�PY�˟g�j�Pb��.�ω�	�b��b���al�� zyg,*�w������챋6m�׿�j_t�&j4�+��Ip�X�;�U�s��Ρ5��zO�w�����b�}y�x]��9��G4��iy��3��ʝ�Z֊�-\��.^�ROh�z�c�< ��w�>��	1�x�p`~�+��@��lO W�cx�����%@����޳����0'��6}�uw�z��O����G]S����+7o�FOo�F,d^��C���A��� �Z�c!1f�R�Z&I��t�^�SBQJ}���A"��5X ,e�q�'�`��g���^��XC�E*��G�7��]?��r��54R
~v��uf�
`F��k��ď>��SX� )�\�pŽ1��$��X�����R�@W���X�⻙����o �����Yx�G�`����c����B8�TAE<--tx,&PB����|���|��=��k��N:�X�B'�����bժt�(=��(2�O~	%��p�\�!��}��]�Prܧ,�����m�\ v����x2�#o��1�Yp��x�|�G��:V1��vIlǥ����546:��x���L��њc��1�v�{��Xg�#��! E�ܹ�O��}��O)f#��_�ފ�~�t:k�r��_J6n�$��%�Y�P���x���\�Q��$fG�/������|�j�:v�0j&�l�H��w��H-;�~Ľ��/`M�'#�y�hL����4�O	V����O`T�g��C�\(\�B!��{�sN�v�MwW,M�5��bV.Pf��_���f�^>/+¥m(��J�*H'~�c`�B[ <E/&wb�v�c((D��'�T��6s��`����G���~�|�q�>Fk"\I�y�Y���>:�x�G��������P��{Խ���s�9@u�X�܋��`�K������<;�����m$���`���^������ه�� &��]��K����]`aSo ��V����X�ܧ�`5����R}�����|�uJɽH�X|����"��y<�2�B��NUD��2:(+!�G&�;�
���/�Z���b��Y�y�P~|�u ̞��N�9�'xx%ހ��g�������ؑa͢������~g�w�9��g�s^΅7�K�ϙ�	�ּr�	ڧųy-V���,��kVZ"R�����K����[��l��(�� ��k�A2�����Ywoh�ٟ�YC*���?�Y����ƻ�~��+X�q��T�b����p9���?��;��1���>�Bry���UJ�S����ӯ���ۿq�Y���>f>��������I��Ix����CB
3�$��E��
�(Z�e�B���=�����h�W���p�'Mg�Jɚ���)cbx�-���v��[gW�����q�6f͜�Kny����Ț�Z�p]!X���y2���r?�G� �~��@�y"���z��"��ZM�	�D$�H�TJ4��$��p�s��¦������R�<�)�NV>����<₹GY{R�pn%�q/Ҷ�K��O%��̉�p���xMx)xP��TO���[��?��g��X��t�L�����c��b}:��#q�Jc�w}��>|/�������,�Jy5U�Z����� ����dB�(�J�8xW���+?���*��s�8~����=�W���6yJ��k�>��@\�x}���{m _�δP�d�¼L�k#�u����.������7_�ޗޫ�5׍���Ҽ����Պ��q��/���C"#�9*5�ϱ25�*~̐�w"?`���c��vr1eAk�c��p��sw=�t2�I�:���e"���y���
*k���$9�8MMf�����V���aY���:X̎v���V+��Y�Z�bs��O0y܄�6P(Z#�,zXT��/�ksg��C��h��`�t�LƯ�������
P��1 ���Ƶ�>���'H�*�zЕ�㗼)q٢K4Yd-�2Q� xn���6r���i��z�N�,�kl�V�����{l+jMV��1����_sl�A��������D�������Ρ�J\ �
�'����*��#N�	����,f���pn-bl/���#!�/�E�k�Vc;t�X��˟�2�C�"���7׌5;�F<K��<*�w$�oȦ-_豄ap�,����2����%2Y�4�;����N�����U+�iCRk��ݻ���@��\�x�I    IDATt�E��>��Ϻ�#��K��]=�%.�-�m��ܠQ�o���E_�~P���m�q0���ij�X$�6�yG�Dj�k�{�m�Y���}"0�e�9h��e˫��=�iC�,/�� ����yйm�|� ���-�1x .Y��r�ha�� ���@�i�X����n--��ˤ=��#.Q��g�Z����{i2�I�d���ϛm"Ji$��m���+� ��T)�p<Y��U!�wՕ��U�&�����_]� �_�qh����\T���������-eYr�L��D5Z��S�|��k�z�K+s/J���U���[�eK֠�x- <S��v�8�<C DupD;r-��� d@��>X������N��I8�Ȇ�������u�ߺ�)���ϖ�П���w�x�AV���<h3f�t�b-��L-Z\;�t�p��"������}�!�����G�8O�:#J��,��v�U=�.�i+V,0�-���܍��GgL�n���ם�)�B��x���/�r���h����-�_�ީ�o��g�3�����_≃��/hl8��lC:�S��J��?z����$>��9�*������?�Ο`�T�o �믻��]�B��\���bu�o�ץvP��;d�q�A�z��]�jչN��8TO�>��q��yˮY��Cf�iY�X������c�w?�%����)ƶ��_J.D�aGfB*8�X�ҭ;���{����e�>D��,]�O&e-^�ʗ�{�uC UqY�ҀkR`�����5�-��N �`. �w�EO�k$�C�9��L.��J�d�s<b$��4��c��*�>x����y(%���Ȋ��X����5h�g�q�d�s\���E��hav�2R��χ*��Q򉡼�
��=���r���=���s�<�V�ȸN&��HB��3����1u�+��s���i�?�i�S�Ѕ��r��p�5�x.	���)�0<��S�k���Vڅ�s��{�� �$V�Ž�������K�a�W�������@<�"���&��1�������[�t�0����cbC����pA����d���t���93��<���E�u�ڈqv׏dw��c���b2u�4��?��$y�V�b���NϘ6�9t&���|�2���O����x89
�o-Ł���y�L�@��Ǫ"�&:���@B��A���B�`;w�ԺzY�B����>�����ms���^�9�o�J��}O��W,d��:�Fp�[Z��D:��2�wJ2 �h�YXP��FÄF�$���Ft饗xP���}��>� n0�8X$ @*Or,�E�)E���J�.��a2�h��"�Ċ�o�&19�2��*��;�����-�<=p������Ce�M��Y9/|0E�xތ��	 �x�я�t5Ǉ.Q|����F &c�w�@8cL���`�h��x�=��� �\Ƕ���R�s�����B��9��do ˟�� 7Ή��kg_��k"������c�?��յ"ϲ~���=�l�?b�;рıh�T_ۇX��z�{m��e��5���v�o��J5n�R�Ə�l6n�r%�u~��{�0�w�g`���_��7���j�f�t�����"��2��x�4|g?1��1����@��qD:s���y��<[�>�e2$�%����=_��sx�!X>f��N���@�	N�>���o��V�<�]�|�߶m�x�>;���z��2$-�M�.����3s�"SU|6���4�L8L\H2 ���f�Q�< �Ԯ^�[��b�wv�ֶ�V��F�5_�5��%�wo�=��v��F��h���7o�!۱�h��y���C\�	�\'���@� 90�lQ��< ���H��&�{��# �dâ�\,,,"�+��)��YЋcb9�|Ѣ�3�X�XX)�`Cͱ� �(^H b�}�+Ã�<o
�2Ӹ~����ɽ��&.��<�7����ޟ㑸�+ә�)S ೨�����=� �����G��F���2�E3��L���ճc�O��O�y>��V ���?���?���YE�?��sƻ�9S��g�"I5 �3�(����wd� ���q����T<ԓ��k���˸`Fyĵ����YWح�����X�V����;$�H�$%�B�����l��ɶp�
Kgm0_v#�󧼇u���4��9d/O�1������w�B�\�2.	N���sc�+��{���x�믶���pgg{�=�����S[���7j����k���um��3�Z�y�����{DQ����=}u�[F��|�)�b�6n<�^�ZR�y�kn�k=|���U����)���Ҩ;oG���ŗ\��\}���I��Z�b�P���L�s�� �﬉	0a%���j�hR��ԋU,?pܞ����
��Ɇ�Ka��UϿb�X�-�P��U�f�(�P��)H��|Os��

���ʱԙ�ߋ�@����ŁkYu�yVX�,�,xz������aq� K��,(���� ��U�p�u�Pٖ�3�Ylx)�6,8�EZ��]�=ۯ
	���\�!����,"\ 1�����0tV4�b��d	�+d�+נ��|�'��C]���b
Xq� sWO�{9�a�0f9.ϗ�Xt� �� c��v|xWlG�>j�o�y�8�Œ�(�8k.Ԃ%p�ߙW�'ȳH�����1�����_��������v�R۰�����K��l��6}�|�0~���|C�8/��s�_԰�+���}��N����*6y��B�x~����R���7�)��*��n��6��?j��6n|���Z��>5{�寰Y3�z����vo'�{S<��8�7����nX�����k^s���a�%beoܞ�Ĭ����=�2J�R
���{��y��b®������L,'��QCrԣ�k_�]@-�D �Ky��'�?n�Z��F&`��e��n���\*����=d�����w0wsm���,(�H��������d�2��` hi���bun�`u�`�tx�,�,?��9�� �����>@V�,,HJG�i`U1��o��(րE�D0��(�@k��%p?瞻�3}ѕ�;�Z���k`q���Y�w}V�g�ǀ��҅��?���y�O�p�Tw�= ��
� �Kޢ���G��R*	L�N�g$�'�<��}d]C�K��s���ȣ�X�޹>���'�%ZJq����}�x(|`����y�#.�{Q@�,�������3�k#�>��_���y���J��n՘M�:�V�y�������c晐��F!�9i�|Ǽ��_}��LG��l�Θ�)p/�:�Zq<��^���&����֪��m�Σ���v�Z;�d���Eڑ�.+C2��|�M�8�b�?����n��.=WŉN��>�7s!����N9���=�o�tܲ��v��mͪ������u;ׇ
������:�TN���.���_�T8@�)`	������2�\l,?TG�v�$��W� �Wy��
�Ճ�J�j�׬��նm}�ʕ�gf���}�?��J����"/��?�#����\3Vu6��4�@������p\,y����m��� :�29��������"l <�?�����e�1�U�sJX� @̢�����n�kp��_q����{-N�3�[���11���\/ �W�g�f%� �b��xlâ(�7V?�f��9.�ͳe��&2��3U��.�lx7�[ �Y����<S��8d9��c9��J��$�,2�I-��s�/�c�O%τg�"ʹ�r@�f�xx�.��=��5��X$��)��:��Q���@
,�ݜ����;Pw���\�qKe�֬Yj/8�b������N�l���h�:+�Vȗ���?���{Tq4zG�I�P�ǎw�_�t��� �����^�;�`Jf��k�^�f�C��'�s��J���wYC֬�1c��^�� �:�I۵��i;x�î��[v��K,�����[n��C��zE`=tZ����C��>Κ1����m�R�;c����.�� Q�:��A����~;x��
Ť=^��3�z�D& /k_*^
r9^:�@%K +x��+\Ѡ@�`�:`r�^Փ��[��X��a{wo�d*XU�.����'�)���ޖrΜ�/��~��w�&^�g���w�4LN�^Ԅ�f�� � 7 �}�Sn�����-]�@��W2S�K9�&�hY�R�̤��z?��z�����-����{��e��j{ (1N��Иj��9�ԓ�e;%[j�^χ�=�
���?��8���zO����;������ ���H;B����kd_�)T(q � �Y�J��}���x��w�޾�6]|��Gx'�>X<�b�|����g5����jW4u;�x{Jv`1�	P&��P���%s��;)�����Jm�V�^b�?�;y�����'m���6k�Y�m�b�A�Ū'|�H���Z����j�x�c7�ڇ�>u�L����s��0�0Jx&�R��ϒD�K:l����lŊy6u�$�����BE�*I�q����=��6�i�����u����.>p�e��[ Nk�߼e�{z�Ӏ�1d=ׂ�ꬕ+�k�bM�������wϝ�i]�r�==]��SM�u��:b�r�����.r��������I�t�r*2��v�%�A��h��i"^�R��v�x̺��z	
� Z����t6z�Vk�h�"�3w�s��:��_)� ���I�A�,T~�"����lϳ�X!�: ��.e@*�\���\+�	@5����� �&%?9�~��nط~A�5�'p�3Wb��Zt�VO���X�ܯ��h��4.��K�(J�d�k�X
 �3���g�������pmx-����XR���Y�Q9�!��>ʑP�-4���1c��9'@�5J��R@����� 8cZ���?~�����&��H��Ϙ,
����h���N^��_��=p�,��VZ2�j_�z<&N�yα	�g: �C.	��D��D�% �?�2	�֗��dhlø#���Ž��c�|b���!����c�����b^��ҙ��ݷ��w�_*F�J���iu�����U��� %�@�홝;�ٌd�������_���~$�'��@]�t���~�*�A��;f���U���-�(��C�^��C��y���Z�Z���g����6zEJ&�� "V�^:?���I�$���䤙|���0A�(�������jǏ���������K��V�V2�4��t$�t�Yͻ�-��_��{*��k�v�zB�Aq���J��W� ��7�&)��ǩ�(IJܴ&���kW�W�e(p�'V1ϟg+�M��.���7ā�� �R�7�=��^ �u ���s~�'���iw}����u���&�/%�AaQ�=q��C��/���
���g�;��' U�`�B�Op�hX\�<���Pw,4,.3����q-HCG��Y���P2caN��;���KGa{��?���\7�� ��{�_�����i��Ӟ�5`��.�u�V���Z0�bi7q�e'Z63��.\l�Dƻy�H��:�hL��;��En��a����~���Q��������;O�4����-����]v׿��F&����{�b��Z�P���n���$;�v��{�?�J$�r@/�ݿo��3#����~�-'��t��9:�G2���'؟��y-�L&fw��5[��L����4�Vн�VM[_o�Z[�Y_�:��v���}5g��+c!��y�v���p�X����#L�%˖�%Ǥ����'���k��y�+���[��m��K�,c��7j�qaSm��N���G��)� �Zd���hI^Rp=^_<�:�Q�A�l .�τUr��tU?���J}kC�� 3�����A0y�K �v��n���@&zH�E.�ߎ��f{BD��[y&m�L���ST	���y�,�sX d��3����8�8}QW�^-,</>���#cDIO�PP�= ��P=�G�t�{#hK��uk�V�<<��<c/}��\����ze��3�ga�������o�UW��v ��?ng�\��@_�_������PG���3�S�$ׅ���_F�F����?j�dS1/�p����a��V)S�'��3$<��Kem\�D�p�ž ���&"����X�c4��'<N��/�ߺ��.@`� �g<d�~%��%:`�C�}�uw���i�N��q	g�}��/=a[��D�юu�lٲ���o|�Wm?��ϲ�H�s�� <�
�}N[��rOo�5#Y���2Y������k�s���-�(Y>�c�����e���LZ{�1k9�a���]�~�Ox&�*�r� �,� V��) ų���z�5��f"�J�+`�`%ԫ}F��#͖��,�1��u��ke�;����;N��e��/=|�J��fd�g��A�@8��]���� `���}q,I�ا�W��z�XT�J7��?E��L$a���(��}�p���H��[uQ�e-(|�8�hyql�~,`��⟵���!�h��`�����t�1��la�S��\��L��3Bm�3c�I1r�w<L�	),V+�`qs�LxD��.q�ߑ�@����}<+%)�W"�}��@��(����9�#��|���'�u�E��	�s�:?Q\1WD�`(��G�?���p��IXn��6n<�.8��}.�z&�]��U�)ˤ�s�Eό�{�^껇�����n�����qp�����]>G%&��ȳ��"�Q���=r��j%o�>m���HV����/b�4%-kv�h�5h��#���׽��]�֟ŝw��^�H�^������vǭw|����O��F������s�J{ӛ�h�j�*ł5��}{wz5O:��=�#��r�j=}�6}�"������PP�0�Eo����pR��A��2q�wדg��T\B$�N�T����	���
Sg春�p�Tm+�O&	�M�&[��#�u�;ޝ�Z?��f۲���*.$����җ�4��s/Ǿ��<���Tő��JR\���x,I,�ƢW�5��Q������U�< �X�Pyj�V��%/�-���5�/����i.spc,�47��.�l�_5� @Q5���m��F=D�`�J�����򈤢��&�a�g������έ��/����L��e��\���[s�7;�Y:��{��)��Z>_��	�-��X��={f�{�Y����<��cV�e0���e/}�{4ܣbP,N�w�������� 7�Z)X��xd�7EJ��
0x�i��K���k�T�]v�+���,���v�w=&�4~¨/�����?r'/+�X(���dMM��7�ٖ-[�u�a\�~j�g�>x��ʅA�t�B[�f�-;k�uu��D�7+�8I��ݨ�8���bB�
���:�k��+�í�:��y+7e���C��eqf�@Y@��i���5�B�xͥq����Ŋ:�c����_�Q Ɓ�J�~�,}��Jn+M��U}(Qr�)�p����+�l o��@ � B����j��n��nbN@�a�@7�v�;�AX�쫚F�2�M&�
}���L�;�ʊ����y*���o4�w�'��b1gMM	ה�� �{2���Ǜ9e�91h�Z�-j�`�s���Q��8S��jN�U����_��1<}�J��ŋ�Y�R���G�g�v��<J�'����Xn��]`��&o���Νv�Wi�EU��˿蜧5�o޲��{z^?���A���6A�3��3,��Oˁ����a�r��Qyoά�6k�\+US�8n�[Gdh�ؖ�@���ѷ�V  9'.9|,�����p��s�d+�7���ܼ���v��ak���L�EI�1c��+�c�e]�F!������ٳ�����\�,�_h���A���׌Sh@�PG0� l� �
Œ�Øb�3�P����L�|���Ǌ���)!��Ʊ��}�    IDATd��3( ��İ��U<�le<���ù�sa��	��"�˜!&�, �$u�D�wά���'(�V��8�}K&ʖL�l07�q�b��U�����d�r��ͯ�T��K(P��A8j��"������e����K�͛�h.�u���dA�3���빱p2�7����	�m��&��hs�Tow���y��p�*X �v�-c���_[{�W
�Li�<�Nk�r˕�����G��w�R��8m���nx�M�2q��T:�rp��8�b�W�����\+_�=q���FH~�}�IU>���KC�OQ����/�=��ּo��ckjL�@H)GFa�={ۮ����������,���&U����_�q�}d�364���+ �$hȮ`3c��R9 '���n�ɍ�N5�H������C����!@����>�+�CX��`�X�ϖ)ٹc���5�qCG�m)���I1?�@)fS�aQ]R�)����Ϝc�z����n��B�l���v��K�j�ު�bE =��gΘo���׽�s,Ny��d= �M�
�>G�����R�7_�V{٥���"o�k�:QAAeW�9�]_�}Ӧ��W��M�8ޚ��=������;�=��*�g���]{��-u���V��
ӧN{�i��9�埈k�I�Ʉ���7a�xzQ ŭ��D1Şsv׏�vK�~�,�X����[IxA�̠Ɗ���2�ؼp�1b��8J=�������ÛTSԍ��Ɔ�[X(V����~�����4�F�������w�������w4�7�lKD��ĪG#KRk�)����θ����PQ&v>jdþ,���>�O���� ���9�Z��k�W�q��^T�T�q��it�*����?�w�aI��
A�#`��QI�[�ϭ�Op7?�kk�[a�6��Ze�j�UJ9$<V��l��i�f���ן��x<.J>S��8�;��٧����3����߱��\ڍ����9F!:h6���ޕ��w������gKsY�	�%�Ugj�������:ފ2�k:ʍ��QhdS"�ͩ��
Or���x�R_�\�[xJ�����U���^�X�r5>�w��f����/�8~�%Q��!����~ ������]��Ԑ�d����Z�&O�a�w�;|���2^�%Ȃ��NYc���Ͽܽђ>@A� �C)�\X��we3��A��Po��Fߗ��#� f�U�o�Cy�Mݤ'�x������Ko�tz�H����]��M�<GEtǠ�%	I��E��C�t�2�z{{���O�
�# [Dȣ1�؎E�Le��� z5s)נG�����e�ןe]x��}������U�I+�)�7��n��-��>b��������K6��9-����ɖ-Y�^W�ҌA�*����爸$��y���z����&M��m���m���~�۾��t����à���{�0u���{�m_;y��:�o����a$ڇ��In�/���χ��^ld��ł�=n|hP�T��g���g�a�A��EF�/^8ٗL&0A3,;t�X|(%+�a8�?�붣GZWW��u
�T������.����>cV,T��3�r��NA�i��>�\�G���� ��3�c��&"��J�%H�$ aٓ�Ż���[(E�( zz����F���L#C���F���#m���,]�؟8���N����u���f��Xx�7d�/@!�9�^��zw�(ܛ��p���}�h�o���]�ܥ�I�?m˥�%��mʴ�6q�6u�l�x�Ű��U$�<W��p���_�B腲m�t�]w�[\�D�B�c��k����T]&)��d�޸=HxQ��B��,޾�^����8NC6����YG����X�V�O�>��;n���s>�=��ӨŇ�������+��O |�{h���Ui��cM�	�y�*�'����PJo{��<Y�	"����8zsg���K.۳w�l�ci��5ҵ+f�-�v���@�!��4v\R��5*�h�_,<�r��{V� �]C4���
P5R�0�@�` ���ᝳ?��{d�����V6��ˌ���Q�A�@]Я�r~���&su���A���m����!����9�z�=�}Y����#*U�^ݓ��|�袋�f.Á���s�]bm\�%�)�H�V:3�.>צ͜�u�JU�� �Hy"�'yEy,T�$�듟��Z���0���?�C�Kt��xv�R�@��˳�=`4��;������a1�ܳʐC�])�ĩa2\v�� ����Sq�/h�8��Fo�`�EE�"-���x�dM2y���O�#� ��=Ǻ��Ο	�d���YC*i�b�R�=vؚ�m��`�/T��7�������T,A�o-�nՓ�<��>�k��Ac�?i#�O�7��L����"D% �ÄfxY t�P<:�<	�m۷{�0�' ��l��>ۏ�}��ӄĵ��2����#���k�������V�^�F���G�g�>x&j��v2���`�?��J����͘�6��[��x�b���[��9w��SU/���x�Y�h�Z˗0�2f���d
'���)�h�nN�,��������k|��dqkjhp��8��uq�м,�F.�� 	��àO,h��GH<�>p�ӦO�����O���WC��?XQ-���>'�?�(E��cM��S�f@��M�H&��Vw&21QV0iFj�k)�,�IXS6fmͶw�V���9H`iii����r���' �MM������g�M�集
�R�@���ˇ�i�9��rI�b%3��� Q5O7�zD��*�xa�3V��?��%xw�I ��A�'��A��5r}���#g?U����b"��}@k@y��T
פ�o5�q��lq��^؍���f�zB���yk����˽��}@ۅ�δ�γB9$m�jP>)W�d���[�fNd}ui�O}�Ӯ�w=?%�*�ސ���l�G��u�<���,D;ɲ�1�^�e�{{z^7��_�h�jH��S��:�w���y�b��X`\`�9$e�äQ���n=�:&�Aޚ��{��J���"���J:?d���	�f.�梪 �<F���������󢪍� &F����82��� b��f���j�˂�*�e�Ŋ�q��1�����R�c��/-���5��kb��9�x
[�|�&F%�|��O�Խ����	>��I�+���E^F
s��(~W�!�9s��U�<�Ua�lM�[�֮4��:�SΘm˖o�L���-Rޝ���ۆ���%T,��{�ֶC�ٿ�,��bL<�P�d���r�(F#�&>G��O�8�� j!;�9Nw��;==��}a�����q��G-�ݯ�h�l3a�S���	,��ކ��U��D�z{�[_�u��Xww��#��-��v/�ݢf.���cD��⎁����5۠�/���2���]��ϻ5�A�hJy���Ϙ�8.��sw^���<	�r\��0�j����� {�(�r-c[Mdؗ�p�x'�cK�/V=�\��U�f?ߑ�����:ߋ#�~� �[��o�?��:Q��|�]x�9v���Z����x����>c�M�6߲��4N�B������s*����v��_}�
Q������K�+�K�bj�=*3S/�74���TOp��_��� �#�8,	ύ��~�Gp�Qd�);W�
c�KcA�Ť�����H=�X�i���f/�L[8�QjU�L������9m���#�왡�`T�v����?a�_=�cq׃?�E@I!ۡ��~�; %�q�ō���
Ń��lT�)���u�b1��(v���B�*�5J^T/�"�����!�W�R�;*�W)��Iu�D ��y~G�I��\�ߓ���������S6��a�
۰�\�T,���Ӻ�h�����V�m�}��P%���뱱Z�z�����?�s/��s�e$*�������Y��Kp��8��:y[���~M<�8#��u��~�7��O�	����?/��	�	��9y��M�ădo��*����:�8dmx�#}be��4:�V+)��l2d����0�Z��]���W�VP��?�\/]�����ON]�z�5M=�C숚0d�:hᡂX�
�dT�w��'?�I��_UQ�i�"�KZJ-@��2b|J�L�d�q��|Ϣ��,>��1�@U�gScP��XD���Ăǵ��S�d��x�������[����U+��mݚ��s��a"Q��W�	/�R��m℩v�K^扑P?(�<W���Я�q���J*��� ����<s� )|FYw=#�-C���Q^G0>��"8�;n����Qi��_��
�ؓ���xl����Rɪ�U ��B�8��� `��j��J�L��R��j%�V󖌺a�g2m�f�����l�R1���^�(8c���	�����>�B��,jh�C��G=�g\�DH��Ģ3�yM�9s�G?��� ��t��\��e؇r�xxT�e�����g�{�g(���8 ���F�-�	E�ꇅd0�?$v�����im����4�q��\gϜ�
�� �TUO���&V��m͹Km��gӧ�ɚ�g0���\��,Y��ZjF 8����[���|�;߶� �er����Ӟ�v�~G�GGY'�.�8��<�>����0����N�~�wo���O�濽���|�K�Ї(�@������Z[�ڑ�W���;��L��R�y�ZD���D3Ed�{�1 ?g�֘IX�4�HH�'R���ޢ=��6�Xƕ�R�-Yl�����Β�����&�#g�� /T6/�.�'W.�A�( ��Ή:��/2QJ%3�<}j�6���>�5��h��泟�ĳ�	�B���'@�<�*����8@�)>`�J��liJ?s�|��͟��,Z�9ǎ���-Y��ҍ��:	�C� ��c�P�͚��s��k ��j�����p�;k��P�V��,�t.��۝v�����~D��'��'���=P���l��[-z��x��>�/��)��܋�BA�u��[&��� �L����+7o�VOo���|�V��54f,ח�j�&��uM'3�
��i��fuB�����ِXLLJE��sTkE��+�<U*T��x�6����'��9f���V)�)`Ԝ�,W�)�,NF �A-n�.��s�vq�S|���:$9Tp���r�)J�׬d�_Mh�տ* F�H� �s��l���7Nd)��T^	�C�|�!���`��}��c�(���7��M�|�9�dYTH.���Ch�hu�W��NU攬��J��C�������?�����"+�������k�xUO,�Pճ��[�f?@���V)3��r������M�5T��S�[n��ٌ?��ɤ�ko�굽h����\�/u��� ���}�S���� ��5G<_.xŀr��� �΢LǼ��;�rȪU����`(I�ChH3�紶�GO�%��j^��R �d<e�]�R�;g͚��D�]R���b����� <���pl���冻����RkA&�5���C=�t"�T��;����l�\o�%1KE�Y��L���~���4�f�'l޼C5R�����I^����=�3������>��Ɉ�x�_}��սB%�i��JU�D*�ႊ/Z�e��y�O<���a�w��.6 Q�3���M�8��А�_)�d�B}�������F�-�xy�{�;$��PB� ��Y.�Г�8�k�
�˸Vj�qȠ`,O�:���s��	���P#��ڄ	Y;c�xKF�J�B��b%���[`/{��f�z�X
��q&�F����t� ���T&��	�x0ڔנX�EmK�Y�P�!es�Rq�l;�앎3fd�!���7`;w����l6m�R��r}��~#Nk�r˖Q���p��usή����y����'O����ϼ�C�����(����i���z�������D��FI^���5�k$��'|�l{vo��{�ZB�M9����T�|f�>{��m��M㖬��;g�-Z�0���b$����M�uY�xp��p�yNyB��ū�>/�	8������s��P�����ࣨDIe���ܵ���n鲅������;�UvA9c�����[�h$,S�%X�x��G>2T �kW�k;�:�Cc�{Q�,�(��w��]�HhA#>k�[�p~���퓌�N^_Tm��œ%[y�"[�z�{�rɒ� �4aǘ�4i�m��+㖈g��o2jd�blE��찏�|�{|�����k��z1�H
ʜ��G4\}�r	.��R���mΜ�^��Z-{��kjj
yh>X`����8�U(���T9*�=� ;����ͷ�t��i$�-jw'�Y*�����W��[:2�r��^%�h�;����O%A�ep�t�'�����A4iy�������+eȜ�J�����^�:.���������'��6�f� )��2��Fk9p���!���[&KY�͝7�� �.X5�s����������n�C�!X��5�d��A^4��;�6���+�:E����=`-�d���J��������c���a�(XI�h��D�W�,U;�Ia�����իz?�C�� �9�K,W΁�c:�V�7d�3�Pq>-Ķ��\%OX�Tϟ�>sf���z��r��֯[i]�֬�w�'�(�X� 64N��7\��o��P�Y�3��vx��ԧl0?���^L���8�X�'`�G4�(-l��+^��v�K/�d�R,dq����~2�T��=r=�rr���1=��\!gY�Y��?�W]��+��=o1�KE��)o�r��+�寸�z��z��c�;���O?��4M���sV���o�q&{���R��LQ;��XT
�s�Ԁ?�1Oaokuݶt�X������;P��С�ֲ�U���(nc�ۻ�m��O*M ��<���#p	�U���e�SٝJ�g0�z+d�X$FRA��x�3�:�S@ �PGG��h�W�,��� ��w��k��G=�K��:(�DUZ�	�sϪxn��f� :�?��O|���:������+�Я���b�@f���y�{���.��8 j%Ā?qU�9�S���D'�@�b��X�{�!����q[��L۸q�����W=�Z�ĬTIZ���I����.�rm?}|�ޛt�-�,�RZ�����+(m����K/���Z���ډͰp1Wd$�w��K.��z�o���J���ჶ{�km=d{����x�2[�t�-X�ĦN�IPK�����py���S���:�����v$�'��I��5kV�u׾��zl\cʛ��w��F�L��'��JO�\�
%���앶x�
�\H�ԜEY�L`$Ȑ���CC�[n�ś8��-o�^��eM`�SO��H�hW��9ܺϊ�ǭ����./�J5���mv���Ya��/���m��%6�l�Jb	��4�*p�:!����� rq喳���LX���G������f<�A�99�+��h
�!��{��?�f{G�, 	��$� x�y��\�V����Զ'}�R���BQ3$�\=��0d��/@H	
��P�;�g[>�}�˸b�q}����%m6c���|O�H�J%)��kk׮���W�%9+�l�3�-�Lv��3M6c�\,Z�`p,�^�i� ?���t�v�H{�;���hx)\���h��s�])�':�wB<d��q��gv��n��ͪEK7d�!��\>����	S�׮x�M�1�E���Wo��:;)�w*˿Z�>u���e���-�����s�H�IC��7�卶t�|ˤ��Ҽ�J圵j���nO��S"��.Y��{,W0L�;���>�$�Pޕ�����?��ݪbB�!�]�U|��x�r&&ނ,�z����h\�l"c�Z�b�۳o�:�-I]F�������m0t�( �9�C��e���^|-
�LLx\]^
�62��    IDAT)�~>��[^��ƌ�� 2H=�(� {���3^X��,7�|�?T,�_� cE�)�鱦q���0��Sr�cqn�	 �o.�.�?��<lG2�T;�6~�lG�K�$rn	*�RK��@�cɰ��Nr��^�YI^!˶��$��D���3g�V-�������Oٔ)Sfۜ�l��Y�;��К��\�`�����B���s}��G}�p�Ϛ��$Ç8���L(�{���X�R��Zﳖ�v����k�X�\�*�:��*��3`�J�~�^ms��̦bw|�{���ĩ��-�jq��iם�U=7o�bOo����}�M�b���7ؔIM�L���߿��\��K&:�<�-&D���6�׬�Xɮ���p�&����ʇ����qH�-��ʾ��/����E�B&�it�gܬ�kZ��l�� ]@��a���Y�<��Fk����1���@��X"fK�-�ӧX�B�PO|4�_*�MLZx]�E�� �	��k��?@C*�1�O �!���W�@�<C!z������\<���, �&���/�=���|q(��3��L�c����;��qh
�V�����".�^J5z�b���s}�A�ߡ��XCn�)����e��"2v$�4�<�-�)���騼�WC�
���r�f�2���s�F"d<��Y��L���<��-_��E�]���"�z�s�>������&���?q�,��' ��w�.��?�q��p�)X���m{�^K���>|�r�3 ���í�֟+��`ͮ��7m�y-��؃?}�n���!I�H#,j�~����+����{ð�O8�lz�2{���n�b�Y�h�����K.���B�k��:�&����m�uX�����}�h�
w�x�j��B3��Q3������2���Y|�!��1X̸��h� ���Qy�ᥞqK[��ʃ�M��%����`��R�X��w�p-��%K��i��Z�I$#�?��kf�cyj1�u� �[Dfn��H��ol��'��d|1f	��H.[� ��6xdu��c�d�m��$��.ՖȌe���� �l��N W	d=�U`��9����A�qY8(E���������op�d�K3Ͻ{eT�_����F��T�_�تs�؅���E�Vڂ%묯��|��QD�0�jV3J��	ć�|������
���44��ʜ��	p�k,d�Y ����v���k������w�[�l���h�-���<{��W�kw���nhN�6׮�������<������7�w�g%*p�G�X-��,^do���J9gG:�O���]t�:ˤc�ܼϺ����N5Z{{��,�h{���k/p���!���Sn!/��c1`v����,g^��s	(U��p�O%_��q)�{l_�6;ұכ��h41n���y���	�Ƭ\�[�Ry��5�KU�$����j-�&$�- �1��/n�I���ǳTޅ��#�@��ի�k �xW�?���G��]%�i!����'�!�?5�1t�E�w�=�`_��j��,V|ǘ��e�3 #���^ƍ(%�˼`�S������v;��ɤV)����K��ɂ�x3h�E��;�S*�J�l�������
R�[�\�_�xc �Z������#�g��'/�6�������@E<)��]��kw���v��sl�����������;h;w�l�dk=|�*��}�C��K|�o>c{�����ؕ�Y��)U.����J�~;��a��/�`/\g�B�;��	L��%����n���m��|�*��UW�}�{ߐBCV>3�f�r�X8X>߾�;���HT�� ���p2��|�FI�����юfk��g��#8U.��4Xs�ѡ�/��ր�,/ i�W��(	�[t~BC�09�������H#�?������L� `�2� fx}������E���w˾�U�vޥ�����{}�R�����'s��{?��@/�P �ԩ��`,b�
�]�{M!�
Y4���!�,����ˁNT�<��Py�(���o"^�b��֭;�6]��9�|+����ON�e�W�5�ĳKZ*�`�\�
v�P���'>����V�<ө7����@"��C���K�Ƶ1���b�o�������s�^lS�N����T��d!_��{Z�\IX�^�TR�я��������ܼ�KL(��>��l�o'��e�L�2�>��?�Rq�R���v�7l��U�y��փ^���?�tο����Ÿ�i9f�6]����kM@V�5�U7���7�n��@D�`yPPj��[Ա�57?cm���ԓ�.�(Y�"�Z$i;p��ԓ ����A�|*�'�%Ǌ��U@˟=E#���(����� �����qw>���ƫ�3�/e��r�ԱFh@���>���fl�p�, +`��z����?� �j�����[�@
G��)����˳y��}�f�6@kB�
�#��sqN5p�����4~J�gSc�����V�E�y�ԓ��J-m�M��i�d;���V(�,fiK$�<���ϸR�8������7W������%�Ur��ϝE<�tv���?�|�\k�fl���n8�����\�v��o�x֎w،Y���kǛ���:p��-��8O�����n��m�}���߾�ە�7���皑�>h�����h�_�-�?�j��=��}6�����`_xў�D���l9h�����]w]�����C�#���G��d��gR�s&�{��׹��-�?,(	8�H%���쩧���foW�M'���Ja��	z�v���<hǻ����=���z��8��8QG��:	�"Їw*�s#�`� :�Dy��~���=	EX�H/���*�ޱ�6�S d��R��&���]���O�'�:��O7.���E��wj5�1X$X��s P�]��(s���i�GM�J%cV��_{�'yŬ`U�7$wR�N��K_a�Z��unt�X��ڇ�\�Go��3qy.h x��_�5b)�7�����~N��G�w�0�bǺ�Q[T`qj=�i�]��~���k�`�7\�E�ܺ;��o<'�o�A�?}��n���[N?��r������e$��lX���]�Mv�k_k}�]� h�mmV*Z&s�����~/�0q����W�����V(E���o�;n6�~Ǫ�A�U�� �.#:a���z���E��re����b��sO!1e����b�<��-*b&̛� ��%�p�r�#���)��U����*E��$Y�����g�i8�
t�/�MI� �(�>@�"�o��+I^�Y$��*����0N����2FQ��v�w��E���)�E����N�`'�㆘eh<�c>@��!p^<%��1^��s�Z�	w,Q���Zb�֞c�t�*ł%��n��9e�6s�W�T+�ư�Qǅ�8���˾���9�so�L�ʰ�s�����S�#۰�bPʥ�#v��>��hsj���R%����H5X�T�;�Y2�`�����S�{ىo~�[�ӟ>4��)�v�������t�y$�@�/�\qk捿�z�3w�M�`--{m�Χ�ۭ��{(U�K�Y�m�s-�j�����N��Kd3 x�b�o�8��������@F�dU+<�QGh�^v�*�56em|R��%"���$���Y�N��Q�ki�|2|�zEQ�ꑤ��3��=�p����τ�?��Á?�*�1h��-����1E���0��'��z�� ٗE�W�I��%����3�n���߹�[N�`�(X,%��������@[��)��?�#��8��L���;�4*�2�K
�z;�9�ς���ȅ�&Mj��&{UO/�Xt*��05����T&�4Y���c�]In0���Ɛ����3���:���-���	�f���Rgh\6iG:Z�8���;�����^8C=�����%�^fM�B������/���	���- ���mw�z�WO?���>^ځ�?��^�y筱�_�?��?���zmǎ�]�s��O��d�̚� �R̃��H��%��ÝE����o}k��?�4z����?��?��L&ܠ�����?\�77�k��X�T�$��(Z��)�ʖ�d�>�%�F�^������j�Q����_��M�ZU%�>
62�Ƥ�?������v�n�±������^x?P����{
��E� +@�g�ƍC�d��J`c1�P�*���n���;h#�9 �𦼁<Z����������Ϙq��ba9C�2W 9�sB�: |����I%�CU�t*���>������:}W�%~=.�%K�yrd� �<�RԎ�gt��a��_�eμپ�>��%ܻ!��c�!ཽ���y�HZD=zĽ�'�|��Cpl�˯Y���=w�M�8œL)�����ǝ���t=aQ�$�1�$M
�8���T�/�d��f�&M�	��Z|����n��
�H�����>ॺ8r��ċb03�xXE�_�YX�d��
ϯ���`��m�3��b��~�R����
�Wl�S;�)�b��*D�����$��(�� I�	񏴃�B��`5�� {��6��O@�Z@Ř�l����h�js9o�5�v�\�9- �D�
�R��*�'ޞ�]��Ї>�/Zs>��Cm�c<��p�,
@ �x��P�?�$I�i�H�/c
��j$�
�k�܇J���Ϟ17�}�'qkkk?��1i��?g�$[�p�UJ�fR�P�͛�{����W���L�T�L���.X�Qt-�W�5&Bc�8��x2�B���/�`	�=�1O$��MQ���\�%j<�����$�
100�`WO�3�|X�K���7�s������-�e3Pqu	� {�ej��w:�,2q,fl+��Fݐ��=�)4�*U���X;z&��%����ޡV�];�c��<�Db
@R�/�g�a{��^���>��͎���9O����
p���ͽ��[�'���;T5��0��?���ͻ'Y D��0�G<3���w��|�� 8�� ˛y�1�'��Up�xrP�Gq<��}�W��@P���W�wE�n��ÜQ�"2��:��Mg@s�>G�mBL�RW�y8��k|�6h�Zf�_mF�R�X"��$ǁ���k�lm�Ԭ��B	�Z��嚢��2��_�����Qo�y}��/�o�>扏0���
/H
 ����3\��c`NJA�*�2Hهg�������JMwZ���-������Ƒ�J<�1Ȕ.���dnP&/������->�^kؓ��2�M�'��ŢW�� �%�TUO��F����3+ێg���P*��Y&��~�P���Q/�Lc5���._�$<Y��OF���k��^|X���\7�/W&E�d���y��7������ċ�nx��HOJ�y���&y%t%�_�+�|��R���U�Y'=� 0���1��X�(�THF��J�
Us�1$�Bu�6� |�L�W*��E�%�W}!�����چ,�����β��g�b>��wN���Ujq7�[{�7�
�@������y<^�Q,:<G����s���<&�8���Y��>�яz��W�A�<+B<8�����3��𼠿XP�����d�c�?
F�
�UISJ)%���jG��s*���ZH���AY�|��h�نA�W@�Z�u�	��*�'��Xaox���4�8ٵ;ةZWW���{z:��U:��������w�O�y��b��-^��fϙZ�UF���LV=i�%'T"�\�z�y��' �V�, ȭϺ�������"eч��pT�$8q (G@� c%�L>�ˈ#0�⃪�0��4�G���ƈ
�i�H&�W�.�"���o|�ϋ�EP`9]ŠU��/�|^�W�7��%�CUφlҊyJ�������Z]�>V1yz�O�4�Θ:�/^:y�)�q��>$-66f=��2����н��w�*j')9��j� �澸O����IU�ERυg� .�=F�:��^��H
���P��JӧN��4�z���K@%i#��˲R�h���|��>�C��,��n��i!�K�Ë��L�b�xSVw4�cB�`�H�y���\*�-V+Z__�<�ú�[-�E�@�Ѥ:�e?��a��H����-�g�fOwz(^K�j�s��X5xUp��&`�*�� դ?�e��A����eA,�n�
���$�D�;�� ���Bg����{�2/�`̊Ҕg��\΍�1������,M
����;D���3��x%|8��Ca�V�N^�U=U�٬X����t�rܪ��%bY�5�L�4y�54��L��
%4��~PBC�[Ro<ݛo�Kf�ӷ��Z�0i�'�a���H���ûG����_�Ǭ���L���^f��,m%~1�����j����������#�<|�i�Ղ ��� �@�`��~y���$��!@�Ń�G�n3����眀?n#�q��[�qo�ސa ����Xs�6��h������;CU�\�b� ��ϵ9s�[ie���*�~Z�4�����;��k��P>����C�/�%�幊g,�D����AF��V�!N����ƽ��Z�%ٔU�1D����ǖ�,�EsPF�"���b�x6m�<T�M�ζ
rj���=Q��,OEU=CI��4%ɻ��ϱ��?Ǫ����9�;g�^`����Tz�W�-�V$^���{�*������O9��
������|�	�X�h�U�n�h;C�.�AϙsS�D���/�N����2�O��W���)e��B�W�/\�.^�"��Lhd�������Y˒���-�4�xMx=h�D��;����IKO�[oO������>�S��w����'��b�x谵t�"�3w�U������g�
xVr�5����+��|�O�J>�
���>��{��� HW?��g��ƶ ���q���b�y����U�K��~
��#/�G�D�Z�W�2�D%�k�˜k����Hj29�P=�J)�}NJ:��a���a�ٖL�Ӄ�l�|�*�:s���d�s����H� ��<����3_[�a���}th�s}����
��QZ�1�Ƚ@�To�K�g�g�©F:||���UKގ�������M�z���?EwM���������{��]������ٚm)�R�Bh�iIDEE@D=��S�v��;˝�������"-	M@J	%=�������g~����g��eg7!	p�/^����Oy��y+
/?��4[nHic�nt]j'��Uf5��aM�N9�\@�� w:@l:!k������+�d ��;�c��L˺\�@��ƣ�-EG�Yˮ���?bd�U��D��W�o_��&��q�1P���������\9�����K��AZ�\RH��z�=�G�,;eq�:��\~<֛�#���La�tMi�^���w5�rƿ�y��|7��9�����!˘�ƌ0m�1���H��4Ǝ��c&��D7�`"���L���η.>�hU��c���+ĭ@�����r�����%4�����+��!���z�o�Ĺ���_�O�s���b��kim�����g��_B����
�� �ߵ�\ʙ�d�b^K�T�F͞��c0}���$0��Lw�:y�N��G � `qa�{'�/�+��ͨ�9�#�X�~��e�ǳV"�g=��7n����n��O�lZ/|~�����C7�+��G?F�<�2�Hu�J�R��7o�|��	�.��8q���-��;����m�ē��r���g2�T�Z:t��7�+�c왑6b7�Dp��(�,����� �����u�x���0�F` ��4-2���T�沎���5��w�)�OO���D���`�UW]�g��>����زy�ݻ�ݽ����Ne՘�葿Z'�@0
zy�Aq�V�Z�Jf,��9��Q8ɿ*��/�3�F�Ў����-��M�g�-r�PUgvЏ�3��S1�e:1c���1�D!��.�E�4"V݈��&6�    IDAT1�(+���l�p<��+s�y��i޹RKU����,k��x����R.������P�/5p|�n�zj����+-_�kZ���埓�HDҚ��f��ڠ�!��Kn�~�ݐÆ���m�J�}�D
ȧ�uTU7`��Mx��g���ΰ-]�ʍ�EC)9����R|>��[�v�]mh^��څ�
_��&Rq�T'`nݺ�������E6݁3'�S���O��"/�;}A�
Q�3E44�⤙���u�+M)�ƸX���mZ&�=͖^�[ɋ  *|����O�'�F�P<D��4�!�/�2�����|�L�S����ez	��wU�������_T�qoLA�C��XA��Cy�K�����|%kS�2	���g�ƭV�L��9�I�X�v�Pd�����ӳ�z����,�s�F�P�@߱#?�k�a��V����g��������i��=���'��O�fl�(0��3��"��aX�p+�"
�(3�`+��n$q1K��\�$�:ȏ�y�6V��4o5�SXB` �oni�~p��/���3jk-2oZ�I�B���r��l�
�޹�<_ח�Gn%	 Å�@/K�)������?�ً�h !���2�Y�C����6nي'�z��$Ba���p���1f�XdҎ(�ii,ء�G�
��:}h��v�Џi15*�����ػ7n�?ӧ��I��ǍǉӧXrD8��c*r��,�ٜz��5��+����c�f(ȇ�A��`v����H�6��x ^/^�{����'YR:KTV�>PПn�A����+e�w�V~6.,C�)3%�W1
�L4��*�#)�;p,3RE;��s"{��2�'p�e�_�p�u1�U��#�w��|���j$��رk7�T�Y�R`�Xv�:
�T�hXiL9��<��޹ۇt]lh�c�W?"!Ge�HvPkl���k�oτ@����$��#hjn@.������ѳ�s驝�Rɜ�|(���'];Ѩ#g����`��b?^��!JQ���tv5D�Λ�"W���4�
#p�e����"/i�^
N��i���J[J`e��xj�fJ��o���6y�
�tM�k�tHiJ�R���S)~��?)����N&��N�F�
WYos[�� �H!V"���#hjj���G�豣1��s0bD�-b�&�@G�������7~S`�����%1O�����r�e�oP>eA^��ٜ�1�Ҏn�����|��cu�ً�Q�8sYa[�q�- ���:
� � >�w�gT����}O�K�\b	�D��*{/�����`���x�����N��[
W&�᭭8��3��:�t��+-�i`X6L��u$n�D�P��ތ!	����{L�����a@�]]��gFO�˸ TU$�t�?\L)�"4o�SE:����k�{fΘn)r
R�`��,Z���v�!��"+��O��%�,K�x�����%ȿX阞�;R;��[�>�j��x�K�;�t�"38x��딿�wޏ�+��5��3��Vz�W_w��������RN��}l��4����Ǿ�ml�Ej�|�|i*Ϣާ�x�/���ۘ��|�����t��c<s{�g]�[��7��,�h�z�����wߋb!`����(��DCat'2�j����t�"�[�]��j�c����k��I�����5�� 8��;X<��q���G	���~N����>��!�����b�ݟE^�-�7J��܋L�t�����(䄾�k0m�q�1P�3��}o�ހM^���b-�T������|ģ��r�x}��e�9���(��ln���<�1�&q%���D����5�*�����{����ꫯ�s�������h-��4���f@2�s�������o,J>�6��������]>�t��b3�ѕ��3N�[=�'uD >��7(��u1h�̸#D�~��]3o~`�!��?l�� P(&m3�Ǎ&R1����#9ʡ�;��H#�A��n���Q�,��:�*<O�ŏb!_ dϗ�q���E����X�
pj����ek��Ϗ"��C�_4�y�	���2W�sW���S���Q��A�g��@��5*�2�.�r��vr�}�qN�
�f��h7?n�
șu����}d��d���B
���(�Jb�I
�5k��?]��_˥oz��t_ݟ�{��ʲeϛO���G��$`�u���<�����������u�7p�N�gL���^ U��woL�g��{Nq���8��_@??c�n��P���TWע;���K�3�i�%@K��>AG���5҃��?��������\����p���"��D0����²�F�le�y���	3����)S1|�([l�,�]�|�M
?�{��Pr����j��U%�O~�S��\ ��4P���'ٙ
*�i[���Ի`D~CUHrQ�r���]XR��~_+�+R+�
sA�cˋ�H&�6�Q�E�y f.8���,V/P0.j�N���Q��[��aaN��l��,'��;>��ʆ7��;>�}j����̆�.Y�
l6��X�h�)�%���6z(2�iS�dQ���&P��p�B��}���s��2�>���RiLl1�$`��������i��tPd!R>ւ�|V��/WcB���B1�N�0���=8ͱ�w���~nŜ�)�.�bP���kɕ�ci�X<���_����w�{�:��c	jn�l�*d�7��dZ5}Y�
���W�p̵_��A�We�]����u�x`*~׻�X���	��.{o(&�z ��^���fR���O௩�K9���w���a��عk��SScƏ���3N�~�������sK���O������:�ނy?��;n���,���8G�>��C���LC۲e�|�Q�;���0�����ο�ǉ3Nø�l�R@��G?*7s (35졇�x��i_�U>w�\9�L�,�O�� %�kA{ϯ�a5�8��6H�Ks����ٳվ��B*܆�a����5��!g-n �Ԇ��#	
�S{$�dm�>ט��:�l|SH r��M;��A;߹-r(�]@�.��.�Ի��&
�a�%����	rL�%�����/?r)���!�r-q|d�p,,�C?p0�xe
E
K�E�\|��ˢ�,�Hԏ|��K�_��~��s`��Y9� >Q�	U~���06W�sI:�Ɓ�E&�:�����
~�r�oB�ד
�s~ow������(���|�w�C�	�r-վ�/A!�GkQ�@�W�C��*��Ԟ�P9u�)Fa�����Q�����2�g�����g���n��I�Mwa붍xq�2�]�Y�c-��s�4kƑG���M�X]$���7��'�3}5��_0�����gZ��ITǪp���ٳ�J'��Վ�;6a�ڕ�XҜ%v����ޑDC����ך�g����g�d�YH3�.!���z �+'����ȇ��\���'��``��kj�Vֿ�x���M��9��,�ȣ������hf&����ȕ���g�,ɥ$�1A��1wF �l΁-�P0Rr�el3�	v��c	�sHf҈	�A��	������cڤ ��|�H0T�hx�Q d�����~ݿ$t|�����YՏ*ӈ�'��I�܉hU�	��6|���m�Fb�:��Y��C�e`�-����y}Z]�R�!��v���>��6�����|_�o�~:>G՜-�.����.}���o�G�����/o~(ʆ�xȚ���ۓ��������X�E�l
��*g�����4˂+Q�H����)�bj-���B��/�Ӂ��ͣ���ǐ�¢���g>��F�F��R5Y)Oz�����>S>?���5e>�B.G���ذn��چ*r�\&�5��b���v�L�s�F�Θ�/�+��)=Ͼ���1�����ߏw�o���S�rݼj����$��a4�U�ww�S��d"���6��&����۶�D2�Î])\r�[q�Ygوs�٨�����G$p���[���Z;"�Y ��w���hCie�@�/ ��UN����t����H�ՍƦZD��X~n�u����[�)u�+~�3��O],�@Е�s��s�s��;���Q����(Z��I'�� �pO�����\�֚�F��Ӊd"��a���]�W@�#Lh�K&��8] 4�0���sYz�z���6�;�C�lٺ�R[Z�͔D?���_&ldb<���	�g*�A$\���v�wU�0������%�3�``n!]
9���v���)�ڣ��khmѰ�P������u���;�mn5���F��b$�j�N���o��xI(Ïp��d�w�Ecc���e�0Ǎ�fKZ?���\�,�0v��_ l���xD�Ae%E)�Rp�n�Z?X�_�Ϸ��(��8��5Z4	>7��I'��/����g?kV�R��\<��<r�n��ғ�2��y�F��1���-�͛v"ѝFWg�]~f�<�((�)��寑+d�)B�m�q�n�_�����U_!h��Q�F�s�������v�0��S���ֶ��7�`��lټ�`5V�ۍ�Ǟ��~��f����]�(���G>�[lq�zR(�˿��� >����~��D*gn\o��P�}�9�����|s�<'�e�П�!�u>��[�@�B۷�㩿����{pͻ�j�'���R�r�_je��H����K�੿>�a��8��3Q[C��TbOp)�-L�n����~[6n�I�gb��1�{b_�B���{�X��R˪�d�YhF��T9�aAD����]���>�V��g�Css#�:�4C�
`�8�A:�3Mه4�LWdp�
�x��'�Pi⤣q���/cq(���A��OR� �q[ :;�x�'�Λ;��KY#ΏO!@߹��KMxؐ���������SO��L���5wV�*��P���}x~�Kv��SN��)cM ��a�@�IQ�_)S.��aǮ��랽����X<����8��	���o���;z?,����5F�C���s}�k_���>����Y�ϦM<�^����FMT��ɿ�c�D;���?b��ᨭ�F�Ƶ���0���JᕗW!k@[�5v>�w��^�;v첖�[�mvsPR�z5��_0�{������E��TL8f<>����V�Z�g��N<a��v�؆T�u��ՙD[�&���qL�|<>������I���B!S&ӹ����'�P0����C�Z���Be���J�/]��WҾ��M�.-���@��-"�9�~��Im�\6��/��IG �ڃb.m�j_>l�`A�b�B�y�`;vv��G�!���/��p��@�im�&�F�`�|h2S���kVo�#�=�au�p�[/E>w�}�8�R>f�d���?��#X���q��:�(�3=�{�=��.��L*��}��q\�΋P]4�`UU�4g��JUz�e_۷����?��#G��K�"_ �e-�)�r�&�g9dr��b@�����59n��v�t$��P`��#닙h08ZL�62�B��r���9gOGsK����Dssn�S*��*I>G�y�V�}ϟp�)'cƌL1��ǥ�z}�.5�M!�!��%�-�O<�3�:S���v H� A?_�b*�|ϴ��c��v,Z�8�	��yfS#�Z\����^% � �� +����-1� �����d	�%��#F��v�l��n^��L����-Ƨ����OE��?kּ�'�N�6MMðr�ˮ��AgWk�lB&�N|�����_Cu���.������+ʬ�ڻ�̟!���>Ǖ}��q���o4M�ޭ��Ow��9�M�ݲ��DW��#�Ύ֭k3�߰1�	��7-^��� ��M�� ����ċ;� � ��A�3!�23�߁}��\���Ո�ʄ���_�/�8��Y�8�� ��c<D���M�C0�3�~[�ua�%Ȥ�����Q��ȹwf:�e��4Sr�(׬m�c�=���:̟w1�$KrJ�����ӓF��j<��X�b5��9�?�l�U{�h�tG������,��YtttᲷ���z�I�O*�	�ְ���lX�>�c��/:��=�D�˅�D2�@$
�$�r�0��V<��X�v=��0	g�5��N��R�9b��~?��\���6�����~�aÚpڜ��:�� �RK��y�Ɲ��_1>�c6mڂ����8�sp��Lw�Ͼ/��K��{'��!�z,_�
�?��<�TL;a<ry���A��qə��4��wo
-z��.k=
��rZA�V��>�����Q�>�W�J%�����X)ۇ��~T�W�5�D��/Z[M�a;����wYV��X/�y�[�����N�3@W��5+���s��!d3�\��l ]�Y��E|埾�`�ʺ����?�굫LY�{�/�������@d���#F��|��e\��n��4�8 ����TPƢ����[�+D�qs��x
n��F����n/�2������6,\��x����9g��{�5��m�L+@���[�l���c�+8?�@)n�]���Z�3�8�=g6��X,�7��#�4ͬ�1�7RÆ�Y�ޓ£���T2��_~b�r�����ϥ�Q2߶T+^Y���|��:\�ˬ�]u. O͛�T
�]J��F��ú�m�5�$?}�{}�s'���'�s�JK>C|o����i\z�h���=�����/C6�|�e�h۰�-�*��r��"�NWe�u�.����g�o7���X��q�_�f.�c��|�k�1�KQ�b1��N��f:+5�?���w���0�1�r�-K�.'
�_v�"	 �>֮Y�|��~�N�Z��;����Rx�o�G�2�=�|�
K��h�������cǘ_��DP�G�>�y�|��?Sx���ٓ��E�ބ�e0��;�̨W����װ�����J�+�{*��
��J�KqM�'�?�f�2w�ҥK�eFk��t٩����i����	ذa�~�^�7�����/ K~.�zC�wc��G�c[5����'>���aX�n#~{�-�M���R��b�����A��e �`J�>������z��]x���8rT���]�{M������љ�捛�i��j/����5r�Pkb^��f�?>^y�#l���W��c�a��ٸ��������M �8L�
�-i�}��p���bx��U��3�.�ɓ�@0�u�UV.����o �?ņ�x�ѥ�z�;.B4l��������X�ڳӹ(~0E�P����.A(\�K.��/�p���L��.64<�ebVK��۫�x�_�~�F��'Ok���"M"/�P[_�\&��D���5�"�L��������s�%� VC-�Yg�nT�� ��a�0RE��*{��X���3;����ٵ˄K0A6�<�����ۑ�&QS]o.��x�<�֬^�Y��a��V���teutbյ��l7������*��;���=6�����OPW?��2�v�4����~��]���?`ƌ�s�$:��]�1���z�5$)+��T�a�O��4������ǌBw��(��6!���+�D��h�hG
�0v�N��+���E.�L(�]q_��G�sޥ��@�k�B��ʖ7[HnQ���������R;ŧ�=̿�׮]kץ��Һ�3�O}]�~�>�.��`ێ-�%M7�ջ�CX��{�ص���}�1���Z�v�e����^�=o��/5J3�|>\r�[p�y� �����e�b������2��>�5u���@ۖ����_�N���~��X掸��կb���fR�8����$��1����shp�H�e��.�/ҫ����`��-XH��gҤ1Ȧ]Jlk��6����G�Y��w�!W̠:V��;�X��Id3�u�y�U�H�hEZ��Z1z�K�?�^�;�	�PUU��k���Ï���W]�6�	�|Y�=b�}�Q�ݳq�F�m���mZT8T���[�5k�aΙ�b��#-x�L ��Mhmn�豣-��qs6nX_���~�b��O��@����CJ8A���    IDAT�������l��=;�m�f�X��b�Mx��'��P�K.���_,�b�w��13z��֯{�V�������I�m؄�'LŌ����k���c�����Ƙb�q����B(�@���������a�Y3��\gV�)�5c��񨮪Ǯ]۱e�Z���.�T�~�I1k��Y�`ֵ�y�9��˦����-��=Q��]V���Ą�c�򣻫Ú��6��@g�[�m�Ν��L'	נ=��,B<�,k�ƛS*D�AyU�W���ڂ��H����}����?|_i��!�s�e���[�j�^V��|��!�
N?�t�T�g:�n�Kصs��@���Hg3�ҫ�fV�K/�6���W����܉��.,\�PO�Y���P�oni��������1�A��uj����x�ϓ���ш�n� ���ȫ=��>�4^X��Ip"���>� N�}:&N>U�l����I+A�L�d03D���>6u��0b�H�[�� h@����ޟ\DFJ��~>ܜX�:m�����X��l���w�-s���I��M��L<u�����8ַ����]����)�w�"��_�֋�P��a��5b�䩨�kp�7�70f�<�ϊWV�i�}�jq��������Ǝ3�j��Tr�Y�ʺ��I�i�},��U�0��,;)[�"�ǔ��[u'��\N�֬Ya��-�:;�x聧lc�����\�8��駝�|�o�[ca�%��3O����m�_�����!�O�=Z�����Fw"oEl�\�����+m�؋a��Eذn=fΚ��'M7৛�����8�����b):�v#��Buu=~��[��쬳g�e�0d30�9u��o��@8��ӆ�<i�Z���W�5n���'L7Z�L>�qG���e�3Q�*ڸa-6o]i� �b/,{�=�8�;�\L�t����Ģ�8y*��u.���GWW�7;:��ol.|�l����c�1ۗ�1�_�ֳ��c�o��,)b^k��\KS�Y����T\��ϸ�<�v*�&����F��شq=�a	6mjC!�A�u�˙�Hkw���8��3�٦r�=��w��]�v�ǧ��?����"���l�5uHuw�8���p�EZ��ݝX��9�̙����S�Zpgډ3�3���n�����ؼys��YY���������"�b�Y��O�w���\D��SS؟�}��I*Me����ތ �s�������QG�1�3���N9���
w�옝ǚ�+L㣏���E�6��[�z	jc�( �#F�ńc�������*dy�]���=F����ex������dc˴A�-��`�6ړD%ScGb/���æI�U7�~���u�}�Id#�5���N2_��9f�6+W���V��Dx���gA̿�\��ģ"N:�TD���,hcЕDy��6�>��ۆ����g�Gĳi��@um���#�M�,_�ľ�Фe�K/c�ɳp�qS-B��ة���[���֬{ъ�BA����n�bU8�hh"wL#F�������+���M'���{v�et�btIΜ9�O8��+hI� qԨ#��A�H8�]�����9 ��^Y�Gys,�j2��4Z��q��i���?B.��/����L(�^��>�{v�j���z�`���_��_���Z�5n��3���֯ ��?�9ۧ�����I�?+������bP����n�E*k֬r�D��{��ZP��9s�c���1�-��H$q��oǣ�>�)�Km��A��@�@>��?v�����;�\ǟR*n!�15 ��ј-�Ԁ;w�4ʆ�^z��wS..��'L�����7e���5�QV
NБ/Q!�����ӹZ��)!3��4o��g��|s瞅Y3N,q��L�oji��ˏ��V%�k�V�?����Y�=�l=�HG��Bc�(TU�ώ���S(����c1m7�{���G�Ōf��u����BC�00W���8R(sh߻�,��K^�Ë�9���̓���n��I4Է���,1��Mw�5�hߍ��^k�I@۾5�+��#��3�c?u���kh1����WU��u[����2�}̽�|�9�]{m\he�@2�t�w�EZ��oCw�?��ο�0a�DTW� ��Y�OK�&�
E�2L�d�;en#V���;�c[.�w	F��6�U8X���ᨎ58�K��H,׍ή=�h��K/��SO=m�o޼y���2¶P���Z˰���u�T�,���N��)�w�h۸��c�%f�dShj�Z�2;���YDcUH&��s��3	�}���a�fd�yK�e�?W����wߌ#������Be�y}��3%RhP�E�u��FL�"�Db��(����V�y睇�有h�4�R�o7� �G���R>I���Ltw㩿>a�E,2WR�׸�J������7���OM"��t�3�	J�?�S�֙��,���0�E��1N	ݨ��}��f�o,�Rր5����rQ0����9MEf�9��/e��g���(��L�C�|&n
ˮ�pՕW����@w�����K>Q�.�?�����"���M��M7b��H���e�����;j�Q�2�̾����sK�����_8��0�����d-��M3E.gi�N�8Ͷ�{���m�މ�-Ɨ��O�h�oFu55_f� ��U�1��&�Gx��'��_�����U��,!�\��L��0��-%0_�r���
��w?��O8��Ӎ��2_��1�ч`�u�rM;�&���g?�)V�Y���w-&M9�h�K�D��'��j*(X��	��꘽c&�ړ#F� �l�s�C,,еBM<C-�� 
�<>���z�U��{fO�n�,��9��S���4r��ձ�(���o`��Mx���c��wOյ5�˰��DB��,��*�4���;��o�4Z#�DM(H�z��yy����ތ�5��M��%���ܫ���-���ζ�<���x.����*c��!Z�sΞ��g�RBp�%����?T���1�F��G{�^hB��6���"��ń[r�z�5���T�~��@.�\�}�J��Hu'��@��#�iy��H�B]��n�fA�%K��ɕo^t�ܨ��\X��9������^z)���
�F�lق���[#��G���V�'`k�_����T�.����@�wް����ry\~����>�qJ��aʣ�8�'�p���6[�KKK�}�{1bdS)>�F����N�s��r���x啗��}����y�7o�c�$�u5+����L�|2���p����w[�ͧ?��3
���8��
8*
Z�Jv�>�X˖?�[n��=i|�_G��<�d(�ppEZ�7[�TM����p�w��{�ԩ���>`<F2jst�T�/�\�b������ ���obÆux���o-6	�|_'����	���eEV�`���}�߬0�C� �Zb�V��#���F,G�P$%C�����L%3֓��ʀ廮yg	 E]"��3��T�Θ�
�mNw�܍y�.��g�m��9����UE1˭�.|�_0��B|?Ο���[kwO/�����@� �G�2)OR����`���c	�7\w=�=�XK���c���5��Y�O���B���U[[o�>y�dL�t&M�d������L�,e���|�)l޲�h������
sO��7���6s鳙��L�&��<S�"�*�U'�{���䗮.�<�6,w��=V���=��w��]��f�� �3������q�@�[�8�>��{�\^��3��mWX���9�b�JI�GkJ��|7f8�}p�u�YIw�l��Vk�n�Oƍ�ϲ����o��/�%��s�W}�@��>��������+�.�m��vwZ��EpV���Kˍ�+�̚�B���j�g̜%��	aG����\�Ɍ�p��Ԟ%�պ��b�����������1���q��e���]�������|�Q�Z]���C�z(�'Y���*3o�k��S�rt����OBC6N��Hi�^0�k�87]ݝ��׿n�T�gS�S��"�ý��<^~ �oޗA]���7�lV(Ӻ�}*��r�������q�l>}.�G����ɬu� ��i.g�K�?:W�cj���|�u�p����-U�
�mQ�g��"���MWcN�?��?`Ŋ��;0q�D|�S��2m�iS�I��r�G=L�mj.Ϋ�~��x���ֳ�y�6І��o|Ê\�r:z���p��ӜB�*�a��͂\��R߄J������c�Y����3�\ݻ�F��X����.!��\Ι�Ȕ�}�=����fw��ח����	Ǣ���^承���5�	��ZR%�/p�W��SL���8{�7���\s>yi��p��'�ۇ
�2U*���;�k��`3�>[~WIx����S���]��z���>��h^��Ũ�A��aP�B���O��O��3œn^
5�mR0+�G�}�kMy�0SkC�$כ�޵��$ �����n�����������p�X������<����޻��x9�,��O�Q:���X��O~?��O��SO�F�R���9ܸ�ٕ������fk���ݍ�����J�����GW"� �]�����C�5�����0p!�s�y��>�7�s��Z��2��k�E���6��s��eQ�gq75�)U��[g��q����,S榛n*[w^��2}J\�|>+7�O�Ss��M�Vp���y���l�|^*�&�k��XI��k��(tLP��Ҝ�7�T|f��_ti��#KV��+i��%�3��?�߁������@��>��WZ��?Z����g̭C�g̎���ts�QY���s��ˊ�Kq�
Y�"y�>�?�'&X��N�﷍�~�Cop�?4��c5��4�}ьg�We�X�/�R�����4N��J��1�!^��z\�W_��JD�'�A�K.
�?�;Ǉ���$p]{��S`���ečB<���E4�p"ë4 �ݧ)N���}�ƍ+��qC����H��y�	��ɭ�}n�� �����bޗ�?��,i���:+Ҳ��$���
��j�^W�B�"AR)�J๪ %�����r���T��S�j���eM�	{^�;��	׃,!��[�x��i��)P�Q��?;����˕ƹR�W
��k����ה�s|��x�	k�Ƚa�%>�]�F���ԓf�U~dux��!���h�aY =-��&m�m����F$['9��`�� B��w�X�e!�}��ɟo��?�ϟ`Lp��T�s��I2���N���DN�����G���l�C!z��� ;P7[������U_U�����X�?�~��_ۦ%��%����njC͟�d�,�� .2�ļ����PY�CAI��c���3��4Tj�^�qf��`�K�}��Oa���,��֟���1.fi=��~��aM�XZ���������{���l�e��ɱ&s's�Y��:��)��b�.!�w~�N�JH��Y��_�u�[��������i��X�g8���?�b�0��H>����%U/�MB��� �<=���^ӫ����ͮ�+�Y�\���,t��(��뀚i���$�q�8�Y%*��1��]�a,���{��/~Ѵ4�T��Wr2�-G��[���	qik�*cD�A�=5�z�i�H
��n.��el��.����O�����e9h2t7�閠��?��Σ�e@� F0�Ї>�Oo�Jc��p'��y�FL%Gn����z!�݀�g�u�i<^�Z=�i�󹔦���5ſq�8�|g�>�@�8	2�Ko7��u貚z ^kDs�U<��z���޷T�{��������������$ؗ�X���:�O_2����4.
Uj�	�<N��?hr�?�k�߻�}B��]���]�8��N	�D�f�]�L��ޚ?��c�l+1��tKP�_J�/95p�ɾ�8���ÏW���ڠ��㩽3�[�L#R����I��k��V��S�3�ր����o��4L��ILŀ<0������7O<����]և��g���g�	c+�w�
����TO�+��FA�Ɨ�Qh0���)Gj�{��eE����_��=��y����j�e���d�p�6�;� �  -J�,еT]O���'MS8#�����/,p-y*���#����;��������.kS��ڽ7��w��˔���X  AN��Û�9�f��	��
�)�h��)��{z�!����� <� ����W�}�9�=�I�A	������[np
 �'��&�O�;��;��\��'�+��c$���}	� ��Z��b�6Xa�M���!��@�^�KS�'S>ǅk�V����/�嫴Β�q �+~�ؐ��v����x+��9�Z���)�%O�'!�w�6�h�Z���s ����pK�'ô!�D���+�Sօ6�ib%��-��e�-�|���8-N<���� @@��`/^ %ׁ�&z�M8������;�_�`����C'�D��Sȹ�G����0G�����	D�M
�@�a�����5���xǍ�4i�;�8N�|x�� �%Ùw����j��O�^vdJ�q������'��&L���H�Ф�4���Y�}h�|@#0�4\�+�b�=M|P:�,EU��v�.���T��J�r���6��L-���W�Cg�qo�NU�e�Τ'P3pK�?�2Y��L��1����5}Q�������a�)x�
�x�J��\�C=4C#``�(�}/�v� ���<NBA^�O��z]���zPk��R:����'Y�7ρ�Ţ8�9V� �	�B�-غu;�[�Ě�����M�''�Z�R�zg�ȊP�N�ƿs�9���|��ch��#P)���׊�oJɕ�/OS��3L`�8@a�:��޲�z\�.�Hx1�����r�m����W�]��C{�O7P'�t��'������3&FNYɛ�((Ĭ���>���◿�\r~Om��}s)E�o� �<�N�1���+��Ga�
C#04o�(LռJ�^��8a�8��!y��*Ͻi���1]�B����Ć�ͨ��`/��^{<��J>�P�eeĢ�_��y��s�8[�������	bfN9���햮&>
o~/'�����=�R\4��L�!�#���=�F�Ў �CY@��`vi0�2�|������V�R^�J�
짟~��՛��lP������nG{�#���2诧����_lz-M��7m�|���Y:#'���	��g�2.wJ_�U2��Yy*�~
^�a<��y�����GB7Ѿz��eedV�e:t��������U+ �Y���8�����U�KE��_��f:,DzH'���Xu-�i�4�J#0o���������3�k��Ϩ>����4�]��h����O?�-�6��C���c��)�����z���D�NV�R2쯺�*+���?h�b� ����}R<f�7o�;5~��Z\�P����8�#0P���7
�*������pԘ��
ho߃��_���/�9�$4�c��4u
N�>�N�2X���F&�c��{v��;��U�b����>_|!�?���GG�.lټ+W,C���+״�]��/��a��=hj��_��r�.��S*��6"�<�<I�JA@:���;����Yu$�>��
)�W��C�d���f�J��ߦ����o����ys�	�T��=���d��*b|�ᇍ+I-���,���=�C�,V���z\'������L��p(�DW�v�1i�4�{�\�&�F���� 	#��b��f'����y�e�+��6K�[�p��cxk3�a/�#G�!ѵ;wnF"�i���c��{W'��rؾ'���0>Jb6V�_�B�yK���ok���3 i�#�7}�C�."c%3�xi�io�3�t:C��#vx�W���2�L��� ���q�����yZ���v�a�
;�>NN+z��n�_���N��X�a!��g�KN6�ö�q$ytv�p���4������� V?��R:iI^�7�������s�W�y    IDATq��{�����
�|�tn���s�I�6)������=�شq;
�0�m�c�)s���Et���R N�.R�ra0����[p�h��j����xQD��t�!���n�7�Շ���5+^��N�\�l\3��#ͺ��ץ�;*rO�Y�7��Q9���?���[:gW�<���3��uQ�X�"
�����](ॗס��	�mÉ�N�o�d�ܼu�%�l۲���{�J.�\sK�����m��o������!��z�أ�~���nj[���g�9�|7�n_�L*iڸ?@n�6�����6�cܸ�֞Q��_���)[L�z�[�b@O���"sz��E�����:(�;yq���(��\��o�i����5��`P6�ܲT����O>e��dOe"��(���iՋ?�$}TIHw�S�ߋ���ں6mZ��nrd�ΐD2��ϯB0P�ݻ��|���~�2|�E?��f�Y���D^E���������f{{���}�l�Q��cƖ��W��p�ٳ�Iw`���Hg%��:;��~�&�|�X�������C�`o�(jt��[]T�Ϲe���i���L���RJ�����������P(�����P=�`��hY�1N\<ܣl���6�ai��ʑ���I��fNl]��Mvu�����˟��܃N����jlܸ�{��J��o+WmD6�Ggg;v����/C�%�o��k�������#�Jc��1����4��R�N�~��p֜���Ѷq5�.͓����q�m؂L&�u�:p�)g�{��y���;��'�D3��6w����L�`�L��9*4Sw�����{���{��4������¡r���_��/��]~�=Nk�,����~���]�� ��><f��x|�]�4i4ZZ�a��W�˧��`c�4��+���Ua���5���n�����;�������imn���n�y����������-�i>��`dK3��<^� F�jB�Ѝ�{�!���y}~?��3ؾmv�N`��$\�vK�$�3��\4�.�"q���ӭC�9�	�����;	�n��~�LM>���c��^�(��}�ڱQ��.��7~�������;�q�W�ޥb���g�q����E�̚�`i�3`���]X��"�TPc�捌��G���;;�ص�\x	�=�D�bx��p�-�X:���+e�Z��/ۇk��<A6
a޼K,�3�Ma�m��ٻ{��B��k��<�gG�6lC8ڈ��q�;'��o�TOQ=|�k_3�gF�z2ݓ�AGaB���~`1 /{���6���A�zd�܇�y�ߐ� ,�_���"�̦3�\bꕀPU.��ty��M7�d�B�5l۲{vmEGG;�9�����l�p��֬݀t*�+���ǌ����nK!��������o�����?P�o��#�3a�x��w!	��&���������Ĉ������Z1�ē���	��g������ގ���:�������N�nQ{V������K�ސU���uoٹ����j@��U�C�痦"�h/Į��^'KJǊ�[)�bB��\����MT0���(�v��y������y}��N[��Z�I[Ԇ��[���?�2AҎ�W�H(��TO+D�5��i�0F���K�E(��3a
O�/�@L����;��{Cc�&6�{;�ʚ�R�����uEE�)�j�#�@֬�-���zy8��_����g�{S{ϻ�1��w�m��T\T��I��S3"V�~���<��/�͛6��/����ծ�u*�A8�$S̘q2�u����mہ��zK3�{�R����y��?���R�7��ۀs���ݍk��N\tх��E0�����F�����{�PX���b�'a��3W����R5YuG��6	]=��ԧ,��_�2��f�i�`ж��|Ŭ��������ڜ��`�^���q1�	U`L�`p�L��t}��4����м.c*e8H#���ܔ]t\3���@J B�,��+}O�ϟJ���Ϟ=��*�CA}�(K���^>�hx{[r��#�c����	�us��GY�p��[Q>��_i���t�h<ԉ�?���ΝkkQ���i}�ƍ��̵*^)i�<O���֐�U�\o-���i��IF6Ї�s�g��SO-�K՜j\U��yb�<��wT��~��`��E�G�/�������'5s�?���bʔ)`;L�'A�}�9�=ʣ�c�����D�f�j���{�j�
[�&p�>���KQ_7d#(|����Z��b��c�����h�hR6g)V�lʢ�'N�n�܈�H��,��0�� ��"",��Հs۶mX�x�i��(h+ �����җ�d������Y���H���j=��{��*Ս ��w�۞�@��'P��gg��-p<�
��g�8Â�
��$�%W��o��o6�2��o�G$�]w�mD�e��w�	�����a��s$�x�)���i�eG3��T�Y)ܴ|Ư��e롯���~̸��n�^��nu�i~>�����M���c�# w�R$�2��*�'����-�%�sK�X�I�����2��J�*�4Shm{�y9�V����&��@��~�T 4�R~x-u�b^�O<a>u�[i��`�`�x��kM��t�R�df�=�̳x��l���
�����[��_��_mdAr<�'��'L��"�t⬝R��'.f���/��K+�;�S(�����/�ws<�q}%�_Ҝ�C!ׄ��/���/�	<j�X+��ĤS�=��ng�Z�Ҹz�z�ro�>���M���}C��Y=�<�pT��i��]o��4�ú���4<��;��P�������*�Z
L��XȦM���8�K����c��/8.�P�|�[߲":�6��κ�����y��n���sx��|�,
�����YL,ܡ�ƹ�Vʟ�'���P�'����:Ӧ5!W�c�����'>�ѣ� ݝt�鴍g>Wj���~�,zx12� ��"��&���4�\c}��$׮_��~�����3�
	�a�?�S����Ϳ��q�1��nPo�y_뀱�5ZT�����߼�M�b�}T����*;�DkF��K�Fp_�z��w�'�t*z,� `��:�ݏϨ����;�-�<y2����@��2�@��d&��h���x�������y���*��d�m�w���?�wį���<�M��/���b	���aĈQ&�#W��c�m�b�H\\�r���2k�,�`����	&4��{���{����a ���X��k��|j!��%���9K}-��	[�)]e%u��i����oV��y�j�/^���{���J_ڧ�Ҕ)|9����%
�4�e�!����q�Hx	�5��X 3�.����b4�K^��||^��8j��}w/��9�т��z;Ə��ꪘi�Ŝ�1A�߬�l��N��~�%K���b96����80퐂����y]�?߉���_X�̲�<<_��֯\�\���ϟ���>�ƕ��j>��y���J»�:��B�2d8��I(��k�YY@�5 k�d�RYܡ��^UV�u׾����rl���%v����*� ���SӦ��jL�:3N�i����Z�\�(�
ؽ{�Y�_|˖/�`�Yxp��IH�ߧX,f�[Zo���^6�����W�` l����h;%-?2���}���b�č� 087�|y\�
Ԋ�� C�+]�r��Փ��:s�L+�b�@n-�}�C=4K���"?�Lpj`|~� ��ǟ\���h�`z%�g������ K��UV�5k
��AG�$�;��I��97��xg�mJ����^ם�W�����1�t������T\O�J��}!�PЇ�G�D,Ze׬��3��s���Z�w2�l=���� 	���"1#���lr����u(5>r7�
'6$Rq��Fg/�*�D����1�y�ǖ ���WZyA��N��8����\^|^^��*/[��x���Z��ť�����.Ɯ9s��X������~r�0�DE���U# ˓���pMM-fgry
��)���q�;�]��/ 
�?�p�T_�Kk�����{��_d�h���v6n�w��:l��6`�~̂�a�	|4u��5�F޹���h\,��c0�~UnP��e��dpL����IVgi[�78d�3���M��Lݔ����H3���+�?e-�R��@����~�^KMA`>���	�y�,+l���u��y׊e����r!�{�����5�.���u�}|��<�"Zʱs�Nz|���[��Cw:�T&mY�W�;m��#����!!dq-�)�l�("UQ*~'A�FD;�#���Z�^7��-ŀ�:Ї�?݈��y��'��\^��)6����-�,^�1�Ә�8a�Cʅ�C9�P�"�����82�ɖ�,�8]|ʝ����&L�0wkIY�4�C�_I�/2G��l	���}6�����28_A �w� ~�}9�o�<��XNjE�C�'5f|����P������O��@��p}/_����ƔF#w��@��m�k�C��8�jb�ո�	�x/�W���'���=�Q�,�L��|yms[T����+뽏6�4P��xm���_
Z(���x�Q�o?y}9㓊R������w3Ѐ�(|�XЕL"�ݍ��%BB>�57|F>��G�{��=��Wf�U��?�nP�}Ya��������;�0J���T�Lk��O�TP_{�{}	cY\����|?zo)�^+���|q�r��w���|���:�ڰ���,Θ���w�Wpk���ܰ�C�8>-�XUM)�9�B�Y���ks�u����@n��>���Uޏ_q%߾>��O����j>.�o~�.�\^��b�t�wmmm��HM�	�|z�q�ۥ�b����w>������c�F���8&qӊ�n|����&PB�2���9����
��	��1�j�����	_�ц�������]6P_�� �E#`?	�;ݎ��,A�� ��է2�}��V�[��|pL-1@<��2�4~���ZEWy�5�׼{�Mq�}
��ރ�Y�W�e-����y���t��Zpoփ�8�R�O��SƞR_��y�A���[0�g�xǵ�|�}�������k�k���11��c��w �G�r��R��w����'�&��f���iԇ�k���m����*ȕ4z�p��#����������Q;��W�ل�G �{�B	�$ zP��i7�_6�����{+��9���WC�����aN��{�B���L!fŰBPy��'�Ng|mK�������b�U��S�0���@�����;�C��k����iT����*��c=އ!Ϳ�ٚ�`�/�����^�/W�4x�b�?X
ZQ�C�!�]�J���K�0y}d�݆����}�f=�s�ұ\��E2�EE��"X6Iݜ���S^�}	�y]� �==ǻ�D>�5��o<�~Me��_�����p�L���h{�Y���8��K�;�w�Cm^��R�@~�ײ��!�?����>N���t���b)�3�C� ���>�`	&�B5����|�S!69���A�?�~_�P�˗�*X�0�$ �R�	�S�2�5��e_4����!�?|��/*��}z�?��l���3�K�O#������p.������e�x����W
��J@����A��3o@Ϳ�p9��.�n�G� C����uL_i}"�� P���ؕ�/����^�UX�C����:ʜ�ޚ����3��f���r�i�o�n9�{[O<z>����{�!�<���_(��1��7����qzh�;I�$	 �M)�._7d.Vs*7��+����a��}\@]�CK����+�?}��Z:�?h�>ݩ��;P�t�!�?p�}�a½�z����U1�� ��-����[���om��`��-X���x��*���A��9_�:���W1o��0&�������h
�L.�M��������G#~�@��+Ư"Q7�U���U,���7j(e�0E���������"P�~��������ZB���R�?��q�|t�Z<��*�Qі\i,2�Y6W��Ze����y.�->�ݔ���1�G�����0�^�z-C�S E�9s�(�O�U9����nx�p�d7�錍m&�~P	QV�����|V�6���J�9Q"��p��*k��s<ʬ��b�bU^
�ǎ���X�� �k<�TZSz{+�5��ޞ���Y�益=�{C�Z�'�jo�^Q���G�\�-aV\>_N�渲��\=~ �h����=v�+N̻b�e˞7�qWp6��?��y�"���������q�?W��E.m?F�����zm���>V�=�B!���&-�j`�&K��k�8��*�i���#��?��% T0t8��\�L	�ci���w������n,��R+T��Whv�L�6���U9����K'皙x+O�!is�oW8�tm`iS(�"/���=^��J�������E�+$^���������r�����@��)巪^�hir�Q�H��.9��8q���lh̩�X�TI��
�%�����sz]���~����|g��8�t�QPp���sq�xoS�I��kk]��������)o�s/�'��Ϥ�=�i�ڐ��U��.\GV�۝Fsc�1�2|ذ$Sd�u䆉�k��V�$�[���9\�\M<�p���/��m,G�Jt9���g�y.�{>��r�O:�4nFiuiv_�۷�4C
m i*� "��F!�	���w/�x�B�`��F"�i�RW�~��/�1I�Tۻ��	��	V��x��}P���N�J�7 ���#F�w��W��ss.�R)mb�8���;����x
x�Yc-�d667�S��ל���_ȣ:Ve�.���pu �Q4��
"�c���Y.���������:3-��E�,&	6�#��(���	N	X�{�ݏs�{h�Er�k�;����Ha�߇�E��,-	j��Ƿ��ގ�=^
/��'��s%���g���0�Z���ӊ>aډ�����W�.�h4�ؾ�:s���T�zV�X���q�Q��-�@�ɞ���/����x��>�>$v�3kcU��e�I3��oKS#2���X��Yk�F�-.��ԩS1i���k���.l�B�a.|.n�#�<�ƍ3ӍVB���M$-�C�?�:��~ ��MWGg���h��_<�V�	ۻ����{r3�1������ �U�oV��m�L1	g��ZB��TE@o�W�KSK�Ϳ�CZ��xe�\�Qy���w|G�]���Z���ޝ�_Ȥ��҄=#���]���=w����!��RG����f-!���Xr\ml
���:+a*ˇ���J�)	yZd^b;���8n|w�I�=	��LyǕ�	]�	bY�K�P�{o�Y�)���:֫��~N�:�����~�s����r��9%(�F���q�U{đ�DB�fRض};�y�i�w��Z�Ţ��;|�H{�h�Ŀ�?��'k�h�i n�A����a<�qc�oմ����q��ދ�G����(���c�`˖Mf��������Gy��v2b���nH�L�~�7qQ���<�_c�@n"i�2����5�v�����˟1o�E��H���|�I<��2[%��ߩu^xᅶ���
8R+	@���&�Q�)���x��)�i���8q�]OZ�W�P�}�=�II���^b.�#�l�C�^j���e��r�xP�����;y�P��B-͍��c�8��+7倾�]1�<y�]w݅�/�����F&H��ƙk��#8_����[��yK_x�>�h��D+�q�e��36GlIK^S�7ޗ�p�w�y�)Di�_��O9���J4^��uE�C6���l�Ə,$�}8FrG��ټEc��,Y�[n��L�,�X<F���1a�8�
i��	,~)^Y���&0�!\g��L���3g[G&<��_����j��F^\�7�s���?h��?�'�S�.����w酸���+f�N%�f��xa��,(GL�O-lW{J��s    IDAT��������r�����F�L'����6�}�Y�[��� �!7�c�=f���J�����;�k{�K�5Ea�9�6��K�$���{���\m�����5�\c��X�x�cC3�{��6m�\�*�F�v+-��8y�d�i�r+�Y�.
�qd�1���K�N�/�7�bw,cW,���s����c�<�쬪��N���IH!	%4�]P��2"��"
D�*���S��\D)6H �t, ��i�L&m2s��~������̙3%���'�̜����~������Q���ި a��}6��{�=���FΪ�j�p�~����4Z>��#�;�����f���Bs�8���2^��/Y�T[.ug��Y�|G�\g�64���˵��|3~uS��ڧ��ֲ�Ro��#���4S�Y����9R��q{)��T�E<�|����i�(Bt�y;J��J>�!y�'���u��qo(�\p��Cy�S��?����V��{
��"�3�.���mr��G��%y��X��t��Z	8���e$��� �l�Pe�w�o&��^q��2k��2]��c�� i@���Δ��6Y�r��tw���<��w&,�ΐ�9�<6��p�X�[@�Əf��~�i�%Lb����!|m�r�є�i�����y�W�blsr���qPbl�{u_ɺ1��5`��f7���D�E	��ۢ+��h�ԼV��i��9�����g��5��� �W~�����C�h۠F{�6|(���i9h� �O`�`lX�?��������t���K/��ӧ�����k�W� *��oֱ�/���	L���s�Ygi�l���1�e�*T��9��́�N�lNۏ�X9�kZ��0��DkHU���|�u�i���|��k�T�� �Fu۫~�k�g�ش{�=���|E׽�]�y��=~?��hw{>�=~�}③ll^,�T�������˜#�X�(/��5M�$���u媫>&3g�.�lA�x�or�=�H,��}n};#]��~[2��J�j�O�� ���ڨ�}�r�����r�rI��f-�M�NGd��9��cK}h�������	�S����Р��CM��S���3��r�����8E��̵r���1c�>����#o�q��hO �i{h~F�������K��u�P7���q�  |��6W�k��J1�b�?�^54f�Q������yJ4E��q��&(��Z�v���_j�E����瞳w�/�P��t����E8��Tł������ G�q^�*��;�MPs ���35�ߴ}s�+�Qp�6��)SJ��	_w�y�j��h��Dw���t6�6׀?=|�^0��7ø�m��+��_���9��W���UysچR���i���ӟ�eie�yN�w��Hn�g�zHƍ�˸	�d����U��tN�-]-�\X:�S�����sϒQc��ˋ^����_��͙;��ɶ�+�?�3,�ٻ�&W_�!���ic�<���r�GK>�%MkWIgW�ĢԨ��斤4�k�l6&���d���Ҳ����җ���'�E�hٴ,$۴��'NP�0-�4EӺ�Kܞ��s����cƨ�vb �wM�t�E��pԨ�ȖIH�ײV���h�f�"�\ )���`416\_Z�?�/�B�'�d=�����E��s~��|l�an�]��/��8-LШjh �1�t���CF��o�k��8�]��q2f�o�ͥY<G��9}���ic�o��8KN�~�X���J�w��-��x�W��u{��W��c���uO�ߡ�� ;��{��gk羦&GU�u��O|B��|�+�'#���3F�,}��ڰ'��c����"�iiMI,Q/����$D�I.�ma0{��l���G��?g��&����G��s���#WX"�����By�O�!��-�XA֬]�m1�
��l��.�6�O�F^^�V=�(�B�(,P8bQ$��pL�����Xx�Y4A5����4__s5A��-n�O7��1�	Rv^�����67	b�e���>��kn}�ôG]��xWz�:��1���� b�c�����>����S>���'��ρ%,q�\�:��U>��/�?��aB����� >���O�z�{3Kz{��Ӭu��>�\N#�h�������{�.8}�~��l}A�]q�J�-_��<��{�G�'Ə����)Ţ�ĥ�+/˗5)�l��)�Z;��o�Pԅ��䎟Ȋe�J}�s[�����j�Oz5u�NS��k>.�b^��.��m��c�L�]6nZ+�=�.����d�4��$�y�ؒ��{�E���*~4>�i4`�J�^8M8P�p���;��1���Ȩ��6y{.�j�f��Z�@�`*�8L�y��}��7�EE��iަ���>3���=�����;����Aɿ�	=�,�����ܒ���(�&����k�v.��]���+ 6���o�3��M �
�	�Jc���߿��*�����s�������2����� ������Ϗh(�2���X�PfX(��׭�'{P޲�,i�8ZV�y]2� ?#��lFd�+�K$Z/�YIeC��]'��Uo��fY�b����R�Ap�������i��}��1r��?*�u52nL�,��Sy�>�J����u���ۥ�G�	i� �[��+#k�&��S標�Åޙ?~ɁH��SN9E��Ǎ�R��[nѰP��\t�F[����j��&f,o4�������L0��i���f��`?_�5'���K�F<�}4��9���h����(�Uic��H����l�|6�v�6�c�='��} �4�V�Uc��߿����)��l��������}'�/��y�fY�M���j�f�� ����9��w,,z_��X|��ΎM��ӏ�N�GI"�ի_�Tڕ�A{OO^^|a�D�d���r�ۏ�y��֤?��w/���������3�gvĂ�i�7~��-yU%ڇ�Y��Qrּyr�[����VI&7�����"�0 �➡~��Y׼Q�6o�T:$W|�*}`<�[o�U����׿��=1�h�\r���%�m���.�C��k	_��,zc�x8�/�\��4/_����/[���[>0�Z5�� ��7 �/��|喏��]������<>�җUe��K8�}k������J��ӷ<�}_Y�����6��/��p�z��Z�׵G~��7_�~"��?�|����͊�Ә��@���j����ѾQ2�N��R��C�����BL򹰼��5iK���^";�<SCA~�a���%��T��w��u�=w�}{����/���xC�=ye%�ϓ��T�n��v�X$������MR�Nm���K!�x�N�;�p�m�=�D7�勉ǂ��K������w����%���A9j��x㍚d�S_���y0���Q9�].��V3�r-��r@,�0 ���%`/&tʩ!Ӽ����W�����������2��}��\�3��e�F9��[ff��c����W����TK4�ݗou���r_�9�4}�����$`����Ja��l��K�'���p?����K.��2I��*���חȚ����t9k�#TN$��ttfd�Y��A���@$:.��^eFՎ���77�a�e��Ͽmā�$/�_#k�9�t֙g�	�'�I��Eem�Jy��G�E�4��E���C<DN8�d�0q���&����s>��'1���Q��	���-Ġ_w�u�v]�j˖-�gc��e��+4��6������26g_Ԑi���� �\s���G����1����s�F]�w}�5|����[�3��)��@����?._A(�r��`�mǚ 1N��90������1�[}��h?b�W ����XC�w�;\ߊ��Ӭs�s���WK�K�dlD�� ��<���}�{�+�|��c��j��_�����4�]��� ��g��M�9��s�}$�/j��G{T��կt�`�/pM����M��p����dā�����f���*���k�/��޲�d�i�0�����.kׯ�H$�^���Q�'���x�F�v{�-�76 ��,��,:�a4��{�q�>,6?m~��w�߷LO�2��6�m�j������V�7ЄmL�¡ڵ�|>�����7�-_p�S��P�Y۹lN�D2~8����1�9-⬿5�h�Z���i���ߟ�r���{���)�}�A���5���kв����w��cʬL���a��E5���:���.3w�x$*�|J�I(]�\-�J��<C����Db���勲x�k��L:���Ek)���;�~������)h	�?$17gyW���c�	z�n3R,��ڶ�X��H\6lؤ�(�`8{��q�<c
�>?1�"�.]*].�Ӿc��@o8����w�\����\��U��>ܱ�����w���	Z��\)�u[i>�\>������KHM8p.~�4q��}�9��{Hm]��pF�Ơ�s���W���ߟ����w�a�}/����
`���T؍	r�TzB�ϸ����d�ӴD ��<$.��W˚5k4-�� �Gc8�st!|�ߔw��r�W��C�_��7!�?����0��l���\~��-^~�9c��(�.�n�3���1��3P�ӱX |ƌ�g�$.�x�����߯`mt��[��:;z�V>��#d֮��J��m<�%�)����/��ؼ~�
����:�{�
��Xο��kRa�]c�b�uM@��3g�t��ٔ
2��E ��n�KI7��'�"c��D�|�T���p��iZ������V��b|4���YMPq�JiB���m5���1�n3`����ӸSj�S����Z�T�%�+�}OUU�^@�6|��h9�F���)Sd�3�&Ӓdv�x}�J� l�����ߜ���\�ol�)ٞ��R��{(��n�� ЇM���+�f�?U+�j�HfK�e�=��h��=���t ,�`���{�Z��~D~��ȢE�Jac`���l�d5�,�6����T���lc�{ ��ߎ�7��~f�PoW"���ֱ�O=�TU��A�ɜ��`��?�h��|�8w-��)���}��8��	ܾS�x9��jUϑ��6sa.�9����s�Ľ{ci�����a��s�2~��7��Q>�yv�Z�.b�����'�"ف<d���z�qu���ʬs��E�7i\���6�q��ގ�w�j��MX0C���Z�r������O�'�?��u3�9W�y�1\3 ^vL$���G��� ���w�+�F��?w���d���4<��SIO�>�$�o�]X[X ��kSP���9UM�дa���Z�2�V��pJ>x�AB"Na�},���!}����i�&��~�-.,�-��������������3��g_X2�%l�!��\����J)=y���{���U�H6�@�I8fmb�*KmM�*\q�Ǚ�^��M;�#B��#����xK�=yI%��|>� O{�z�Eh◭T��{�("�|o-u����� ��_ViM���a�QŐ���'�/�o�m�X��p��%�X}|?���E2X�J���p���;f��},`¢x�ꯖ=nܻM��('����5�q���Vp>�f:�v�D��������Wp/��\��B���,��3�4�������8�*�O�n,��F D� ~H�0���F�
���j�Y�u�c��'�.�����c�@����]�\��Ec��p7����#�4ݓ�s�Q?�EE(p,��M��Ꭳ��{�՜&D���1#��}y�m��a�zO)ʡ �bX����tc�z<7֓����	u��w���T�����g�r%,"N�{�iڼ i��^�Z�
7
��7�Is��G��d�?tE���\�4��
��.�;�R��Pi&�����c
"L�N2 ⺨9M\�GhX�
 ^V����
)dz%�����m�2�/+�ZB�{�k����Z�6���4�+>t����Pi)���L^���9��SUU_4�5Kry�21*E���D����x4��H��Hb���9��3���MH�<�Ũz���ϲ��֞�H��	�hB�Ǣa����ϥ�~�K졭g��o�˜�VEV�� yʀ�֥�_�)��o���xn�G�>2���
Ղ2S�d�}��P>4��!3�%�0.	���}O�\�v��sP�G6�W��#!��b��$1�,�6��� �Y�]X�E��D
���F�����-��s���?f�I'�K�w�y������ӱ�5	m��|J��X �>������n2�`&��8Z2y���$�1	�3�tHM�[:�֋d���HݨIR��%��c"9"������ϰ�Q	SS�%ߛ���l�N
Q�LT�y�Q+�ܲ^6nZ��^5-�C���~��d�`��VdN�.�ϱ+�3�����7!�X,��>��-�ʔ9W&ȸ�j���;����p��l�Y��`���9����0]��J�*�|���?�aҥ#��Ϗڒ��*i�L:@��C����a�e2���������g6�.Y�����r��6�Z�v�g�;K�O+8�
y��@�i��o���f��_��u����/
�c)�$ �m� u6��SN9I�<{���Qb##�IL2�uHw�
y��dݚ5���mǾSƌ�(�bA�E<�0�XC �<�
��Diբt��k$'��8I�k$��H1&ɶ6y�OԒ݉�:�Td���/p��̙��YT�$�Ȣ�,�k����O�����DùJ��	'����{�Z.e�s�b��}�����e>=��h��M(���zA�%��{4H�T+.PB��2A����_-��'~�i���k�FMM�F�(؇c[4Y/E�� �B�F���˼���n���P�M�I�Nш��e`<�̢��;��=)��Iy��h�#l��\;�l��Xb���!���*�l��J�G
R�I$�*��:���Ț�Kd����ݍg�����y���6�m��d�*Z�)���J6:^�?C�z���i�I�������vB��'�r�c�� @ȳ:�3�$	�>t�	&@��}[so���$f�(�ǀ�$
�q��aaS�B��������؀0N^��P= /�5��C�R?fQ���2�SJ�?��[]�o�4��YҹZUOʹ�)�ȡ���ۅ[9n������b��L������+�V�i�,Q*%�˨��F]�Z ��S)�ɤU��L�H���t���-5��&"�#t(
Ю	����{�±Z܊��D� �\���I"�"�^p�lްF� O>�Q����G�F���ry=����c�}$"�P��#�$/����-H}�hy�EjE�ui�x�s��{�� {Y�y��2�47'�>3���g�f ��Y�Ͼ�i�n��O"��XY��7�կ�ϱ��@ྍRV��r�Vp�ņr��ou����J#	8��ܵ���c����;��dۇ*�>,>�4��:�ҮA3�#�6���w�}4������
h"h&hZ<L4��1���M|���|�v��U���%�؈�	G$_�jr�Y/�x��82���wu���qN`C�`��c�f=|�J���*d�.���P��:W�}w�"��keڔ�2g��R;a���Tt�`�/�׹�)�~V�DX#��IE�J66Vr����b�F��H��I:�s�x�|U��P�7��8�h�Dv�\Y�4�ӟ������cL�5���&�:�,�����k������?�W�u8���-�����d���RS�ڻ����h�
���~�D\B&�SkE��׈�j�����N4�|XT�pL::�d��3��w��͘Q���1Rp��ާ�|w�,>�i4�%����Oߏ@���Q*��%w�_�K,'s&eD�D��gs8<��Y%C;@�0�H���p����3��)��&��i�f;%�k�����n���52i�$y׻eB�N��I�)��I<�W�@�O\�֑��|1,�P\ґ1��-    IDAT����Lx�d���
jRc��7|O��Z�B��r,�2��G{Qd2
 &<�֦�����G}���e�����G�{${�,n��u�ܹ��'��)K�B�ׯ�iJ�P�����Q=%� ��!��|��r�1����SU1����ē�* ��]J��T{�#��5p'�V�,׏�M���#o{�12��4M��f{4�C��_A('��P(��1��'�����vg��o�|���a����z��|Njh�I�i��pF�|�'`�!�i$'E�hS�lЧ ��n����@ ����,�^�7~�g��F!-�BJŤHO��������2m�t9餹�0e�tt[xja����POH�BB��h�9�	�M�j$����z�>C�߰a��薛�E/�0@�V�۞ c9! �瞫�}ӊx�-&h�ϛ��|� (�ƽX3h
�)��Q�*f{=#��L�(:m��ɹ眧U=�����&�F՗rn ����0�A::����ğ�T����j�/��dD�>��������G+�>x���h������|@b���]'==���+�i�Ji�h�D̳=��Kf�ds$m�f�7�t�.V���o}?���4����[5I�c~=�<��-�J��R���-?Q�?����Ȼ�}ݜ ~�����$���4�����w{�?��X]7��#��vi�u-ᨙ.��%^h�pz�ܿ��Ҳ�I�N�*'�|�����d�]D$L@��7�gP?�����? �/D%��tt�d��[/�P�&|��ٞ��������R�\���@��̔+��s���a�DЖO9�Ufx�[���<s�G��5i�ja�>�VC������k�[	��4t:pN�x��ަ�N3���e���I��J(pN�)@�˚�����YH�ͭ��ZP���=r,����#{��C-r�N�;Zeٲ%���0y��m�=eԘ��Jgg(�L��ؔG�Z.�F4��il�v�=��J����l&/ӧN���u���mw3v��\�T^~�yy�����E�A�%@gƴ�e�}���;Z(���z��'���]�t��g��P<���L^� <m��kl����a��5�7Ż��U	�K����$�RISP�����XM��p��%W�v���I1�)5�#��&��*���Ҳa�����O��:�cͻ0ϡ�4r)� ��>�� Ӝ�I&2�9|#��KǶX,!=]���?��!I�9�a8�>>�E��U�X8"d�J$�O���0��#�=��$�
eb˾cc亥���w;�ʐ�&K�4(,�p�PO4� }�#?��?��pn���_�Ĭ{�@Y�2������n�:�h��y���?��J;�C5�1�M��e��瞑�uM�A��tugd�]f�G-�춇��.��GV�m���9��w�?����B#jf��lZ
��,ym���ҳR(f�.�~�$�HWGJ:;3�����G��
��w��]u�(؄���g��?��j.<0u�i������g�yF��玚��x���P���L$H�l������m������s��(��P�S��Pf���[�e�j����j�)�?�揀��Z�B��֬Dk�P�JN�%������	��p�v�wȝ?��<�ğ�TW����۠% ����I�����wb�)*� D��c�t_����+Y`
ʶ�~�������������}�$Q��c��|���dJA�B�/0�J1�W'k&S����䢋��C�=�~g�)�����ַt�~tc����_�4l�����^��^]$�m%�^'��:I�����#�~�z��݋P��]?W_ k����0i�#2�s��9�J&�?^I�g�y_{����.�fH,"����"�F'��e��l^/==��$��rE�ܒ��%3r��)S�(x[M��i
\�f�Gu�nD��X��K��అl�}�-��K�`J����$�$ �A�
��)���}
P��JZl/��UMG���4v��%����������e'h�������0��|�o!\�"Ų$_�s�ђz�6qٸ~��z�O��?�4�m��e c`n`=����k����g�r�Ъ�<+V�(Պ1+´c�?h�"4��-4gֿi�f���l��QF	��Ϛ5���D׻��V>�����Y�k�>X����(c�D0�P�$��{�{�k_�����8���.�HA���p��4��/�X9�I�tHrs���6˺uM
�(A�C�>���^�^:���K�a�Nz����k�#�}�'ߑ�z���%���l~^�N����5��6�{���v���e��W��#��_$��u�7K�ڍR��,[�^�9��ڸ�M�"�����d�����f8���|�C�/}�K��iM)k�q�8���CY��!��d���z-E��8οv��
��2�k���u�����餝�{�	�L;%Z�,��*���M��NS�?N�'c'L�t7��f���߬\��a�0GaM��b.�%%��d���ʈD��i���G?�%˖J��m�/�P�`�_�������X)�A�Y_����΍ՊF9m�4}ˀj��9�ǚ��?������6 h��Y066�T�S&�	]�N�6V�p^&P̪�s��u�]'+�-�4�cY��%���|�;
�P@|n>����o!-}��2u�x�PN^}�F���¡���s��2v�N�t�j9�'ɻO��x�Ң�jo�,ݻ��_O;���/�s3��,���c"��l��$���r���b�G6�4K{{��c%.�iY�n��sY��]v�uO�n?��M��/|��ݢ�������8�8|>�я
-�xX��o�߰�]�~�W<�ޠ������Z �_5�=�/�w����U6KK���c]���'�3�����e�r�#�|U�'��������t�<3q��)��eu��3;Dy��D]M]��Ʉj�G�K6<J2E���g�f�*��?��Mͮ�S�(7��_�y}[�?y&֏��8��;�	 �~XVn[�&\��� 5����8�aj~��9�� ��bV�YF��=7� �?zf��뚀5*�_��<��g�^��Nj,z�(=�Qj�~�U�Ę�@��n^/O>z���,;�N���AW�?&ٌ��Eˤ�v�4��$u���ǯ�V��FIgw�^kŊ�zn~�����h�l�0�k���CW^!�pQV�\*?�k9��äP��VKWW�s��jd��ViZ�IB�zY�z���!�)g&�5�\SZ�,z{8ַ�
��ޟ$R��8�m�9}�`���s>��� V����5�	p�u���o��匇�EI��֑���
:�!
B-f$�k�Da��3����&�}��ɪ�O�?$!AcZ�?�H�\J���7,�bL���;!���_�1 v��%Z�aS[�UE%t����mƀ&b/Ӝ�Й��|�R�P�7��zt������$8z˜�s����\�	�q� �����H;�()s��}[�:�F�"�L�.9�i�t��gȧ>�)u�ҫ��k�U`��K�B��&�h�x��e��k/���J�<r_i�4V����1���l떥˚%-׷KgwV��m�caٴ�EE�.ݲ_���Vf�h(4�=gϖ�\}�Ĵ�C�����;�y���]�~�jimkQ隈�K��NY�z��r1y}M��e߃T�ǼE�n�Q�>X��ӊS���Ik(���g	/��@7�v�cK�qmAT?����\2W��?�}�� JNi����^�+ڡC�������?�q�u��LN<��D�K������|�.��?~��h4RD"�!j�Nϗ��d%$4 ������}����#	��(1��|G�l��5Do�������M��F� �ti@���}�!��1^>?�uW~,�e�o�I����_�m��˵�"0G��6?�o%�IO��í�i�Ҵ}_0r?8|���<��#�<R-�;�C�.]�S��g�(�����<����̖q�G�kK��K��D��saye�r���ٕ�L6,���:=j�tv���C��0&?:�����n���5�5������~L�j*f����ˡ�'�b��Z�B
���i��M����뫤�#/k��ȱǟ��?���8�j4R1G�q�<,6+&�]w�UJ��}����M��^��m?k:R�R�4.��k`rSBAk�����x�C��崺'��2�
�E��ˠ����Z��K��#WKD���f%�k�p�E��M�o��u�d��i��O��JW� ��GjS�;res���Y<9��\l���%-=��C5�'��W_����/k}�����WU��d���b�ͱ�),�}_\������[Pۦ���%
ڒ�ݞ/�K@���S��,��^������Fa��^��P�,��PV���8� �gs�Z����(k��a��iz]:�h�p8"�]=�|�jIeD6o�:\�8���+�_[.w-�/�5�m6���ܹ��L�]]���]�F�{�{������ukVJwOR�6��\�Gyr�$ź��U�o��Y���רs�ŀ���4v��v�J�{�WZ���A{D`��㎅R��s\s�j�O;.��JN Zd,���u�>���xc�����Ւ��q�:)3D�E���u�jA�l6%�t�$�Ih�g�Hj�<xϝҺa�L�� '��Q�O�.�T�GE����{�i���	z5��aL.2Z
�1Z�!-5"�z�<����_��������C���F�;��sh���r���A�<���a�>5����l�}��6����oK>M��K��l�K֭}U2=mZͶe�&���n�hm]��^�$[���ʵr��W�����p�N~��?�/�KF�%����m��8���m��+���ƙTJ�._���$P��d媥�|��QL*,�t��5������3%��V�1swV$?mq�qN�iF�C��x�%n�E�B�s˜J��ETqkT a�泙��:���db�5;1W�=�5�kj��'%�Z7��U��?�u~��-k��1�[�y��w ���F�eR��vK,��!�l����r��ۥ�y�4L/���4��O��H������<���2�4²q�a)(��B�^r�1*z
1	'F�g�)��w�-���Ev�?�����/�}i��Q@��?��X8u�@���9�9���/��ژ�3�����M��A	%�GK8�q���7ȸ���N)Ƥ�'#>�;��?�s��~��ɫJUϠ�b>���cG�YgΓ�;X�]�m��i���7JG[Ri�P!$�h\�L�*���Qv�6K+C"�)��׿�����x8�}48U� � ���4�����kU��*�O��q����Z0*��%�i�OKWG�߸�E����$	�Õd#;���@�/���S��f.��{�w��х|F����%%�L����_�*�Vj�ƹ�d���E���lZ�ZVZ�IT{���/��/���I12Jr�Z�)F%�-�L^�Q��ǷH"�V�v���b���,D��2F��GI�)�����w�h�믿^�=`N��7�B&5��x,,�L�<��S���OHw��E�g����Ւ��s̱�����3V��^�Q_KJ���������++i�tɱH���0I�s�<y�[���DL��Z6o�H��+V�����HmM��7^r���?�L���ø@�RY$h�˖-�Tp�r%j��vq왃W��ΰ��_� s�r��O>Y#���:"�Y�+�fZ|�UWT�z�5�O�1��<�v8���N�����*g�{��I!��P!-�ѼD�ݒ�l��~�lni��;M���q�$�FK���Dj���ϕF8�5��/Z<>�0��:)D�$NH�>��:���R����)��H��ڧ�2�w��ه~�nԜ�D�QR�`�|nV?�d��Ib�߽�ҋe��	l5��sҶy�,Z���\�R�'64(1z�X]�������=��qB>��_��?w����+*�?tN	�pxf���w�q���{�)��u����%� �ߵ�u��IgSZm�����-�>Rn-��+��� "p�P��/�+�A����í����ꩧ
U�Jt�g�����|�s��д,�?��I�=�y}���~*�%�&M��ft�m⡜�r)I�Ҳ�y�!p���S����K��ه��O5h��<��#T �HB��I���ȑmIm�M�em�j O���Ù�ߡ�7[o{p��c>9����M�+�y����^�����l��o�8�!� ��sl6�ў�T�em�_9.��+��������Sa��1�uw�q����46ޔlO^^	���IM����Ak�\CC�w�}�|��%��C(�鲓��K�_��,~���q�\�߉r �k�]w������H j��3����@�[4�j�A�ᆪq.�K��h��VD�B�}�1b���E�S�`�M�X9�� �j�ѨjN�\A{&S<-��Z^
�n���G�R[C7��� U"q���?Q���$��Ȃ���91�XH�X����G&�W�N)�"�R	�X�n��/�},J�֩	�сo��/L @�@����~s}�].��6N�i�2(��f�TAA�US����fy������N�����r��i���8����HX,��.$+���̓�8q��;Fv�4YƎ'�LQZ[��ҲY6on��x��f|FA�h���O>���illT��駟Bİ
 ( �~�����G/m`n�DS����@�NA��k]i�����s�nL���D#��N1��
��pQ��٣ɴh���ҔF����fc�*�e�xI�Y�G4Ɯ>�Ez�F�bk4^��c��3��(��ZKH��[�C��ܕs{i���\@ohhJ5`�*{��k�.�{([w�y���`_�P�~�����t�"�&V�J�n���"��YY�v��X�\�֮�J���Je8�S.���z'�[�gNc�-���%�4�^�ؚ��"�J@K@� +@`��"���ʩZh��l~��Ԇ�BVl�c�.���`IahF�{ktMY7��(����B���-�6���)�ઍ��E1��r���"EpÚ�[Q���h������x�P�P@e!����I|ύ��U*a�`�--����`q�V��O������'�Y��	|�����Lk-�vMS��������5�<[�4i?1��k�߯Y�ܧi�(Y�� ��Z�~�i����I�$w���to�M��?�>�����̿u]3!���YG+\�a���^T_#�g����Ȏ�N^CE��j�P��ҕ9��<@��tJ�o���n&Ο�Ë��;�s4������Jv��	zr�i�Gi����F� ��Z>����| �WH��m���!� %�+p/}��n��p^.z� 	������%V/ޢN|�|�1XL��s~9 ��FeP�pŅ ���=h$��mnݢ"��Kz,�B.�^B΄{�롅㿢�N�����˪�Z9
n5���z�)���u����_�@m�@f��,q�G�PG�:��h�֢p�X������2��:��]�����ޖ�����ی�i��)�
�1���p1@ӌ� �@���O'Q?<|8?٢p�֤�<�[h^��]��Uz ���瀻W�@_-�-^[&ܠǀ+��ZVV��IT�e-�$z_N������c����7��'�O�:a}�R��i���[-״{��
h�\ֵ�t����,b�Y��+_<�ׅ�|���z_`��û���,�J�P[�(W��qƫ 3kz��a1�~��&J�T�=|���A�?�A9�c��K/U@�o�x8A��"G�h�Czq��r0ƔI���}�`D��@i5�Kt�o�M;���(�JZ�3�\sj��X�l(8@�l67�  O��
�ق��P�[]4�7��0���5|[ݴ�ܒ�\��`ӻ�x	���m�KTSp�����?98�X7Dy����~&����5��E�JQ;[�oL)��>��iHBt�����n��Ÿ�H�p��j���:�4�H    IDAT^6�����2�+�5�K�'9�zDd��b��c�ҺY��j�X�{3��"�'d᳧���Ju�Z}.:���#��t�9x�G��6�6Wt��+; ��`�=[�}|�|;��_�K���7.��V`����n'��3Yՙ��d����fZ�{u�Z��>ڲU[��>�?X�zەuc�����7x'h���m�WI�!ʧwc��p��1�w[��J���T^Vc��%�k��_恵u�ŗh�M>���&	���
�Ma�3a@EJ4U�	pn�QiBd@�Fnf������)��oq/�X�:��t����S���1�����o�� 0��>y��'T`�z��h����"�����E�Q{<C+�`֎�OF��C�I/]��:sQy�·o�c�>[������ι9�l��o��  ���X���p �x����X,�.O?�^~��׭ҡ�c@0��g�}s���������ӁƯ1��a�Q��������"��G���;�('�P��pf������b@�o��
��'��¾l��Y�uiA�Cz����}�l ��?�x	p��d��p֟�S�'%��G������W��͌lo��Qg��4wb�*X 4�D�'���R���_�}�����@@���9��}� v@��G���ZtE��� �~���V� ���<��C=u�IL�s&�h�����O����eԉ/ }��Ea�ꄘ�"8,��L��/��m�;�;�T���
4P�Y̹:,:�D��:�0V;�؂�q�����cJ�O4`ͽ����;�*�"
(� �D����o�� �w`���h����?�.��q5˭��ӈ(p�B5RR���&�O82�o �y-'d8�i`��O�:���&*f��U}���n_����e��$�@���k�6�̀�5��B7�۲�}F@��7��+&<��nA�8G��=VYw�y�Sm���f.�&y��O����������MJ�b�3������a��LR�ke!�>�lQ[g�;�/�7���J����~| >�n�(e�z��Q5��¬%��Q�1��s�å�]t�}�o����}I\  ��唺/�pm���������ș���?�����_3A�s�2<�4�<V5λ�/ � D���0�(+NL: ��z���� ����4\	i���V2
�ǜ�|��?���J�H��!��A�x��O�Sy��ϕ�f����5��R	���uNc�k����RþeW
�E����?т������RN�����Bä�.���-�@i��h�ij7�l�:��6�����@S��z���s�/�dN5{�&�M�0��ie�)�f!kV�m8���n������r�>���pL碆�=���%[�J8A�4����0"�BX
9�/$R��L�Dc	�*/mW��_*'���B?{�y��8.?���8����KNK[8�c��I?���eo6�EI� �|��@ͨ�lxr m�g�]�����a�a�s�lH�9�#HL�<;~�_Z\�{!�s�� �K�,�I��Ϲ�[��3Ӳ`�Ͱ�Z�e���s����d7�d�������{F�1ɦ��Щ5��Q����̿c��y��:Zp�ߪ��¤ɓ.Zpׂ;��q�)Ù��w�6�ؖL~�R�'fN"~])ˠK8 �q��a��ٿ�]�͇fO,���k�+������Y�0�!��6��5Sq[��@c6*��}b�)o}Ѹ�t�d#͔%k6�I(z	S3(KW.%�xL��^��6Q�VsQ4�ׂ89��3ʩ�.kkH�rBݜ{�xUt �͒�*<D���^[� �  �Y�+%Rm|>���-j���c�Um0��/~�EȬ*%�t�Ȕ��B�t��̱���Z'�jWe����Y攥�.��Z�|��֪]�,�r��k?��1A\$�]���ح��+	�\М������`�_�F�;����4�JUOJ�(_t%�'D�g�M�2MC��؝"o�����^�|�K^iO�F��c�Μfl2�M�}5���˂�Xk3K�a��U[�&�q���������E1w��VN<���6�̉d;3RK(�Y��$U�H�X��E�%�l��Tid������u�����й���F�VQ�8�m��Tm�������Ǝ[�!��	�4zh �V�U��������)>����D?B��¬v/}}�=��A�;���>��7�!�W�����#6'��Bm|��9Pko[���y�@��+,�#1a�+f�k�� R��y�{�5#�a� $<��%�Y��VUJ5K8Lq�ٜ�(e�WT.F��?gn?��iܑ+�dS����շ�dRZ���C��8P�O���@��8��^xi�����Z�ro���ݚj��y��dr�jf6��a�Y�C9f8�����gt�J!㣥4!~�	0*�����͇%F�|`!+��uP��Ϡ�@��_*�a����p){[D�k���ԓ�V�֦t\ȅ�moڠ�|0a�٬C^�	E�0%b�V�l��O��F#ڇ2$��n����%�O�ܼ)A?����2����]ˌ�,��?^3�V�����h-۷v/%N?k��9�� ��w�]��{�}���N����K{{��{��e��Œͺ^��TֱA�J��

�]4��;�R�:������ɫH���l*źb�Tr�a�hݝ���S+���,6߲	y�񚄴%;d�UkBR[\��mE��/Eܨ���c�ir�J�/	_ֻ��6����K�υ\�����.W�'�L����3Q*#񀟌�Dr���t�R���|1T��C��Sh�oξ��B=K!���&\��;�Nf��R2�ZD� �q ��0����Yw�%��Y�J��+b/+����/9��O��yC��_�B�q�R\�똓�|ù?C��ZG��w(g���N��\�=�9��bn8�	H�S�_���޴��#��|*<���}�q:��	���K�6.�tZ�@&��g��U~�Qio�T�ɯ5������No�^{[�>9�F�Y,JM<!��V�={7�䒋�e`&�a����SO��5�����{�m#���J6_�g�yFc�-ӏ�/��6������A���~�3uH��+����d��@Y$�Ql�u;�SW�P<�j��#����	Eb��B�I��IM� ��aɤ�$^�L!+�X��c����A��6*�AK���� ��j�J �2g\Oڅ�U�AM�f\Tyd=�X�o%��B��k�s��À������Q�?k���,4r�܉'*��7fv/�`ʧ��	&��#)���.�0�����=k�Z3������_��SOy�~�!:T�m�j��e�/��!3f�R*ߘ*�_������haT�LGt�W5��9�Ǝ-��8]<h_�(U(d���<%�$�6l��-�ƍ3Zv���t�2e�n2f�x}0����I����9I�[����EL5)����~�#��6-�8Zs�j%V9x[V�t���|ø�J#�;^K �0��X��ĊiɈ�:����W��nA*v�[e��骍Ȕ�M���[`�tە�_^x�����'K�~�9Wˆ� �-��X�o�X�<C�A�`=0椯z6}]���A�@�ˢָo�Ws.�{�t���1״y��1׼�s-���<�߫��P�����|ǯ����|��=��x�;$��X,$˖.�GDk9%;�5󺶾Nv�<UN>�4�y�LIC�f���C��o������=�h�3w��$�mWW��!T��#�K.�PR�.)�R�ʫ�ŋ$�s�(�X�����1ǟ$3f�f	���A`a�7Z�O<���{D&P��/��7߬ܧ��i�Cs�����W��j�_߸^&�oP��D���D$+�LR��V��rӍ�	e�x��g�#;7�(�Z�,%����JqMV3�W�O�GKw|�d£�yY�k哟��$�W�����b� �8���"�|筽g4���Eq>�j�6&����9�~���ܿE�Yč�*�;��<{��A�ܱPp�c�0�F��Aik*���D%���+�ʋ/>/�������b�����%��%'�����Y�����mwܮרV�b���<`R��!�/�lJ^[�P�lX�$�74�:^�Ԥ!ʆ��;���TH����j�Z��#�<��$��D�G ` ��Oa��ú�DYT���+,΋���b,Յ�^{P��x^_șF��& #�M�0n�\����œ�	�%&]͵J��"�L�����K.OrRX�4ΓS���h�q��_��Co��~U A��B��;�����l^���~�����߮�0+��
~���`�E�Yh�i�vߦ)݈������ޤ������n�F	0�ǀ�w�o�Է��<��E�*{�֬�t���.��Ȕ����L�SR��e�ڕ�a�:Y�����N('�C[7wʆ��RW;V�zϹ2k������������s���P���&7\<"���̝��d��#�45�����U2��F$��_��^����%��U�WH6�rE�����eg���D��w��o;^{��`q4A� �l(6)�>�Na$:B뀈"��"��h�9�q0��Zp�ݶp9����1OY������Z�F5���)��/I�8zIB����N�����&���ߓ\�[�Ѹ�i<K�M�-�|t�௢�^yu��[��u�����L�Fƕ
�1? ߂{�|p�U-�
��=���QHe����{)�}�yM�X����	���P��Ox��vO&�8�w W��r�a@���57Ա�I��snj#A�|�+_ѐU�a��?�����ʻ�<��?�S���'7���>&���$Y�f���V�p.$�tNV,o�H�N6nL�1ǝ('��?���^��%��O�o���Gn'�*�O�B6'{�>[���5��꒮���}�rһ��b�G�4��Q@���I��KV�l�t."�W�ʁ�5�y��8���Э�;���A3@ۇ�4��6���
Vv�8},�e.���ð�B B���{���-�&�T�B�����w�!����$!�?��$V�h�E��n���}�����eΜy�ӌ�%O��W���ުm~7���.+�ՐK! ��=4C���R�4������]E�WP���]�#6e9	�4���O�X�A�'�0���<M�)ꏡ\[5�2aPm��ތ�7�f�0�i���s�Y��y���/jH)�$���sP�xAa��p�z�ed�����
��M��Ϗ�J��wW�0a�,]�DR=���LQ^Z�D��'JSS�4L�.W_�q�������X����-�����G,��vz�w�ے���+�
��n��U�R��>������C%����HGgR%,}f[6%��i��N��h��<T�z J����}�Ta�nB8By�L`u6��f�F��z�D�+Ui�V�Tw�F�u�Y��EW����� ��8d��xp��J��qh?G����-�~�
�jK�b!,�PN��E� �o�����wϝ'Sg�&Y/%~p���f�'�lU�i����[=k����W�������@ɞ�Qp��E +��h�*�O^�L�[��� ߄C�1V^v�rJ���E�ʩ���R�-�g��k�Q9����?�i�+ <�[Ț����<Z_�җ4ʏ}�g�}�҈�y���SO> ��L�0V�-_,�T���;�e��ՒN�ds[��������F�+������?����YC#��46~;ٞ�XE��Y3f�G���$�QiٸV�ӯ����p8%�ׯ��֍J1Dc5���)�[$����u�2}�n��O~R��L�u�]��ll&�Y͛7O31�������$n�\�b2��-�8�*��9v���{�:�D�X�����X% ���u���)�>+�ʲ(Gq�Z?�A1.���
�;Ϳ��N������Zy��g�ԝgI��;C��5���6�}���F�G��>������9 �hno����`�?XW<����)|+�5j����JM4Z���T�P��}��0�V( v���j�;������w�Y��'��	�TA�Pv��i4�F�S���6�oʔ)�-W�Z"���>��ݥa�hy}�2I�;u.�+J1&���H�^��9�������_�DM��(��?�ח/���✹s��L��/�W���ҢL���|���H<�h8/�T>ho)�es[����ꦉ��=���5�d��Y��SNx�)2w�\��l����'[l$�8�I���eQ���� �-����Dk��PIh$�;��R!�l�тF�M�O}J��7�������DC���v���$�����rىb���-7h=�p�^N��?���:�������k���Y���n!����X5�j�3�ʱh�PD���|�V5�&��	�ٳg��F4~˲-�N�Ž�ڻ��HM�����)(6vߧ�y�{&��V���*�p� >N_,gzPn��n�����3��g?��ww��SO�Fv�e�����U����Q'.AX�.	�H��69���e�Y�HM]��Q�z�J���y2�gräK�ϟ[���__ح����E]S'����-��!5�<���2vLTZ77K&ө��<�I��d�Ƥ�i�,m���+�Y4���n����o����6.)�d�ZV�ղ)����%nX�E�P�j�x��<����(��s^Uƅ	K�x�.��LP��f��a)�sr�)'No���OL�@$=��&�)��o�;o�A����i�g���H�8�Ԟr��^j����4���L��1�޴ȵ�u���/�Ɂ8�yA#P�� �4?+�փ k�5J^
�4� �|fl����~&�����m�������Z�q�o̲���e��ђ�X4��_���g��ǔ��N��%��l�[6�4���O�|(!�6u���kecK����d��p$"x�O�8��t4A�����_����k�q�G�|@ҩN	�Ҳb�bY۴LB����0ц��	��²is�L�eO9������Z�������i�?� ���E��ԤZ6<����M��$y�:O�R_W���7F��DB�r���fiK[�R�Ԍ��lA�����P$�)鍧�K��;S�uǥ�3R���-���;�'�ߩ3f�_2�i��6C�M��<���8uU�7���c�'���"�L���:媫�ڂK�@8�s�_t�E�\�SM3C�T�4p��N@���~�ܔTF�	�ZQ�G��xs����(<p?|�����%|Yة��T�d��l�{����\z?� 7���ɼZ$�|�C���l��j> ��;���
�Y��"�Բ^
���ջ�n�V
��,[�$;M�.�x�I"r�P�k�dR����'Mn�l�]~2�4�j_�,��y���������)�\V�z���<)���	B"�e�<i���]�!���S�5�
����o~�	o���_ %z��g��X���e�Z�5�bc���J��U�I	'�?�X����
�!g*����"!���:[�q%a��J�q�����~����K/���~�kFr����3.��?�W-�j�<��s���*9LK*����os(k�ݾz����o��,[[*��GT��M�lx�>?4dӢx>P`���_�܁�P�cn�u�*`�Z������`%� 0��iԈj>`e̕�c@��8��s�OV =�q^�!�,ɑ��mfB��"֞�� 2V+��t�2hå}l̾���p/���P����?�Q8�n?߳,`��L��1}����Xs+�.�t�GǬ�%^#uu�d�]��#ߪt���O���n��]�j�W���{�����2|��O�E�`�Q�	چ����>��j�(6���n�g8>���+��( �w���i�(����v�M���ok� �C�fX3�j�OooY�h{i��U1/�HDk�G�Š-ڹ�x)��AP����+�B�h��$H�
V��z��,ި�%���K�mG�Ux@��Mڹ�y��k��Dr�r�-�ӌ騂��2}癚<d���9T����0�PL��'>��>	hWW	.��-
�����@��>p�* �mp��    IDATk��&���7��u��h��#���/V��^Z�p����~��G�g����̾"J��s<[ȭ�B�%�k���?�#t�$S.^�Z)+8̧�|�߄)
������gF�|?sl�c|�#�Ep��1��fT	&��a��B�{3G=Y��~�3�j�ܴ����~�z�Eۣ��+��$��3�h����c,^k�d�Z��駟��k��4���� ���4 "X�x��u��jR��BAM�bT˰����G��Z$�m��R@A-�E������\Ahd?�O���_*Gu�V��������z���yN��M��p�$�����&��j/_�g-SX�4,M�"������ |��!��ZrbEdQo��Z�L������7ARm��ל��@?�1��/|A��=L('����� <��K��I�:Q#,��s��!b���D����b>+��wh�}�@����\rnY�����!���uڃD�g�P���<�W���=�����X�p�V���������ϗL^�\��ˊ�tP��zݖk��|Nj�Q-���~�.�K#-�)��`�B8T�����2��U�����S��4���4�7;�w�v��ш�� ��'N{SK�
�lp� �� �X��}H�k�������v��m|f��� �;��wܡֵ�a�<����r�[,,�
͟(����O5�`��Y����f��v��V<�=> � ZWR�Ǭ�� ��������:JKD�]�|�w��P�
�C��a���Ϳ�#���1�����2��Ĳ�X��e�Y�"�3�m��u�^ܯ�c��]q��p���,�j�8�~40�3�@,�El�j������6ܾ�����I����4&?Wt�xE��=�?�գ��}�A���ϣb�?��(�(�or����F�F�� ��@��}~�NZ4UA��������?c6�Ф��*Y�80�o�k�kXn��?B��g�ؗP��?`Z�6��傈�s�'؀�H����&�/��BIq�Z|�%`]�u�����1c�j���B�h>~���a�U:ۻ��������t�Ι;����k'��Y�.6̀��$eaqF�w��O:7���/	���-|�-��P�;X��@�-���>�C�@؄
p�QI�H�����.4w^�܄�����4�j௙����>�8G�>�������i4Ž��{�/�9|����g�h������_\��v��m|�4���t�w*M⃿s�;%��
6͟=�%C�ǣ�C���?�����/ �|&��M���m("�Ц��1v�V� ʤzJIZji�M���ʭ����b)�7�2*��N^#4ο��d{�r���s�ol��i&��AZ9�ɷ0N��i<��o��,�dq�!��ބ["�z���y���8���P�װ[l��4���?�q�h���p�M���������5ZY�h����\+� J�2��?������Qee�.��(h�O�~}Я�����?��1m�/���"�������1`6��2>ބ�Y�������-�������7�Z^6V�5�r�+ױ����ƹ�?jK&/��&�m���<��o��k����w{�v<��Y��%qY�-t~�>�[A��Q��ĩ�B�9�q�.^���M�/Pp_U���}x�,h��q����ڧ+:]��1�o���i�����RS|MD���$�ֈk�u���LR"���3Գ��7�Ǣ}��њɏA��e��r��ڱQ2P��	U���t�6����iS�6�xߺ�Y�$���ri�����m���9�y�ʼ���{�
V�k��_a�̝ss2�~i%�f�BA�0p�T�຦hT���^��_mCb�
̴R]_/y"��!J��x��L��X\2��d�"�0�D�.@�8�[A������ΔS�}���E�@���h��>��{6.n��z��WK(H�y#���'Ml����`��U+��'#�N��f���LHl���3��k��i5�xȤ����󀳼����m�vaw�]��A��A��A4R���&Acbc��I�Q�`��&%	b����ԥ���l�;;����{��s睻s�.;�J��������k�-�9�9Ϳ����!%�kF}�9>�|QHϿj޼�_�I�%����Fm��%�5á�N�ܔ�ɿ}S�?��6fa)Z@בE�@�,I(Q��H��Gs:�cZO�h�,喖���%ʫP*Z�R5�������Th6]��+������V�v�ε���\�/9|�}F@�n���M�(�v��~}Y�M4�a��Z��V��h� �Ƭ�F��|�
���袋<�h;!��C��j+�o&|xV�}h���F�����^� ��x�o4WR:]	{�4ք�s���;�����O@��Xf7��ȹ���6u�5����%�R�m&uX�Z�l.8�� ��p���eZ[lm�z��h�j��?_1�?�2�P�bs:ϱ����8|Pr��ܣ}����O�������<շ��� �������LE7L�?�>ǏF���u���B��{z�����%�ܾLʎ7��	%��Q\X����FC���9��������8�I��;z�	�����J>�s�x��~��i#��8�CŞ���yS�X���T�/4�UOq�\R��l%��$y�����Z�>K�zp	���A��������ߠue|�AAP��R�j�~S'�%��t�3\�
ȎMm�;֚���v `b��5Η�#�#��N4��*�������3.J��b�wliku�u��Ͽ���xĴ�"���hA�s9�3Np���|���M����#m&6�M@<�����,�ac�h�x�����-����I�!L5�#��*��[X5���+Y�J�}�m�����3�i�Bۉ3�8��r�EV��]�_p���C=�?�Xdn���_�MH�(�E��P�f/�'M>�jDT�X׏�n�{������Xo�C����
��cy�0�^�Sۭ�lh���'2��9��4��E���/�����V�o0��t��5{����ҠK�ġV��q���P~G��b�+�k<�(MχD9Gswm-�,^"�Z��ʹ�{6��įJ!�����]��L.���J�5��H�/UҞLv�)'�e�����3�-�"�'����"�������6���o�Ǎ�}���B�KȺ���M]��KqX*����v��I�Xv�B�u�l:���0�XWZ�)�c/�J���8��ⱎq=�SO�	W�Y6h����x���� "���O�6X�B�|5m���D9(�wSP3��뵃^�*;������L	��=ے��׮��]���߽���x�0k�h�T�|�	�ٕW\��>p�.<��q|yv#Գ��R��/�'��M/���2��V|~�p�1�"�?�"cZAʋK�/�����h�$�G�c�����5ݍ�JH`�C2}ϦS��M}�?�y����4��1���=��Ϝ5���o�����O���Ku��\RB�0;@����o�Cʈ���`1�/n4|
�Qȉ�Ʉ�@M@f<�F�?ׄ�)��v��ϲ9�����Vs�fq�fF���Yw�z�����z��{�����Y{�X�O�y��!;��W�UW_bϳِ!\-ZKe����J��s���iU���W�3�c���t.�B�� @A󧄂�q�#s�5������(�&;X��W_I֬(�p�\@�84�,��]2ӳ#l�7�c#�����*����>��@��G-�O�'l�$�������R0�s-�P	<�/`
�#h�0�ͪzVK3g�x���fq��c[[��f"r�
���a�v�y��C\���t�Ig�t3�����͛�l��LUi4 ��>�!|�{��@�j(e]��ߴ������F��JR<�1{�l���7y�>ז���j���3\qՕV*��b�h��p��d�z����r�Q���5=`�r��U�[� �f���v�yo+��V�T����A��0���Wӓm�u��KLOp�ui���5�`�j ��8�\o������̈�\2�4V��I<�l�/�3~��j��b ����<C��#A*��`�
��8��C<�u��h�D�� �)W��#���O<a+W-�r�j-�4�
ax)��G�q�-�jub����}���/*;Sj����zՁ6iR{�$
�ļ�y��/U���@���뮻|�dV�V5o�6<1�h&D� �|��ޡ�?	;���aƳ�Y���Ѵ��n�lB���>��������L��'���כZ ��
Dۭ\��L��J]I3�U�͛>����L�ٝ�ێ����?�a��L���nV�NVP�����~�%�U�g���0vZ߱,v�}�9}6ָ`�r�r���Z����EK�BG&�;{��9^�eŚ��R�8��c^k��q��M�p�Jh���6))8���k�y������B�`��ϴf�ђ,�$`+�'+fvg���=�kE�Դ�JH��q���/����5�b�`}��}r����͜i�����=�2hȿ��/] h�0�u@���c�Q����3�\��뼪'�%,b����Q����k"ph�'�P59�c-��P��Ѿ!�����nSuJ�ͪ�3+�Ղ��^Ye�b�}�Ϲ� M_�ﶓ+#�[�ol	lP�2#�9�����VjٶֿVB�
�$����,�3A."-?��a/J�b��aQd��5>�	篨(�Y�V6�����7	%�1�|	�gǲ+�{Q���9ԭ 1��׼�Zr���������f*c����,C:CK؜�E��O��Z�iߘ����Z�К�9�v~��;}#��}@�6�LV����㏵r�`��m����k��8y�n!���v�񯱝v��
�Р�ʄt��s]��G��u�8���?{�w1��5���as���FĢa'�X8��gu���6�O��]v�e��?Z�g�j�b�r�\��]�Q^e����͟�J���?{ι��n������V��ץIR�: ����.Vi��c.m�1�����V�t!.�\�k]+XB R�&i��˾�}�q(n������jo� ;�}O�q�o\L�Y4�>�o|�y�˦-C~M~�=�Я�_�<�T��ε�Ge��q��N/R���ݾs˷���V�X�q����z��74�R1^��:�����k��bi�2���X��~�z���V����S��p¤�מj��� ������pg0��'�OO,�R�Y 4p�q�<���G�g��g<�����(�+L	�s��$��IH��ў��
GWlֶ�ؿ|���:"O�5W�\����W��o�w�� �v;g��t�s�5���9�T{F�y�����
�l\�5���㙻?�s�*�k��M�Ԍ^ �Ϛ�?���8� @q,���ԱT����:�q��g����}�����}�q�{��l�vKW
�j�2{�
�5����!�r��'Y��SՌ���cg���aͲe��%	���	�1s�w�z�����O>ڧ�����ο��gҡ�+���;���-�.��yOY_��\�Ժ׮��g@�kw�Zg��e,d�]7��;�Y���ַ�A���B�w��S,, �9?��3������cNqS.�)KRB��#�,q�Ҷ8g��CSH�,�m�N����-�	!��R�Z�U�V{-W\g����߸���m�s:q������sd�R2�[Ç�s�HX͍��
�l���_A_������l ���j���O���O�aq7����D8Wt���P����3��~�;q�����?ֱ�p��ҬH��"�d*W���Ъ�O�V�(����~�"5g�;�Ӭ4�o�}kl�����m��.�e�����T���ݽ�v]���~v������6�c�}�;߱_����'�
�fw��9�����!��������v���K=�e*vם��1Gf}�����g\��j�[�.o,���ڲU�v��'�\��ˤ# ���ڦ�zϸ�hw�Ue�}��x�����{*�&֬�����X>��a�Z�)�-�O��uLF[Iy��ʖ�>˖�Y[e�Yq�}���Y���X���l����
�i���Ӹ�뱗�~�ӱ��Ib�{�i~R�:d>�V�}zZ��W>~2>���W��ǳ�F��Haoq��gu���-$���4z
�3�{�����k�j����7�[�����i`�_|ћ��4�a���3�K�=kJ%,xƏ�㾮��2��㿴�P�͜��=;�i[���{�
u��E�ʴ٪�n;�����ϲt��~��Cv�w��@o���hkuBk��tv�SOO�Ɔ�5��*��]��k�=����k��w�f�q���Ru�E�\_\���A[�d��*��pq����������Gc����8X,��;��}�+�WZ8���ŋ�O�bO��9�6u��<E+(tT��4�X+��Q�f �3,��ђ���Gl��휳��JѲ�!K�z����T�Ǿv���S� ��Yi��W�~ɴO<P�ų�ʈiJM������g��d�>���[���O�����'��-�y�3oФ
z�#��z�OIg8t-��3Xԛ#�^�Bk��b��
�_vɥ����}v����4�~��&��k�-�6Qqt\�b�=���۾��bS�L�矟�ډS�ٜ��y�b-ֽv�v�y��򫭭}�[7}�f[�d�V�o�@fϙ���|��������o�\{��Re[�����e��z��}�յ��z{���U����]��?X�EK��+�;������c�|����BF+�ē�'��{�mT6��O⋇��vl4��Q��{���U��P>�=e�4����Wmr[���!K��<�kš>+�)��\K��������v�G$6BbD�n ��,0��|b�Xf�+�v���RSt��h�/��'��3k��o}�7>G�˗��%�?~�����X�ƲҮ��Z;��|�1o����󛥜�����I��}��uk�zT�BTIY�?��}��i�@��g���{�q{��w��G�	��>���Z���Y�X��O����|�������g���]0|��_��_������HMh���9��?��������Nv�uW��t������)'g�L��?����>�����l��%V�v{qI���+݁��ô}���_Kؒ�/���ooG}��s�9�Ezǝ�s�@5��&����n���8&�%�9kC��p�'�(sV��j��բѰڥJx[&kE���]3�y�b��h����I9d#Rd8HkDZ�f7}9O���F&I:��Yk�e�6z4��6�XJ��v�o�.�x�Y�H��͟��3�я~�Aozӛ�W�j�*��>�яz����>����m��=��o큟�eG~�M���-\�B�0��
Q:�b�>���E��)�G>�	�2y�����׾�5���s#譭����sf$����F�O 6k�v����`�-4#)��}ێz��V�5kWY��5.$hX�b�J�^���dE�q䱮ɠ�,\��#~Xtj�ƽ�T� |��g?���{｡v~�����?��c��@�r�nC���%� �8�˰��L��28d9��V��{���� ��A���}�a���w �7��J���d}lrix<�k`ԉ���l#P�(X�P5dU�Ҋ�c�?~z���������� �F�O�s�y��Y�{���_��g��P�(r�]v�;�|?�����O�����U���w��{�lmm-�l����'!�<b�Z���t��s�}�ʫ��z����^�%'�JK��Ϛ1���n��k���'��L�omi���n����暫l�=w7��#�����Qجh]���W�T,�C<��s�z]��YW���~�����;�?��O4��tLS�s��n���������8�R�c�m�m�Qj����Kg���њ��gCW,GR�ӡcX1]���,%�	�䟁2���ޗ0H�x���@'p�c��lL��
(    IDAT�?�K��(IP58}��f���۴i��+�� �i�8^g��e
�D��p�^~�e��>��5�>�����C=�� �����<��`�|������ͯ���cOe=�z��d�
�Z���/��?�Ֆ˶;�t��_�tv��CMY*�<s֌+o����N@����ϤP��M�o��k��%m��?c^��&Y�R�����1�%˺l�=��#�<�@L0Q"�/���F �����O��a2zz�{�v���/Lڗ��I�Q^>!d�V�+��P�V
OQ�7�T&e�T�J��-�.g=s��?)�7raK�'{m�[�v/�:�B]% ������Fxr��(�F��;��ֈ�C�� �G�����-���W�"<�M������W�}~G��-Ͼ�� ����:�i����V�E�����˭l%k�d������)7c��csm�=��O>Ͳ�V��l��η=wH�ӈ�JJ:_uǭ�~e��ء�$y)
I~������ra�Vu-��}�y���?�×�a3��̘1�Nx͉����y�;��mh�Lc���=���k5u�5�M����s��Ga�,.%em�8�-��]8UCMO���:�4 w�d���0%����2�!]	UC�-���U��� Ц`3�x%��Y�>�^����7�w���h�?�n�Z9
�e������{�5׸U���8�������> w�ֶӦ{�t
5����ş�/��gS�~A��;ﴃeR%[��E����l� �@w���[�~�Pr%e���n��ez�m��Lo+:w�\��׿�B�YT�����O�{��n��KG��BU�C>8Ak�Y{G�
�6�3������h��Z<�v�a'g�;&Mqg��������}4�~����JO� m�����;(����3�BMSZ�c�+N�x�>���f�j�rմe�L�R�lE��+�%}z��L�J�@-\tʇۖ�!Z��X����q|�?�S��ڐ��8|�͛WK��8�4���]w��0_(\�3ڇ{�\[;����+.�k�X���G�M��߃F����[
����>$�N�h�\.c˖,�����}�����w�o�Wڱ�g��S���6~�B͠�R3Z�B�����n��扨�&��~g#�'��5�J��\��:�.��"kk%��6���`)0�CC�E��~�Y������MQ�C3!i���������'�͉G�$i�\��@ �s����e�� ;��sN��g��-!]8`d��cx<�f�kc��|��˄0OYX�ކ-��Sx<�����7Y+q�'mN�$И�Q��Q��X��v��w�Ã)ثh�(a8|k�S�u�a�0c�������l�#��Ѓ���q��5�чɞ'a��5�F��cO>�d;�3\9t�X.c==y���m7é�.ϱ��ߙ|#��p�w�(����5���sN����w4mve��7���W��N?�4�o�}|�x�\��0���g?�(����9*�8d�}�;���w�B�D� B��n�{đ�+��	5�N��6!B"u���8�{�>��zp��h�bn��]�A�(�{0�C�q�x���E��C5��y��������|�=
�9߬m�c�B4U(�~��b�ࠏ?�S�[�M���:1YS�t�]p��3N����˗���w�=����/ae��^�����l~�����ӿ̐�s@d@�f�{5ΤP$Q=$xQ�
�5a�� PQ�
�i���%��jqL��S�AN�Ϣ��f���f%��d&�Ae��H	#������R3��I�fB��_��q���7�x�GQ'\?���ˎ;�8��ǧ>�)�&eQ(���I���j�����{͝�WX7�^������K��i��B6��c�?�9��W�P"XZ&?E�H�H�h�7��?�X|�T��k�w�fD��b%�ȐEA��T%�ap���KfS'O���V(B���ڵ���z8w|�����w�?�������0gP:�~�pSwE��3X��@�?ɠ;�s�?ȸ`Q<�����\����, dBs��s:�Н�_Ӑ�I��2�Z�L�6�IP�1���D�9L��E��R������{,�!�����D;xꩧ�+$���U�g3��lsn�|ˎ�4j6�ֈX'�
bwGwRwF�z�IO-�=��r��H�DY:^חe����P�?�u��x�Մ/��!*����N���1|�����M|(� �Bӥ\k�gl�L/��a��R���P��U6�����w� ���W���܅	<K=hk�@�ȳ�?��FB: c�τ��sf���K�O����1���dVk3q\\S�8h8C�I��\ t&�s9����`
@����4:i�ٜ[�ݲ#�<K��Se�e����ޱ&)������� i��ט=�u�{�4O�?���xF���El��'�7 �Eϥ����R);�f�I
�Rb�^�ʞ� 䂕��A\K�B��<#�f��c��N^P?�>��k�P8��b:NV"��t����*�^o�qo	�۪���zgwv�G�'U#�_�Y�˱V���:���L���f�5_���ٛ��f�����X0�zg�y�Kw"pTq�"�bw<�s�[vb͌y��-��ZІw帎��i�zz��@����k��aL�H`p=S���@?J�ñ��艐 H<�8�`�q�(:=��%z�����e�och���I��TEb�h���/A���~'YiB̕�Z��,v�B�� ᭆJ� ����@�q�-��c�T����9�������|��F��+��A����8�J����-���\p����U��9oٲeN� �!�.Ƶ)���q�18�ڪ��,�X��Ġ\oQp��W�Xv-7)A�/kU��h��2؎k����^8S�����?9��e�d, ���N2Syf(�M3�SVl���%tmů����E#�ߟY���3�z�į"!.a,� ?��\����%@�@�1�<�����K44�+bc��j�R�5c�U4�s�����+�����$ˤ�yZ��Fc��i9G|?�7�o 2��<��^d�����Ƶ����t�s���L��?~js�4O=
�+������
����c7��c�����$\{C͸�Wq@��_�[5�O@[��="K�-�t.�P
NU*߃�	n���H�}�e�fp'�[a(���A�j�["��'��MLw���O�_�g�/xA��V�ϱ~�Jh�M�=�;��'�{�ܱf�9k�շ�r�M������9��Λ{��7�Xï�~bs-6W� P���4����z�������2�!��Ŝ�Kۖ[��C��@JA#��M�	L�f���a�|�$J� 䑲�7�.��2�Kg(^�=���@��R&��c�C��P*�|3k�3�y."Ɉ�"�&�l�X)�G�Z����˂�r�eE�;�b���.1:�g2D�T��	�-������U�����������a�$�Q&�%uJ��p�4w)�RP
�R*bZQX bc�Z�VgΚqՄ��sf%�﹬����I�b�I+��%�%�X�/�q}���LҖ:FZ�6�ứ��� ��5�`��e�b�S$[j�{]�Q��1H�;�����k�}��k�����o�|�����p�KQ2^ԣ�40׺�K줓Nr ���?�$3�9AԒ�o��,$� ��K/�ԭ	���.S$���p}�x�l��WG_�E��T YB�d.��2XE��Z=z�(DT�0#�.Z����fB^����ɐ�V�G�Y��=�St�ش�x׎Ώ�0�;j%D86���SF7	�f�w+������6��ɒi%@�F�F҄���8@ I��uo��ב	-gd�o��&�Hi2����^��I0ΓbPԥb�/��͌��o��o\;�j+N~4�v��������!�4.�2 ���_���[n���Ϗ���	'��?�>��>H� u���E� ���p�O�k�B%YƙZ7�?k�+�&�LLKĜ����α�pl�O{q?��P�)����$�>]�L���P��l]W�RI�j���V"O �V[���L����������>�q.�D�
ԳC� ��19��=�QH���o�1標���My�c�&K��)��n�$��H���Ц_AIk,8q�rR�f)��j�~��Ό�ų�ŕ�"��b�������B���ȣ���[G�Gk�}>'A�"f�iA�@Fc���/�Ў?�x��hŃ@��T傡���}��j�r@�0�\�gĪ �\�k�h掁�@�� �i��Z�B�2�����
1�N}��A��k�b�\R�����O�aKD*�%$ejs9B�O[K��9�J�leچf�ҫ�}(�b8�w��>7e=�t����E!庶�:�M��Jоe�H�7��'��ߌ�g�\�M)�C1�|�{r�2��M6�&De���MY4�����G3�5Y:��M��^Z���2XEn�`���_�4�XS��>����$���_�����������?� ^P6��������~F��: ��H�BB|�_p����x�8�K"!��x!<�}xA3Q�W~$i�γG�/��WrO��O �Bk�H 8��K�-Yh��͍Rj43��y����'0K!n�+�)�y��J�`�,��RVJ����)���Vk�%m���-�
���rnsC�s���hj�Y�(D��f�'�\&`a��Λ�=��7���1��] /
��/N��z �OR\[�!phf�5���~΂���#-8������^,t M\&�g�ӟ�4l����e�������C�w�ԃ�'�ZOh�O>������
��K�U���hd�}������՟�ٟ�` �n?�n�kB��~���=a�5�r��w������G<;U.���K�q�G��1���=��8���m��b���L�c!�fU�y��UI�80���2N	��%�[�q��L%k-�i+W
V�!KUKVv�?g�
I ��M��$�������]{�uȍDM)@@J�h�P�"D
���w�ڷ͒�"���?g�PO9[Ўpx[�qlB"7(� x��is0DV��c#��2ɘ�\�SE��h��=�G�}��~#���黥5YL�hƸP헱!����g,�k�Y���a��)����:��g� ܧ�z��J�_�0������q,V�b_�tVׄʁRB�#נ�V�@2�9�nR�@<� E�i��\-���W���شO=�C�S>p�Y|���U�k�Vm��w�=����V�B�bm�f��Y;%*I�*K�:�g��a�w(/���=g]��XO����2��;d�y�1+.�D  8?q��2va��M�3�q�C���O�	�GYh���~�8�B���0���L��Ϙ9�	�̥Y��(&II4H_6ٹ�ז� Px�����pP��<��.���¡x�E�L#8�-�x˄	�F���_^�/�;�28cΟ���
\��g�6�r�\1��5'�Ua3�����%*ǠBݯT� ��b�E5ȹ����|�r*� �i���7���Z�f�U���Z��O;��8�Dˤ����Ҷ�������3@\�;��mP'h�:q�А�,S����u����ڊ]�կ�j]+��Zmw�'§�D�T�X����Ж����c�r	氖���'�x�+�̹B`����Q؍a(��1}�hMh�oV�G`��
��s�:�N8�P��2���n�ZK���|�,��utLu��{���2��Ln3�̖>���駟��R, w��WOc�_�U�P��Sc/�L �����e,�{�t��
�Sē@_}�.�Q\��=�� 8K��zNC&�8BD��d�i�şK�������_�Z�c[��5�nf2U˦�V.��i'c�{�IV*�[*M�i�Ǟ���@��5�O��Rٜ�R-6T*�50�+�T�h�){��Y��+�h����k��?��m�]��J�^�)�9��4�VHyd�Lr<�p�y	N�W��?����;��k�S�T�U�,m�&4�7��$��*!��s;��o��P�![�b�����قE�\.��D�;��C�SN���lk�v�B��tcΎM$�_�_ٿ΅��A��sbPP�q3���P>g�vz��{�s���|�Z�W��}B��?�K
@����]*�������6�4j�6'?���:�F/͚��lTzAsͺ��(�4u�g���/����@kF��^ti���(�_�g$� A"Kgx�|=#�'h��n �{���٩'m�j?�>���l�v���<CJ�t��Z�m��1�Z�H-�ݷ��Y�n��"�m��Gm�o��RC�*g���h���w,ߛ���Z��=���J���-Mt���[�i�C��d���Bi��j�+�B����ʷ_a���a��y��.��ϡ�at����;V`�����#�w�Cה�P��'4�7��_�(��g߽�?��&Mn��U�����Gg��5�kQ1LJ�[�v��Î��:�'��&�0>%6q<�t��ALv'-��@m&mQ��EM!d����أ'�V:p�4,�x����	��T��c	2�
���" �!�/@�˺�8]WB�ϤM*�?��ba�k5��e��Z��H8�&�6���&`��1#��!�3�ϡ�U���~�s�k�ԓ^m�r�����mmڶ;��`ي��M���e�mV,T����1c�M������P���gh͵Y��gK�κ�.�j��ҩ�u��ؗo����X�rV&��7��g���X�g<'�G�[Y� �A�-`]��>�(��u�㼟5c;kɘ�p|rr�Z���Ckٌm��L{͉����z�C_p��9Y��Yi�����|���F�>���ʦ�6{��v�i����=��k���^m^x�z{{<b�D��F*e�Ww���C6u���_��ӎ	��~DgP���#D���	Ĺ��o~�I8����I�
����ϕ���S+������|ST�P��w�ѵ��w��a`�������@1S8fY��.Y /�'*�*�����
J�=�/��"
(~6	.�d�����xw���NT��e3��}�k����J��*Ռ��v�Y;�DҥlҤ)�΄օ8|{{��\�����v�P �{lh�ZrE�Z1���4�c)k��]f7}�[��b�T�U2P��T! 4t��=6��Y/�5�
�V^���}���3J�J�s�8�^RV���.[��{�鹶�7�t�?T,��@�֮[o�춧�~���ʹm=��[o�x XF�O'y��}b�z6�͔I���iӷ��2���w�=��+v�R��-z��}\S��ށA�Z�e�r�-�׽�ӳ5�8���-��ވ� �����pCy�������/x���!�|,ir,����j�c���Oc.���{hl>i��$��<v�BH���c*�O�P�S�0�"�!v��z�N��K� �yLO�7�*�/��{Z���;#g�$�3���<�4E�o�R�>{����I�=���>�fZ�c�^��nX[K��������R��P���´��&O�/�io)YO�E��/5+�[&�f+��K7�a��a��"�ԁ��y�u�A	c\Q���%������2��>����m�f�>�kKY�e�[�x�w9�500d�m�mɒ����V�Yo�\v�t�V,V����[n���h���&4�7��K�1lםw������X�w3�?�y����c\SX�|�5Pu�?���/\l}�f�W��~�b�z׻  z���Hh�LL6� �٘�9��u�U�\킀�!�nEn����8uƂ���?6�v��f�c�޹��6�w�99J�Ҧ 8�x��f��`9�b�&���u�����t��9c���Ɗ�QB1m#��A4�^]�T+���X�H�q�;�3�v�%{%Zt-����
���N������'a�r�U���.Gٔmw���oZ��B�J���th(OC����X�0��{��Y����׻�o�d+���7�ak֕\�SF�	�    IDAT�����_�>ߓg`�E0�\�`�PY�ˏ�dt3�(x0X�KϷ_?��}�����Y��s�u�;x��l�=�س��vؚ�}�������v�k�+W��<�ŋzm��"�W���s���lOw��F���Z.�>{�e�|�u�Mm�������c�y�ў��l�"����	�d�֓�%K�Y��j������~�����v !�����y����L����H<�y��>��x�v0�C�9��scC��[��r�4"J�F��{��>��̝�hb*@�W�t2_
	i�Ҩ9^��|��/��:�,��U��}E=��~=��Gk��R%(�N��_^1=U�p+%IЮ��Y �h�T�:�9�N<�(�z�Tm�=�:�Z�gY��/:��	`$w��������� ��YOOޓq�����Ֆ�-�j���{�k߸��v��b��MLmE�RԍVI<���d=u�Q��o��6/����C^y�^}�}��f�n%�Ս"8�����_�mGq�M�:ٞa��*EwDS�(��g/.Xj��$[ݵ�֬�O��=J�ZM���{���|<�-�a%`��o������c{���X.]�%K_�_��#;����R�ŋ�@G�˶8߿h���ڳ/���~�Wgd�����?\�h��ꪫ<��+�q~��pΟ"]J�  �(�J�l���q�V��ǠG4�Nr��$��o�� �l$H�o,�w�e����˚a��S�� ]O���|�)��m��@�?q�|VuZ��)�ɲ��� _����	�RB���[b!��#�w���W!�
��5�,U7�v��N�לp��J�VI����l��if���0�=X�sV����RgK�����2x����P/��
C�V�H\%m˖���[�ۖ-ﮁ����o�F�����b���_�c��O~��W�r8�x���|�#���z �������~�=;�l���J�h�\������-���Yת^�d��>�i++V)��ӟ��-\�|�*���X9���\�p�V1C�Y3���|��V)z&�7�q�w����UK�o}o����D^�p��*-�pi�~�1^G�����(�t��l6x`�Wac����Ss�=6��Hӓ8h۪�7����? ��;@2wp�l�_��מm)�Z!���UV��b����/�ιd��X����,rBD������B8��X��Q X[��v�\��ƽ�YOj��#Z��F����G���R��R�;o�T�,�1�Q��]��l������9�
C��ɶ۔�{Y*=9������\�t�ޝ���{�X9+���0���a�������
�P�ǭ��B��5��ׇ�|Ya����{��w�XSO	
������^W��f�c��"�W�Xh���ǎ�Î3l��'j��Ht˶�ܧ�Y�J��m��N�go�¦M�i]]��N^�腭��h
�L�J��I�f�d��Km��w��\������Ͼ{�`��]���4����x�R��Zo��%{Ӆou�`C0�ԭQ�8����cs:/�¹3��h��).��7��V�o��f�% H7��T�C=T�×FkYr�rGE�����
@0 ZD�!���zj�E`��gb>w�K�)�A�?k�{B'��  ��L���r"J@�kp�]w���p-��~yQ/�u�f+�(4{ u�_JX������W*���%����jf��b���#Z����ed)���@��U���r[�R��[*I����c�D�� 0N15w�Eفh�W嵳P ?����R���B́�&��ŖIlĽk�&������18:�l��նx�*��ڜ�7�QGo�t��>���緿S��}��U=u�J�&��3O�׿�4*���}���l�e���L*k�\���Zg+��m���|��j-����"�ŵN9���j��{�q��a�c�N��x��s����#(-Sa�lZJ{ �R!�����<�N�����bߍ��f��W	��:�ی ��Z9�ro9��q��g���# }��|�߬)�G�>פ�3k�sE��i+�D�EMd\�H��C�C�1]�G�����p�|�G+/�<>�R��M����J���H����B�E%�s ��f�3BI��uPM	�I"��$y�9GFio��G�n���<R�A@q����q�E�\��o�r+��.�[e�kW���-זAY�5k�=}�1y���^o]��-��oo~�%�݌�\J��w|�~����5Дc���������[�\�?�r������9�_����6�×����O�`���ˎv��o��ӦX�2d��=��Þ���i���l۩����w��;ʆ
%��@3d�C�F0��DBew٤�+N��墕�!���G����?����3��(hȊ�Q��;�K\U1���#iD1���hq��@������ơ m�K���h��%A=)	`�U�
�qM�����x�y���`�p" ��{�zR���� �zQ#	3W�+������'Y���ݳ5*��y�н�
hᐸ݆'
�L% �?k�U:C�^A�'1ܴ%� �u��ט�g}0�c,E�$OB�����c0�(x�;��x㍶��)�^�d�-x�9[�b���-ז�l*k�C�6y�6��:�;�H���N��jU��t�Ͷj�jǯ���`fwv~3ߓk�hB7����N���>�.��ki�X�z+�����'6�U�8x�A�ٱ��i礡�~;X�s���J�\B����4O{�����'_G�� [���S�WR�X�������U2��#�H��[���}x`�`�5��.?�/-PU,9� �@q,稜8�����Y[�8��(%\+Dk��*��{��f]J J���)��
urj��֨k�������Oi0�.Y�5���(Y����ܡ����h֠Jl]���U16�����7�D��+�(g�X� ���1���1c�Q
����lp`��Lj�+���w�e�}yW��:m��6u�t;���m�]����^f��q������En�F�?g��������S0C%�8��'���:�u6���z{�[kKp�6X6ko�_�Y_���P��~�;U�A�x*��BaC�,��niܿ�6�2/�H�M [��9�3�w�^�:Ná�V*��ŝ˪�󷦕FmE��7���}� �F�����UF'Bց�����u���@����7@3�:rfs�"~���q>���ǰ�P�$X}���.r�A.��i��qkP��AH{�ɰu�ţ����M\���o�;�� �[7RR�sr���Wj�FM�4X&��J�HI���t	�ׇ~�)�%@��B@��(��ߡ�O?�u64H�G�r-T~�vE��E��nc;ﴫ
���p�i�{��ahO�I[�H�k�WR�ab�>�;;���ɿ��.6}�v�h�y�v�i'������!U�g" 6�SO=�� ~O?O��)ڇ��?�����W�£X@d������
4I( 4:O|�V����<q��`ߏ��=+�s3�6���%�� ��ﰒ�S�$��|B �D�p/�s� 7���zA0�9��>` �1ψf	�@ @'r,4��s��\�Ǳ�[օ ]��m�X�xP2�څʀ�E&?	��9�j�2��ƥ��$�zR8w����	�>��B�}���������哀���� M���>hN!!,K�qf?3�8��8�o�� 3?*���>��{��z<(ԛ��z�ɧ���g;�8��|̳��|���}�1i�Sy��|�������Γpk�ʷ�C�'K18�B�謥� Tڴ�^g������Kd{xm�G����9�=�����#:�J�|1� <�lhLB6�/���������9�n��?�(ʹ*�K�s42�wM�R��ߥS��U`���%��a�3�̭Z�1�k����3� ���h�h�QQ�P�3����7�FP��$�?��5���M&J���V3��Ij��+!�)���q\g��c�<)����M��Ki��s�GO�I9�c9��4�kS�f��u��(��o��M4��$%�k��օ�O~��v�]w�~���+Y�{V����gM�A	P>�"�v�q{;��cm���9�-%�2tt��=��S^.~ͺ���*�vL	��dF7��gΚq���~S�q��s�t~�'��htͿ���R��b�r�!�'�=��͂$n�P�+�8������C(�����a���� �Kj7�=4�K.�������%{lb*�[aS�V�{�D�H&|�xw����"`�?��^�Xjr�h���������@փB|�+*��կU{L;q�k���N"����*�W�e���RX$|�'X<	�'�S��寪Y9��y�������0�k�W��^�`��0��2ou|-��F-�3�{l%�<f��|�U"�'^'�k2uk"~�v��; ��׾֕;4*��ЩJjd vS*>�
��P<4���|~�uw��|�$	��o�R[[(3aqo�Q�����C�XXmI|�����n�9fk�xQq��c�ɇ2@�3���dx>��N]s�5�9�}��j��7׊�!XDlLg@��������29�1�[m��ix��f�% d�|�S�rK�Yw�$?%�c��p��E}��qȋ�q�^��ω鎀�8�Ѓ!�������6�~|l
��>r�J��X��1��V��յ�@��f>��H�c�%��أ�:�kn!9�%P`В#�?���<QK�a��k�BeCoK�w�]F]\�}��KC�N���t������S�=����'���E�/�G�F��<jxѲs�׆j��˨�<��4�S �w欙WOH�������{.l���}#0LƆQ	A�	�b�VE|8Y�4�V$��=I��?�s/��v�2��Фah��Ѧ�
8��B;}���~����}�V�lGi����Р�0Nd�G[4��� x6At��8�3��˓���Q��J�s���$F��s��Xq�����߯��$�����f���b�������D��3vs.kF��a�0��^z|N�L�� �5Ф���y,(�^@>^�̔�4p�Ԭ�@Ŗ����)f��P�m���9�=��W���$5�j͉�1V@��/��-��ZK�
�|L��~�(���u�?�/��{Ml���%ߓSc�	>��l��R5�lD�Ol���i�M�?N36p~,���ȩ��� G�L{q����Eb
a���"�t4&(�[��-�������8xd�5Z�5z	E���B>c#�̜�<p�18�2!��)�'�G��<v��3L~��㇫e>��蚪���̋gB� (P�����<�� ��j��<E����B�9�lt*jJI�y��x&	]Yc���"�D=%eFV!�s�@"`�.���l�40��1|ox��Эk<�Ϲr�K�I�3ỏ,(~���o�A c��FBIyc��U�c|f��	���,�$�����w�ynRKsd���]M��9*-K� O�F��C{h�j�)Z��Y����{�:�+j���F}��^2�"P�[���E��O�<�|U"�K��><�B$�k��]V  �s���K��gNI(㧴a���9����"�T:��	8@�8��?I�=q�a"���z�B�)K��~�[���Nn��-�z%×h~P���Pn4�MDՉ�A`IS��r�+p��\�����O���Xh.CUP�:��Q*&�w5=���i7����+ƞ��	sc����x���6���k��fb�'0�"U��T��C�Ģ�糁y����)h]C�����1l�Z�i"h��67��Xm�,
QͿV#q��Y]�.�q/�+ A�:cD������.���g^T�pt�o6�cO/�7O�J�:J�����	o���d����Љ����Wq�����6�����B��f��y.��uyv :�s�.��_~i�Ϻ�'M�x�y��K�9�Mx�����j���P~g��x.��b�C�I�"��zI�F*ž��y����8]��>ße��Ev�-��s��4��p�&���ԯ����#+T4m}C�F����'�7���Fm��i�	���8�e����E68P�����j�-Pa�0@4%�H��8�
w��y�������/oX�Ζ�����$����d��Ҥ���pH����qrj��\[N]�<7��	ϕ0�W�) �f̵ J��$.Yrr��LkO݋��YJ�R�g	<���@�����}xO<;�������d�] �:Áy�A����ȓ�@�B�q.�o�w�8i�|/�Cd2š�Z�::s�G��"p��-�_*�C���}�(����3O�z\���W�%���4N
`.D5SNF 
5�^�~�
�1���wD��(�A����h�A&���K�!h�ld5��si�V��1��,l4=ř�@���V્΢��rP�D�/�7�m��N�F��ܺ�k��ъ����_��X����c��>�y�<�( �U�8D��&����̭曹��&�Gh�P9
��oU�Dx ᙹ'�����e��s:R*��15%+�u���R3���|b��L3�C��,7�A�<����^�7[�zUT	7D�[ �Q#Ifq�ŦM�nm�>��W��/��^*ݩ<��o��/�#���=}&z/����b!!�b�<c,0�	�f�~Bk�c��7�z]C)[� �5��Y��@�4|i��6��r�rY ǰ��81�R{��K� &��.�f�� ���t�fZ�,�!@	s>�	����|��4n�A�.m�EEc^x�>
I߇����?~�[J����o t�K������;2����X����,XB�S�>�g�����EY(�RJ �
�s�hA�N��O����`=���f���F�'` I�c>�`��#T�>=!�*�)8��Җ��l֬�m�?�Ψ����CJ0�D���t�8�'"�_B_�@���W�ޯ��	��[���sD���#��3g͸rb�z6)�6q��e-�ZN�@ҦT����X�\O{�簨��T�M���a6�;��@1�2'��M!}'͟��YX�i���኱�"EkH��Oir���U$��;]W�%�CTB�T�ȱ�N\�8%����Xm"}���T=�EK��E;4N\Ka|�uUs߿��Dhh��H�_Y�������xZ���3�|�s���y�=.��g ;B*	���yF5o��ǪDH�"+ �
���!�<3>�I���M��g��)�Ce�1��\b��GF,%O��޽��U��Ο}Ʋ�S4��a�n�������-_��È��?/�j*��p��֐�{	I	,�X�|m$ٕC���=*�r<�+�=���`�(	o��Em������v�Z@����`�y�v�I!:�J�k�V[Oo�ggs�����]� ����=Ĝ�&[�D�B� �-.���Х�iaJi��ڸ�X4A��:_Z����o�K�u=	�%=���_�a�kSmI�g\��3��c!!��g��������7��q����8t���ԙw��́"� w���#׵��3]	@�g�p��x�N��ܗ1�;�y\�.^�[�B3�;x>@��Pj���0� @�X��VD���
5��9�Ѓ�"o���5��D	8�6B�p������h���RY���5��/<��e8l�����<)r�'��%�N��qh��E�tl.�q���d<j�Ak��N���'�n,0�5�1K:�O��ϔ)!�pg`��AK;�������B�z�lhpО�;��1[�l�ku
��s&��?J��̣.���"b����\��h���c ��౳Y�4���-�A֎61 %kF1�S��H ļ��@�1�Z	��'�%�_�Z�w(������[C7�p|r�z��H 0l~QE\S@��XY<��=�9�q��:1�$�Psm>WY*�z    IDATG���{�
�^d������r�yzO�{��Eiq�rR���֐��|�;�i�|�V.�?��*[��n|����Y�~�lR�?~��n������~'���e݋��w�:s.g�[#IiW����X�d�c�M�����[���γ��	߇	��������������s;����_"G�4L-D��������4�a8��C��K�l)i�yY��i{q���/~�i��f�$�� 	��l^6*��hhp�t���'�$j��C�F��~i%��ka��9Oe$TZZT�֭�$�44rT�P��Q�]�s��X�m*�I�%�7��g���6�(�ሿ���2�f���ҸD�	����%�%,W�Y�þ��h ��<���`���@�7�Q�9�&s�0S�/�Pv|^�!���Hg:��k�tnSN;��3N���/a��J��(Mc�5nex�V!�Z���:��J�OL���)�-L�@N��E�*a�g�k�0�<� ��|��x�=QVX����9���;����K�ٝ��/W )c�أT��n���s;o�i��15&�EO���k�w���� �k�Hb^hlm�9+P�m���Z�}{��&d�����}�Cd��qt������I���
`�|�1�C(� uxӄ�Ȣ��8Wi��% `�'ϮD��;A�NDY+�4cA��&Y�L�"ekSIK��-�������L*8�Ѩ�bQ�A�4�ҋ���\BUVS���$ 4��?:���I�g�5M	%���<�E�i���!�_V�)O|���xM�9�N�_����GZqpȆ��e	�N}�j��p-�c�whiks�v�i~.�>p� g@��s�~���}$|e��j|�\%<�ȘB����y������,��T�M,L��BHպ��ح��ns�>�nO�k٪�7��:�t~�;�����ς����3N;�.����Q�`C�}�����?u3��6}�ǃ��Cl���I�C&�x	�㚢C(`�$#͗ʞPI4{x��_�E�ЬT$�x�����$-� �+��&���*G����Ǳ,T�?r�/�C�ݠ�dxg /��4�wBy):������f���{�]J���%i��1"��R
�$�%4e��/1� P�ঐI�ב��8�l�(M_օ�Be1�>��/IIF�3��
VF-���-?�,>�S����:V	d�{�Æ�/�u��3���.��?�iT��tu��=�(e��^Ƶ�oPl1奧YcJ�"�������z�2��;���D��ڿ�Jnd�xF��`~(��7_dS&wXGG��9���#�sK���
;�#m��l��P��>���ZWW�_��i2����3���|�Ս��X�l�]w�ٮ��Z�2u���d����<�+[�n��n���f���vԱ�ٌ�;��S���;�9~�T$��� �f�V �y������W�8�BZ��IҒ�*s\tE@�pB5�fA�*U�J2c��3�8�s��� @������Y���L[�c��Q�%pR2�l~� 'c��R�8�oi�G /�� ����ǪSct	'#�~��$��;q�S�=��+��se��)*��ay����D�`n%�@�DH3�Ж�Tm Y�(i��ro��i0���ޑ�QLX�N�̏��1�'��e%�]Y7D����;�_���w���e�"o�@�&��Y��).^�eoi�GQl��0��'ƛ�ZI�i)����m?s^=�Y��~���z����8�;�'�:�̳�^�T���h7��U_͒$'t�������{��6��-�gLJ����O�޽��=��\[�����`��q�-����U�l�̽���Z5	 �� ��(��g_�j�0�p�X �����E"ڠ�O(��Y��}Y4lp@P�,N4o>�"�cC
X ��h+���V	�(-�c�X��!�@)^�s���@ı,r��x>�%@����#��Cyj���A��{S�Ǽ6�(t# L?��H(�
!� 楱`��L���C��Q�r�ATcƘ2�*Ɔ�e�'�n�B���I�$�D�����q��K�zi�+	�f���X!��K�j���lHn+�J~����4��������ʅmʂc~�����Ip��!�G`̭, �7�Ǿ�={�����Z�E_�'�>�}A&Mj�� ���i��������v�gy�����q���zH�VͿ�̞3�������?�&ɤ�ɮ�Ϙ���������]w�e��l��EV(�ͧh�ۇU�cU[�v��=/��4��6��j�ڋ8r�E�_�$���~^r>k���=�� �?]����\� �hҮ�[� ���D�R!�A�@6 �6�|/��84��4{�� dXPb
��9;ƞ"� ^X�S[�����pGp�Mw�N^7��s�cm>�͙c�X ��+~zG�LƵDQ-�=��8�ZB�p��5�ye�r�1��!�$A]��;z�.���X��C�^� -
e��7�x��h��2#5b�t�Kb��\�ԓײ����y]�J�p]E�q���z��}]?��5�=뚦8L���/� ��Ų+�m����@����xɋVA�kZ�RM��E+��l��e���o����ו�{�C�6#�3ʺ�`���ȴ���OHh�]��?�{�*%�f*������t�1V.��E���\�i[���V�\g�b�.[gx�;rj������,�йP�3�I�������<�T�qj����7�KCf1�)�bt R� �~�3A4n�h@y@����;�	���U5ZK+���}i��>���3��{��#\�c�5[���ϳk�а��F�g\����b��������v���:4�l�XQ� �;Vt����M��jn��-?Ϡ"p��^ ��h�oE���s�K��N�g�o�%̽�L��M{�S+o �y_��~1t�
�y�.`d�# ���
�'%��[ ���Qx��|w,����σ:XÊ��3����}���`�ux��3ԟ�_��m�ݶ�i�;�g���"����\���y��*�zM���>��K.u*k��.o�l��Zص&����	M�t���\w>��F�?���g�W�{nx7K�.�g?���䓏�je�V�Zl�{�C͕T��u�ڲ�]68d�t���+��pL�����ᣄ���S� `Cv�a.���tg�Lhmti��4mD	iʘ� ��� 0c� ���f( �}�'��Nc��A��u�h��f)��}�B��0���1B0�q��b�Z�}b�I��-� ���(ʉ����k�D�W@�� ��;B� ߈�r�s)�|��=� c0�Z<'Y���.��� o���%�'�P�=��C���R�����o&b������{���w��?��2����p4�{��c�QV���>�яگ~����e�w� hտ�˿�� ��1��S��<�����;�C��Y�O�y����\���6�_�g�Y`����.��N�����������������hNa�U�o��Wv�y7{�{n�L�b^|�~�����c�R�׺V/����\��n]�-_F��6{a�:;�����x�ob6%�ڕYy�%�x/� �x�|h����O~�V��E�H!~ ���E�p=��j�9*��DE�<p��@y��@Bh�@(��P:�g@sAh���Z�|T����#@u�<��=��=TE��Z���O�TV�h8����|g��;D��S���`��F�W�NƇ�� Tm3QE�0WC>��������o�9繘/���،3�@x0�Xq�~�G�Y�ԍ����q/jN�Ys��P��=h��p4��p�ui��ǅ�t̖Y7�s��Ϙ����v�[|%���͚&G��o�����H��8����+���ڡ�c3fN�^���2�A2W�����-�r�Ŗ/�[�P��|쟼�iw�:���sYT�4��̪��c��/t���4�Jp2�������h��>km�ط�u�w�V.���e,�_k�����Z�Ζ.]iUk��K{m���eeX��,�h���7|SJ�C{@+���˜&��i�h�z���XXrk�� /�f� ^�L�C!�h���"U��o	�)�����������[|��Y[��u#�5��ⵡ"���~���M,���c��������\Cxa�J���-��y@H�G9n���x��k��V��Q���S�;j�uy�)kQ�g�y�x��!�'�h8͕H)&��-���	��	������ܷQ��%�K�"?��k���~�aW�k��C�A����(���J�͟�_��9{����C���۴�s���P��R��E֞|b�����_���d{׻�<��*��>�9[�d��q	>���c���ZҤI��w]o;n����`?���e��T���k=�~��,؋/,��]�mmw��?�-^	&$��~%K}�c��s�=�Ԣ��E�H��;��/[��ə�8�F_�`��I���|��L ���EI�i��t9ͅk�q	�Pf�d���Ikk-bHQ@�6����; �u��I�S<~[Z��{���=�??�S�9+UVL|��P����!h%��c(���z�}���a1��b���Z�2����\>S�#Ń��`�<��(0h���j�!�>t���H'	������׃�蟗r�M���;͹|=��1�>ڵ|.�h$���ކ��j I¥�3��V*�����ȦOk3��k�J�z�j �,�j�y�X_�Vuu��g̶SO=��i
eOo�֓���������[�\?^�tG~)C��?�Y�/�]�ٙg�n��>�z{�Zo�:[�f��^�Ԋ��X�
�P�����ޛ��]����Yg&$$B"�B�w"�Z��IP����ź�o�׶�����V\��KMX���(UPA@�%����6g2�Y��{?��̓Üs&���f�����[�����7R��n��$���]^���Z��c�5�h��[5�Ź�lX�9G�K(��}�r6i�*�`S�v�J<��^��xnv�h�C��܏�b�'�h��{	E#I��<�T��V��'����u	%�8�ǻ�X�����L� 
�8������	�J��w	͋�8H���w��%�]�KBw北�:�����d%j�c'&�AQ;ʚ�w�}4ǔ�@��Dsƻy"�~Z��0���N���(��yz���������/E-V�� ���Z��S�#ʕ��E֘�%]P	,ٺ�)۸i��ض�JղM��[-�����lp�j+�Zk[���eo}�͞}�U��~�;����l�#s�h�,��_���
��w4�} 6p�Cgۻ��v;䐩V���y���l��uT7������������C��N{�2����>�X�;�0��+�ʿ�Z��7����/���f��6��s�Øwf#+kT$�H��"�A��7����'ϣ�mi�Z�z�84��^�v���6)!$s_����eE+�~��������VA���&ca0�H��#�� ��3h���w���u�ݩԂ�c�'��X�`.8^�ɵu��+s�υ�������<��k=h����]�G�:��?~�;��W ��E3����������G��k\Q�����̄�rX6@�Y�YG�j+W-��+�yC�O2)UISV���u�y��c����`9���o�b�Q���V#�Ϝ>��ŋ_�8G��5�|��Px[3��dj1�ɋ^h/y�mBg���)[�z���w���k���-�-��ڬٳ�����{�M�p���¡B�P�MY}6�e����͆)Φ*��/�C�A�C+��6��ٷN�H�i%[`  ��x�7�V��.��K��I˽����J�����o��d���w���v�W�X�I8�z
���9�o��OE�$�~�Lڲ� e������" �oqss@�#�j�K�wZZ�Z?z�V��-�+Y\�x�Ю��s��Oi���9�_,9^����Z��U�,z�}4�d$���9w�(Ǘʡ�&3��L:G]����Ю&�p+�?������}Bg��c�s#��[��=��mdN����E]d^�r�V�^����,�e˖z1��g�9�y����̎:�y�7���w����Р�}=�}���;7_w�������P���f�/P�=U~�$���KmE���P�3��߱���cƌ�>�^�;���l����YX�~��}CSo?�'�E����rE��B=y>ORK���QYh�W���?���;�/?@��wh�X�y�X��CDE�rs��CWI��i��(��	�h�����|_�?�'n�g��Ϙ��V�Vi쌯Jr<mc%����s��BSS�Ɖ{ro���+��9
�9��^s�8�.�*	X渝e"�wAc幜���I�B�B*��y��Z	�X IK�����Z�\��|βD�O,������pP�J-��0�����)۷\Jh�&�ߘD��.<�T��h<��ݗ_� ؃zn�(� �v�*�%�O�l��vt۔��G`��#��b`����Z5�wt�����?�����B���'��?0�����.���)��w�PŇ�r����7�ѝb+4�����+&tǎmo��lHi�L:M+�� 
 ��[��V�U�`3�~������4�j���b�1�<<?��;�#ԏ���R���� Y���Ȋ xV��h�h� ���(�#\ �����w��g�TbB��8+�������e#K�f���bR�f=��k��}��)u\�1㠕ƈ�!��3��zH*zǆg-	LCƖ�b.9��C(sՐ��J��J� Z�"Ɓ
�D;�7��:4s��o~SO|��P���t�Ӻb�.������{�΂mZ��K��ё��M�b|�?�Z(��1ɦΘi���\���~���m��-�t�I�3����+h��+%G!��Zan�3{�t��"����c��;|/֟<�Q>x���e��X6�	�lGֺ:����R(��u&o�����?��;�Q<;:r������>c��nY��+��ߦ�c�[� kq�c�R����?����d�׿*&�����ʖ,y�^�%v��G|�]w��ݐؼ��ԅ��
��G�v�-A&�q��N���zQ�@�I ��ffa�0
��w�$#�k��.@Ģ&I�Qug ! _�HBR�H��
�8��1�t��3�q��V4Ҿ�}ėJ����:V�q�Xm���i�����T�&����g�4�'Y��	�)T�XT�[IZd�2~܏yc���/��a^G�S�Z;�Gt� n�e/{Y�i$��G�+k��^��C����%!�(%��sϱri��{�~�*���\&� �
��ZMp=��'b��Cմ�>�X�5k���6l�b_��{l�A覰,����#�u�%M���.�>s'kPY��Ε��P�s���<���ʎ:�9^I�=�N�c)�LV���ݕ�L6������ZP?��߮�;#m�IS�~�-�|���>@cp���*Ւ�\+S|q���I���|�	�I� 2|���x�� ��-FE ({Pe��w���� x��&͓{ΊL@!	Iڦ�F5o��`I ڪ������Pb�Ҍ��І%(��c�S<����Yisc��|��u��[���-򪬲H�)�ڌ��=O5c�Y+l|��f�'ƛ����an��5�B�C �@�ɪD�o���܊���=@���*�����P������������[b�u��V�Zi�6oXo}=֑!>�b�r�i4M;r����J[-3ѦϚm��j�j�
�}��k��ǟx�)��4���E	�� ֘񮪃$�]>1/���7�@F@��ɜ����#�������p-p�`��g�Ppq�[\�#O��m�f�*W��w�C�W(��UK���������B���>���F��
�;�x�5��    IDAT�B�g5YV_�R�/���2�/�i(����O�����^;Nk @$������rN㚊��Bi��(0�f/�Ţ�z"��De�*_E�x+��H�q�𾀓|	��POT�~W�6ׁ���2�5`�;C���{_���~�O�u%�>��@	2_rFs,Z�֔@a$��Ɗ��'|�o*�J��7��]&�c����r�s����]-�s��'�Q�xY	����?���=�[�@�M�r���w����趘���Q� �TyЬ<d�V���7[�Be��[��'/��CCUO�*��Us��9G۔��:�wz�_�p�=�d���!l2��.��b�Xrq`�LD�%�}�}�K_r˝r�u�]�E�"u�1��͘8U4y���o���PV^�*�?)��P�A�w�'���#��6�g���)�����=>��t�~ܙ��ģ+ X,�P��j�] ��OX��~��C��Omj 0a�Ӳ��f&���}��"o��3�i�5�U��X%�(�H}b�q�Qy5�V	e���`��,P����Uw82.� ϳbEȼ�;@�s�O}h?5$G� �|��/�k�\�Uc)*l_9|���i�K��&驿��#��
��8w4:�� p��\��^�U~�VI`Mh#�S���3�|�u&ڌ�#a�Ԏ�Q�'ϫPN �P2@|�ִ4����J�h�D��+���s���{,���Ƶ���c�ufҞ�J���~���8 תVM�l03��3�&M>���i�6��_���VZ'J]RZ=r�֚���|<ק?�i{��<�| ;�r.�k��}�<� d�3�Y
R�<d�X��4�D�|N�"~��}),�5�ã|�7B����Y	h���}*�g̼�L�j	��M��W/_$9,���31 VtO�P ���*�aP����������y�Q�i7oݭ�U��I!ڠ]��$L%TR �������� ����DkDp����y>��B&�@����;4Gq�,`��g��:��Q)��V�R܋��Se��K�_���g�]c��͏S#�q
%LT*�;|(�h�|���YT[�8�����P�*��5���fYc�J�MF�h�N\i���M��%��=�X��
�][%z�K�0N�Ԁm��rV�5�V��-����Ւ�,� ����TΪ�iv��ϵ��DK島e�v��k׻�c4�����?�'i1�j���O~�֬Zm���7����~ʂSߟ��1�Þ}}�k��D]ʊE�ↆBX1��I2����#���Jz�|�O�V�̘9��o���_k<�}����,*t.Q�'��	��K8�Ɨ�$c^�b�[ȥ�l�i��f��|i�, �8\����1�i���f�������s��sU�+�CX��N���1����E�v. �'@��@·
R�H��X�*7�3 ,q���� � (Y ��u�w���x
��DК��G ǽEY�V�C�Z�[\9U?U��Z(���������{	��h-1?qKF��|2��sJpKH�* �IDOi}J�ig9�{Qh��yN���i'�`��+C�~��c^�����ͤ�����A���?q�A���i�7m�k���=��S�'YJ�kY	�4Z͟{K@�;DΡ�S���N�(��0'�7��/��/�-Z�w�Y�A�Y򱐕BJ�N��)�(7R�5�T
ڧ���ߊ���-�I��a�g@��ed��ؑ�zh�f�6rp'�����l
�pπ�J5��]K�KE�p��.�f1�%\����z��,�&��k�+-��%
�N�)�x�[	1Q^zY>\[��! >��w�j�tہ��~��k��ߧ6.�)G�@V`�؈;����A|/ �z�
�JK���{�ΕI!�����R�RxX#G=S]�%]��.�x}����x.5�܃:Bg�q�k��r�i������W�N��.Tm�6�τ����߶�`_������K�ӹ �{��+�_�_
��]�� �1g�ׯH;|Z̟�nY�Z�4��A��9m���8vi���@5,�)Cs�j�[p�8O ��	bT �2����F@j�6��9)��'<���:�Mh	���L;�ԤM	|���:|/� ˃��9��:Ց��Ε�(^�Rڹ�M��Oi���j {����3~�����������v�Y����x��4F��"S~[e
�X��Kc+kP�1fXr
�%̹����@V�"��%4W$F����<�-��;�z� %��8�T�Ҁ��l��ֻs�u��CA=�\����;X��G?�&O9�JՊ;|���km��-MYD����h�I�/TJ{Y�1Zl5s��B�+|r��}:L�p�D��ĉ��aǡ�M`(��aއԑ��8���n�&�H�x�w��'�$uК[���~
��EݼM4yi�,8w6���ht6�6��G��1�h�I𝀸t]I,��2��'�]i�a�,:������������g�<���qכ���5��[�RG��(�4 |���d��=�y���%KB�p�rbK�yD`-p ŵ]�I��@?^��;vr{�H��²���Gkݶy�-�ԚC����gX�<d��۰v����p���X�])��C=�ռ~��6��Éذ-�wؿ��ڒ'���	�] ğ�̓�	u�g��-8hC�����+�H{/�S���Byaܓ(�B:���q*������<��7[��}�å��,�$��'��A�%����Z$o0�[�n�|E���<S�x,xb ��'��Sa�X[�5���y��Z��b�ǀ��γ
D���Lև�_����k�1xb�ƛA�I ��0�y&(�_�>�<�1��V�A�q���X�J+�/f5�r
�u� S�R $���� ֕����K1�wAP�+���V������4�����M|�YgZqh����n�`�};]3�=��}�zy�9N��6���6}�LO��oL:\�f�lϱd�j���)�Z�{SV����֘�Ա%1]Sub`!���+K�-�,�$A��l�q�g�U9a�8�����3�N9�6s��I-Z�9ߛ$X���]i��9�L��� TG(:=�|/�1��c��5�H��4�F��X�-Pӂ�~Ah��&-�V`�0��5��Jck|T\_QJ������#M<�}bMZ=~e�s�6z��^��K�Z!v;�hT$�֐Rc��<�^��敟��@9��)jH�C|s���ח/G�+%{:��x���8�=�7e��;�s�\����?�{$��p~���/�L;�&M����t&�͈z�	�{y�x]�oQd�?�B!�!<�)T�$V�4�u�<���%�v2I�"ǖ� �#k���Z�|vu�����g�w���74����h�6�_s3j��OU��i�!Ty��uV��qG��	-�����v�g?,��Q �w�7���s��cmN�/KC�F ��,J 8�2����%bm/�$F2y�1�Ij��D;�D���p��]}-#Y-<���B����I���S��4�=�UP�B0�!k[m	�T�:귣���+��w ��� �t,e/���;�Xo�7$r��wYd�����w�q�\�g�6�Xu�O�g��?����Li7V#}����֑�oϚ/-�U=т��"�R����rŲ��l��e;�Dh��YB��aa7)B̑�]މ1�
e�Uԑs�N�_�ּ�0��lG�[n$l�P��;r!����CuR���X.��a��V~��X�o]�!h�>95����7&o޼s��Shf�8�7*�*��v����,&Q�>ͦ�?����c���wo�Q/�&-J=�x��ħs��?QA�P�֢��(��ck MK�]G�[�}�����^���zҤ�;O�2�}M���K�$�s��]*$��*5�ԛ���n��;���@����_Q�� B���o�ݣ|h������������A�A��AV)돜2K�l~��_y�!�{��_�E�PD��d%��q�����T����	��Z�W��Z�����%�fRV���9��V�f%�}���Ý�MI�0GP�t�J���aI瘮��m��J��+E,Vd�/�r(Um�DҜs�Qv�s����&L���*p�|�
[�jm��9���wtUUh�ߦ�[:������zgʪ��o���E6��s|B���r专�R�y�Q������M�;�(F�W6�w�i_|��� n��f/�,���B���&Y
�}L�H;�ƌ���v�V��"���.��G��o�L�*$H%��]�P7)������J���4�%#� Bat�g"ڧ�;P�3�$��'���_���l"Q���44�v ��ݾ��o{���.��rX�4���_^_G�]w���34a\��^�'����?�����ČG����g����̥qݱ��B���̕j=i����[BC~�u͘q�W��;�8�y�t�|����{����k��ҥ���w��a����;���g��i�r�j�Z�>c�{oY����u����-4������P�L>lj�ܜԩ�_-��n�L�^��/8ߦL�T�����n%�~�͆d-Kel��^��^���1@S�����\k#&�l?��O�/x�oR����ы�Q�)iӇv�&;�H&c�s������Lp��( P.1>�`�w��OL�	���X3���{�񓟺P�v)�E�.�&1�M{!5���a*���E�A} (����J���??h�q�>�nD%��CH�������3n��F�S�r l`U��J(X	���Z�b$���7�#X�?J�����|��|�7����b]q��y���BG�&�\l5ǁ���������e>��H�ճ�/^�:[��'ͣ�"X�V,��Cfx��'�Xj�/�D�\G�	�'	�#����V��Y|�^B6oC��v޼��k_{�M��e�tնm�l+V,�%�?b��l�,����c'�x�}�s���ȍ�SA������/4 �۩�����}����Q��+��K�,�ו���
HY,&z�"@�8P'�W�d%����v�F�l^�W� �>��j�/0�3���[ns�U��w,�Z@���)��wн���)�����[֯��3|G#X��<�ǀ?7E�����}>��	�#�i�A) ���0(�} o�h�����6�( (%� ��J,�������}3YN#�5�w���Oh�.���_�}�dK9����U=|QT�O�-t>���4����VX/eֻ�y��m[69��!3���͵l.o��Xg�{j�*/'�z��?�h���j.��_��?
=�����3h,@*xN��f����J�1}�UJ}�}�f{����򧞰����iV�x��!���?��<{� 6����
C��_�����|�+�G#$=�]W\�<-ş����E��i�b�̵`�7�E�l�V�C�����_��o%)�`���i��Q�	�"�~l�[n���q�u�G���FZjD�#m�����?vFslɆX����G��\�5�wu.c�Ӵ@F ��W�(� ������d^o��G�G�W�.���_K�g���w�!����*Ҁ?��I�0N����D���O+��{���"�u��g�������÷���>�N�G9 ��Cq���g��H^c=#�����g}#�K�?�7�\�Ry�{�a��{�9�Dp��6�?ds�e�}�͞��x�G1��n��P
����9���M�r�8��T_�k���۲��-y�!{��-��zQ|fY�e�lgϠ���q'�j��z8ߗ��e�p��{�s����I�OU@z���	ƥ�H״-�F����"t ��5�q 	��f�NL-5�rů��*���B�i� ɢ�;��{�}�����K.�gD�yN��IS�ZV�,�}�9`�{�+���gV�Z�w~��c���9����p��O'1�D��{����h����5�s��� a��������s�T��5��;�cF��so9|��C���D(?�e8yk�>��p)#�1�ozӛ\������[xXq`��z%k���\���sө�elȖ.{̖=������i塢w��첁����؉'�f��y�z�,�,��f_3���4�����k�N�6Bg>o���]��c��T�h����6uY{�l��^��R�����l��-60h�ik�����y�?&�g?��kq��1� L�/~��&4ϸ�7���dS+$NL� ��9�|�T����88���� ��^롃q$�H�B�����1@?|4e�#�U�(���h	!m��8��m���?��'��GGçp��>����zVǩ���G5�YNz�/s����8��P GB�n lE}iޕ��#Q5�&c�H2��(tX�c��q�OE�R#�۽d��u�gl'5��u��CNH ~rB-L�o��?����������h*X�>�j��p�c@����f������8�k+�z��%��ښU+Bu�rj>7�֮�d�}CV���-o}�<m�<���d?���u!+ 큫����U\�3�����:<�䆯~���O�\�+��_dCfҝ6�_�IJن�v��'{�*@ʅ	_�0A6����*@,�0A�C[ToV6&�P�D���׼�����PWg�h��.\���V[�xbU��u�<1M�E��_�!��K������V���p�bR�$9���x'�h�h���sEg���
e�. �xʿ��}���.��r�_EH�Sf�d�i����u���h����^q�hȝ�P4}r}��a�vCͲu� ��m�\��5s��w|0�l�ga�`�C��/ Jڗ��%�A�p~����ۻ�CgL�I�'چuk�FQ�u��r�f+W��J5c��vۙg�k�{����k�-]��n���m�������T�s��q��?�c��Q�~۸a����;l޼S,�.���Ox�_b�k����m��V�u����l�	��#���&���|����	11�x �-�_����:�JQ�Y� �Z���(K0Q4\0@����<M�@��qBSi`������Y�ȝ�q���]}/��������D�ƅ�u��1�{�IJ������<��T�����d�ǚ�(A���c?.���j�����Bz1�-KNV�֔�Y���؃�����E����$vՂ �4�g�c���aܘ+�p� ��ĺO|���u��,p��"�/���l�#��_��N9�h�1�[�أ60��� |��@��u�u{�uvM�_�q�wM�����ƛlŊUu�����p��3�������o���>Գ�毥v�s�t �Z�V�z�~������n�T�֭_i�}=I�D��-ڪ�i�m�/�`'�r���M6�wh�C>�4z�^ >��?�&'�mTB�LR0L��E�z���d����q8����Z��Z����+�tx>�Ef2���P�lFۇ�G�W)�v`?ҳ ��>�J5ǆ��y���P|�`��)���� 4�틠m)�E�)	7Y��W��9�k�B��6�Iܞ����z�XP�^��i�~��n��KV��^�*[�x��k�c_@���o�i�J��;o���8�>x��Z�<�zz�0 e�=���Ga�v�����~β�N����o�b�r�	Qy}Y����?_ڬCg�'?�1+�,m%��o�h���ݶy�:��� S-c=�A[�j���Y۸��iej��ѫ�O�����L� q��lp���7;��������ϙ��)�ub�w��A|���3�n�k9RZb+��H�w,_zH1�#l�/>#�p|�a��d
)������s�|�|4�ǳ���c�Ɖ^��k�ɇ}�u@���k�|��������5����N��`lEi�]�u�N��'�G��6y�Tۺ�ە�U+V���	l��������w����1k������i�{���}�v�
+��i�N�mg^��v��m��m��ګ_�jN4    IDAT�z��=����N����F��w^�.����)ޜ�"
ɹ���8��e[���L��4g�� J:�xB�	x���?BVj>��Ku�#�>�x�!�G�/*N91����N���������=�C�8�g�b�;��{�#f�Y�kV�p �8���oK�\a����M������ezh���k��j�=����G��V��τN;h��v��U�Cֳc�mߺ��wo�Ri����%ˤ��/tÆͶb�FK�&�;�����~��1�h�$[a
����O,�,e������׻U��H��J�#�x\��}�
b���8rM� I��~��	��磈'ێ�!
��V|SK��n�������ڱ�{L����C�N��X���O�Mq�*CQX(~�;{�R����l˦��ݽ������}#,c]�{G�=��%ֳ��.���6k�l�T�v�O~j?��-����)��%cx�:|���QU�t-ms�εw�������[��=��a+�l�L�f���@����c�©6�9�8@������$ƟJ���DD�"5֮_��f��0��deӡ��H����?�m=~�31�p��V�+ �Xxj�  T(Q�s׭�����G�3!���c�1�X��V�]��ʏ}���O}ʁ���\'J��N�qQ���8�@	�_�q�h�V-�e˞t-ʇ��\�_���`�N:�t�{�)��uX���]��=� \j% �8�VU=�VO6D�,���)S�S����V��k�����k˗=�WS�5a��z�iv�9���鳼�@Ov%�J���D�/Z	�-���� ��N�V����J-s���7�5d�9�q��X�l�+�EV �1�OTq(t��1M�HłA����9���,h��<�x �XޓwW4�"|ؓ���<��x�c#G0>u{� }@��˟gR4?��=^t��T��Ѐ=��v����+�[�J^HH�<a��v�ة���5���<��gw�ү����s`W�lQ�_]��JE��5�bG�������Yg�n�Ҡ�je*؎�[��[��'|�t�T�e;�X���y�ų�0�lU�'��/�ω'���]D�ȩ�yh0,.�>o�1���h�fe�h���]���3kmK����=���TB��b�e��T�#�u���Z!����eK��iU��ݳ����Z�]�I8�	�&��g�P��������,E��	=����ՙ��ނu��ڵ���c��>X3gf�"��t�._f����~ *��Ƚ�g��o��Uw���(�J}��|_����/8ߛ,PB�hRJ�ԩVC��޾�����=U�/����W_�@�ǂ���+}�X����_yHQ
,���ĉ.��9�� �������0�S�-�]�z�gvS���P�b�W�H��0�U-�N۱�k�$B�<���z��р|�cT�	P�ު�p����+��Q��`�<��Hй��P�^������_w�[t,+��~����o�B��G}ܾ���Y���^5�\�~?�����
݅KGN�ҿ1��o�P+�F�&L�I}��W;mCyg>��eaB�l޼ս�j������1hj�v���A$;�ݮ����¦�|���f�����u��E/��pdƺ)Z� r�YH�m���RI�K~��a3C�ocl��Iy�V4��s�єw`̈��Z�ot�kG��hL�	5T�ߎ���l�ќo*9��7~/@�3�UnC�[��O�c��*˺1���F�&�4@�������Y:������<P"�s��@V*�uMԏ*�����^U�U����Ο��:"��G��t\��ڱ`b/S��w��l ��_Ia��vK�N^ټ���!�ε��&{73U�,�"���3"���==Ng��O�������3�?�{U�er�w ��9�|SQv�֊ ��kA�����z�^p�c��G�'�hB=�N \i��$���MD��JU�z�J�1h?�z���ΧV�C���0S%yQ�ᐩ�F��5K�P��| ��H���I-s6�j��o�AJ9��y�X9�v���PVl�Vr�	���v�h�}�{�kK�� 9�5*�9(*I���<�ϕ �2ʄf?�0�}�o��"⪣�KZ�?� ��GQ�\����C�k:�=y�s	�x���8Fu���
#�{���zdN��\=�����I'�uE��1.���}^��н3��gýR�`!��F�w;����߬\����!�������`;�Yw8�� R�l*d䖂êqQ�����'���� e`)���O~�K1P��k0���Ь�Z����uY������/��K<;��z���$�8r��w�'�2��1�uI��nu�������f;��X*!R��#�*!�ZD��9����ƒ{��۝��R�S_'I��:�\IJøގk�{��%PdQ�Y���M}�����E7V�˳���R*����7�(��8�X���r�����%y�w�q��ؒ�] ��v��|�a�8�9����&�KR���_ʹ`���Ă�n��(���;��2�j(՜��10��hh�����©q�aځ%1��W:�����& ,��iQG�k�$��(
M��.����n�4��q-� ����S�3Lnh�^L� %�<cA�CM��%%,Ne3rV	��B*Z�#-���H���i�����4��y󭷸�[%k%�)M��c���;���Jƀ��&�*�;�I<��6�~�r�&�����+n��F��I��=�w�y� �`Zq���)�����gkw�-��땠Z�$9�S���Ny �͟�J��/>88�'�h�=�H߫���Uq,悬b�Q��P'~R������:��4*�uKh'-i�T�d/�I���z�p��`�9t���c����[�a����:|��)�<�n�jA�G�
�t��b4�J�ĭ�r�w&NG/��D�o��w�Q�4p�	��4B)8~B�`�?=}��\RW��O���P�v��1�ƢVm�F�_�E
��@ʂ�7l,0�	��ӤƋ�Ն�����8|���t�Q?5~D[�n���$� -���/�_�\��o�y�V�֧�㿧�6�S\��)�d,��1��3>�C��D���1�ז����+�Hc0�wP䞔Q<�p#t>�񏏘������j�!���ZA$��t�M'�%����.��{/&��?��S4vj��9�ƨ~��0��̹j%r �p��TI���F팉Ŝ��o,s���v�]�a3�q��D#�����y�E���c�G�̹^��_���GE� mC�&	o��%���9|o��mN��;�GμUO�}|���ռ�, 61�<
�y�ERu�&}�1	�?Pn�~ 5�6�Nh !�^c���7���X0�bJ�k��%81VXI��sٝ���c��Z��<vXJ��6�ؖ���5��s-���}ޑ�Wt��>��{����M=���s	����#���[*%��L><Y�h�`����j�P�8(��c�lοE��k����HӚ��L#�j��PfA� �Cㅴεهs�h8��f���3�T�.�A6h�Ī��x�K_��_o��ݛ|���}ڙ�.���K(�H��_�����YG��ӈ7'�}�[�����Z�%�j����p��&��r��`����(��7�_�`ų���ʺֆ\H��Y��]Ig�� σ��:�hr�]�!a˽dep�7��u�[k�v�DϠL�՜�=���/���Z�7���/ņ[�ַ�o�(�MhY�g\v��۽����u|/�E ��Ou���]4
3)ij(q����^�B8y��� �]���B�'��F�g}�}�$�V��6(��������J9h"����kv.�E�*b3O� � Z���j*���U��lp	��h���z�����k�'�3s}@�{�N��h
�-	gv�Ӝ��J�½�������v��L�,��rSI��	-z�	��d�k�	,�m�=�>����
��y�K-�f��ˢE�p����ޚcͫ�|���3��:�_|�cu
E���<�p}���{�ܘ�z�K]KN/�����|
l5�;�m�Gćs��#k(���k� 5�w���5ͳ�}�� �@D�����}���,��U��4r����a�N�c�}��Ĺl	�f���]g�aV��%���ש� Z�j�qԹ,�봇4�X��$���ڔ�`k3K[��N	��G�^���":���7��ɤsP;�m�X̭>��X>ZԊr�i�+C�N��X�m�ϭ1ֳ�����Ƈ�cݐ�G�a�k���W�q>
oe^Y7$���_ �O�'��ց�ќ���F{���H�VS:᮫� �(d�1�K���G���{�ð��OJ�H�5d�"n߮��j�����5(�_ᥚ{Y$z.�����)+V�\:��[�:��0aP�p��q�R���bZi����Z�UfN���ŋ��5�I��z\��n8\(�Z�f3!<m?PA�
�d�<p1o�9d�2�����[2��P|���^��/ ���r���AlA��'`�l�*D��e��iNc`޳��c�T>��9d:k|��~��e����{�U�k:�~K�.��2������C���x:LUX��|��zA�v�/���g�9����E��e#ϥ������+�|߯��u�^X�-���W8�j!J��s�,)*��%�yX#t��3d�Ha�<�Zk�fَP�'��Tj�vM?X��/���l` 亠t��������fQ'�_�iH��gsA{��ET*A���	�삏/�dtuM���m�G�X��Y��5�"r$)����`���18�`k�O����o�������c˪����6
���v�?��ey0/ZC�B(���ؕ@˩����X��<�@D��Ɖ碥���|����xʊ�T8��=��كs�!��}+�_o-�.�ZPb�v�':_�[��["�CG������mw���g�a�C�JV�r�k�o�	C·"ɔ�r�c���OP:�Y�Dw��f�h,;�����eѢ�5��[��2�vH�pS*���<ҙH��#����zz��9��*k��2��7W�?G����i�P���c#$X���A9�c�kԲ��Z��z��3vJL_qSi����3n� V�\4�.n�'�I{$��a��r���D	<	t�ݓ�.}�.�5XG_�����+ϱ>{੓���[N�Ш=|����,���-T I�5�kX�D�L	����eB*�sR��E+A�č�[�#�	в���i5t�#�PX~ �O�?�"��-ʸ��Q
�|H|?�2�}*�O�4�'�@`��P�	��3�-4��#�wIݓ�u���{����I�ä��j����+��+_��L�4w8IY�h�ī��� E P�����P�Z�5H����t�Ӥ{���6w;�2Vڧ�{����힯����^f�45�9"����ii)7ɉx��7�R`�M��m6o�E�p} �� W��}^J�gQ�I4j�l�r���+�%A�t��(����^���{��QC�lҫ@'as׸��e�r{�q�^lq��aD�o��*�u��-<�,�o�%�޵�M�4��e�E�S�vJ���B�ּ�1��=���g̜����{�N^0<�=�Č�8a�k�z��k�>}�o.����pg"���r�
���d3�������S$'}�{�sm�c�S)��G13�Ac�yGF�D��]�����H�c�v�>���>#	����{����Ώ��;�M���T�t~�����Tkgo�"�ⵡȣ|�^AR�	?Q(�$�Y���a,c[n�3��ц+f�|�.�G�A��E����vy8���o�����w� ��h5�/zE��
��=Ĺ�o�g��	����,a���7��N�����3��a0��7�a}�\,��_����w�s�K֟�w����s`g�.���B��f�?���W��Ͽ���/�x|_�I�>�>��p#�-]�G}ԋ�!��X��$/!����!d�&�DkPן��4|�\���`m�FN�QP�u����p�÷Q���tO�c�v�����������d�b�1�lf=�z�{��^=�}��6����@��8�����J���k�j?Q���U��N�8-����9RO��:���^��:�SW(v�c�˾dL��ȇ�ͬX���	����n���d_��?��{�'��"�:�'|ods6y�A�y�6�ݸy�w�A��r��B#���m���5c�R��l޼y6�E^�&��o�f�
Ϛ���O:�4;��6g���2����#���7��<>���C���?����?���Ԑ4 ����E�&QO K��'5�ݱƺ�������C�'-p_ܿ�5�PX+hb�����x�����$�v�s4��2�&`"��}�)?��=V�����}/�Cs�s2Vʒvn��|
�#<�2�I(u��'��4y�Y?��T�z[�:�X�`1P�ΡW�%랂����~�m�C��W�%σ0�3��/���z��1����_�Z;���B����mt��rQ�4�����$�;\��Kig��8��3���[�F�$��Ϝ9�.y��v�)'Y�4h=;�ۃ������>!D��P�{�̙��9�γO<�r���o��v�Oux�I%J���ϸ��`��ٞHu�M7�BQ8� B`o�v��@��g�T�)vp>s���TH�Q����k��ۃ*2{�;�a'�=ޣ[{{lӆ5V跮���xJ�V���� �P7%���s���I���ȭ�
�쩕��uBI �	��s+�K|=���uS�����\P����~����Q�KKz(����g�A4��fO<�����_ن���EG�;����K_�J;�i�����3�����X�Ԟ|Mn5%�I�����=2gh�^���eo~����X�V����Gy �Х,mIĠÎ�ݶs�l�}�)�����d|�_p+�L�^ij�	��B@K 9�@	"\G�9ƪ9�������h����}������ڶ?%�N��J�^�nmw��|���:f|x^�8�qکf����{mӺ56�W0��)�x�\y��@瓊VLuج������X:�a�6o��v�=��ɤRR'��w�e�)���UI/|+�X�m�v����*��d[�s���N���?�K��m��'l��mǎm�ˇ���ض�������/p�'yq����5o ;�������G����f�?!��\Ʈ��]v�	�[�<d��M��a=�M�a#NU���P�6o�j�r�zz����y�{��o��>�
�BCIJ�FS�o���1�X�,�}�����4�i\��7C=�=�Cy��}"��Ya9��Z����[��P�m^�����[6U�t��QT~<�<4)��>ڮ��N�YGk��l�|�mܴվr�W폏>�+�N8ޅ�nr�%j���|�9�9���|��������+}��"��p��|�	�ʨ8�g}=�m���l˖��}�V+���O~�P�f����[�k��v���d�Ϛ�>GJ�C5������1��/�����U���#f٧?�I+ؤ�v����K_�+�ؚ�O�P1�Ϥ����o�W���!�������h�+W�ts�E�v�$oȞ�/QB����x!��(7I�g� P̡j(5���������)��=j
:P$k�}�{��u��V+Z�<`�6���m�,[��UܑN�r�g5�\��8�	�TƊ�)v�Q�ڄ�S,��t���7ڣ�?|4%v�ǘ��2�����g�����'?���wB�����>g���o��(~D"  �t�l���;��C��	9[�f�����~����mɓ+��s�-}r���%�_��I�z��-[���4�.92��`Ⴏw
ok�1�s�e������%۶}������i�t�֮{���{��e�����    IDAT�b�o�������csO8���	��/���o�' Iߑ��kV{$�LH�\�7�����G��J�ߛw���G@�}��Lo�P}6Γ�3��Ph�r;��ӬZ�L�d[֯���sT���x!!���:���9G[��If�[�q�]�MN��5�p��c3�PO%g�X[�k��N�o��o��ˇc��K5�T"�pN�İ[���_���v�I���i�l��%68je��R���\j��D�)XG���G>�e�=�._���ڨh$��f̜��3���7�oo��cY�l�a��UW}�2���Y��������ϰt�h+V>i��`����m���f�&K�'ز�[�O�+�����p�0���D�Ш�Xl��p-8@��r ���`e	s��8���z����N�V�K�z����1���Ͼ`ݣ��š�rѶ�_i;�n�|�h��̥�g=�W�x�������?�c�z�6a�:�_����ǖZ&��������/'� ]�^�erxN�{��]����T��}��\�(�|���=���7?��O?ΦM;Ȟ\����RC�\IY���Ǘ��J��ne�Q���������W��ei�z��
0�q�o���P��c���|�*������n��[���e��N��i�2����W�uk�8�j�v;�Գ|1�0�pH�R"���p�͋�uHn�{��_zM� ��Xi	q�X7����f�����5(�u�����1߯��S-�\�߲v���������<�����pNJ����MʩSژ�+�.;�����I9�a�6�{�I�>{����w)ɐDټ�U��K/y}=�����Ɗ'�+�6��|���n�Gp�Z��~����I'e3���_,FLeϜ��Wm����M�ի��f���_J���E��v�?s���,^����1hޅdls��9�=퓵��{���Gl�d��J���l��2��l����D��Sy��9`�W������ۼ�^��=1�E�VOU�X�Q���5k��0��;��]w��G�@ H�h�1~�����2�u����kd��x&�M[�0k^e���f���_.Yy��6�[e��[-�*:���s�?r��-D�0\2m�s��	��t6���W��	���h5�8zF���ڹ��m��]ٓƯ��4���>X���Ϗ|�#^�{�f{�ޟ�ԩ6m�[�&��j�O����-yb��Kۺ��N9�l{�%o�l��Ճ[�n��>�4���E��,DԠA��Mo�y�βJy�V>��OD��MV*S�+0qZ���wز�k�З���>��?�~*�+�-�_ř ~������淿e+V�p�W�Iu}�Q$������ZV�B��~�8�$�U�V�+ئ묷��&�3��]��fB�$J?�Pޡ��Z13�fqdh&di���o�����%K<)ʅ_�#@�Q(�(�W�J�ñ?�[��Ź������bG�9m5��F���gj�fգֻs����PiЊ��z��T���A{b�S�}G�]~����G[�����.[t�b����w8���uj��L�,X�B��n,��90�9�ܳ��^�5��|�=����z�2��-���UB�g&�����)���'�EA��?��?{B��_u>N?�tC`Q@��G> I:J�V���D�rm�6>��`��M��@M���ζro��};mݺ5�ӽ���L(�P){�j)�����[��pJ�lαϵ�3�r�fk׬�k���_�[�t���bv�m��b��GV/����|x��.��"O�BK��Q��i��fW\q���u[G�h+�z���1��3��8M^x���6ڑGg��=զr�z������
�Й�f+���)��Ќ�'kNN �-o~��ܼi��rY{쑇��?�gO=�ܵ
�M�2ɘ�SO9�;�X�0�5��~����U�a��kQ��E/z�O>���'�}�l��yZr�&ܳrW�?���bT�=���-��sfϱt��e��n�s��8��R&�v�5ۤ�����̆�;x�t���ٯ}��v����Kg3^<n,���Rv�BV�s�ᇻ�O�{��6n��A������ܕ<W�pL)���~�I��mp�����>۰a��{P�3���Km�aG��I[:�����{��7%� ���?}��?? ��/X�`qw���f௸{�e�v�An��>���b�y�F۸q�k�8c �9�g۔��Z���Jռ�%}�"����,t9�X8,~QM��n�A	 -�����Q���C�G`�G@>	��؇h��K�������i���JRO�`;��7�{�dC� ��syotB��2Q.y,�P^Y �[��f/��#�K}�TЯ�kO��
@�Wƾ�J���[.���'٤�]6��ok֭��[6Y�@�G;utu�o����������sg��46l�d]��R�|���h�\CA&�:�d�⬁�g�,jF�Y���-W�w�������ކ��rI�Z�B�������� �-��1�ݻǘ3~�d�� �>�F8�N�T��x~��E���?OS~� ���b3�\����/��k륤�m��nr�q��#y@�=��I�1��:�����_o(٠�`a�D!,:)�X�0V8f����^!����S�W��6�Z�����Qb�4y�$��N=��<�v&v��8�H�K9�t���v�]��D-R�	��#mGf��'���\n��Vw��!��}����kk����
�=K���c���n��ִ�Ls]V��U-nըf.O�2��}��| ��<��$d�f|o��q�!��)��B�k���.�GA��=��c}c��@_g�	�N������>˻{�96i�D�˱��W�xwa�=��?�w�����������颜�E��¥M����E��rJ=`�Qga@�I'�d�6+D��.e�n�:{rٓ�uTke?��^����|���������Iǜ�$���/}�^�{�g�������Ox�F�9�:�Gh݇it�x6g>��TÊgv�(�\:X��%}�^a�����pކ���z�*�M��aһ���b�Ja�h�T椌QK�ݶ���H��[n���<x(�SԮe��1Ӟw�q�QC���ֺ����I��� ��Z2��g����i��l���-�wh�B�K,��*�)$ӏl���W�&Y�.���+�K�I}�At!�$�aʱxT/����Z�*?�7���l���z��T���(?�o�G���V�F:sU)��M��Ϯ�<�(����@��Thv��tٓ���t���l�T�Mq�q����.��K�ѽ���5�y�G��H>�},���>V�s�\.o�	���A�� 4h3h����i�jq����=P��Z:|ہԮK��z�g6U�V�d�0� h�w�����/�ܣ}p�7 �_i�m��6����ydA�:_�$��03�}g��3�v���iQw��=I�zvvҌCᇲ�d;�c��c͓�"q"���n~������s�]H ����[�s��J�(t����9��\�<��Q�~���Iڵ��8nMg��Ww�ۃ P���H����8�"N<k��W�pfL��������t�v+��N�'�^h�� ��&�|�6�I�Rr����gqxƐ���
�5{�Z� ���\(t_Ҍ�i�hw�4�H�HׂD�F8�QC&#�i�${�(Xh�p��?�� Q�8mt9��=��,�F�R`���H��I{�������ꫪY9�Te3N}%�qR��"����ZXm ��3�;�Y�A�|b*�N4�D(Ś����8b%^+í��÷��0�`�?���`j�T�H��r+�|>�A3ޟ���1���F��q���u�b�|��i�E���@0r�E�m$�4�a]�8Gxb�oT6C�]��� ���[
݅�5�Ȭ�al0����ݵ�P�C��&l܀lB�b��y� H�ูs��_����G� ��|����ځ7k'��c�s4�����"��H���6����|�p�5J���F4��Q	u��Fo��s.s&
A׌��Aɛ	��g���]@0))�b ` 2����
�9K~�z�9=����]�曗@������/З(��I�S�%
�5��`sW���� ܓ�I�fb	Z=�����@���v�q�Ջ�)��y���k��U[�8�!�����hB� ��ڰ�$4^��a��*��:̀?~�x�Ŗ � ����b���;��š�qmX����M.����7��4���f�Цiw��o�}sd��j�Q������
i�~�H#��$:�g?��Gy��G�^"�D�i�wը?잼a;���w���e/�g!_I��Hӗ��"�#����<)%Nt�~��H���zaTJ��y�4�yXL�7n��S)XJ�ЇW�SFN-�^EK�okĺ�?�,�?��<h)��g�����������w A�5�@2v�{�����o���/�0��X��'�ä�$d��7"rX�h�Тb��Do5�rI�m#!�nc����O�n�d~�k��'y�]v��#�S����6��V~g�5�׽��노诊3��)ϭ�h�Q	�=��9</�Bx
��1S?��K.q ��C�(nY<�֦�T�?�C���~�v�d����� �IɆ䨘�ј��\���`l�I�fi��.�b�^`� Ƣpȕ�В5m�����beLc������0eLe0�g��Ɋњt��,��c�. | �u���8�9o�[���mh�с�������<�MT&�DX�p�C�x���x�Bk�)�����8�+�h�l��*i�!��NDD&�z�}����uɌ���{�J���ҾΫ��"(ش*�G�Y1���ַz��O��]�W`�����2�5XK��r������}�c@V)���F��H0��#Ǣ4} ��������=w�W�����Dah/����� �m;��Ԧ������O��ݿ�m�C��<�( ͵�K��i`}�=��z���X��t`�f�i$�W)_	�0t)��`ķ���8��bǵs����G��kk��%��1	!�D��eq�~� �`���h	���e4�M8���&�o|�;��m5L��Ip�o��q��(�y��۳�c�����$+�ͩ�
�CV�Ýު��/j.Q�Ma�d�V8����g+A�O������$�(,Z
�9Gq墴(6ȹ|�(�z�?���τE�j�b��-�,}�CH'�a�/8�����]�v��X�$�R�4��ź��[5�J2�+��#h_+Z,�V1��E�P�%��1pBkС=�C�sW�u'n�^
�<��$�HB���{��>M�R���Q�X�������^�W,�i����6|aW*aMS-����r�4�7���A,�4��c�\s�5u��V-$�<�?��@S���Vϱ��٘�?�,�GqB�G�d��%4��[h�1u�9n��G�ٷ�v�����_����Ų t�	�(�9�:�/�_>Ɓ�~��փ�����pD����빗Ʈ�4���@K��%��"��=�&9!�z�g���0Q���[o[;	����FzW������*9���`Q��^ba*�w�Iiq�I��	��  ��
H�s�o8����U��g��[-�z�q�V^�_�G1!Lrp&��X,{�	���PC��s��`��g��!�h��ڀ7�i;N]����5r˼����'��x�R��OPS����$υ���UO9���M�vϾ���%�{wzI]4���6&sR.���&��8i�Gċ4�Gy�#4H�{����2̳��4ƌ=��C��/}���������;�0w6�p�����w(,E��x��~|��O���1�� bE��p8�'��P@x'~g=b!���3���|���e;�Ph���)�(;�	�q$�F�_L�2�ڇ��~��J��E�J�c�j�;�9�5�����go����6���˓!\�s"Z����!<�����۔t&Ҋ�r�'"FJ�PցZ>C�%Ky"FH� ���&�����L�R�Y4L;͢FHk�f�x�21�)���SO�%�i���������/: �>�E�
`����6I�wؗߏ�1���	E�0?�6m�wN�]xw
�Q�	�j ��Z][��\@IQG
���s����������w��T<�a�5G=V���U�6�d<��z?E��"��(�����d��iR���Md��L�X 9���=���Xʖnų�7�F�  �<Y�R��(Q��bv}�Iu�l�f�:��BL���'����o�g�e�j5/���nj|@��k.�vO��&-.��Ҩj� ɏ�3�K1�9&d�i;�?�6W� k�5��/X
C#BD=V�XQ)--J�G~i.֕�;@qJh���Q@��&����m���x��Jh|d%p<�+�z#��kd�����w�6w��	�JCܟ�'���?��d]�����|�󰁪0K�ħA�1Q��X�_@��KE1�5[�����+SV�q�s�����$�+P��8���z&t�_U69�DU�a�Y��,+1�z6����`A��C(���<�1Yj��O��u��'�d�7���}VhKz����P�֮]��@��t��%���'�����5��o
=�5���i	�_u���PaS)��c�����;;;|a �;�&�@ ��O}�S����|w���b�V%�BT�P�0єp��PBVB+�'II���Ɛ��p*�P���'@�;�/Ĵ�H���Q��9�Je�����@,����yVE^�&y6Y~Ҋc�E`]�I4W��8=UW�x����@�gx뾚�v�'ZNjY�. �!�MTǒ3��;�·R�>����{��)Q]�J�:���	?D{��V,���yq�c˹����c�'�k^=�GN=h�K�^��z>�jmE��AQ!/��$�9�Ƹ؆�@�?p{�.\��B����?]S���>�>t�,��9ȗJ�t*�<hK��o����cB1�f�~�kV,g-�MIF/�a����;�vXDT�r�Lf���|:�쳝n�)�8	�j����P)8Y耇��:�
�m�}�}+���%s�<� R�x%�(>����Gs]=�"������tc���6lp��:{�E+��*���=���q'�^�0)p�gfM���;�Qk�[`C�a�H���`1T��o�����$��������;�$K
��X��O�AEO|K��z�~����y�B�}	ʕ�=���x��9a�u��N���s����~��۶�p��k���7
=�l��Z�ڏ9�h���WY��édS�`۶l�%K���֯[W�+���	�og�=Ϟs�qf�഑FF	g&P ?^��� ��b�U&??L_��|��\�S%P��]W��fϱ*���<�Ѱ1���}wa�h��� پ8���Kt�������AQ�SY2�c-V���~��� �.�v7cރ�NxQ]{��㋢Ě�'A���)�/F��ͧ?��\P��}R�.�)'i;�G�]T�:��3�K�����T�Q�W��(�/�fmA�~������;v�w�̛7�#���k/��^z���O^lV�X&]�'�\b�V���Զwo��`����{��v�igء�fCŲA��w�u���e���.���Pxw3�VC�c�:ʮ|߻�R�l�҂%[�~����{<�'�	�#^,��P���*6�������rV�~�eJ��� Ŏ?�|(�a���.�Q���h�8�����Ƅ;��,�����Ak��׿�NQ�nc��o��h�_c�@��;�ck�x�V�_�-�-V������>h�$�)}op�Ҁ�����:'%p@\8��'�Ē��西�ۿUVk���4x9dꣵ�e��4*ψ����x�b����ݲ�#��+�^�w�(B����A䟀�j��Wi s��W;ː��l������ۭT���N�J�N����vX��������3gz�2�/}�Z�0��8�7�\�](�yS�'ڬ�=�������:�+���G�\�f[6��m۶��Ѐ���&��d�;z�ڂd    IDAT��3`���]����ɇ�����!M�@&��w��Zil���\��_���9�D�Q�5
�=tl� #4�$q���}Ќ�Iʂ�F�_ ���}����[�h7���z?�񖦪��
9m�c�pH8�.ມ}�M�7�_�'
��E�ٗ���z�s;p��g��1s�L����.�3}b_M;k�s��wQ/�۟�2�4j|"������]���wgw�}�7jU*�? �/�B(�.������3U+�6ԷնlXc+V.��[^�D��l6o����y�����\iO��x?�������:���]��bw���f�_K��G�9�>�����@�M����n��.��� ֮Ya۷o�\��:�]�u�[�n�Y���o��N8Ů��
7�]�Z _� my�ƍ��H�yի^� �{*zB��g����*}��z�ȗ�ǚd��T_ ��
�����w6 �Ɔ��;���X�o��}H����w�+�BY�� T�h��rG]+����D�z�Nq��G?�dAU�P�E��u��FT�	�ڇ��Z��������o�AH�r=�&��g��%�g̘�5���|ͺ#T�dAA��X8c)��	��ՙ�O-�AC#�3FPP#3���07�&NX4&�q����d"b"Q.	J�F�^�`��@7�s1�xM��#q�Q�iA��޻����WOq(��k�jY���t�W_���<��>�rP�x�Y��M�Jc�����׭5~�ayy�ik��wW�o�˫͇��7�1�w�W�A���u�Ŏ-M(�i��H���<d��u�d���_�5eʯb��݂?�燆�������M7�p�|���<������Gc�MC�G��9f7L4Ti6|LPg�Ix�f����QGO�- ?�E����8Ё�<�P54 {��G��ի�Xx��J��^fF
�;�?��?}�o���Z~����[���Y�%��:�d�fu䘳>p���� T�8w�~0J.@�9h"�S���"X�6�M�EO�%
ȋ�"@1q���yꩧl �@u��$��3 ��/�Iu<=�("��RC����0�a'ث.��0����7W��>5f}çf�A�������~����ֽo�����bQ[�ߚ:��-��K��<�Lq���/2ш1�]e�������cL<�l>��cӴe�Ow�+LӖ6��ǟ����yo�f3��/��.���0l*�@J����ۇKI:"`y��[-=|�p3c������8���,m�S���R�A�C�台�.����JM7�dG���k]�G����g&���M�TI!�"�'��-�.�5� _un��<
q�|�X�d���Y� �|����_wQ>�f+�y�ր{��,��^ u��M56����9r�5 �V���QG�6���}�|P�.�$a�zM�ii��-M���%n~>w����kk���^�j���g[�IS&��m�$�����u�Af楗������d=�����<�$����47��`h(j�������ΐ���Ō8� ��N��\s�]t4�ܹs-/�;L�>�Eê��&��c�)�:@P����\௳ v�
�l�����MK��ϢH*��1��m%�FA�����V����hH��	2�~�Q�Z]Z��a�����~��t���C�˳᧒8�X��2y�9�G���;{Z�s4�C��|��]��3G�=���>f�wM{'����6�xȼ������N�HF̜��7Ѳ*Ӵ��zZ�Ye�?��UԖ��)S��/��P���G�0�~t�ikm6}*#�ŏ��i���f��LssS�(��ټ��ԯ�Ĵ�yf]}�w�?��*�}p�(��h��1cl��,����F�0dlD5�Rj�
Tz�i�/ �2�0Ȳ
��eec�0d|�,l
�y���}7�ߵ����Oh��;��Ϻ�R1�}�]̅hy�<X�Z��]@6S�Em�C`��N��@_���&�y�1��c�W��۾� ����Ƽ��-�67��_z�x�P3`@�z�*�mNUl�������۫L$��l�3�c�8�_L�>5�ݕ������?>h��/Z�����s�zZΟl�2���!f�W�f�;oϴ����+�j'�j~Sf������6��Έ9���e��T�e~'�kN�'5��xW�/]��*e(��\bU"��r��)p.���
��B�jN=�T�{饗� ����L�w�cU�?�%��^��N�F���_)��.\h���gk���m�R5�Kɳu��s���=7���+��Wz-s��o��k;v��������%ւR�<���iv��u��0��m:y[{��:&u6���'����]mZ[�滧�iFr����k���^��C�t�a�Ǉ|Amm�}E���LY�5����������ϛ��C�d�;[�����7�3ﾻ�������ܞ����io��ƦN3쀃�q�Oܦ/��Y��<��ݨT2rF���*
c��	E--�=��rnfDO�?�������W���(��{l�Z��(�02
�10 #
��5R�]�$'I����V ��G�=���v?`��;Nl���nO�
	��||,g/�g���b��b?ślX��Gٲ�Q�jAk
2���V�����u+͇~`�;�MUE�54�imQ��xɈY���f���jL��l�����y����r����Wjݱ�/Z�h�=���'?�;3�Ӷ��:�/�O7t�����g>��`ֽ�����?���z��N�
E��Qc̸/kF|�M�b��T����c�*Iכ�'k%�e �/!S��Z�͛2�}��kv����g`������m����ݢ�l��a�_Q�����R��B�?�F~?Z.�>���2(���X��(Y�
����qXQo��,�G��œ��>���Q����I��)�FԨj3x�D���7&�n�Z���_�����^5��wXs��:ZU��|��c��8ҔU��:���j���{MWW�Z���2h�E���w#�?�;=��O"x�3<�\p�~��6SQI5/�.v���&[�a��>��4π�M(L�0����8}6���S�G)�Hq#�p�|�@_���������y���!�s��P�}uV��J�T���ϗk����@���J�
HRTUc^�o	��S��8ܞ��M��U6�/�`S�|jW@}��/��v����Z,0�o2�ԟ����~ �?cٝW�-�L�K��U� P*R�M`�ޢ�T$�B55�S���Y�<� ˥I�$ݓ�l�w�3��N22��0~"}er��*󅹄��ء�m�Y�V�N���$9=�Z!�x��}��+�@�t��d��P晲s�ռ��u��4�4���I���|����oжй7�p�Ut�r�<yW�T�Ϝ��Czx�J:��x|���wW���B!�|�!>������U���o[ϊq�zy��4x��ŋ�Ut�����EA�Sy����T��iXm~��L�l(����k�͙��A8�� nZҲxO?���JQlmb��ֳ��ci۾(�d� o] +��o�l�w�y�n82����¸d�Ӧ�	 �߷��4�8Nm>�	��N�� �%����Lj��	��1Gw��{��ލ��� ��\�YʖM+�W��������)���.��gP(l�p�m�ؼiQ��ś3^��s�̖R��e� �|�?���i�(i�.G
�"< [�3�Ea�1�ָ [���@V�1'F�t�_����A��}��-��J�=�5/R��Q�F�8cE��9��T�=k��>�2{Q���x����I��}��r�`/
��!7_2�Z�Ƚ�KH'�I	�=��y�P��u��9)e>�{)л��@3n�eW���d{y^29dА鵵�w�O�2��Xl�iYi���^r�%i�P���2�u��p�b&GY�dA�B#+��E>���m M�g!N���D�p_���{�9��]ֆ�g����V��:�'VY���o��;����,O&���%o�k��l[��WXA����[o5����=�@�a	o��
�@���)�٤,X'Z:c�1mf��OA-Oϥ6���U�/`�����R����n�=2!0���f������<�J����?� �?�ܒ��u?���+��s<2���;��sm!# i��3�5���� BN~5�����IgO������H����)����d�k�0�k���y�f���4L�N�b-�Ħlz~�Y޶�8�:s�J�3g���@>���yF}�����K?��/�j`
Ɣ��xd���<�U��~;>�	�i��HnZ�<d����u�.>�8��b����2�m(ֵ�N�,~iu*��,"`ON?�}�m,hr�9T�ŕe�=%�,�[\"�c��h6n1�Bl*�q��������m2��ҳO�4�o斲�mO��
�;u
����S�>m��WUT����y��l&)-�k���x��h���r�=�	�]*�g����q����7�^��\��Qq��ѥ�v�`�x��z�H�\����SbN @��w_R�Re�} 2d�,�=�.�(�~���chqrޙg��>7Z�>K\�b�-�1�Ϥ�d���[6����c2��s�O��g��{}{�F)ɪ�QCCq*#@ԩ�J~b����w�� pƃGKJ7��Fź�]�}������C�e
Ƙ3)>�xP d��ٯ(�[/Y���d�Ew�O��(��N6�P��&�_ZWՋ�����4��>�$��92a ���
S�xJ���j�An�� (
E�k�IG�*j�T	cM ���u���J�rS0ڂN"nA�GQ����d|x"<'9�|�R۸�@UHV��R�6������*�Y��&��
�G�bL��8����]�Ck!��뤸v%��'�LjL�����di�&s�����҆��|����7�W<+� ���E7OR}�1�wJpd� �6m���3-��d	���'�p���/Y�ʣWF�֒�g�jf(�M��?8��,���3�z�V�T�2�}O��`��KT{�q�x�������^a_��`�^c�6U��Ŀ�E�fƈh_�oK��simm����)S�b��og�d�Xx-� �u�]Nյ�e�sf�YH�G��ʱT����D\�xg�ϱ�\���?��u��a{k��`|?���|��M���?�����pc��bG/rL���	@]�������������B���y�~ �>�:[�L���}{��~}}�H
R���񂠜Di���������"�2t�;�ȋ���Yw����nv����3�N��q���F@F�*��z(}_YW�||�Z��|?^�&t�,X))�����:�w��7X�^s�g��W�j�	䛗xz�${�1��Dɸq %> ��)) "�^Jo������/E��3�%Ydb�0�k֬�^s X�c.�,���7M5)�[ލp@^�"�H{^�\�EJ�>��-�������ű��)��_���@�)��N.g,�ׂi)3A��I�
�[�wJ�k�
tt��o}%ҁ%��r�c9� �Ud,���J�g��R XԎ��x|��tM�����/ZŢ͐���O���>���
��e�5�@���f���l�o���<3|�a�2���gPX��Z�?�Q��8k���ڂ�9����z�QGٸ��5�*��}tϋ҆:ԚBy�(AY��R�2p�K � |�M��K<��ISK����r�
�?�D�7�H�~�<���=��+�����9k��e}\�'��ε��KE�6��c��갺y�|])��xc�l<�ﴷ��(�[�F:��N����b���g~?����Am?s���a�R4�.nHaK!
oDm2���d e�=�Sy�:s�E�*>�2��X�qj6�( ��L����ܝ8�dIZ,�A��U�h)��7�{��J��od�5�CX ���{ �@��թB.m�*�Y?�ļ���nu8d�w6��!!�6c�!��象� �x"����������,}ι��=����$_���e+�U��`3纲A�lN?�ck�[��c���UJ������������V��D� J�C �~D��PV�A�+D`��3Go�����!N|S�f��D��p�}Cn>�$0��(*�/Y�X��/Xʌ᪟α�*'����d��k��"� ���������s.M+c�k�RgϞ�ND`O�	�-ݚ��d^dy���Y9��h<cP���衇ڸ�G���R%�̢.?�Y���\cEϡl#)���Z���amm�m%�O�����d�?�kd �X��d[ @���� ��ȹ��z:��H�:�`�m(��Q�6֩
L ��+Ț�Z6�F��~b���2b�� d_�m�@�����o�_)����Y	xc��I ������Y�� .:��� i��Rb�����X۠5b�?�я�gB�(
O)�xU�.2$\�����s�A@A2_o��Ft\����͂s<����{sv4��1��O ���� ��/À7��IW՜s��f���|�i^ޡ�͟k�H�C�"�,zf�����]��+Gm�0�JBI
�ˀ�U2��}��naݭ%����_�?V,��SD����
�m�`
�@�2��7����s�)w�7%%e��r�-�2"�!P�����L�����Oa�����?c����k���8�kg���O�1,�Q�F���41"����ǈ@�g��W2�I���\?�D�Ld��Vy�J]���|3>y��_��k�I]�O�N�VLbW���<��kkko):�<e�c�����h�]�0;���Y�JU�u8F\m7G�;�*�{e)�9e��9l�N2��;�;,�s@�Ԁ:Ԅ�����[+?�����9Wm���l��--�������Y��?��mV�G����W�})�".!�������H$}�D�'N�'�W���qO�X�7_�����}�`�h���В{����ߕG)�P�W4����7{��1�}�����̪[�h^с����o�&���O6�w�'PKJ��q�A����L�/ik��A�?�?����4���	 �^�������F��ˣ�>�\q���anPrk 7���	����s 	����K\5��B�?�r.�$�W@� .� �,(�ݦ8�b>�d�'{�TfёPrx-J��	�fƸ�3;�������\�����(�Cr,��Y`C�� ��|Emm��%���h,#,������
*+�$|�ff�*���m"~�}6ΟTO����(`� �7�'=��C���( ���PN��p}��e��{���x��,��Iٜ�����?�NcA2�|i��Q`�!��CB�3$艵��@�9c ނ|)��A�}��'�M�m(EdIVv�\��v�.���)��w.�_��x�����(h+�'S��d���Ʒ�ͮ[TwS�P��g��ם���5bQ��[���& ˆ<���m��
oد���dc 초����-��!(�!Ç��j��T;2������g�W|�8X�>A�6�_�	�����	Z�fX��z
w&�KcA�'���R�$�
���^
��"�f��W�&�C��^�_5��,�w7#&׶앩���Q�x��񳁿��w����*~W��(�ނ����S&�6�b�?�>�( ��<k,,�P�Kr	�6�r�*/I%�|h@��*<�N�Y4�8)u�M��1��M)\+�%��_�J������@�o	�}P͕��Z��1!�MX���?��r}֚���Ɂ�'�/y�Q�ɋ葇ӅK�c�C�4oi��#d�'�T�jŐK��ݲ�1n�I�t-�\��˂��*�E��mo�zO�[��?)��CO'qw��;�_�� �y��6���m�6�v���KdEʢ=��al����w��%ݓ� R���,.�
K���'e����w�%�{˟N<�B�?�?���rD$�Z6`���`i�    IDAT\j�'���@J������@ܢC��1��P.j{�ߩ ���s�1��d\1 ��y�.��<���������ɤx��D9�j�He��.R�ʣ���Ӥ��Naw��z"�-j���w�9��������:X�8�^X�p��9V/	�@��ķ�M��|�K/1���;����{��M/��\�2>�_U��L����](	��9�\h���� ���-rÒ�(K=d ���v��W^wwy�=ɔ���{s����3�.�e���R��t% ����yE:F$��y���/���x��������Yg���/�˳�7z�@^:�2���q�SEn�<�WM�,�'�|�ƕtɹ
����E�6��M�8hGɂ����ރ�Ҹ�]�]�y:�2��E�a���)Si�5��
�_@Z՗�'mjDux�(�Bȱ�iŠ�Mq��բ@-�y^ �9�?�n @W]lF5�S/��x�0��òǺc,�r+���/@�kh� �����k��w�A�(z������]EQ��/pI�d�駯yU]�LGb.s�*	? �,B㩫+S��52R
�x�z�W��ǖ&t[0p=�} i��B�P(�G� �T�r����}������9�w�F��Y�ъ�zRT�5j�o�(V�+<���0��������ŗ�?iꔇb����S�?̓��`�=A���b8u�+��T� -B(���-��O��=��-<?����<��s����K��d�;�?@��/}Ɏ�!��q�3�=\P��ML�7���;�$�K��d{�m�l3CRV?���~�^
@�� ��?�{���ώ�K�S�bs.P�okB�/T~r�F��5u���]d/�~��;�3�?��24ħ�� �mj��R.R&:�:�X{C�=�<��C:]L��n :��>�߿�GO=�D�w�<e��i�5�!��)��V:�
P#����\RH���XHV���Xx+V�H��U.����	����`s2ר���sp�ƹV�I�5���a�A?���h�"[�K��P��#&o;�KV��)���y��S#�<��؊����c�  (�����l�[)��v�gw����u+b}�I����#�ܐMƩy��� pU��|'ʜ@$4�:X� ��c� �(2��3BYI�!P=('��w����'�H�v,͚�{f���O8�������ŏ_?��S���5�Â��v-��@3�� K)�XH_��K��B��*vt�M��f`#�7���j�q�]�p �i)�����e~^�� Y]�8��a�Gi�P3:>�s��w[AwG��T�BQ���Z���P�� �m%�_�M���m1^x�U��T��ۄK�/V�w���a�J�����j�u��\�C����:~�Oz����O�|�^ �뮻μ����j��?��F���;ڲ��i�9�5�a�o�
���{�N�U����S���"�V9D�v���1"`|]��;����g^�0����|�]����O�')�vO��Y���*�d#�	A�{6  Ϧ@�-�ʝW{�̞��VIc.h"��s�Il:�uF0o���ҍ�Ld|6^p�9���`vu���#��5bx'��k�eA��I!�݄�/��T��\p�����r� P���S
�>�\|�V�*O9h� ����i���h g.�I�k�	�gm����?�Mx�4�|��Nu�d�-|��U�(/Q�Ɍb���.����j�����l=����x�s��a>�У�)B�r[cc�=�~XX�x(����mm����aWf�,���7��T<�VV�{������8�b���ӛU�� ���X��lB62uӗꇱ1F�1��6�!���(*p��#�1�?���R��ݼ��<��)N�˟��g�.���,D�e<sQ�r��$)�C�s���{�N�H .OS�G� �oϝG�U���2��N[)-Q4���߅|�{d\j�#ߜ ����I���]9�U.�x�u���u���o\��-���L�n��ƫ�T�OgJD�v#!�X�X�:��M�S>����tK7��0!��'���@�?�B}�y��C۸��5�Rg�jL��;����+} �j����Ac�Z�j�Z�|k8���-�K��6P1�?����0?�?��%�-M����8�Y2&o��e��d��1l|��	��t�WkKO(*�m�>�g�)��ؖ�Ke~rO�_^��+Y��TRyԒa�0�H���>���[����4�/N�k��������oO���'�3m~��!�m����K��4�":(�'V��$]�]s�VѲ�]�K�#��Apw�M��`���i� ��z��d��]#���Wq�֦n��.�W'11�dz�y��f,�yF2MHC$3��J|�Q�TO8��LJ�J�eZ�C�馛�x�����9Y��b1�7�с�2����x~h}WZv�er�g�X�(`e6�5�<gbܬ��;���^����w���a��3>,h�V�#{���O�~���z477x�7�y�O��7��Ͽ���^_������W���Now�Vs���Pv9V�<��5�  ��'A`0��O�P��݁��YY��=�!��( �� :�Qx(�8������K'�i��o(�e��pjn~
��W�=�%����g��y���`���yꮲ�>��������ᕒ�C\�s�Y���1�8Lf�ܹ�������J����&g��w�1�ͳ�<�[�w�ڢ��|�G|������l����=��]s�����ٰ�e���8d�����)k$},A>� �H��f\46Sa�t��`�ɂE�͘1���~hSr�� ]�E�qh�[Z2�0�^,h�rt=�B �����O�Q����k��?���y�I�ĲG��ƿ�� �W���Jnh��}d��k�i�X�6��mW�|D%�g�d˟uW�+��θ
����e7Ͻi�	�����9��˗G������۾� ��"���D覻;�+�(>�wQ�*+Y@'�7����lyv���H�� �A"*�`����)� ���;��������aEqo
��P��>H�$�"CF']1&�
�����߰�I���u�.�ÒgO�g.)�c�PH�A� J���w������$���o[o�އ�=�3c`Ȏ��x����.Yzaw���3��(��O�x����Y��P�]*�W��-vw�����С�d`(8���Im(�_�)$��͟6	��un��RN����c����= +�-���q= �L��Y�����KA�����Һ@ֿ{���f���8ԅ�o>�Y�FoZy�V�?��5'�S�H����'D�
�WZ�^$��?xg0g�l��T�2��ֶ�	��y��=[���5׌[��s�Ps�ҽ2b�Ӽk����_i�n_ײW���b�\|�S�gf]�gm<�,�Ϳ��J������a�Pm�p�B[��D�?ܿ2F\�E�|ƯϺq(� �5k�=xE�\�	TP,��]/��C� ߮'�{*� F��d�`TA��8���6̤%sp
��<M� 
��ۓ�}���7��Omʭd��.���rS�Y����7/�q�)�?㌕E�<��c�}��~S�J@���}������XG��4Qt�jS��|�3��<7cb������%�����8M�Hl,��*�����Z��w?�Z�����d4�����¤/�I��yEQ��"Њ�̳g�>n�:�Qv��?�?@��!������Vz+nB�k����ϧ� 뎼�P9���s�I���7��������@��ͦ�~e2�s��o�{�-�A�����ڴ����sX��R?p�z0ϻ����`��"q`!���Q
�R�5�LlO���SdD�/Y�
�a	`j��P�?�x�Ny������#e��w�ːB�'=� N]�tU~RYK���eZ�x����?�wPH�h���T�>�ޟ������/c�R�������<��axfd<�_�}��˵����q��յ�k��o�qyу]]ݨy��-����6 �pQa��%`^�޽�孱���&��f���t?F!�k�Me͕5!J�9���LOr������ٹs*��wS%L(�2Zb�����9p�pǀ����Q$V>Y.��
��J �'#��cUc�B��=�>3�a�ųJy���ݺ㡭6�N��3�����g�bW�G0n(�y�7Y���(�"�L�//]�9�O������~H��+
�2x�Iz~�p(l�xZV����]�.�P�����z����s���:l��t��m�1�c}Y+�*�tXŠhT�{dUQ�-���lsR����~�UH�b�T�j�\�ϧ�rʧE�L��i��[�z���x|�N��F�
���%m.ޚ�G>7�c[��[����'�! �r����>N�K�\��75nN��"�)�&�w7�����E_��<U�r����`�*A�� ����'U�X�|�@������J�T1���Bʏ;ܟ�S��HhO���<�h�J_Ei��g�� �')�/���y�駶i얹�p�s�J����!�#wj�)t7��w����m�������-P�ޙ����
��a_�l��+��<3
�y�M���O���ȅ��HH(�\tw/��XEvvvn3f��{��/Z��*ڇ�_�`�~,�;O?Myy�; ��E�v �F�:�r�7�Y��>xܸq铓�LP�tEU��˃E(�Q��m�UQ����L�|��L�cu,_�Zuڤrְq�f���yq���.��Kyq/�	J�MN����g�B�j�\/���t��m�V�*\h�p-v<z�C��l�%p銟0^�}��Ȋ<��s��3�ِE��SOn���sJ�?��/�0�̧*�W�[�gf�Y�&��-CF5̽���ho�b�ʬ� ����q �]�_�N�S+y��DQzmy?��dXN���k�O���O<����\~��ǿ��˿�ӧ�H{�meEZ�܉��s7C!�����r]^�,0�!��e�a�;6����Ea��Wm~��_Z^V�"�Ue~[]������TAO�M�>��yYm���㓲�d]���D҂?�̼(��!&`ѽ�,�^�	�wQI���O��z�(p͸�QQ�'��L)@�O�QAA�>���m�E�06�g���4ߋB�Y�lN�G�b�#c(��z����`�R�G"w�� \zO�\4�s_��%���}�q M���p����_��| �����U�<���^ߵG��Rm���rV�?��y���)h�����'�|mCC�%����9�J�]��K�4��D�ȍg��:�hk7��~�3fL�e�F�eVL������}��g-��� ��<w�)�9(gS��~7��sdZ��m9� ~�6(�Ϻs$��C�v@�����/����(%'�r�H
Yi�Fۙ�5'|ʊ�'2�zi���~P|tO�z�q+;H�,E!X�����/�} 8r�a3�%�Sͭ�S���_~W�T��p�G4��h+���kC���[�-m��ȋ�^d8�.�K+|ݏ�j��.�3k�Y}�n�<�ӯ_����_��#��ܓ�/:�gRx��!,��L&OE�宥�����=Y�\׈��e��a�6iA;��@����<����"j�,�_֢��I�ϊ?tw��y^�Τ�D{$y��M��pĔWT��]��d�+����w�G���a�1?�ݑ�v�$4�X�:V��x�_P�T�P��QO(��K�R>��9�oX�dĐ+O!�㓬��c�+ݏϋ�p��֓�c�/Y�����z��B!�G&�%=�C�א	��UUU՞�<���:
U$*�=�]�s!kY�e\娹Ҙdd�������s�(�C{j,'�A���sT4/��Mw�W �L�%��m�ng�J�gȶB����%���W]u�'N���^E	�����_?lٲe�&���P(�E�Z(�mƠ	-��|�����
�d��
���cҜp�rQv|7����wb���-mQ%����/@K��*+��s�Y�9bd,�G:;;�^�y�U�!Qc�6lذ���/ZB����,:ml�'�S�G@�^�������ŊP��6Q^����B���M�Pn4�#�5BqṸ���nZ�ƪ{�l+V�X���}�z��6TVVvvvv&����x�kkk�.qsss��7�<�����D"1�ϩ�R%N6�;ǢQXGY����E\/%�idz�?��}�dp���ʢ��mŕ	'�Tb���;]z����P�+���TC�ВiӦM?������E�L��W_}����vk8��#�b�Kg�t�����u��7+@R���h�vԑ㶩���=l e�P����Ӡi���.g�qh=C�����)P�(-��O���֯|�+����y���jmm}���	�*|r=9�f\�R:.5���)��,���<{�g]�s)և�9����Ҧ1�J�m��u��ׯ���c��3��,Y����n�<�L^TQQ1P��F@�m�P�R)))�LP����nR>�����^����I��C�6�#�S��{K���!X��V����>�Ogg��&M�����/;r��&j�̙_x��7~���|Ruuu9�� �+���L�uG&�7�u9J崓�uhS#c�y�\�6 ƺéM���V�����ZX�x�O��o��/�~�ĉ�͛�yPvwwvv� q�xpV�y�mv�����92
`� `}}��	&��\���5���/f���\�D�)���K�i��5k����WJ�QG�{b�����I�V�y���	<>eE�{��vw�()Ŷx^e7��ʮ�3%N#E�꥕����&L��ùs�Ο��H����Y�f�O�YUU%��!(�rPQ��Ke��=hs�|)v�J��pD'%���~6S���
���s�euf~�P��VvGJ�mPS�ȕ����1��a��{�wP"�x���k��/�uQ@o�fv����R�t�u�]���N8aNO���g���[n���h����d�E��Efܽ o*����\��mI5ֳ�AEe��� �:�*���������'��(9A�O*J՛H$:��˞�������:�����&��;o��§gE�E�0�:g��M 4�S���{�.gs(Sg�j�i�e���E�p�����M����8_�?���W�"�HcMM��ٳg_s��Gg��S���1���NS%(��L��<=N8�閿K��A�,׭[��c�=����|�w�q��yvuuUD��#cU��������i�lRY�/���˭�p���|�S�Ac���x�{|�ғrPFolll8p�G'k�܋/�8�>�5��;����O��������G�WS3`BWWW�F\�@�|a�I�m�P�����o.�W.�v  �O�}D�d)��H��~��UJ��Xuu����}͸q��s	��yh�%�+�1�(h+�_ ��"sn ���[���	A�$_��*풿�8��L�0�P(�p�'|����Λ7�Ɩ���*��?Q�W+N�o\HAle�Q���ԙk �2ʌ�� �έ�����O���gd�RJ!������C�wڕ�>sҨ�:�z	����n��sK�~�g�S*+*noo��!J$H��6o>��g�N����~�K�2H[�X��&+����t_��� p"[���i�a��[��kN:餜TOj\�c�<�+̯,~Q?���xBA��~o�_���;>7�@����q��{�8��C�P���:��˗W�r�-��dӧ�VTT�+�\oS
 �s��Bge	+�!��������A�G�ic�{����lR�*ڔկ،�&����k��j���5gΜ���^k�&{�=.���#V�Z������-+UQQQ#�I�-�Lv���l�&�|7�M�e�g8Qy6B��>�΂�$�������o��7��>�z���d2�`8>��� �G֒� ˾'߷'_�&��A/)�mݸq��cǎ�rG-�ǲe����_ߵ���*p��.�+��̜�H  �IDATy�C�T���>��/�V�	$v��Lr��^A�A�	��h9� ��ۦ��������:�����g!���=�͟��g���u���S�x_����D�	�BeA�Y��=����$�t56�/碌��L�l�dM�B����S>�+�r
��M&�=u�W���O��ӹظq�QMMM����k����,)
�h��+(�#�z{���9��3f�V9�1�S�zÆ�ǎ{��X�����ȧ�x<>����wSi��1�}�qf� �A�c.�WO&{-�4�S�D�o���}_�-?m�p�)2%����Æ/=dԨe�_}������%�߁�������y�o�f�ڣ=/1���r0��1������G[_���m�c������X��l-�d�+�F)���(�!zuvt�C�Y��b�!���dk�,GnL(�[�!i4e���I�?o���ow��ߞ����[��0&��x޿W��{�ҥKw(?��������YC��h�H��СC����&�Tjoo�ڰaC���2���E��]�,K�·��gw�}���9C�2g��i�������p+	�{�����[B��F��^nhhxvܸq�������˗W�����4}��}C�P�"��}�z���^YY�d!C���}��uo���߳�dS"��������(e���3{^��8����Ic�e��m7���D"������5;�Õ�}]���m��n���Vw�X���i�<�-�յ%�%�G��F�<��G���СC?�6mZS>k���R��Ʋǽ�dɒ����������6m����N$�
��D8��ɤ�,�3&	A�d�/[�掻�q�{���F��x���a��q@�1i<�Θ4.~2N���O~�߾��"a�ya/�¡d(i��ԘӲ��1&�������pg(jO$M�H���΍w�}�_�������w�jjjD�����Ӳ��pWWW����-�d�-5���ye�%�ɴ��L/0�LF��p��<����T�B!�3�L�<��o��S���z�k����9��K`�����RH3�]��u���d2�Qc�t��y�
��P�q'��L&�{�GH�1���J$�Ϝ�e4jMd��:��h[(�t����9s����px�>}jR�r�|��i��~�`���/o�{����>ӽ_����R�;]�lV�<�8�dKE}��P�}:��%�:]��ʪ_���TD������ͻ��]�0s�ѿ'.�{��k����m�lI�w��Qm���*/-��'X<��j��/�Lߗ�~N�Iw��~u����Q�G֩.�~NU�6t��Fc����q���K<"y���!��ˉ��g2ټ�OJLI[`��j���A����mP�C����X��9�?���cfAt��S�b�b��_)��%��i@k���1O=$���&,� ��~.�� PK   vOX@��)  /   images/b4aefdef-6992-46c6-bd27-cdaf728c7c35.png�{eWM�5��I�� ��w�;�a��]�kpww'@���;�>0�溟?�~��յ�ԪSGj���Qj_�q�(�p�|�@@@"  �`��롭���w�t��熀����1��
W�,��sރ�ch�!��թb���A&��A怳�>���P1��c4�{?�ԗ̈́�p�i�7�o���q��'Tj��7��+ ��x�t��5��@�4ic����}���R�&�%��_�&D�]���]f3�d�Z��4�����H�Dc��K�j���]tЋ���2������o'*�k7}���������vF��*���g�u�ҴR��FR�(��y�J.���{���>u-y)��ȕ̚���7���/��L�B^��Yz�v���~rm�$�=ھx���%����$�p�(�ێ)�b�d����RW��#|t�#ge������&$5O�v}͎��l�<��էa```v:_��(�m�Xd��!�wgKG�}p�9��q��Z����*��Qp�!S��r0���t{�M�����/*��s�OV���1����3�eȃ0 C1�H�1��Z/[,V��c���~h�~��y�o���}��!V0oڦ���\�#�<��n�����E�v4̥]���<@ �!T���x�ف&dlJà�m������b���-�Ɨ��u�(#x��)���Ŗ��7|x�Z�j�S��(u�2hU����Y��W������ݦ���Ԁ@��Ga߾�X�Qm^�{0xy���pg����w�ל���/[��cu<َi+�u"��ʨ���۳��I�#�Uc�&�[������׉������ܱr����X�rAĈw!��/��6I�˻/Ty�O�R�0�,�8*ɽM*�}�վ���?�kV4ʷ�%�Û��1��[��/uzM�g�P��_a�'y�|�1���!�cQ/ے��恑�x���w��0y���#j^�gX��n�DT}ҨL�@�"9�=H�y_`�~/*�W%�L�kH�3DB�5,�W�@?{���<��������ѻ��껀��	��/b[;��W.�܍d~UI�o�/����R��6�P�wWа,����T�^Nw�A�֪�����%����t��'7��Iy�-�r�|��cC>�܁�������k�8TZh%嘙�k�,lV3�U��{��T��}@���旜�4ӏo��g�.��Bv���sfK=s��:����ʷ���L�1����]�j���1� ��6��uj�[~|�eĔE ���^���/�O~�бd��v�z�7s�2��L��xm�$dr~�t��������L��E4O���q�~�k�9�C$�@«��
0*�9�A-p����"���A�ݻ�ޜ��۟�6�[t�s~U��q��x���}Xń��y��m2ß���É���R����[�gb$Q3�AȆb���$l��TDl��4�m���NIͰ$��te��S	�)��>�9�'���B�Ѐ��k���vgCFt-*�P�ط?eg�Y�ny���N~�
�57{zz=���a�	�ãNݧq:.�"G���-D���e��'7u�\aww���jk㷎wuj,8˚3�"�/?*K��:�%�����v�v2�1�bf(1?���4.�I"ɍǬ��^��k�N���ɢ������"�ථ�T01�Ѝ=�ꊟ��:&2��f~��P�O�Lq�?���N���r��`l�e��ܫI8�������)�,����_��K����>J��r�9Ih~yC���)!���5�н}������[����T�'�-�>*0��ʏwLx�� ���8?�|��PK��O)�I/W.�v�x;�0p�R�l˘�)ո|��,���/��'��:,�d��T������u�b��
��%Br���w?���iI��Q_bu���qՑ\�#���#��(a�t��qeg�� z��"H����l�D���b���.�ө�n��\{[A����a	{Iq&��K�vGm��c��q�h9���
j�h]��<)Iw��q�U����դ�倛j��^ ���������\���D���->�ao��'e�讛���K#��L�FPJ�p���/�_"K0v��5���h�	�80�kw��t�y�V�����U���O�Gl��t4�ʱp�ll?%�!7,5:���n�(�6�,:��F�~��%��OVfJ�z����I��P!�����'�A��F�3���촗��p�(�?T�E݅аA�F��snA�
�ϥ�=�̴�#�b�gV�-�g8����;��'*.U{q��  4E�~���N�I'���P�x��A`�*p���C���Kښ�'��O��A�/6���ކ�5�-'_dD�ۦF����Ά�()��]�KLjQ�E�~NMq* @��5���C][���pQO^x�/�-�&y	��� ���e�lYfʷ�iߝ~�k����}�6z�{t����͞ �N�qC��:;1���ަ0��)�U���vi��C�s���W�C��e�C�t�4��zp�X�_��W�����|�C���Y�å��h,q�W>x����q�������Q���Q%|u� �� �!lg]���i:���x��0�2�p��Trchuy����^@�xiy�+�Aa�N��7���]@4F�&�e��Wl��ȶvu��4��J<�_�a�n���^����h�3� V�ɏ�0����f�N���;��iu�K;~���j�۱�
���	�p�9�����Ew�'11���>{�� ����Xi��n�^^���H��3�@� `���п�jYY(��A�tޠ�������S/�:c��a�l�z9�51��ǡ	���.�ɘ23��K��~�h����~<۹��c`��.-0�`�2B��Ť��M MH�c��2�동k=��y��4ع޻Q�S &&�0����f�~�Dp79y���b�2��L<~�/״���Wz\y�-VSYؓ p��y�5�m��(�uq���{��1��c�ɓ��Oԝ��CK� �4�q�j���Jt�ru��e��c�^�Ӗ��󅤋)�����iP�rp��������Ѱ��K��9��L�����l�J��,����@j�z؀�8��)�����:����P�@��Y��+�;���?��1�p�F_�ϟX����s������>s!;�K�.��?&F2[�i&%�,ߧ��AE�o��U���n'8���?.pr|��~��"�9������Be��t�0��Is��^-�����V�k��]�������~�2����ԗ�\���I�p��Ʋ���0�_g���)�t����N��SR��O�A�O���� �A�酵B)o�&	\��ᖨ�q���?CK)f �����}�Tz�������-wfm�J�ʯ��&T{Y3�E�\r����8[�O�����:L\�A��.�
2���N�;&�i�Ut�����s�e���K��C�
B	W����n���~��NM%�����Δ	[��]DG(9��(Hs0|��T��a>����{L�d���H�ю+�S���ʅ�'$X���P��k�ζ�iS6�huI9g�TݓKև�=�w��$�o����''� �;̽��������q������أ��}�GnȨ�D���Eϭ�z$�mv��C�C�e��a.���}�î�d�"��_:|�y�,4gZ�L�1ɺ�z7P,�eT�_��h�Y��;u=�A4u�U��A����8agF��!�@�� ~7[��k!߷Qg����÷�Da?)�%�UZ���=2X��=o�5�r�+�j3y����s�$Ʈ�}��������*9��2�p�[i����~m�(���n�g��Y��v����h�T�ɔibu�3�T=}�"�MZ�:-6m�_�>G����Ↄ1�C�����Wwt�I���i��f	F��P��8��7��!z�Q��Y䖫*K�_)��z�C�r�;j��v�-�%�%�XNi=�a�[����x��Dww�Ϛ�h����Jj���hQZ�;�|����ܭY��f�
=y�ne����ֽ���X&t������.���t�@ � ,�˂�s�}M8Y���!�� �2"��>���
]��b��@�16����iE���fO��Zz��61�Dg\F��,�N@� ��)舞J�����Mm�O}ɟ�C�`�}�!�7���5it �dC�lL�$�I�@0*`Z9��2��`�x���bM�=9��m��:��?���N�X��u����Q����;�#�ï[�~#Hqi�(�O��P�w���w�����"	���W8�@P�&�u�kg���J���;�z3����{'�&.�����zT^����l2�>M����!UG7>�o_�{��r�&w��/6Ey��~��<kB���׻�N�I�p���f
�&u������C�Ǧ�;����U�1�������iDJ$�w���v!sT;K�=Տ{r���Gj�{hN����q$���ͯ��X#)aG��Gy�^��	�4 �C�	�^�X�&1�O�֫����D)�Fg����S�L!G}���ϼ(nq9�2�tR�+��eF���#؉ey>�NR��g��?��tBy�L�}�Or�:\K��t&�,GY?M[q+1�R'S�Μ�4�G�oֶ`���3����|���d�H!E�BΛ	��.������W�ɪ���!}{q?ڃ{�fl�|�J΁���e�8�ސ��ìs}J_n��R��.���ι�7r/쮎}o���=���0��B4	�
κ��ez�Pބ�O+��MMf�һ����I��3��O6����L�?fn&�ٹ�I&�)�z����= �w;zm�)�'��'|�����\���~ݚ��������>�� �=����L�o��ę�r��{�#½�o�wm�?^���]�s-7��0�B�����$���\�D�O�c������&yG˓���43�6Fcq��dUK�:4����Z�X���(��A����wā���#H2��BLΔ� �u~� .N9w������o�^�u2i�x�5�5��w��<ay4�˳HI�/��y��X�׏�II�D,���Hė�>����S�����S�_䬺i_��'a�e׎3��f�֫G	�?Kо0l$�2�4��,���wItN��f��s]w�=ےqh����o��x�@�|Q2CX0��*o(��r_^Q��ֶ����2vf�=�6hu�B�M���U��;=���s���~	��z8�B��sJ��W��w�Db%�������{��2m�ݗK��w���R����&Q,����U�UL^|�Z�$�%���d�GҫwIC���.����~u=2jc-�e-�U"�mo���9����}?�Y5��8�K��~��b��(dk���#&؉�A2+��4�2��&�(p#�u���^b��}Vt=9�M�q;�u�����S4�9X���N�A�ӗ��(x,'�.��r�j���n�\��K�MI�T�W��2�����u��uP�l�����ّl	K���a҄X� Oc%%�Ж3���J�Sd����R��Yp0�0�tXF����0E�Z�T����� ���#-�B-F�܆�?�]�<�K����o�	�$-3</M�_�N�f̊��~�x��)�Q�En��k���?ĥ9�ZY����x����Ìi�{��d�W2O&E��_���'*�N�
6�+<�.R���S�^�G͊o&BT�7���3K�����ݍ�o�0~�0���Vd���48B�Df8����ƾ��Ѻ�ʑ|r~'�"Bm����wK�lN��b�-�37��:�������h:`h�t�2}���;��-�)
6}h5���LY�� ̓^Mj{����6}�:韬�sX��е���'�W�P�g
�l��LI��g"�P<A�9�a#�w�S|��1�H�8@_�����fP��qQB<��6��
��T��I�as��!S�����S#l��}�t������P�a�蔏���un�(-@��{XV�J�@="��u9�f��6]�8c�π�n�1mڒ����d]�^�h��c�M�֤�8�f y��} ��Q	���x�^�;۸���L��ܢ��:f�$/�駭��B��,��/!��g�cۓ7���:	�%~ �J�O?��������X�sG�</W��Š���f"�
�u�t�fC�s�������4�;tڇ	�c���;B�dF��3F��
s�U���o�KE}�|�	=��9�&�Hs��|�C)���	c��*�n^� �S�y6A��/$=�N�1&K��i0�h����ߩQ��L�\�%ޑ�I�u+'���U�U���/�A/3� :Z�AY#C�{��:M%�5�-�2���h`���B���fϩ,�f�K�� Dc���	W�@'B$7i���#�yDh��IoFb�&��_B�����4�� �#�\c�aA.�%��ھn޷��UjU	,C��^��=��EU�($bP��rq�℈�?���BT�Mm�)�Gj�d��z�㦨�OzG��|��U�}�т� �.����������wb���ٙC,ddD$�hQ���q#�� :�9�1=#�Ȑ�X��Ǵűo����B����v�X����S%S��!�g�VrLo9��/��:}s���~�<���j��h�`D=W�g�������|~\��<va���|?�=�ď��٬<
?�vJ���M�C�
%�� �T�h���>�7~�*�į����ȵ�H($�
�Zn���E��v��g[�?Ĥ:¥L{�Af�b%*�����3T������G�i
ߘ�jih���&��xY�O��fB�,	n*�×}��?��V��NeV̛ X�)�S�';*:�2<8B���:&5��їf+�N����=�V���2��/�)~Չo�u�&��N���v�y*�'����&����޽�\}��O��3�ןf]@��o�VA@�<P��]�:P��1W=���k
9�����5�o���~���b��J������qpW^�W����q3D��GX�a
���9����������d�o�S-|�>KU�@/�J�t���������x��
����shu��}�h���_�����|fv��o�M���I�>SD�K��/]�P|w��=�	7U�2��mv���٢�I�D~���z}��	����g̻�a�&zF�#u�F:��Ʀ�<CHJ�����m�{�|Э��Y�f10z��W+��C�]�Qz@R'a��]/	Q�O�����Gv�k�L~�x�Jn��ʻ�[��y���bI��H�lۗ�8)ώFnE�P�U�[cW��q�y�t��S��9�"�
|X��:[��J�������O�4���d�m�7�q\K�,"y�=�T��	C��'��c�J��ʕ$�&���į��#����1#X����p�E�.Mw].�K����1���	@���87�N�'Lw!6�ۀ�5���=�?D	��F�~�	ن�y���<9f[T�	1+�b+8�m�R�JO��Ũµ��Bgw��?�F*�.\��$�x_#���7��;Yn3�j'�����=]&϶��D��ID�x��>k�7�_c |af*PF!@7S�� @��o��]}i��f?�"x4�IwA7�{y���nwȆ�4�> �.Io�&�p���kަӢ�֌2VبXݘM����X qJ������Z��=1���q/g*0{YY����;��d<�/�����_R���*�[��Vݤ�*�ڜ�fS��O�ʲ1�)N�CɎ�'�������5�bc�s��ID�Ή	�N�u�\����7S�kM�"&\��2ԥ�^:�s��b�#�po"�V'-#������Xkz��^>������FR��Ν&��v� Ix7���^�Cf�� �H����|{�	�Ce2&�?��׵��l9�^"~��o7���C���/K��~O�w�&G/��qvm��(�&uv����7{��Y|3n<�#�Ɂ�Kl������v�X���(��{��!0�2qƪ��\�C��D	f�n��_4����Gx���^&���|"�V�-�N�����/1v}ŕ�����oӉk�]Z�4����_��t�}J&��MP�G�h�	�+��4O����Zy��m����[�^�RXi7kz9��\$v��V-�>�_������Λhp(��:;�{9q]sl��wy���x�	q}���EGA��+Sͫ͒D����A�Y��oG��G5T��E�]-��D�ep/CX�H�QY6��0�ة��hK$���J��N�Ã�C��k7���ON@���,2����l�r�����p-�'J�\���9�����a��e.
B5I���â�s����.*����=�K�?��4�f;�:�׀��B��B�aJ����1V�O�)��/�E��Fmcڟ��}��_��t�l�2��.����1��g������6R�������lN2,8�
�]�S�����S�}U�@X��Ɔ�Mve;��a�0
$��P)}��7#.�T��G\��lp]	>����%t.����V���΍%+[J� �D��h�li��z�X�� nw?�x@%�>JY�x��h�VP��l�Sw~Eji��u����|�M�6���j�^�n�JH�ؿ��dbMߋ�̬�����F��U�!�k\��O	˴�͌7T����r&�m10ͬ�:�j�����ז3fU��Ѳ��W����������E HRBt�U�(�}f!�JBN�,km΂L���HVӦxG 8t���h:�A� /ɒODO;���;�zo�;".�G�,W����%�D:�C1C�5Ŀ@������z)�Ɍ�#�2���OR*dҞ:����ıd�b����t�q���c�׏��q�s�{��RQ��+�ж�mi��s	�l!���UͿ�!�
���)�;�;��Y
c�)�PCp��N�G�_�E;Wh�̲e��	���̲f���56�eV%���e1�~숆�գ��[�+�������R��h��R'��F&��	�@��8�P�'H��E��KX��G"rr�[ZHK�G)�c6R2���=n:�HU�@6��{Q�f�aAb���<��װY�O�}Q6�w*���3��#�����I?I�f��>�%&>4��y� ���VrCｰZe�|x���'Wj��i�o8��e���V��2h}���=�)O�Qe�F2�!�45�L�4ՖuVj�a쫓ρ��j�+$���L�����BU�{�^���T�� :��vYI���
-str�gv�B{t,����kk3�hƃ/�I�'�_%߿��j�v�M 3�ѓOM��D�%�͸N�������z�MD��+���z�@�wL�5t2��_~�c�E�7��G>�w'*3\5�kImt��m���~Oq(^�˘��W¤�z��%7���C;�j����p���v��^N7	a�cz��u�o�j���'a�$��%�7����fQE	6c�c��|Π��|��&� LD\������Pu53asE���z�[_�&�W�@i��D�%���Q��kA�_�4m\��T E��3:���ÄGZ	�@E�YdF���-��>?s�Iz��b��m8�#C[�-�{�뢢!t��!���R����g�1�z��E\���Qly��1sF�;/
l2��g�(e����2`�����H�Bl/!� ��ޏ��ǘ����M�c,W�|��8d0+vP�]$B�v"��GO�����+E�a&$���ћ�P:�>K�P2kŖj��0ߘi������L��o��4�Y{y^t�<6:�V��\�{�}9I~@`��;5�W���o���j�9�ѩ�Q��t���]���k��ΐ�M�7�D�_8�<�C%�[<2��� q�J��ڂ'�B&܅1{�h�����pg�-�^�Z�����*bA�ʭ
#>���+��Bn��d�bksx��x�#}\֜q����|m~�:��'U���A�V-���8=�P*���]	��Є{��9p��Ɵ\�m�ی����o����|{x�[�h����k:�h�f6�>߂����j����<�'�(k�p4��V�I+�$���L��K�5ʿ	��J��l4���t:e��<�9�PU6D\�j��m?[nNp��)�7��.��쑙Q ��uA0��H�Lm��P�ݰ`�1�ixʧS���\a�Y� �~����i����.������|�ɜ��V� �tJvLv=rq�EZ�0+�R�b�nE�G��S+o�V��)-��жx'W~�>3�_[�x�����}�}�z~�ʃ�cQ�C¤��-	 �"$��"��5h���K����g�k�e�$Cjk*�XE}�>�~����וVBVk��'UR>�S����r6����8u3�p���FM}�ԟd���d�n�m?vR�ܼ;�?�~!�l�9�������Ti$�	�vp�}�����>�CөP`�^��,��]�&=5h~�O�{G�O����[�$�G�r������:7Rv�����IF^���9%�L�;���l���&�z�0,�Y��-S:�$���f�	9�)X����8_������O����9�O�k�塩\S�m���B�+X�9�ylI0k�����C�1{�^�� ���-4�8[��8�5N���I^J6sA����ʦ����j�QY������硖�k���M�(���_/uu$#]@�>�$�!�!����Ea��=����fw�>H3�94�Q�]!g3v6*݊4������ǥ)����t��T�_�P���6��~�a.���7",�U�K:�|/���βڶ��]�y�}*�?P��*�~_1�y�.�<���%�L=�-���X���>Ҷ��*M=9��P��od����ck%��x}�ȒMP�I�]	��1mS5�Ҧڝ5O�`L�@卬F�
�%�����7+Pۣk��I��,�G{4BI�0�1�֍�.�K��~��h0�4�E���;˺�~�{����,S�Ѵ��i��=���.%��o�˹�A 6��Z펩��Í�ݿ[�q���9�$M��<q侺ň�����+���������=ʐz~Ffu�X�|�?��}o��K�!p0���ur���8�lD��g�T�>�P7�����a�"3d�3{�
g�������J��%�����|�_#��N������f�j�TO��9=+qT�6�#�L��vf?Rk��|��g���qm������O{�֦<���K�ڝ�E������(u��տd�!�ӗ�A�vi�d݇����f���i7��тG��C���eCX0�h݀��A����'^X����'\�eP+�θz��J��A7�K� u����S~�Z4)��p�W6 �����$�+p�c����`&X��8Q�p��w����Ϸ䠊9�6���A�H�ӗ�u�pV���*}���F���x'�ssd�����1c���{�L�z��R"��o?E}pA����򩓲��Cʜ7���*G_���cv��U%[:٣����|��&��y�|����C�w��fv~]��__�F7H0���$��p<^$��E[BM8�NEG^&�ht.�C$�Q���l�uo�޺��`�4iM�w�q�j���cN9w�5u<ǹd'Y:��n�����.�m~�}S�֥���������x5S�-K��y�����5]G�_�R�-��x`P�8�v�(O�>�n�ݣ,T�XQ����w��������� yR"Y�#l5��`_��ݍغ�G!��f߅�jV��+�����ƴЅ�����
����=��޸ �*
Rj:m�z��>�XS���=:��uy��}F (@�ɽ �X}���p�&Ϩ-��a~'��J�'�:�\}NP�U�&ֽ�m6�n9B�����Z��+�V�[�=���:&���H����ʄ����wR--VX'����kT�g/S��*9 ��T�x�r�L�����J����#v�j15l��H��`����07��gQ-!���@}U��#ƽdL�6Ά��
Ȇ5��?�k�2C�r\`q՗]��b�w���t���yb�h�&`�!�+��k0x�í�ϛ���J�{[K�x�(u�J�Q���j�8q��j��@]"���z�8e�i!�#�Y�Y�1[C�u(��| WuFR��}�S�-�ƹ�0���Q���.�6wm[w$��Z��C7FMЙ���o���ZTnSfv�-a��i\7�φ��_�v��i�u,�eV�;�'ᶔ��B�	��s�a��5g����'|����%���2��\1v�Xk��_G��!��a��H�`����*�41`�~�u���cɈ��t<�	�b����a���0�$��e'1ί���e��c���
���fjg�*�c-z���m���ٚ�����a�fV��ߏ埞�7��-�cfN ���ˊ
��C�+��a��Ѧ��#���a:=i���ݦ]�W�ú�{K6����*�%��d���.�7�y3����-�ʸ����G*��N�Ѳ^�����}L�[��
H�9e���"#Z<��
�F9�6�T�B�ix��P�_�3�̪���W�f1[(��O�|�S����|=�$���b��X��٠�f���:{��J�p��j~��,��-ST�z
=C���+��}�?����X��-�H�k�~�}��XD:I��
�q�h��Dj9�+#D��Z83��På��{��K�?@݂�uq���Tȟ<���J9�!l��|�3#́T�T N_����"�4?���i������0���`����1�n�=�����r�(j�!H^�wp�e�<���\����haBxPXFiY%�Sgd�����f�*�ZH��ɩ2����tƩ�*�(RU+q�h��z��h��/�)ݳ�P�c�SPs�H6���i31�~42�x�Of��l\,���\���x}Y��>9=q�ґS��U�.����<jK�l���l1�#�������m̲�����X��u��Ē�)'�Y��G��}�e�����ū�b�3���n��o�\�G�wį�/m^��P0n�ө\��r�(/~�=4,��.�姚�LCn7AHB�٫~�#�y��cl�qt�*����ApCZS��.fe�s�6������{��BO�<ae:6텖S��:��N��.�Z:0�ͣ������o�(O�����'��f�y"��8���M��q�U�<X�^���>�!R��q��<������z�V�2"���s0�_�5E�HJ��ʿ���P�,5O�!��1��X��7Fq��̔$��j3��w� ���k��[
7��<�E�Ӣ��~��x�B
j�y�I�.yIl��}�-ɌNR�?�$�
�����&LC�DfP��R��J���݆�׈O���Ά��/���,[k�R�yEaQ����3[Ҕ�ڪ�B�l%n�k���@�K��fT�
��ٗ5G,H�ߴ�6r4�id�LB�O�[�j.��e>��f{ġ���@�Ñ$����'���䱳�yl�sZY5��s���5����k���7{� �c�Dqn�C'�q���Љ��S+)1�I&�4W����+u�8D���w�ʴ�s4�Dse���;tQω�{!H��$�����n��P\��n�y�m?���Z.�
5���%���+������/�"Q����K�K';�0+�O_���fpm�ֶ蚾C[%X�Fǳ�	��k��p��/ 5���Ge�K�;\�R�+��2)Ʌb�S��&�kS��R��%>Y�'�M������"��gֲ�����j,���<�K�p���Lz?���(�h���p��X���[zeON��B���J���qSZ%�;/SSr�A��RO�>�g%*V�9K!�����,�M���F�� �ね���ѱ০8��r��wa��'g'���km����G\�Z�Y3:��#�Mp��I��)V�f�֨���ˏ6�z�<#Y+�3�=Z U��Wں��-2⺃��>Ur��|֩^n��n'�Io��D%	Nvr���f2᪣�L�!JÞ���7����[����̖�����SL��tGy��i~�Et��TB6��O�Bz�-V*�A��o�Nb#W��J�,�W;�EZ�h�~-��:��
�H9��i|�
��󝾶Lw(a�x��ZG�(.��<� _�;dּ�5<�?C6���[�D~p��ep"P���4\a<�|�E4��CLT�Gz���P����6~)5�^R��4+�{Oc�m!��U@��s��~#���Ygw�Q:{ԄDA�Hǔj��`�l���m�z�T���^������(��y��yo9(^<iJؠ�X�D�H��~3{�Ze�hz�A/��ܬ&�L� �q�} �#j���U�ea����m�~c��J���l�
�R��3U{��a@ej������7��U����~kz�j���vi��&�h胃F��%=��o�ETYB��&F��l.<?�-I3�t�'aV�D�^�$�~ř����闧U�p�$�d}!q>ah�Ă��~t0�jn����#��)��Uqs���B�����	RH�	Z [��������U�;Lq�t#�*��9�#gCp�mX�B��bj�U4��ݏgY��,�}PZ+���OZ�YMh�l�dH���c1�]�tP-����
�jQ JAq8��|��Ҡzc�Gh#��p|����2�b���QI��H���;
W����	[�e���ALK-є��|�L8Aqrp��s岎z�B��5�Q��0�b·��5�X�H��w�~f� �i�p�Y�~�.ஊEH�4�/}�J�hu�[��1��k/o��|�ߊ�d�cf�AcpWq�M��oJJH���t~u(]�ݚ��F:VV����GL����4��f��'�������G(=Wa��?��)7���`{��P��s5b@ɠ�4	�03��+�߁�pߔWH��^�M%A$^9�>�L�o�NEt8A+�=�?1M�}a���V����ϥ���l�'@a�dI#����h!�H?�M�i��Y��Q�m�y��Sx�%պߙ�!�G��0m���ɓ(�B�n:#	ڹG��$γ q+�x�Ɋ[dO
�)�@y�>yS�-8.:�=�W4�k>�f&NWtO`�^�57H6f25E���vi��4���W��Th��� ���eۣ�ub��h��U�7V�7j��kc�{u��M^Ou����p��}�S�t��KSf�`+�5K�F0��G�-��ݴ%q����2�P��I�D�����-��?�i�j��"�lqln/aQr��[���]�d�XL�B�O�H�F��ڽ�ϣI~�<�H�8�q�9w����-pcRފo�5W�����6����y�_������yhiu/�pS�(WQ!�O��hn�@���r�|�U�Vfٛ��!�㵪�R�+_���6E�f"8�i�)bR�w�p��X�rҹ4�؋�t�vDU}����ΆCo��#���X:#9�.�%��7!��W�d�q�Y�5v[&!�/6�a���&�}Me���5��\�a�$�K3�=�Z��K�y|	�x)v��3h
I�k�8[���CY�9�"-��b��ʲ�8�!�[�ed�Ρ?[��m�gAX��Q_2!�2]+�*�^���_61��ΐ����F���c]׽�J0��;ad��n��|43X�����?g�/r��h�?I�tf���X�f��N7�i���:4�շ���T9�Tɝ�l	�%��5�J�@ա2Yg�t�<ԕL��KO��W��|І"Q��[97�b�;V��K��F�]���}9~��-�
E�AЅ8���e`���5�K�5T�-�J
�� ]��wE���d'�X��Y�{L�Ͻ�/��pd��Х7��ofM�$��n7�n��ƒ�P���z���6kjMx�>!�O��G����D�����do�� �����}v�zﺩᩋ	���=�05s�T8��x���T%`������f�P�F���1���i%�˥�9�`\�&�����Y�s����S�l���k�t�����|rZ����$7���"���C ��	�]ωs+5Nf����0�?t�k:�V�@j5��泥������hƄ��m�"ywc������N+�wa�,��6�9c�%��J�Q ��qx�e	�;x5��������HB�	���$��#*����v�յ�?9"M(��DV~��Z������N�^|�k�S�B���Ch�0�'�	����ŕn�dc|��`@����=���p�NkWm���F+ox�l���@����U=�}�Q�7�I<�`2��� ΑI�R�e���L�J���gA�^��-�ˆ4n��O)@Y.���߹�*���?nnl.���,?w{�e9xn�c�#�g2!�����ԇ�p����� ���֊g�n6jg�ݤ�D��w�k����<B�n�w��ۣb�=��K����O^X���+�.�L͗SOYf�j) �"(�����3��_����L>t��aݭ@����_��X��?�Vv��Y� �\r�B=��u��7+_a�\6�Z����oy�{߫��I�r�����{�<��	A^h�ha��,9Nλ�U��̳����m��fx�^].�`kq�{��y�{6��	���4�!��`��nيSe剧� ����|ꩧ�� ��yh����Zy��U�c2���7�?�,Y�D�z��������؈�E���}W�k��rQ�Ni�\���0����faiٿ�[3xӞm<W����v�1Md�̦$b��6Ԧ @������ܢ{d��sn��`�{3���fdS���s�|<�	�,���eB���mA�&)�x.6*aͨh�����Z���7�n	c
@םq��N*��e��?��I������#��r���m��B%��B���=�a^LJ�l �!����ݽ]
���B\�L�=���fM��j�a�[&˫/�B^{����PA��)�����G��C�ۨO��c��>�6���+L�I'��e���Ym���������a޹���y�0  pL&�(�ʠ0���c��]��ʕ��l�/Z�$�d���+�/��dD.�u{�r��%=��q�O��g�cNF���C悈�2��m���0.S�k�<��s+M�j���)`�`�N2V�"�9Y�Ƶ&Ș]0�7������6�8�E�(x�
�;��m��� �� �XS������/lIg��m���e}gW�(J-f�H�`�H�b��@�iZZ͝�/�5����>�Y�H�U�fLozӛ�G?����|\(8�:H��A�� 
a�1΁�q����{�9���uP�9|ͱ�&n3�!���VѶp,�t��Y|��CK�a����I���h#�YP+�y�+����ʍ���ovъ7�&Յp�={�Q�^�8�S
}�R�`q[�V[�y� �nb�?@��o���<�DW�[锉u��D+�� �mj�Ԩ)Ad�\ 2K�K!�j�Ԩ�ٓ�������S��B���jx>�R�pKoP����s][n����砐!S���r��D%��Z&ǘc;�)hf'�E%�S�;+0"���9���)Ӎ��Sk9�N)�ӎ[_c>3 �$��U�Vi�}��>4z0v|��|@���AK��xZ�ZV¬'Xp��M$��Z����Wf�c�!4�
���`�3�`��orB���I� C kD��=��D�Z]0�0AH�:��4%E��9��&S���q�>���Ae��4Z�ʲ����{��[�Fv��l62�X�ڪڭ��S��؅3�5�	�^1�`Xd�7k��[���1���9q���q�ݾ
��ϸ �}n�}U�c���?X}�|l`ι+�"�u�jSxP萑��\�����cxM*9n\�֔ƋB�D���*�V�}�>G���(u��.>$UyAY3߳f��x�L��@�(iM�V�y��k���Jv��M��.�}�z�ɚ�w/��:a�����^˶`�c}2>B%�c��H�A�������<hR�YK���Cca�F���# Ԣ�_e ��&:M^jVdH�	]F�����'�9�	�&7L=������L�Z�ٔ�4�8���2y��j,�}{wjuC<������c�\Ư��76��zfI�C�ɝ��(�x97�;6���q��Ժ����2p������$L�q��]?�мO��.�A���i�3��j�T�sq� 7��bl���3�q�C����z�TɨR0x��n@V�&ok����3g��!FѪX�3\: d�gRz���ף��F�fQ	����Ý��|Í�p쨔a����G`n�t���o� �7T.�4ak���ΑF��e5@�'��H0X,$�KޠT.EL<ה�����ӛYtA�ܰ*� � ��P�Z�|h2�Ajl�ri�R��Ak��1Q�@��}�?]#��
�4�kt��*8��s5�cw�i����� ������OF�Vo�68:��}��Q%V��;wFnBׂ��B�G�w�n �V�{b����.��2=� \�َ߃\��gD	�p=h�(3 !F��Z0xKbk� �lT�G�؏�DH2/�����*3�Y�ZdAֱ�����ڗ��S�k�PR%ݳRƒ���c�*@��芳�����z�5:�pc�0���G,�`����	�*�q�tsj6oh�R����M�h��z47DD��0Ml�FZ�į� D���8��R��@.�!���q=�H͎.�Lʞ��&C��v,۰)ߨ\�ճ�`��i��/2�t�X&<����oW�4炕S]�>��=�c7�t�n>7�]����;2N0�~UPD���
��Z�h�1F�}�_q����~��������8'��abS��x�-��d<\fH0��,@�0���	����������߯y�k���>C�_���� � 0@�l��Z/A��6��BU�޾^�_ 6
����V��,4�?~��(yYM��֏����
E9w��7ܠ�?ʺCQ���
~���댖�Zfx��s�X��`L`���q�����f��v����L��f
_A��R��B��G퐈�������Zh��k�>{����]��ɧVK�*}���Z�@�YlQ�ޫ�G�;�O"+-��.4-)��) Z�T@W��v�8�Mr�>��`=@��&eB	���q�\��K�.�x7(��+�g���!M����`�{隵�ۼy�BfP���KK��up,�{�'��\ (`�x�5e�b��!��KZT�:��"����F��{����u��S�į�_��g�2�W���rkn�"�g̷E���ݣgq������ *JVٲ�����B�yC)g�E8�T�xp��+�d�a׭��v��B��1*M �����#�礹Z�;q 2w�(�M��Z��+�B�ߥ~!��ν��COjUO�=��%��G�n]���f�$5Ϗ�:�7k�'�#�%������_Z�{��H����6͋[eQk����܋-��$޿�����w߭��:9������&����`ʌS0���Ƞ/��zX8�t� ��f�ƅ@n^������,�×���~���Gq,�����gsv��p<~ñ� �|�I٢�O3v��B��(@�U�u��SOJ�-Z�y��ǩ+4O�e�&��0 o�O����[��`�"7�H�����q�� ���`��S
�M�Av5|��r%u܅� #�@�Ƥ�ZRm��=��<���mL�Nm6�|����n��֐�^2�-���������� ���F�]�IYa��H.0B��B7m,%-�e6=��BW@b79j-6�4��z}�[%�;4�@�k~������� � ���C�	\�0?���� ���r���eP��Q?� 7�k�cG��!�tAo��袱L�U��k|�\U$��2o�+�j�{�N�/�F���	_���%t�Kk	h�����0��ZP�h�q�k�`b"������Bak��?��gRҹq!3�B���es��@n"�L��Ԉ�v�b��ohz����ק@�����\��B���6��w�N��]Q]=V`�B�n����_ށcC��9� ���h���
 �#H���g~�_����0��`&8�����Dt��."ąC2�ߏ�i�L}7�׍Q�� ��pqshE0Ǆ�D�ؖ��h}�0O�/QP�s��5�ǔn�1�u(��^`��5Np�:N��3Q �|}�b�� ǂ�(c@&<��ts<��606��/Aᅟ���TF9wno�C�	����΀�3qӻAN,.|�=>mdsp��:l���.�:V����W얖f�,GG��� �y
}eim�&۷�UV�Ug��:�4�7�X&b�� �(�_{0&OA@���,��l���Q�%��5]j�86;|��3�b��,>�8�b�q-�tuv�0b�<|��l:Zp���5>��I���q< ��d�8����?�=��83�)p4���\�ŭT�ZXcO������9{Y�v=���B9�bE]�%-����C�K_��&��Q����z�9@�C_|����q��P�y�_��7���+����omrq� 6}�4��F.$���k��(���M��f����Ѓ!U�[�R�5&j�4�=X2]ʅ�m�e���Z�X��*�Mii$��w!c���3�ʶ�.���w�[�����I.y�7F�}��`�6���\p��Ua�a��
��[�S&������`� O?1�y�d�T�������k}�k�q�x@�L���7D���Xo�jH� ��J�lI��1
$�V��gl �#Z�`�e,�*af}oݺMv��"�]����݃]M�R���e
J�) "���泮C?���T{���\��J�Pֿ���u��O�r����:��?����#C���T~�\<.' ���+������E�z(��ڵO�=��J��\�Y�[���
T�D�K��֠�. ]L��,uiycMsHd��w�� ���|�)2�?h���oFv	�
����;������#D�v�✘&�����*�87�F���:��lὕ����c�7�	��V!MW_}�Z@���q#c���z�*���O�T�&ċ�̃���@ny�������2�I������c��@c?[��{�V�\�x�\|�%�kj�b����Ui��|�H�P�����B?U�NGx���=��c*�+7��E�h���Z�J���*���\S-����~�'���#��-�j���6Lm�I\<�\��bc�*	Q��N^5��Æ-Is>-My�8У�/� �V�`���m���O���>�}AK��A�:܅ձ����/��PD;L���,Y�9���
,;�5`l4�/���'�|R��c�6���~����y�E�
w\��eR�V���$��K$O�m�����b��\Q��н�w�Cq�����d\L�" =�� �YXXn�9 ��3�0��k����.����|�[���Q������/̾��%G��_)�TE B�GU�T�E:���}�,Eb�=,��P{8�󬲩��la78�Y��M֢�2���������9V˼c�����C<(�^\�%f��N�+t(�2���ɠ���'/��n��C#hmn��^q��^li�k�n)4o�0P<�}�4����Ȏ۴�+�}%�fWC<��(��ۆ�]�2e_q^%b$�p���!�l�fq��$����+��@Ҿ�V�,i�(�b�����j�Ę��4��e�Wv#J�>�'Y� D_4QR`~``�`R[��8n�����׍��w6�p0OM�:��A��q5z� 6e.�U�,m����_�B	��Gg6�j6o�$�=�Z�Ο#���&2}�4Y�dQ�L?%��T��L�h j瀝~�{ߋ~�~�!��@/������#Z�T\p�w����)p\���I^6cW������^�sF;���(H���=��@Qjn�*�Y.��1�A����\�W��@AT ��c2�xr�)��+�kk�Ұ.1��vݻX3hԂns���u���e,�>���eR��C�\�Z]WPf�e3[m�\J�+��P�y�3���>ʲk�G��k��FN;����rQ��:tĚ>}�E\��`B_w�uZ��6�x �IiYpBt�d�1���k}�|��u1V�}�g2ZO�%b�� #�����;8��e��k��$�*d� l2�M��%�nj�����K�:JD��&r���w,Ǎ�!��H����(p�(�+������[*J�P��x�jts@ns<#��<�PD����V	�נ["���-�� ���};d�]j�s6�f	޳��y�	ZP�J���E(8� %��#d�z��}l)��ZO�ׁ9����#����R���׀򁜌׾�r��F��۩ �fË�v���5�'g�q��6�w���$�,��Ϳ.��g��d�Ye��^q��r���F[��"۷o���{��Ӻ�ʁv�9��Ur��ʹ|����>�#��b�]�9>Wl�!�/#ӧ��Ν�d���֔kֆ�U�Zj)ؚ'E���i2�Qb�fj�����H��"p\+����S�fi����X\+�����x��P
���j��j����V���g���XC
V5o֕"���	"���ȃ+}��``��`~Gȧk}��4�9V����B��92T�tQ�X�:��/L�4n乂����VY|�rm�R�x�W�\�I���S5��dI7K���h������_��_���B����&�ʤߞ�EZiHXl��񤣳W�|�qy�чuMa.Qtn���SVi>;���<���Rr�D�b��{�?���̀	[�p��y�*-�Ma��r�}��R� K�_�Z@�`�c`����m�������vO �#,5Lm�f=�7����yg�M2w�B�>m���K��κ��ul]r��À�ϩ�9�?�I�]�>lb�3w�2a$��Dl����1��A7���k-���R��V?��ƅ��!_C��HVz�pu\���� �u�� (�6N�r7�}���h�=��w�c=:�>6n�[9�*���g�]��D�j��=e��*֌��ڦʱ�N5V�d����J;kR�γ��E���S�yGa@X���1�p��1c��-�o�p1G�c��Ռ���J�7��=&;w�0����m�7���O?a��.9�3����SČ`Yt�t`�;���h[�dB��x�J�	�	�g�9�x꼱
:�&�+�}�fО1��+{�w�r�u��	?�St1���2W�[���Ѩ��|�fvw�����d��=�չG{���,r4}�ثha�r��c��m�c�	ƅ&:�h0����5p��D0����̰9Yր��A."��&�t3��Aӊ�@�B��tx0��	 ^�&�L
�=Ρn?Ϗ����ʡ�?�!f{��E�!KL@`�
�O�����H#h��$Jh(ˉ��D3
Z���Ǟ���}.��1��P֘@���f�L6L�j�)����K�h)���z��%��,�[�����1A�Cq<}�c�X���Y��D�pЧ7(w˾����m�Q�ɓ��W6��QZ2���+=����+.����Y�Dݍ��)�!.���'jIg뭫C�M�F�L: l�s�����)��z�̝�n&�7Z��P�����}���
�Ǥ��؄��N�5�&tr��sf1���H���0�L�f�I/V ��u� ��0=TJD�K�KA������e�����S2�K�/� ����7���������N8A��N���ʏ�# ������=�I�e�9I��C����o~3��Z|X�lr������k����w�|��%�i�����uP@Q,��}-�u���J�{�U� x=�����X�F(V+���f�K-�ַ�U_�������{J
�����Z���:�%e��������M4_~oo�TM���^������[.X,��:S�S((�z���@�Ρиg�A�HPH\�S�LW�	S)϶jKy%�:��h�6�J�5��.D�{dR�$ٵ��M���Z%69zw��t�x��~�^�E����NYֲ��im�I.m��r���E�R)!���o#��Z! �XOl6�Q�o�� >C\4�0@�.�G�+��:0Y h���+TS���������|�Ҙ6�]���2�pʤ�
�۷�h�}e�+�����w�B����5�gd)
�qpO`T \�)��������5F�s�O�	0B������
��A�J����j��]pġ���d�_��v�/�˥�2o�!�cm��P4?�s`�̜�D�F�+�i�T���s���SU�?.�7˖/���g�8m�Ƿ��-:�_��Wt�1Gl��?�vwȚ'�ŋ�Ȭ��e�_�4���^�3�=�roi��Ï<(�/]a�grdMn޼�Go�3͢��2P��ф3ƎZ��93�6��l�~�L�fi�e5��VnՒE�Ф#���7��C��\D�?�zܐk-mi���'�o�M�ךg(X �{��- �?c�\'1���h7!���nA5$>Aಅ#}���c������������$8�52W\��MX�((x#@��+��2�� 0Pi��#-���&����wn� �k��q����_/pK��ѳ�>��G�"�@�k%!��6r��D:�@J"�@a�u���%+��_���eS����e��Ge�	�$�d�~�(�j�%~�C!¼3~��}׮
���AX������K��	�פ�:��;�aƻ��ת������̄�
%��n6s>$
�:�q0~�q��=p��A�ɕ�If�E��[�[��,��#BX��Q}���m��_�����;�!g��)���m�ҴԴ�=#T����O�T4,�(�,��%}蔟Ua�����C��J��)*:�p(n������}6wN�4vb��2x���، ��]�	�bW��0��i��������<t���w��C����Ѳ�𾨀pL�}���;��#�{�6D.�����8�pq���RPQ���g�\7���<����p2T#�3�M�6���}u�jv���X�3��N�9k��q����[Rf���=���c�v��U]�{h��Gy$Z[ �0���]�7�e�+����	q,V�| N��b��?�y]������Z�{���}��0���o1������f5�b��S9�M[,9
Be��S�<����� �!͙��f�h�A�*�XHnh
�|.�Bɨܶm՘�״��V|iknU���#!�h��Y��|S����3���G�K%V�g�?d.�r|>��*�4�[4�-pr5f�,1=O&��{@.�хK�̏�w�%�(-���Hp��ܠ,����0��ɀ�c�2l�QQ�x�i�1�D.ѺaN��=����C#�K����@ �4N�ux2Z�1�^��a�a_@1*h�W6g��t^�����+�j6����X`�yͫ��y��A���,�����
���w��	�
����
�2u�qъ�eZ�Q���Y�ip9�I+��9s��!<�2�u�憛��?1��PD7 &�����6���=Ř�U��U4@5%��)��}$PuHW_��Ɛ��877]�(I�m5�!x-$
�ǲ�O|���1Y��t����b�5�͒�޽)�z�t#Д�2�`���M.�����9�x�.��ޣ�&q3MyW�e��������Em��Bf��� *�-��
>gv���;&�1a�P@���ǭ��<�D����/>���?W耈v"S#�g���
5�1�C94���*a�J���߾T��7J��Հn�Q�̝ky�����29mʲn��޿�Eo�EF!	�f�z���h�Y�e]��.C�M�k>���=�ܣ�/�ti	`<�Z'ˌYs/i��gsm��t�î����Im�F �x��3T �,��6�����z��?���v����}{�q�d�tvwȹ�](k_xFt���KS�h�d]f�m�$9jANҹ=2g^��d��ps�Իꪫ���D �����N����(&p<nb��&�M�����}��K�Lj��+����V/�@$bf����"�m�X�~4�u�nj�.4�ڸ���.��L.�P]+­�J���&�1^� �fܺ��5;W��o���� �����(���$өU7&�rqc�u9NC) |>�y\F��	��0Ǆ��Ұc^��B���R���9�|Æ��q`�с���d��^[�Y��ß� �$�L�9��0!�hˈ��4)�w�F�v�ؿ���kUY�AY�9>�' �~��� . ���K˖� [�m��[v(P��y��PpSk��O�5O����j��=,��>'�]���R��~0A�>���<����<��cr��UƼ�&}=�̝�H6o�&���/�*2�\�Yc�Z�ȢE��Y�\����{�N,��/~13�.��ԟl
bLH���vh@��~.:5+添d�ֵB�O�u�����tQ�j!�]MS���tv�� ���ʨ�[��M�'s��7�C�k���A.f�ǻ�DfF�h�E�Z_�8�v���d�|>���j����
@WP��Mܪ�'�I���q��߱E�`;�]��q�R�G�%�g�[!�E*���3{��s�z��^:s)�?��ޒ���<u�t	�e��
��ɀ��Lׅ�Ak,��)Dρ����>��ʧ>�)��~����H�s݊ p}�֚�|�lE�tv�ɶ[e���77	�VI{n4�Q���'���3t��ث(���r��R��_S�!.@�M�[o�뮽Fʥ@��Y �k!V�?��J\$U͘1K��XN9m�6�����[�zu���O�G`����Gsh	`��>�� ��!& �VS{��r�@�y���ӹ_U�\�G�v�����d�
4��2|�h�hM��ۀd0��.�k� 2
��e$W@���x\���s�)��!ƙ5\
W�P�PP��w@�_�}��u�D�w�X^�.)

�q�;D(�-�x�P�k��;}���U���:�@72�0g�8��W(<𗷷O�Y��j= �����E�Sr�+��+�`&�X3��в6Ϭ�q##w��._�ׯ�1�5�\�l߾�X�}�}��������z�{߫�$���]:�)|���_����2c�\��.Es�<����#΀�����rs_S���+*��*R�DP=���o�3���!�U=Sv�L
�&!C���.��~_xѥ�?{oe�Y��>{�]c�IwzHw愐�aPX��̹�8� 
.��\NG�\t)2xQ��W�H!!�$9@�H��t:���w՞��{����U{铳���*յ�7��3��ɮ|���A��� ��l� )����[�����1 �!���x��b��w��k<��M7ڵ�^�X �!�.��m=��-��up�+;�R8;&���%l��Ш�w�;x���-��m�52���aOeSfIZ
�Єc�^�ȩ�6ŋELD�DL�	��]�G�2AYeo��@�*u�T���!b�F���k��*Z�&5�Q(c��)s���i�e3�B*u����F��Ԥ��9�R��Ɲ2���'ռRf�k�~r-��2?�f������v�s.�|;c^Fs��9J���9i:�j��y^��C���G��7�ךA��מ�y%�s�yf���J��9��V��V�c繶�����x��h1oذ��M@�*A��_� ��mp�$�~�sx��\?�?kn\)U\�'������>�r���V�6�\u��$�YPD�	A�B���W9ae�4�O|�U��^�:_L�߳I�� K��ˎ��O�Uw�Z �� ���čMQ
l F�{[>��NMuY�)m����("�
����~"��k��Y���MoT-�)������W�kP�y�G��|�jhb\O��y��R�M~�7�c=T25Ʋod��
�@(�c(�bl<���I���¡�Oe`�!a� �&��0~1.�Ȼ� �^x��)�)�nP�}�	s���'1<1/�m�w+�5�)H4_�#�d
�;��(_�y!g��@���wx��pN�A�λ��]av�����	�2�hS��iw	x+���,�76�s�O�B��u��(M�g�p?4a!H�W\�_G��6m,۶�[�λ��3�mb���pѿ���v�|�8�,*��}���
��b��O�?����ߞv�Ev�3��o���i �$p#M�N>S�3bʂy����ӟ��8t�v���O��o��661ލ��s�p]\���z�T�{eh�U���n��׵��J��C����an1��.�A��.˒b=E�������!'B������pec���k^�':hD����P�5�%�=ER .��'�t!|��_��\�/|�δ�u�J =/{@8�t nDm8��Ĉ�׿�-�})���H��`116���B.?)�?��Ow�������b����"��\!"������'?��o}kW�L5+�M���LEH2�d^ٷ�SjӀ��¼0.��QB}���|����Ks�&��<�&�Q�{�~{��;7�fZQvdHs^g���N��K�p�g'�F)H�Յ�Y8#�S ��d����ǆ�ne��h�n �L��?�|�㡞�x�A0_���&��0¼G���ёh����u_�[o��g�$ʜt-�������������:D��<�h�>_Z������i�س�������wo���ZR�zh���V�~a�F��DȦ�T��ɒ��*t�<]h�v�i�>j{�;<;�\` ��o6�G��=�K��@t�Z��7�Ϋ^�*�w���*�A�%*VyOȑ�F�Ď�Di�H&���qe�� e��3�xS���D8D���!��nਬixaF)E�*ڗ{!���Y�� �C��<�@�#y����(�����B��W�W6\){?�a0A$<${"��#80؊~���=E�A�T?��O�{��^+^bh4�94	4��%�u����&�>�\�T��h�t\C�*����&AP&�ά�C�e>髊�@�`����s��΀�?5d����<}�ޙ[�瓋i�����?������v�3.�y��.4�hƌ���Z��f�_tG�۲�ϱw؇w�xR>��}�s͓���P�%�{�� �� ��D���N�CoP��Nx���uVe��$jB5�i^uhI�i����\��o~�C�!<"F��H�z���F�պ�a(�i���6?;e����>RN�P�s��	�-d?�������AܐH���7T#��T`	6>Ă�90�*ϒ������U$Z�	� ����1�)�"���4���B��Y9�"�����
Q�@s?��ϐ�d���B��{�~q�G?�Qυ�Drg��P�����{��!�H��)��!
��9��ClIj�X�]���ų��r�i�ar�9a�`�h*F������u��z��_�-	��2Ϭ�`42�0P�
q���_�����m�Ͽ��?��cR��kVwn"X�f��:�<�X�AVd��\J�� �V�y�~T���ce]�3�XWi�eQ�W='�j4f՛��꙱9���A��d�	O�����R��O\������K��n�9�HNJ6
B�懀�i{SW����������o8����ol
�8
�d8\��9x�"�mi�����7�CL!(%>��!=��#M�BAuVrۈ(wp/s1�:$q"D)�5�ZE�
��D��k<�k���@���* v܏���X_K���a�1	P�;c�Y8@�t�y/����ғ�E�Y5�-�*/2��nC�@�PY2�DK���Nt��%��w40�>c�Bg.y'��0�Y��~�E�+h|��4h^�	L����ݚ=�c i�B��ǟ9r��*�! a���:�C�AY�琺^�h1�s��w��?�A"~�7~�mx0`L��%�F�)�UB{\�����#f����M��'��N�6��I���I�"�r��>O��xD"/I���&U�������~[D�JQ�,�!�mE��J�ǉ|!@v�j���SL�u�!v"�����|�c�C���5%oh�$�8�X�9��Op,��1�*��sH�Ż ���x����,�i]Fb�R5�hD����^������@Ӑ�esк�/��E����|(�KP!��Ar�鏘&���i��^�W~Z�]9�i���
�VQxDI�k��\�c�b��aj�����p=�DJ��h�p%�;��jt��Ԗ��,��)���t"��V7�R��4Qf[*G!�!g�����<���c�a�s�s����5ߩ`#�I��ƽ���L����	O�����_�Q��æ����}`%?�^UL���>Tw�y��*؛^����R沴EO��/mz�p���ik�w\+��7iK����6�s!����Hlh2��2x'x4� |b��$m��8��Gʂ�+H�Z{f��:�`���,-�#y��� ��Wy�@�U�F�T9�0�a�r�4��B�=�R3�m��N0U�15*s/����+*M��҄�H�Q0ϡ��1m��	舾2F�B"%��&,�Q��#/zFz�41d���\l'$G+I]P%�����t�]�fUA`��|م1�O깕/�܈KQ�V�a�SGm<�{ͺӲ~������u�7��.ɽ���ޑ&�%��`��~�<	�Cc�ӂ>��M	�FZ�[�Q*,�?�'in������{��S�L�Üb��Z�Z�Y����\�����,I��z��m��Al�&g�!�gO��A=B�a��*C��(�=i��w|b�_ �0v�[��C��MQ��H�u!L�7��	B
T!�q��v �0R����4 ��3�:����-oY��h��5���g]B�W����p�.A��	��W�
�]�H� <����?�o��R!-b�3`���	�]f��[����L���O^6��Qqi�3��G�G�W��H?�%#��ɟ�I�����Ea_�y@;0,���3704�R�I�)�6k�=r�H�����^���ʠ�}W�����ϼ}�|�~L$K���=�ަɧ�v�yOw?�b88D�+�]f��	wj�s�6��g�䉖2�4��v�g_�m��i�^z���lP;y�}D��AF�?����L���I�-�0�I���I��,����{�����'�r!��C9�9\(���������S���6���0xB�t�E�$�*��?R5s�����+�} �G��!�Ҡ$#��H	�4���:4�s���Ic]�w�����>C����T�{�L��ES��N����n�U�A|r[Mm!*��� "#kߤ�f��@' 1�h�N{ы^�D��q��I��Aȶ³���=�D�1��Þ�d�D+�ko��-��&��{���	�j�����[��@`Ew���<����&�sS���]�ў}��8\p[Y{�,Ac���pX���h�Ae<���$�)�Ms/�w}���|�z�t&����N�2��Z�W&�7"��7������2���#�
j���1K*����q�/����>w�ҍ���f�o����򐧞&�9��呲5���a��ݞ�-�Qbu��d�4����aʁ���W�b+�'��0�Bd��!���NW�p�ͼc V&�:��Ƚ�T���+!�+	i2��M�7i6��& �5/{ُ{��/�K����9��D"f�䨨bދwRn����e<���K;����L���@��y�ޘc4i�t�w7�|��^S�"K�Y�xўpYe� ��V�P�n�&��Ǳ��C��N6��7�4�3� zu(��EQ�S�KEzt&5\�.��pv��m��aۅ1���^j�X"-ƥr�:W4i`��#���8�,� �A�R�u(!�xSc���_�i&E�=����OїZ���Ķ���V-,8,�CN+���?0�v���61J����*����r6[mXeh�#=Z0W��!�O����$:`y~�w�c+��%ɚ�a
@H��4���"�\)8x� �@���K��O���k�%sL ���X��r��; �MP��e��zJJG��i gA�!���`H�e�8;Fd�A�af�*��@3>�x�≫!^&bN41<s�ԯ�q�T�L�H�H�w��6�w@r0!k���f�5<�5��9Zo���-�
�G�O*��N��bVr�;��/ =@¿��!��5�U��Ԑ`���eƤoT͚<r��AraU�G���i�9?7��[�5�Z$���,��&�E6&�����71��Z��KsHQ1�Ԁ�w�N��\�4��Eӄ��Uׁ�MU���׏B��Y�$�b�z0@��B��b�i���F�-�t�fl�+y5k$�����m���?$��Mws�C��P�š�<����Y��Ɔ����Dh	U�H�X�6Ұ\;S��á�� �a�PA&��5�\�/��H�&pp�Va�;��&� =�@�C�\!Ykp��q��t	؂a �cc W�p���
��3n ps�*��H����0R/'EKRO��@����(݅��T:�9H�0 4$�|��(���YW���,�3<�����K��K]�����ye�06�S��-�CVnm���eײ����92� ��w�C�D@��`E�Z���4�V�Z�l4�*�B-V�Z{7��%�C���=)�]�iHJn(�Q���b� }���L{�@/�?��̘����B#]2�I�,$?lj����	��V�d
o�A`+5A� $�B�� �Ky��c���������I/a�h0B�ɓ��Q�j�l���p!��Ea੯�a4�t�Cͼ@�8�B�P1�H�|�DL��%�mAϒ7�pr��J���c�C���5���x�,$y�m��)���˚DF��cj���H�z ��a,<�Ƹa J�3n�@�8���������9t�'�PAY^���L����B���鏌��v!��k��3֒q�n�
?�Z�y��~��{�\�ϐא�ni����\���{�%�w��J%h;���fg�:׫n�o7��ɝ�';\�nS���$Vp�tzv�Ƃ����Z���H���9̛9��ʜ#����#��,F HL�Zڀ�f�����9�Ym0�r��'�+�<j" *l���o�SŽ9Dlt&�Ŕ���i������jZ��e��C��x�V~F>��}7�a���Lu5�yK|c��#H0�?1iw����34H��`��[��uO%��AG�aH��n8�*�1f�_�-e?_�P�KJ����I�$Bļ*���QZר�[,��3��He��3�+Y�=� �\AT�tǵ��+�>�LM{G��$P�lْ��!�K��Bc~�b�\��()]j�e~蟼E$}
����?0�UQ"�0�sn4.�$� �??����ĝۋ�Z�<����-��� �չ@��묭�,���I�d`rp�f݆��ꗿ2{j_� I�!`�8��k9��R4.Bb3ќ��d�Sռ�`���{f�G�ќ�a���[{��:��I��9�I�b�J�g��CF����F��<0��a���`�fa�	 {���������\�ؖ3և�Ƽ�h����?{�f�7H��M�XS�X�-7���D|�FX�E\�R%;l»M��tjD��|�N��N��4ikj�!M4i�b���I����jj��ׄN�����r��@�"�)!@Wq	�%���(��Ɯ�A��T�L=���IS4{R(?\#_��&�K�&C�[���	�2�,ͷ�M*!��6�[g��M�[�k[��0ng���:�����nrJ��sh8F�N!�=���oe��,�FsL��/�˺p���4ڏ�'R�'�'"��aR���h\��	D�'Xyuq+����˳D���W��Ը(i^�&��Y8�dAA��K���z�-h����>6���06�,��Fk�I��(mR�4Y�]<I�������֞�&	P�H�B�V1K_O�C?MN&)[D��P����B���AjH�O�����.��#@�Z�`�(I_k/��ԅ/��Dr"�i!�t�(�X�g���'iB��S��i��ԦEK������(���X��7�nh.��Rv1}���GK���k �Sg�]����:�ߞ�����/LZ����({-_�.�HZ��3����u�x �/�F|y&���H�hz|Ƴ��F�?��/�$ոE�?|MB��v�����9i�8jRW�I_����_���S�/�ik���[�x��a��3��2�B��B��$���.�"�"_�^WO=�	R�߮�g��`v�У�n�X.��P;�G0~�ż�f����Ŋ{3t�����7�I+��+C�6t��_�Մ��`��萪�ZJ�0��'�OR���Ii),�Fh�����Z ��/%������Hת����;D�b�2슩H��~�@�WذRM�=o�j�� &�k��X;�W z)Õ�"Mn���z�W�DsǵbLi��U�?��_���q9+�<�y��(N�K6>6n��l��yf$;�����ؖh���B���~���C��Ԙ�6H�b�i�.�#��g�g�|Ye�䩛}�Q�����~d��ضc�×##�~�/<�<7��ц�GiH�l;�?zj���	����\eC��9j�>b���ȑ�~�l��9g���=�<zȞ���|�6m�h�~֕��#�2	i�+Y)e��$ &�jË��0�"�b��9�d\��6�o>p{x���i}>�w�˹�<(� ���&K�6��8��_(/!N��K������P�T�m�<�f�K���a���n
��H5�� �.Hc�Y?-I�i��R�R�MR�$i��\wS5=u�L��Ik��9�qN��pa�?f#�9���I$<��w'�@Fa>���g��51�T�*¥yW_Rƥ>�{-Ո�YZ�MPRz����ƹ��J�.���K]>�V7�g�1K�;�-����5:uZeO��Yϵ�G�λ�2�Xw���C6;��e!�;^��
�B���L-�e�i�]�����3�58�����k����s\�����l�Ęu5[�9j߹�[v��~�֎#�7�ȁ��/�/�؞qųm�:k���b/��푽�����,��k�z�&��)��6W�q�.�;�l>�4��O���A;��>.��/���E
%/�p��\�����䬽����D�MN� �]�4G���#.g���(ˮ����x(8ԑ=l�tf�ds�{��o�|�0���f��E|�>Ҵ���#�b�"Rq��FUե6O�KR��G�<�h�B�4��u��_�/Ҕ\H$(��K��Yi)Ϡ����������R9+�Mڀ$s��&�$+�O�	6⹂I$aӔb��� ���������jIpW�N�R!���|�[����J����y���H̓a[���{ ��%���>i�cr<y��E۹�L��-�Çp}��8��`�4B]C�Ƙf�u���'Б'l$���h��q.0nn�a_��ce��_��b��3�+��qx!ur�l#˷��笿��s�*��>��O�5���o�T�u�u����!܁H	a�ڴ��i�z���s׹��<W8j�I��,�^�L�">��J��2�;���Zm��mނ�����unԍ�����OHvP��E��q��4�4�Ţ��;%)�9�fg�!w5<E��sK0^1=S^Tb<o+2l����;����Ѓ�
ߖd)"L���EA�~ˀ�7.�"����~� �ȷ|�!�#C�+�I�`=1 =���q�$6�+��1>b��3�m��o^��)����>o�L����5������	�AzG���uAӃ%K�h�i��3�3�^"���=��^O�G�A�/A�<Y��|�#]�N��-�N�f?���m��u�ٵ�Lв��/"���f�Uw�}����|N��p>�v����bXp_R�nX�6��V��x}�ݻ�m۟�tr�o
WG�=���5[Hw@ �ݜ1|�(	S�n��'�	~+sd/,Ե�|�E^.!}�=ca��0E}���u�~/�⣶������)��.�E#�	��I�٧��޷z=z��SY�p��ށ��@<�ʔ �CH�^�c=nsS,Y�А�R"���W� I�J�,���u#*�\?xa�Q
!�������1����<�f5�?aZ�/V2��� ��q�He�Nޖ�] i�g{��Q��w=9y�6�=y|�M����]�S@w\�O��د��hIr��@�8q%ozӛ|O����M���<�|i����q�w�=g�����졠���]�r�ssպ>r0��z���n\>s�9�o�#�|�=Y���'��N?�f��2�r���b����8a���I� X�����{��zo
�0(=�`.:v�d�=��!'`"n2���4�}"ps-�0�`�>�'�=��s��.�;$q|�\��绑�MWg!X4�#�+R�W!"���!�6�5sĿS<Y�3��P�]����w��`�0r��
��DF^?�����(jᤂ�dw�yH�Ja�A�O],ӄmJ�,����0��]��.�=�iH��M N�ϞZ��f�����r'eS2�e�9�	:_�e{��R5סCm|�~�Xs���(�C�I�x)�d�3Ns;�Ȱ��FAc��_��bm)��w�w]��z��9���g���Ja�y?ϣ#Ѱ\,��~᷂�d���*u�M�l&'<��bXu�
~hk8E���;��[�}�1�Ot�_����Q�[Bɯ$�B����`?s��h�	:IS</ۂ;��Ç�ك��t��@�5N�8!aa��!%����	���$���6��A�<Wf��8Q�[���-�Ik(��B�?��9��t�P����w�RE��P�,�ʮ�g�k�sY��V��!���Agh\��܋�QV��TZ��#��
��&�,6#��;�+�:��AG�ĖD0�]m���ޘ"�~i\u�J���hrm:m�6l���-��~܎�[Z�C���Zr.Xs��C?��:�m�v���\�p{b;�Y�Z�Y"�������:�>��KS�$�H@Nx�?��oL=�rcn�ȿv�v�8�-��f;H�%O�q�~ѓ��\�ŒQ��@-<��o��ou��J�KCB������!*¥�tzϲ-||�}�����+��E��|���/G/�����5E�Bx�f	6.��K�5��1�L��eRq���H�8��Ԡ)b+)�)H�g �@�!��I�yF*&���i�J�8�gTq$h���;c�u
xR�0�,���H{~Aw�;�Q�
B���֑����P�{i��5�N����6�.��'"?��/��~p����k����Ş����u�ξ�w<���۴%F���!������Ǻ@q�{o>h���{�j׭�����S�8����v�#!)���I����F��w����"J��+��:� ��D8�f��Co�Tq�=w��u�z�>���G�p�d�+��6�7����x�8:fa8~֯[k���7o���K�F�8V�z1�R �հ �� /��W�7>�r���� @`��$aJcL��]s��@1ȋԽkm��VµsΚ�fPU+8���2��-Rz�W(u7��`����FcG�A^;���.An�nƌZL���%Ė�����3]b+��&��|� �fL�l��́�3?s�����/^�,cQ�p
��{��Fڀ$��(\��U ���F7<+'�b������3`>Ur�4({��}��r�o�]NPx?������-��|�=���yO�V.U\3��)e�UlR��m!J���ƥ6Jҭ���3
sj��?��n}d�|~�W�ӳ UR�Qğ�E���i�mvg�����u�L�>:T.����mf�������W�ǟ��Uts	�|;�XȾl���0[A���^v�Ka���?�G����	�kQ�B�휟�)�oF�8j���~�E@U��<M d+�X�y�>ג�� H�l�~�n\�@4��~�Xx_���ᣨr����v�H�}���E�\�A�07u�٣�"0�b&�#�0>4��۶�w���a"S%������{đ��q�wv�k����`��,�0����������x�5�$E��������geQ�%�#��<ii���)��3`vc�+̃&�/5?�J� ��!M��������@a�	w�v�=D���`�����e�4�ǿ!H�!�[���"R�1�A�|�(v�2�p��}�=7*j/�-�	-���H��@���y�!���:���hI�'�e}��7��6�=�-���z�LO�ځ'{�#y��y��a	
��=��0��[�U��<B>4b+���B���x�A�ǎ�5Q�9g���89;r8�yb|�7.�g�{�My,���@_���F2Z���	۾�b����c��[��={
svȃ6{[��<i#|�U�� _�ڇ�Py�]��gن��mnv��ز�n?x�8=0���䙢��u�]yՋ|s�H,"��� j x0đM�	�x��?di1x�Æ������TPM�?}4�&�B=H9��7!D#��0�:!�kæ�c%�l�����@�k�l��aO$��Ę\-��9�Jf��a`���^Z�$ߴ@����:�%��7}�N ���b�� d;�w�G���CCX$� -�F^Z���y䅣��`�ߺ¯��n	����A+��F)�~C(0C@�
�/�q��ay.̅��YCT�O����uF��؉2YMa�J��ܰU��)b�zr-�C���E����>go�h<�a��/�@�U�����!�̟� ���P�<�g�NU�V׎]�b1��|5��#AZ�gsӁ ����
w�Q�+K��o�F�2B�Π;��+�)�N	A(c��p�Q�,F�<���)[�R�P_������oۺ+KwrȎNO�����OJ��9��߲y����/��Ns�$���vXj9��v��܀���5��l�����e��l��.xz؈�@?�X �U���۶�U�}�o�ѱxp�q�-`�&iR
�#i��?b�㏹��(V`p������!�'�?�CA�ǵ4l�|ۍH�Vؼ�J �@���ߍ, ��-w_��yA���ɼra�b����Z�x��H�lP�~`.儗�(�g��"� ����9$�)I�)���T��I�o�&8���AH���3���'��a�;�d�L��W-����@Z�����u�J&�� �E����7@��?��%Mr��~��k��� ��?����!���3�:0��"Θ ^0�MK�씌�uG�e�L�RV3/�a�d+e@U<wU����|�}����"G�ћ�^w�u��[�Rd���0ƶvݨ5֌�qT���[��� ���5�܂s�p>��͠C�3������y�u&��'��[�/����#�$�}���+���Mm�94g��k��=j��DOd�ư��watj8��h+���w��[Bɓm'<�Ԕ7}��	/�@�<O�����>������7�����U��x�Y�����-��@ H8<O�B��<3��g+��"�Lĵl$
�R:�Z���5ힻo�COl��Բf#fW���G����׾�]�<Z�T�20����Ԅq*~�"z�c	BB2�o�)/D7�Ad��H��F�5N��HT�$E��Y*j!��4Kg
�(��pPyh`���� /��#El*�k��͡
d�J����GՉ����>���9hE������"B$d� ��{�k ����_��B����a�XO�-��3�
�u0vy.)/3~��++�F�f��"L�70���Zs��G� 2����'�����=�;��,���y�� �ӷ˯x��>���֊R�ds�A����6;�̈V�W�U+�%y#{��d�>�����^��Z�����l;���W<�r+W
����gO��2���{l��=���;β��0�s66�ƾ��o���E���&�_��I[�:���Zu�֎G�M^�z�i_��F��Q鐺0����x��Ojz)l�@H<�Z�y���`S(=C��G��`q_n�]�u�ɥdU��k������ᾩ���Q�)�V5F4�[��3|�˓��≯�����UP�M�S�����T�����Vau�9)���)���q�D"T�C��	���i?��-��`R���ai��Ռ?����>�p�yS9l���i���^�g�p{�rL��F�V��)g�4D�[j[`�� %K+Ax���)�.Ps���N�����ξD�C���Ʌ�w ��H(������.���<��"s��!ӟ�Tu-���H�vl9h	��%Z�iI�?��ʖpO�3Ʒ��Q�Wݏ>��(�@8K�h�/�>�-�~#��I��<�e��W����0���w��{~���s��;�|�^b� �0g��@|��p>�v�eW��݀A��@?#���/}���_ז�P�����-�S�ֺ�폎�I���l^6�E]l�u��9;K Ҽcmn$�t\��$k>C��lⷿ����t����jc�[���o ���d�%��qVZ$�`�c65��L!+��-0���{0x��y2�h��-���k�Xz���p�qGc3C�f����Z��	���F�����!L���<@`�/�\�t_�B(���hi}U1gɨ�ajt_v�d>�V�z��`��Щ�������ijo�zB ���M�M\X3c��)����x��|x���<����%h�w �5�ɳ?��O!`���{�����+�3�:ׁ�C�!�h�q��ٻhPt��|�рphh�|�f���rb��>���_�^D�	��D�zZ�|����<p�9d��4�ݤ~���.�S�}C�!!��J���0��/p)��$���������|��a����_���-�ܵ��5�����2`Y�J|p�}#st )h5c�1���������h��:����7?_��x�v?��}�߿�v|d43�M��$��O]���N�����	���#	pPq9�GZ��_x���� y�J�ݖ���_�5,"y����A�}r�3�T6���_�MsU��[�!�܀- 	��i$�N��,��=�q8D^:H�H�ܧ���ڇ/djoJ,i�Xq��P�t�P5�����9������,����RJ����
�������b���]���d��F�	?��s�q/*���9���n�!���ј�Ӂ�	��0�o}�[�>��@�T���@$��e�<���<�Ϙ3�@��<%~|��0����m�>���o���<�,T�JB �g��Ә+�=�va\.�7��wF�^��=" բ<�A=H���Ʒ�F��uߧ}�Z��@P�]F�1v��_�_��~����(@�g�g�D}RT��cM����;�~Ͼ��[��`�w�3�y�B�A�~؞x��� ��'��rWЅ���C�?����QJb�:����&�`�>�s���\�&G�T�M��o��$d�H��ˠ�$��H�HLHe
�`��y(+d7�K�0�з�vچM6;w8�;���Tp[>���+�,y�k���^��(�'_~�����W�jw��N'���d�|���$?�Y�zQ��?�;�`��.UJJ�f���V�y?X5�1��H�iV��I+��@0ހ�0��� �!�z�_�NEf��yF��i Ҵ�r&�њ~\���\p7�̃�} n�� 8,NhG��U^�����}�<,���F̃
��{���T��Y�����_Q�i-
e>�[���
�×�I��{�5i�*��r�`�%A^*���%L]X�ny��9��zιچ����ѽ�������-�:.,�m�M�؍??�`�\���GJ�C�Ё!���M8�gl$�RΆ��8 ��R��F.�^�crk�0�'���}Z��s�V�\I��v⛷�!*`�<�l�NW"���A�'��z���| ³�9{�k_c?��{�U�q5�|!��L��Ar�4��ԋc8vQB�{�"�JC�q۸aKP'��X<&9���k�{)Q��د F�=�2��G�w�t8�O��?��/��s����{�<���v?�ֽ�E��?j\~�3��P�E?�B�^�Cب$0Ta0i���A��N{�e9)4�t�s��t�0�2�ʯ?��&��'���^{�΄xv���(+k~���p~������u׸0	��+Ulnf֦'��?�
������;��soz�y���/{�;��5���R�.����4׿`(E��9�ŰR��bR~����Zנ9CH#������,;m'�B�K]S)Y��|�����sA�:g��߸�=|:n(�sO퉖��6 GyF�0Tj�Ԣ(�Ja���c�q���ȜH{!y�sWo��`��sG:Y_�8��u�s�棞\�n#h�=+)�<�*|'<��*��R�ۖ�< ��7�������"�}�tM"@��#��
��:��Kv�X���Ar��q������"щͥ�h@jogѦ�7M!�R� B���1�~�����ʴ	�La�O����Z�]Z�\�
&�'D���P����*�U�&L����	J�z ��|8���Z�x"��5�,�f@���ۉ�	GNSU�,$z�w\f��q�N���;I�����g�����M� ~r7A>9;�{����TԆ�����B�Q��%,��[��'h��k���b��ҡ�\�RB�+t�#M�j�
ԔP�����۹��.�b��9U�}�������mQZY�EF4{���#������w��!�w`�$UEH䝣w,�:64��
�p���t�q������L���=�W�L�`؃>C� ���z`��4ߗ�+0�Ft,FDy�H2^v~���]�ΡZ+7��g�k"�\�;6����3��#��3������F��)"��n<�u�!aT��S6��
b�Y�<0"�C%gx9D^�00
�h>��3�A��Nޖ�ow��T�b�� �i5�iz"����l|�tX�u�+�=yȓK�&��z�U�.$)�Cl��[,��ڮ~�����+p>	i��5���c��=��l/q��V�'�	_`I�;�x�V��p���\}�cӶb�u��!�$�S��S��I��x$�
�Z���_�B����=�Vn2|��+����O��r0s�T��SЄl$�z��?(& R�ŝ�.>�&����&���G}�:�$L|�B�f������O��HS+MAƋ�ϻa x~!$ +��\|��/�4}�7Z� o��峂E<15C4 �ߵ���m���)%J��R1�0̑�#Vܷ�6���6b#k�ݘ�̗��A������Gr�T!�ԾM�4��*���qg���V|�O���\�rZ�4�*�*q������+xBը�3/�(�5MӪ�J�<�n�������=V��
.�P6[��s80(��
̢m�����ʃ��̻K'�+�B$�~M����J�P�Ӡ���ru��M��V�&�=-+)�1~�S�{h�N*wG(�N~i�"����Q�$d��]i!t���1�g�����!�4 ŀ�]� Oa��y���7�_���o�t���N�Ȗĉ���j��ٓ�r�������u�6�E^�q�}�8B[����p�����mG�J��jZ�+x�����m��I�5�-��޶ԋD��K���t>$]��<$$��`���\"�z�H�0Vmn��~�d'�y9:L�8E�0$r��<_I��X��c-��@�d������=���2p��VjE4��DL!�Z.�YZ��\W���ؽG�f����!u�@�U�K_W���Y�HN���i�g0FEz��k��%�IWM>LHbh��0ϐ�41e,=բg4�Z���px�N���x5k��o�38bs�i/��C	E?�H���`m�s�s�+Pp�m�A���~�	R[M;�u\M<q%�+�E�_���(:+O�]>�*�-���I�4a������?���\ j�	+H�5��0��b;��t�d/��uJ��!��k�@��-��iv	P��ޗ������.3M��p�r$"t҆�Ҽ8+51NͯR�^pt�,��ȴ&����LS�5a��GYYaH$$�xs��"%����"�a�J��E_�R�UeA��Q%2�gb'o�jQݞ���A�G$.,���P{?�z0<�H�{)����T�+0����ƂI "Ÿ�|��Śq}�d���=j�� �!w�=�1��l�_����?7�����vq�*cq8#l�\ڌT�M��$�*Ǐ2=�Z�4F`%�*� -ō�v�el�dÕ��$���F���6�U83ӳAI
?��Ē��V�9%]��%b�������@ɾ!C�r�H�#�m#WB�C��[IЋ<md3P�v�B�Xk&�Hާ<@b ����$�9�v�
`�$e��+6D����������j��N�&AFn��ߒh�Å?<b��~g �5'ؕ�׿.�x����]�/_tXO��D��|�U�����,Ы�A{���D����K���^e��TX�=y��'�9�_�è2*|;����(����cc1hfzzƯ��"
u4���`Iz��O	�
�N�`~f��w/���$��m�}��wY�Q'l�V݉?Iܦ��V��(�V��%��2�����?{|V����� �:�҂䛾��%>�)��Y�J�����vi��
^i��C��u_��O����`���=���Dwzf�/xL�.5"�܄uMZ'���=�Y�s�r%�ڹX�qdl�|U�ȉU4��n��,PP,�S���i6cpY������������Ҧݽ��w$/��^ӑD���y�7�Ʃ@�d�	O�;�)�^��C<U���g�s�:�FFǭ�P�#A�{�὞��۾��݅k��H��+zR��P4)yO�Y�������U¦��29{#��byh�3��N7챃�V]h�T�(��V�+���]iW�טSb�B9��k��Ȩz��jO��ǟ}��J7�,I<�j 6��Mw�P���oqfn��5�]��O��aÒg�`��H�7�C&c�����Od�cCn�y�[~���B�]8�k\�)��'�
���ύ����$���B��֬�Ds3s���cl20����ƀ=i���N�d-�2�	?�Ǘ�>
?;�>�xW��S�n�/��]~�v��A���K�/���4��
]����`�dt�_\�E���na�Hl�tNۢ��i[�U\�y�G�N���U����;<56���1�!5�۱�Ѡ����)��j+����S�O�w��%ҔN-O�'���Y�EϋB���Yg���m۶%�Ջ���!��9'�F'0�3�\:<kÕ	�K��+�3�,�w�K�/�}�C��L�#��!�I���{�� ��fi��3�lu�����);K��k�(4;�o���Z����j����)[����� �/��\��>�����]#l�:���h�T)Lz�"��ٺ��ڦ�6xpɸ���|%���7�t�둵��E��"�*�n�N3t���C�BP]�^l&o��ݲѱ���uWu�T�fe��"�?}ih��(<<M� ����+��jA[��O��o�|��%�L�����\��᜔����yخC�q�����G&�����\��0⮝Ĳ���l
�D��Q i�3M]�r�'�}�G�񩐓\}_��W�}dk-�"�E�!��l�zz`L[����rm$©O~�N|�?��@6D{��?a�#�dW��S;�������q�0p�g=�6>����Nد���{��'WA��{��^_�`7�s�N��_�e�5'E .}^�7�@HS���FU-@�Hi6h%*�%����s �'�-�������0���I�"���*F���T�[s����ک֧-c ���O�<V�˓�$\�-x����CONNۚ��6::�I�<-J�-����b��b������zh��>�������)�&�lg��L��5��}s8�s6��}{w{j��{���wv����3�+v�gۛ��3�����T��z����G+���2�F)}̉�m�= �nn�ff��;��O��������;�ܽ�v�=v��/�ˮx�5k��!���h�#�l�$�"������?��/�c`�t#K����]��g���v;p`�x|�MO�Y��iFEIڎ���A��p|i 2<���(�S�	JS��%���}��j����	�G�,d���o�6q��������z�*��@X�٥�=�ʕ1��j�A���Hު�Bb�����E�%����vw��l7�3?�3.����ܛ���%/y��:�L��$�i�����曾���,�p�n��[�v�z���v�}�:u���կy�}�3�q&4T����}�|;yO\���K.��Nߴ)l8q��s�MO��O�6O�7��2f����_��?8m��ɟv�<�iH�7�LyB��_�Wx`�?��?9�ă�҂TA��y�ۋPJ��߅Џ����n#;Ƭ�+[c�aL/<ݦ�o��Ҍg>̼Iq�����2�k-����ׯ_�M�G�ŵQ�g���?ӌ���_m5�S�T[�en�� ���'���ݠ�E[0'�F1�jں��v�E�:�Ǹ[,��-[�Q�
-e�(s]�`�5C,I	��N������&ug?F�׺g��/�T<+מ�C�=���vn����v�Y>�n�_��z�|�]��gYex��=w��w�9��[o?��;�ߖ�eY�� �w�9�������~sP�6�y�������q��yN�`�n���l���<����Co��%������~��=Ϸj��+H8���˗���rVϼ���#�i�U�]��:Y�x��+x7X��Wng���Ă��O���al�K��O����P����D�"����$#li�k=�T;Վ��׿��;��<���h�b.���7�5�ގiN��6��;�!Y��?����:��I����|�����{��p/��~�4�=��kҝ�|�@�����پ}{=�y�w���G\��ʗ�����}Ǩ?w׎3��;�<��;��?�C}� �E�۹ABŐK��G�c�6���[�G�]Dܻ���1�H��qr�?��+|s\p����o��B�F*öo�#�W��'�#��^|O���U2���}���X�QQgG�qQ����;X��X���y<��@L~�B���/��W���7n<� x#�g���t��RGS��ޜ�P�R��Ơ�S�Q�������)���U�:Ћ�NS���R�S��K�'_Fp�U�ߧe(�q=�+`KcS�ԗt܊9�8U4F��\i_���VAy	i���K���{�0�]1��$�-E�g�]o�]_���!M�R<���)�{����x�����FYG�N8�`���-Y��F��~���'7jYs��~ʮ��s����w<�~�g��fP����
��D֭Y�$�y��]�ن��lٲ&m�6_������7�j�-�����i���V�Pz�}c�\�R�tϯ���Ŀo�K0~��o��a��}��y��m[��������n;q!��������o��o��s�d���q�ڵ���N?ɿ��� -Tgڡ#���U2�p�dxdµ�4�9�L�D�Q�����PM�1���o�#��}���چ��tɪeL�)��C_S�_DB�S��X��mpe=��V��-ՙ[��{�oH@EXD��h]I�����ا�`s�*�w
��whR���+�9H�$���`9�+�\I�y�{�1��d��4��]j��zi�)Q!s Ƣ@4�W���[�S�I�и�GR�b�$��3�-%|-�豸�Z�1�l7ݦ�Y۰q��E���	`�;G��ƈ���6]�-����� �R���zd}���&����w�<��mXw�{��fBok.���M/�[ȕ�H�=w�m?��W{��*�Ɲ�w�b�y��v��N�d����XU�K�e�����AL�Ng)��г}�ͫ��!��0���P�|����M7�@�\��?�zB�c[t�l���=67�f��#G��<'���I7�E͉<�}�o�o~����ZǦ��m�HSɑ�BL(F�}�V{�������	�KlzpP��L*��L�k��"h�LQV��T�Y�.�g�E]��p�&���̝b,��k*ً���J��q�͈HZL��k|�Li&iD/M�O�h����x��� A�&02��5��B�T�Q��<VR/�TkH�N��1����7Xn� j@����h��5_Ms���'gё�Dl��}b�<R>SWg��᣶���m<:��5�Ǖ�
�7�%Y��esl,F��x�nإl#�?s����^�B�LL^9�8<S	���Ӏ�����`Lh8DB� p"dAspG'�"Li�R�r�'��e�(lT�c�ר7|qt�I��l��hZ,��TԴ�js�Te���{���[n����]WP���fQ�vO��g-��ZN����:��)T����(�ry��<L̉���� /$�|��y����H��d."N_qW}����Z�n��!���<� $�RB��M	�E8���ko*���I��N��4'��X�����ԝ&RK�r�W�%MC�!e
),���1�=�\��z�l�E�b�������� $'f��	��>����^�֐��]bip��A�RoTAEiiG�=e�;�:M�N~Xiv�V�]5�o���/�|�ݓR�M�W���B��ֽP{܏e���ZexT��4/���+?��#�#�c��9J���p~p�云�1��83�%�R#�Sw�6O1!M
B�u��9.��lxP��'��i�R�#�:b��G\Z����uu1HC�l�m$�[��Vk̅��݃�f�N�L ��}�s~ )��я~ԋt �����A��v�o*6�b��Z�0�9�	kRM)l�E�6O`R��3����,�v����Z���~�C�f!ց������)/�ą��`�}I׸Ѧi-B"����酂t����m��B4Io�1����N�s%�J*�4-b&��S%u����MꛘIJt�0oiM��_f�#�Ҷ`+����]�D�G�$~ER;�'�j 
*�I���<(��>�K学��Ms &�{5#����2�*�Ij[-��\��z\n�|��*�z�o3�?Vm���p���̡D���I�@/�������Jս�0���g��?�^���\;�0w����m:}K���@V����"i�7n8�?ɮ���c���K�4�{�C�	O����(�b�*�/�����a��g���a7���xҬ	� 'ok�֨�C�<b��[�T�3t�Dx��Xt<f��Q��~ac���\:TIWS��h��S��d±�y�c�
�]��6��Q�cY�T�f3��ii���`��}�K_r/ ��W��U����&�w�Pe����J�]�����T�?H��6R���C��ߒ��{H�ZYkŜ+�j�7ˈ*$�H嚛�r3����G�eҤz%��1N�2'1�h���~�.�`���UW]խ��/����uBJ�L�((�)�EED^k'����:i.S��bAz�$5�ߩ�Ͽy�~`��I���٠��-�l�t+�Dx��O�.E���ͯyJgR?��x�N;��	;p�q_?�w�w�%�������1�o}�[. ���o�׽�u��4^i���K/��|��#���5�"��g�T�u�6;�z�ӂ���iB�/��밖-ըV�Nx�?����k�,xp��]jc#�b�G��l�c�mzf���IĂ���Gm���v����!����&�j��w��~�w~� �R6��H[06� ))�F�֢�I�g�B;��KʡO������!��Q�����a�b�v���p����GV�č����
cÞ��s�׀�$127�Œ��\�P��Qaih|ǵ�G��Ԉ��#|]7���o�%�{!xz��J����E?d���r�|=�S�O�+���`v��u��������������g0~��7��>I���h(���d/�� �J|Ιgx�D���%H�h�A�i�,A]���>BK
ӉQ��@�觠4�*R�+���;�Rږ<���է�^�Do��p:��"G���O[����'�l8��k��f3��2�g��U�f\Pr�𑊯K�:���^W�o9�1����Z�?4 #����m����{�Vu�"��g:���6w���5�,�5���k��Bb'>��dtc"!ި��}�s,$��7o��[ny"0���P��DKk���?�.}Ƴl۶���1(P�߯l lr�5�4��<h���җ��Ŕ��2$��C��������=?d�F�8�p�5'���Ӟt�8�� �>�|�x"�M0n�'��D�&����F�ĀM�
��� �,�k9�h<HFƆ&�!๤��`2_�.���H��@8a��%!�-�l��!A���]|�Ů�+�"̞���w뭷v��@�!>0<�R�qE�h�It4�����A�!�`�3sG?��O/��wa8�^�>�����b#���@���x�'�42?ϔ��{��W�H柹�H�x L|Ƽ���\�#&s��A�b��ꓰ�ZJS�N�0w��&I?�S��A�EO��Ko�f���!.j�x��pK-��?g�N�jW\~i83hay�T�ߛ�eU2�ļ����3c2pb4�����e��A�0Rh�'���a��O��w��q�96_mط��M;x�q����Ex��v�%�k��,n�Z�;�;��^O�r<e^Nx�?����G������U��~����g_ye��Sv��ٶg�#{�ə�y��~#\x���áYX�S����1|��_����.���ȒhW6��5�yM�����Յ�-�����;ǼH�R!˴i��G�.�wo���^0�Xp:Q*,"� !�^�
c��"������5�saTC�s��0��I�A��������"9qX�~�p��< ��%X66`'y� ������Յhn�
qހ���?��3gR��ŕ��<�	.��ox�"am �H��ƚ2<��t\��[�������#���1?�@<��y6��y�X��w�ß�e�!в� �0�J+��z����H?���v���B�w�O�k�����ؙDj��Q�`r����=��nl0"����#�´��5�����9F�Zj�Z�	`�3`���;��EO;;G՘��J�8{��N��w�+~�5��.��מ�c&����?��.�ǚ�ߘOՕ�f�\��0`���c����]g�sٱ.���m:�p�+�a��kk�m�����H�n��˩
:��ۊg�N򖺖�0H]_���H
�2T�3w�gO��{�F٨�����t�MN(�"/!#��g>��@��90��]����)L��r�pl�E�ߴ�Pζ����*�@���ߎ�����+�(>$���VaqK��vߧ���o��*t�&O���
�8C��$^��A��;�⁔L�(BdyLAFK�ć�a <��z�R��?���l���BX����ε<��5��v��F��Y#�0DBȻ �Kpu8D���BZG��`\ya<���0��������\3��O�`2�����D��HPP�l*�Ë��H��^�җz?���Aq�����{�0�fO��y.�/���ó���jg^�/�m�� `�E����Fgh��"L��+���6�����Y�����A󥆯kP�6�`tl��ȯ7�\�/ʈ�%{��Tm�V�9?�N8t��Y�.�I^Br��������������~�;cK�N��g�3�v��}��b�]�%g���Z����O���1�+�aܴ�Ȑ=��>����j߻�6{ы^�O��G��9�g�a��c7�tC8��,I� ���w��UY�j��s?�sV��!�*�� ��QX�b�= A}��a�MR�uLK�(����V���A��s��˭��ѱ�OYA�ѹ�)o��֬�����F�5}R>s!� �8Iud����XUm�[Pb�D	�n��B�!��`y�C�3!�H�D'C����P"�qߣ���2�;#�N����!�2�)]8G:r���C��L߸��>�9�&3�0J�DzN��p�Xb���s��	�M�%�^�s�0�7�=�C������ɷ_�s�b�g<���	k�>��^<�x/ϓ��o�2��I�	�b�0��K��cXZA������vػ���;h�A�m Q�2b?���zw��w�c4�GZʾܰ!B{�G�7�}��Ky96�x��}�S��=�G^`�}�U~��:� ��e�Ұ�����/	�Ď19=h�Hē��q��A_��t0٬D����|SOL�q)��٨���Y��h2�	��|��ԧ>�Ź9���/����!X�WR�F[�7�����4f\M�b��P�e��@�[C/�\?Nl�O��6���B�|持��Ƈ�-�1C�������i�E�Q��q�H� �����ġ��sИ7��?�Y;�c�c.!�<�����!yq8a
4�H?�Fy'k!�O~+�C���x��$�2E`ƉF�{H�"��i�f �<�>\{��A���5h��E�1a'A��11�J���0*ր~ ��,	$"<�*#3sGc��H���a ����z a�AE0C��z�C�!�\#{�y&��z3_�����1�^�g���y�1��D�4��=���RD�S����΃�8;�By��]=��X7[� Ͻg?�*_'�L��g�9��=	�O�T���xff�v����n����Ӄ���Y��F�<��Y\�"��flx��t9�?��~߳�D󲯔��=;�+�y���^��9{$��#�_t�i%s�Ң
ד�&F9n���F�!��� �>�tH叾옺x}�vl??�3�67e<t�>�ߋ��ƭ�A>k�"����i-Vي��ϟ ,I���!��������!�G��F�c�:$Y5{��$�#�qCp�	`�=ćk!�ZS�!}�A�a�H��%D�y���_����� �a]Xs�v �:�4�OZ	?@9����!&̌�A�!�"���7Z��A�Ȣ%HC�9���� 0�����|���<m�Ly70�"M�^��k!��+���yd 8�Q%�A��}%+c��,����� ��|�o��~c,�V�j$�Ѱ�ܧ=���4�����4z/ۘe��y���u�].���gنM۬2<�I�b/#�gj��+:=2�| ��q��o��k{�A�!�1��)F�zMI��~�)�`����>�/0�=Q;�d���5������(�,Wm~n�\�s''��t�B��j1���/���
G��� wN��������Un_<��a�(�9_@9����u��D���kn��X��H2T��Ѣ�]�ɦ�v�7﹉���7<,�#�Qp���6z��J�Æ�@@88�D��o���Ɗ��R~��4\;-�.�7wfȔ߹����bǏ�R}����ɯ^��I��=H�rߤ��4�X;�ʡ�����s���> �L��&O��B�e`�/�[�ϣ�a�`��H��	s���p�>6�'����8`H�M��ɘ��O���y�x7��0�`5/�$�����\9�3Ew+e����@�����r>�qu��b���bzs~
���s�-�	����
�w=_�s�G;����ԟ
C��>���0/֗�����U��4'y��Cl�!ڂvkC�[���ͷ;�w;��ʼ�|v;���saP!X$r�,�c�Ĺ��&o�}���R	�$|�vb�W�h�4F�_��_�_��_w�3�� )�.�_wBɁH7��4���6:��B��!�p<���hƒ/e�7�"�|���4�q�����%��0u$�P!6V$b�{�l<gy���&�<宙F��^�S������C� ~��ȍPy��8$qy��7����lt��o���~����l<1�5�
L#�%	�@*��TiO��f>%,C"?�ٲ�X#��wA�h�B#A����G3�Y�xJK�z�4!}��ZZ�����$Qk�5W\�����8�vC[��J{��-�xK���.��ՊkQ.���z�������u2�	�ŹG�VW���cǝ�9C b_)c�������,h%��w�P���S'��-���\�K�nl��|;$�%�˝r����+��.^��|�qCG8�������A--�Ghg��)
Q��7�#p�x�B��</���p�W�Y�%Q��W��8D��`�N&DCɺn��B$0�}�E��d3(7��i~������o�I{�{�c��G����R�$u�ͽ��T���b�NAW���{�*`2��s�/��*	Sp^%�:�|�HV%HS����yz�,W;��
�V`��1�*xP�RF������� $��Rp}�s���� �Zl`�@�D��adozӛ���4��3�O����f��I{�A^\#�V�z¨�c:�2�k��'��	��0V���}���|ݫv5�5'�@����S��BA9�b�.@i�n3Ȝ�3cD�~P�.�!Q�����A]��ix
�ت7�}���2�6�n�DD*�?��So;	��V*��({����B�|'���R�ͥ�\њ5��� ����z�U8$�T�����ẇ�k���~w��˳GH���E6�.�K"�px�T�:b��W��'�nY�`�R�s���L۝�H�TAD��0p{��{�ԩ�5�D�%M��Hʥɏ;M�JҊh)���4�l*zF��&��RI�&��&`CW��O>��VD����oi�`�A��-f��c�g�)��h��]ஊt�D����ް��w�>1=��T�M��2"��U��[�-%���_o�~n��-�)�c[��3�/0�@�9����p����~��ֶ�y��M�f{�c6ng�n3˻&�7�F3��U���� cFg1O�W��񮶃���张̢0E��R��e��CY!�N���2�b!~��V��ϧ�+�\�&��Ri�Z�Z�v.&�r�' ���B&M�,Ҍ�:"N�p�5��:�{�����?l䃇��Ƀ67{ت�S���RD�$��v��5,�)d�I[K���?�%�J��Y`�TAT����q���H�H����C��xC�O�囘� �x�=���E�щܐ�	���&?�7ݣ흤�D��/4lt|��v��*hxl�S:S�	�A��k�-�BSFtN��i�i���\�f@�C����w��#��Q𿛭�f�t�
O�v�$5�jC�Q"m�W��w`�O�V��b��XʱPT*��E�)%y��3('�6-5�*�w9�Qj�l��8���x��c�Xo�@�|� �/dϴ���$��9��)#'������ϵ��q�?��=1�����sI������~���o��0��1�H�T���[;&v˵�-aM�%f�g�=�����5/�a�Uv�}�&�gl�m�7F���kڙF�g�`K5i3�UE���������vF��Eo�J	���\����^�|�[�J���d� $��m��A����S�q@�C�OE�e����� -2��S�JM�y��;���}���{S�}+��V��sso��9�����k���n�bwio�ji�I߽�_�w{��٢!(�8� ���=�y�8�Ѳiy6A�u~�l1���g������ ���o�׎?ꖂ@�y��`o��2"�ԭ�x.\y�%>c�����,b�CS�y���t(�"xMj!�C���� ��$E��ԷS���(9�QMk4�b��?�JX(��F�.��U�U�<���^z1w�d7�HǆJq�w2H�c%k4���)�.#F���2{_5�q�8/�Kl��٠�F�c.�[�,�1�[��[¿���{r��{��l��7��1�胱��-���/|ZU�jH(*-3m�F��m.mBY|��ִ�����1���w���ش���5t2W�mgƎ>�@�1����x9W��C���p�F(���K=�۟�7��(J���=J�
�5��}�m����(�!C���H��t�8��B�^o��C�l�S'-�rm��6��=�l߁63�g:�X��ke���BZMk���a�-�6�e�f .5�[/W0���؍��>�Ϊ�1KY\����l��_w��h�:��V ��*^� �8b���.*}�LF
��C0��'UX�s�=ç9㔰P:C�i6\�ѩ�C���J���{�z7kh��K�t�ދGB��&�W �e#^�R)2��Gy�i@��c����<��o?RlyY)=�S)������x��V��xtσ֜���Y��#�{�68�4
��c�`��h��9�i4�jQ�ˣO��c���֑bX� L�3zx�B.�(���p]O��f�GP�L���)�8��ӛ���pH�Y J�І���u��q�6z����\8��H���=���<?o�*�k���$ɷF�:ַ��M�ۻ�����gN�sAX�mf�4�jA1�4(1}l��u��l���^<i�A�GDe��l�m��Yrɹ��+��t�b���S��!�I+!AB_�~���X�ݳx84ۊEu#�a�U�ޖ��.x4b��ʵv�78�?¿X�� \�ctXO]�fpl�Zq����e@�H?�W�ݣC�v����ڵ��l	�DؿȔ}���:~���QF��l)�xQf�g���w�7;�9�(���[��thb����@��P/FF�o�s���դ)r��W�RC�9�R`J�y�K�q���_�u�Ycf2X'eg�t�C�+�q߾�v��;���	+v+1w8�~�3T0Js�(FEX�mW�
������� T{0;?��� d�H��9)��;;��-�'Y�m��Mv�5��=��a�y�aC�5�޼�;�o�s]O�hw��ʷ��O��Wz-P�����W��I��~R�N�_��_w&�^�9�?ˮ��*۲ꐚW ǽ�p���;wy<�{��.���ډ3�+v���x<��z�>e��,�x���꫟f/�����#�7�b��N?A�5:u�t�F��M�(`-$ �!%�L 	w^G�� �����5���^¿ ^9i���A.�?iǚs*!�m,�ȩ��SA���S�D ���}���g
R������?�`8C�sJ�¡��-���6�*�v-�5�d�<=���`��V�����1���E?�9�I�����2kU8_��ʏ����W��X%��9n�	�Xj��߲ҕ���	�ѽWE�O1(UO�ޫHOך>�����T��Y=c���2�^�:lB/�b9X�e
9�� h�M�c�a�XS�x�b"����V���&$=��/���e=c����y���ʯ��i�c��q{�w�]�4z.�����0�i/Ɯ����aՒ]v�v�,�`�o�����OkI�EO�%�Y/��/K��i5���`�o��K^�"p"�v{����o���M���~����.��R[�f�5�mgy�RH�*Q� �P<7}�o�[�3h���^+�����"^�q�	�L}&,Jf�y��۴����=웶������8
����t���Z6"H�� ��Vo�TA�f�k�8m�"�Q	c�$�T���u�W�Jx��ƙ/sRe�)ǉy�Ŝo�!���L\Li1��sD�s�񚠕4Q@<>\�^^�x~�)#Jկ���� .C�E��1�7�4����ž��(w��n�����7��Iqn4fmr�v�jC��-Y
mv;�,ve�k�f�s�&����f�n�F�4�������3�8�c�%;�԰��:���S'�ѕg
/���p���k�pf ք�si"��9j�zw(w�;lF�ú5k�&��z���Лv����W�h���u;~���DXl�w�];�ˮ�:�k79.�u�۱#G�?!�b�r
7^���|�+_��n}�m�h�������Nu,���!�=��]�a������lf�D�\:��6���OeHx���={���g��>�����݅�;�����pg���V���n�
ȕ�W�]��x*P�P`��<��g>�Y'�b�_��BO5U{C�!�̙�1�&('x:<g�X�����wZaxpD�FM�g��5r\|膁渖ok����"(�����4u1?Xo�������q쑱Q_�:?���D��A��uk�z�0�����gW@w���p�T�)�߅bֱ������ׂY�z�:[�bC�#I���Q	�:��kϟCDn��0��a�Řbm.J+�e�8��m���{���ҿ��;��!U�q�5��u7��T3�^z�S~�C��1�J)M 9��_잣�O/˟��Y*XU͸�ᡟ�:IbU�����^5j�.X�<:�z���C��׾����v���C��!��WJ��>��hr�0<(�U~�'^�^	���C_�<X)�ël��~��{�}v8,".��N�F���cq�g��i� Z�<6@���kEB��B�@���?��@3 m3��=z�K^����@�c5!�9��P(T,u���a� ��)�a�y9���պPMVd53W�)�!_�� �Ie�o���qm(+<<8͕ J��v���p��;�A^m���C`p?FǆGFI��������X�Pf����7����\8�ڱm�Si0w�k��͚R��<�_o)*��d�cࣣ+m3m��(�f���n,�,,��0$`�Ϭ���W�Q$cH-�'���>�g�� 2����e�U�ׯ%<�o�sή��
��w%�F���O}�� .��i��o{5��?���v���7����/�3X�q��:��YK��_����Um�u�o�� �&�R�88¦:v�MN�� k��M.��x����8�#*`�QYs����y
Xt�z)��u����EpO���-�u� XA?p��V0���52~���;|�#��H�r���2E��X�m'����~�y�#>���ѹO|���� ����[�l��,�Ga �x&��s%���h��q�5kW9$ǳ�y�]~�����\�q|^Ûcsc��9#����(����!���k�E����-QT\J��̱yM� mjR�|)�n��5ǽC�n���Y?NW�.��Șٱj��{	�V����q7��m��I�J��P ���{�)T9P��s^�a�7rl�F
=��]�z��q�����=��ɣ��r1��k�s�3M/���b�䄑X���������.��a��+��w�;�����/���gݶekx�-k�j�#��7^ikVӏv�ff��=�`eWmo��4� �og��+M==y�~���E�B~N�K��K�sW��)q�b.�^����j�����>�KG<b1/}��Kv1�VӨ)����'%KU�(�#�Dt&FL�����-�"����/ӿ��Ω"�p���J�yFT�JC4'������;Ne2BQ�Xxfs��~L�;׆���t���N�^���nܜ�&�0�3�=2=x�(
Un�lX�^tA @����}�QkD�+�{3J�/�>;���ZA` ,/<��銻}��6;q�S�[(D"8h���aO��ۥ#v�nŘ�O])��)���;��k�u�4g�A�¡ D��*>�z���Ԥ=��=�rŰ������#���v�G�R*ة'��ذ�B��}op^���z�g� �z�_��Rtv���XN��� �N�,����a�@fV�F.�"��v=h�a���dP#���Q�?��?�M�Pb! U ���Xo��|_��d!(K�x�Ҋ�Ƭ�*0�6�њ���ɰ ໯�p�.gt+,��l�B�yh������]X� e��������X�,�f�����P�\;K� �5&x*J�󲱸'p�K�=���~,0��g~�g\� ��g��fR������[�ͥ�s��=�v��
�d�_6=�k��g�ry���kF�?���v%����'̕��@�̵���kc.bC�U3z��2a]�X�W�s�p>�g��1pϸ/jCyn�QH	tm1�?)�<�X�_u�W ��=yb�V��|��6�L��I�pK=���l,�6/eee1�Y�@|�4s����«{��{l��Ƿ:�g�E�p����S���0�B,���W�<��̉���?�y��IY���(��̔oڑQ6����A*�U,Kl�)��iz�f#�T�u
f~����R��y�b{!��c���9;tp���}oX��66^��k���E��@YZX�۷�#C����+A܁�@F��E���k\/��DM̱���5���N"�k������:΋@�;Vp6��c']�#�Ԝ��،��^����.3s^�zE313�XPףt\^G�)~�@�o�r繂���|��Ԁ럘��������Vf���G�P&x��ȍ�qn�w��^
־�1��	؇�T�8��i�FA�5.͖w�b�;~Ć�ﱡ�UaM�[��{��k�#���S�����
��������a�������7����z`Ȩ��Ӛ���ke�(z�d��"��"�@��b,qxd��Z�"W,O�"���)��>7��l�]]Z'���Ց�)~=��K�r��[��7l��%�V��p[�l\�����?�������\y>wki^���e�?l�sAIET�3g	��E�(�"��ur�[͠h,X����u�0����H�s���j�
V��/pKA�2�
e���~b#x�pB8��`��^�ʯ�?~��杺���[�¬1W�k���.�q������#�jժ�֨ovܡAM�/Ͻ�9. 9��ب7�n4��ޭϸ�ߓ"`�dg���}��ܺ���+"$�7�.Jx��5���O~}ܓ���%�l|�F�m����k,���~�w�r|��Wlz�7���;��B���r�����(��[�9d�<Pd���/�y=�Y�v����� EI\��0/�~AJ[M���<U��0�RC��& Ȱ�qTӡX�֧��i���TťF�!���� �뾐d�p�[����xk{k�T�e��1[��v\r��׃< #���S1hɕ��q�Q�����[�?��'��\د����ۯ�����ҋ/� �����)��JT�%�@���Q�t#�X��t-�W�@3�ylx$�g�T�K���R�y���j�W�!K;���vX��9�k�{�iG�����w�k��9�U5�E����ի^�P�0ؼd!�����j+&�Q!m^64�D���>;z����e�*��$T�˖�B����Y�g(�
�m{��^
 �}bO���0	N ��և4����pN��9�Q�/֋Z�?�wP��,&yBx�2�a�s��fD�'�+X��u|�s����C9��zZ���1����J�L�5悧!aԣ4���f~��c)5��B������.�E2o5@W<F���Ҋ�MxWR�D�K��X��� ,]JR���v��z���PŸ���R�.='N�f@�3�^��sL\����(���8y�{�T��'�Z�S��k�(_������B��~Ϟ=�'�'��׼�[���-o�,Ω&���W=ﱆQԫ׭��bSӳN�7^̮ەV���ȕ�e���Q8ݵ�Ϡ�Wp��b�7��W<88����_���pݵޡ�۞���C�e0n���uހ�߰2<Ԫ�;p̨�A����K��y���wz0\�\v�BXW]s�o~`m�٬� kyfz������f��m��a;9=���iD��r\� y�r!�+�y��~C}dU��o>?���`�"�����`��]�U5C�H�_�zsU>#��&���yO�T`�X��6���P�����>|�M�5�y��F癨Z�g�޳�_躽7l�M�1���|�P��96�������ؐȫ�[V����^�PR�Zi�8	"Yв��B�@SN��	�*ӊg�ȩ��e��U�:w���ɭ~>j�����c����W�Y�4΁�H�H%& v
���DY�z���H�W�4��eu7s��\�X뭬��@'�?��'&��|���.�](؀��2��=i�&gmhxܠsvt!�Y���7���}�+�؁�/��灂�"Y\��H���"�L�.9�Ë}߽��ϼ���Y�x�6����AV��]87���[��E���s��n8>�?b�T{F�Ӽ��O+6�!��bx������+e�ґ�>�屑!۾m��_����:x�<�a����CA��=�U���BV�������.�!m��K/w�W����&vh&\#�3B�F�@{�	��`8/�
�C	�0�xE;Q����3�u)F�2�\�36PP0�	e�<H��~��x<���o|�=���Z�(pu��N �{� g(�����q��|�����/��9��F�=�<o�d�[�� 歴����=���=�뮻|=)�V7K�˛J!��}Rn����LxJI�8��RPEw
󤰍��������+�,a��+���-��!�+� �=X{����_�����a��iZ,�g�'�{�}�^����~�����R%�ͺ-�o���@x���<P��Y�����u�:�sb �Y�x��o��M�k��|l�~�k����4�A�tl�m�y�%���M604hS�s����B����g��_  �f��j���ȋ�O|���[���m�~�w�yd�^۵�A����+H���˞f�_y�]|�����qc�k��h��_�W��y�L��E/z���%
�C8h#�z�ڂ�ynz�>��OZs��!-��1����5@�<������`��]R��+��źP���z�k_���?����� <�������T4 
�J�K"P�%������Cyb�*�&�0L���tL�/�D����gȖa�!Xو(���o��m����i��{,8Rq�\?��?�0X.�h2}ڲ�Q"�x���.8���T�F�=YK(���7��9���7�1���^ )��e��%lH��f@�Eֵ�q�P��iuu<y6�w�
l�C�N���dm��.VZg2���{ �y-���?6e*���ݳ��{����A91��-/_�6+mbr�ceP����;mF�����'�vvO)Q�C��d�Gq���+5`X7�x}�C�֭�b���>��]-W|Τ��_�=�����z�&��a����g��q�q��~�
ݚ o?˹F�>��Ϻ۲��`��ƛnJ�{��~��`�+׬���.�e�"��E� ���ᘈ�������rx��a��Y�A!�$��<��wx�w�=_����`��:�!�(�u>zl6���rh!�Se/n��>�-/�1/��Qn=�M��MДkG���6���Kγ 12�E�	�b3pl�G�V$���*����̅{I�%n/
��3��=�H���B/�����;��fnT�FOf��/ރ�Ұ�����`����VQYH̓�^k�B����O��	b�S��Ҩ�F��'� ������[ǂ�u,>�='�h�S���1�*W	qF��W,@�[�B0����Q�<C�-o�����[���ӟc��1[�r؊����ʞ�I�;�=�5�6���yn��K�o�} yld��R*�'�w�?\�!��M�X^ׅ����FQ�$���Xx��֯�U�/��n��[w��?u��2��o��6m���0�w���ѻ?����+�Y/��ֻ�;�T1p��`�~d��ٟ��^��Av���k�k���HŬ�:��X�ln�VA$
�)��`RV�\������tK�E��������w(
B����Y�Oz��T�f.;,�/��S�V_�e1  ��IDAT�9�N[ذ�������
��=��3�&�
��,|\�T����@�\#�8��1Ҥl�(�
!���Ȇ�ް�8BOE���Gys��e�f�R�����h�3�g��E�rI1rY�\�,e:�����~l��!�Y#|��B��s=��ǣ��Ul�$DdK(J Kp��K(+� ����
�+���4{DB\i��e����|����$#�y�K橸�2�4o�)-EvU���n�Ev��WS�y��V���gf���[��+lj���1�|h�X��O*���tO=#�򛜎�is�>g�췗������~��z�Z^EVpr�{�����^��^�5<�<X�+l�E�mnfֳ�FG��.�+~�#=�ȁJ����9w�8v{��O����N�� C@��Y��@,�w������n��6�,V�ɐi�,��Y��>v�G\`i��0��@����q���Y��=�x�;��X��%J�%1#E5(�JǙ;K���
E�}
��_��]gb�D��oȃA�2#�	sF���#\�����pl�9� �V�ŀ�&�{bGDx��;���?`"e�7/�����: ��6B�\z} JE�[�����r~�q)���
��X��^��;�c.̕�t���qߠd�C�,��3PSp���|��ZB9W�U�Pe�p-|�����P�fjy���R8U��"0�#�B� ��#��*��uy|(��� ���y���k�xf\� ��?�A���c����8Ć���}�T����U�"��{h�f�Vۋ�ʵj�������E��@V�u(F���5�������]D�X�y�S�[����g]��-��]���62dM0̠�����=�v��G?l����3�ckiI����6��ހ0�&�ed�<�QK����}&XjP ಣP�G�G�Gz8,��f'���k�"E� ��q6�d� (X<��ۿ���i^�R4�u]YMMUm��	+���κ���wߧ��r�c}���c�C�{���@8^x�_��}�V�QH�D��9�"�6 �S6,��������TF�
������
G�1�!����B �>�dc"�`׽��r.�P%�|�7�e����>��7��
�p�@ �!�U�P�?�˵s������b`�PM0W��'k=%����d�=��FW�X�y��,U/�kn��V��ز ���Ǽ喙0�geYO���{)���=��e8ʑs��Pp
��.�4뽖Ѧ��R������_p��l����ɪ����2͍���)��[#��s��ǗŶ�@��Ś�B�}S0&/��J�X�������͠+ŮD�r��q�����,�L7���k����` pe�{�.?PQ�9�5 ^Љ�]j���
��?�!�{��͌�˩�x��	�]�ͷ4,��dq��45�ZeC�`�������/����O��
,�3�����Mn�⡽�>,�^�V+�>��.w���-.��5d5���E�@pE���:x�+_��닻�)k��]@����`T������T����l~��jV̣��:J���	kW�+c�%��W��7�r�����ͼ��:O5D�U�&�e{`щ���'�'�G��֑��T�(�+����\���&����J�w�f�Q���hrr�_S�XP�j�Ny�"!�'�|��"x]�(3k���W�*2���L��u�
��B��_R؉������kG	����5����J��u�&[�vC�C���F�f��2Z�ڡ����=�p�IH�0եp�����T�Ǌ��=���S�>�;*ume�Vx
"����no̿�]�'�]�5�e��Q24�7>ZT��B:5�� �X>���M�<��M�Wit���k��`�u�b�F�����Nc�n����pz:����H�Q�
T
���B~��2L�`����� ,��?P,@-Ef�Nf�7i����g�0r�<�ShcJ��hKA;s�ֲ�����"!��+y��z������*|�^H8����dR�^�J�F���q}�#c�-%����*^W� �3�,87�e��=��o{�E2�����`�c�
�K��p������\熍�eW\�ﱽ��t���=�����u�����f)�<�/$,��"�U��i��vs>�薧}�+
�#�?I���_z�Vw�����g�#>\��Aq�U��ǟW�]�٨��+k�_?���Ŝ��=�=8������xj���6gJ�Y/����q�t�eeҼ��n{�MۚO�K����nXWX���z˒����K�Y
��z&+����)g�B��Uv`��� )�>�8�AX0X&���gr\�,P M�N,<�U���lp,HÁ8��9��8J`#ă/���p��b�*$��=T�
�HlŋUJ��x��z���,�� ��9�I<�(���x�9�+׎@d���/!�g�G���cP2 �Rذ�|�����ٟn���z3��7� W�UB!�V��WU��2uXlz�9�Ph����
v#��\|����s.����꠆ף �<�����j�9ǥ�u%��5_���+��ݏů�n�#��9�ei�Sa�<��=�z�Iߠ{h4;q��b@5镲 ��t���)���?�'�5�<P*ts�گ��BLKu�"�X��sc������_�a�g�-�j>�E̕@K$K����<�����))��=<,R9��~�^���yF�K��#�û�M-gF�5�"��W���^2��,�Y�W�&��{�U׸ %�K�
��I�;���{�\���Gq�7	���0J�+��Pmx����;��L}�
����h��LP4�B���rl�N)�B��CJ�� ��9�
����5��X�j�5�f�w������,���

�`�ū̚�j5� ����x���� +J���2�!��0�W������7����1�N!�̑�@�F�P�iL(BYJ�-o.b�B�F%��'���y�*�z�b&��B���S
�̯����ql���(ԭ�l)�<���B���VF���4+�LZh���U���`�n�/�p��m��gPP����c�I9) �,��^@�s�e�� �2x�E�����F����������p.\�au<_�=���l�ѱ�3x�:E6E�S������M�/]kl�"��d��ĺEp��!���۵k����w |�4W�늴J,o�K�t	*	8��c����y+�4B����_A��H�D��u��7��F�� w�X�j��2R�s�-�5s�(3���ÛA90v*��!�D_�y�����+~e�(@�5�I��$P|�&�7����hE�Y*�|xA�?���\��E��d��� �h�����Y����\}��2���,.%υg�ץ���'��f��ĜQ�<_M
�i��"�no/6�]=����Bs�p�C��U[�:�̍���9O���Պ�n�� �<G}L����5������T�d���h:��E���0�b�9Z���?�������9��3Y8< ϭ.ƻ�ng<&����Sˀ�|`2D�'#b3w��  �c�%�=�J�;q���}Ȏ���
V!V6OS��-�O'��S�TQ*X �4�a����Z�H�!@����4]EFlz�� .}>�1�TʒM�<��s?e2�F�qQ8X�X� U_^��\�x�;�ax��L
#�J-�\��5�=�X�y`=��B��� �a>QAY�YLɬ vz�h�z�:Jc�+u%���c�O��&��5 'I!��<A�xR�>���m�>�_1Y�xO�o�פ�Vz��I�H��!�J=���N^���w~�b�b[�Jl{X�1��	*����.�r�_#�V#��Y+-��n�'U���Ih����x@�qnJՍ��R��]�օ�g":����3�.�g���������6`NY�-��}ou������W�7��).o_�5�$ L���m��p
k����c�lr☍��j�#�2�}��+͔�gyZ�!��<�����o�'m���%s�_�`�>��Kإ�����"l��:�G>x@-�!�!�KU���e��"�
���!��+���%��2��`05������ �X����=�n]*fJy��kd�xR^�zRПav����L��!��)K���K��Q��k(t�T����������ͣ�"�w���3n�նl�(�����~�a]�ךd.ɂ-'�l)*��g��]����������9���٨ (ҀX�N��)���nVx�S;Ik�">ǉ��{[��	߲��4��h�W$ռ�Q�h�~�w�x�2:a^�v�;�6�E��_7�s�ȫ7��r2��S4[u��|�U�q����NA�,�>���i��$�ѣlwb�03�T��5����A,���p^]y�l"��XlY}���V�v��c��J){Eo!,�f�b���=��٘�e���@�|A#�a�#���������6� �p=�{ѵ�]V
!&]τ�c}�#OP% FL= ��e ����Е)�Fձh��|�ǀ@�~S? U��ൠ����|AF���I� �@m�><M���L�Ac��&hG�>ץ�]�,�@x��s��f�(0�BF��f)\���0�fI	��N��Z�����ܴ�����~�ɩS.\f��5W*�zZ\�
p]k��n��sn���W��� H=)6�Ou�4%��$:����t�3���m;?W̕+�
��O���^~���-W�P%�ً��'B
u����=/�?35�ߋf���������-��{����F*��-pE�9wP&���t�)���9�X���x}��۹<
���k9�D������4#L.ndi�ܞ�8�F�"��z-���*���)>����^B?��+=u=a=zd"X�E��� h�5�A67\�z��Y(s��7�6�(��SgScR��,0	8��.X��M������0{捀U����P�g�����d���je� ���̊���s`�@7���~���>�<��96��<,w	@��T�)m����A�)�ϛ���R�����86�'�+�WZ�80��ԪR9�R�R��$,w\�.*�ytM�:��w���o�-�̇�������yC�c)���3�"D�\�=�}��
�����kIXCs����y�
r�6@���	�[z�L��,jf6x/��%��9/جt�г٘�}�w�Z����>׾��1sϫ���(dJv�R��f����7F�e�s��'O�c���#p���-,h��N	�c��Z�:�?����oΝ��;W����nӘ��3\���2F�%�.h��\�^5k�*?l�Us>t����e' א�'�[A1Ǣ�D��t�?�͖��x��a�
�xF�\*����U6[��M����d����[x��s��s!��p�4��5��'Rl�G*]/~�	�� �W.�R�<�e�I��}��bl�����	���X��A�my���,�f��EX����+�y�0�����S�B�_P����B']_��jϿ����#s/4[+��S�H�&��p&q��<#�%�;�����{�>	x���(���Δ���bAZ��պ��y;�W�$u��IኧI�N�������&[����{eͶ���q���M���N�\��{-(�L�1�b�i�펧���?<<j/{ɋ=A ��b^�������9J��^�g+�@c@"W)Ÿ��̔{Jp�7W� �9o�ĺ���q��Ɏ�_��������j�@�}����y�V�:d�@�w���BD
,|Y<
���O�X�T����,#B�-�������Q;z���;�E,�V3α)�FƖ�l�aC���A��#�U��֏Z��+g�4�X�??�@6�|^�b?�-A.�T�\�Y��LBL�.���\��#!�znj|�"2e�nR�+��\%����ϊHB_�A�H��o	���ы����(��*�!~bg�Nn�ׯ3:����J��/IC�&	e�-`.>����{)/����o�)����Z�B�����C«�d6q^���`z&�D�.�
G�NJM�a^��V�z�s���a��lnf�s����䐞��[6�Үw>���g�
8Oɔ��o�s��L��=�g؋^�b{�[���.�w���5���ZԞQЛ�B�əY?���k���$��Q��r�a�}�p��Y�7�Yz���P��*@���ew�U�r�j�`�\*n��_�����S�G��6��Y��cA�o	Yy(8����`�B�~�{�ч�e0����Y�B��g��{��y�a���K���w=#������x��k .Y^�Aۮs�p�'ON���H�јuET(�l�ju �{�s�*�X���l����`���BX,�
�!��Ț!HŻ�e0J����}�;((6��Ș����ȣG�g��M��S��>�h���e������ �v>����j�=�� �)z�(ޗ!�w9���k���0T`W0�`��������e M��DU8���9��;#��s��/���ۻ�ֆ�T��D�c�i�P�C��p��GF�TfAn����3J���V��@,�����n���Ea���Zv�����M�=�r������}ͮw�r��(��|o�˷9��1Q�P�P�� /�����(C��L�FO(���O:/��7���8
��# �Y�G���|���E1{	:���3��H�8G{�v�0$(����Lx#t�կr��a�V9��Lh�Ć��sa��'�&lU֭�>YK��L)�rs, �@�.)�i�2��j����@�.��V�;l��I���]1��`�ݒ�x��>+@�L���K.��5(���ov�"�2H�)��9�k+%S|/d�|�w=��X7��ʓ�(�����$%��$0xj��UK��%?�E�%@�(YJl.��$��&'<o�2!���,|^�:���%e �;�Y�E��?�"��^�qI]�>�*��<H�Խ��|��� �h,t�di�����}�(��	]�&�&����1��{��E�0_�����U����K+Wr1���mr_�kN3�� �'*ϰV�\�$�/������^h��2������9gqu�C���(���LLĊhkG�\����K�-˖۝/{�C��aR��c]��e[�f��ر�>����������A�]��ȓg���7�ǣ�x��٫^���za�fc�EK~ �~tt�Ɨ��-�0�*h)��1ɒa����E"�EJ0T<X�l`�}ua�9=.���W�,�bݩ��S,�4����\}*K�+�5C;�6��aS�ؘ󕅧�m��s��J[��2�2��AKZ%�A��M�~�(ā��E`Rp%:,Yb(A,"�K�'J!M@�cq.�T�у���TL�� �Q�(-�[j.�0`ŒWz(���Qr=	�r�Xn;�����,f��=�؍�B1�bD0���W�<�j�@��z�����
e�\"�	�4՘!�ε��P�j�.��X�֋��GZ4���j�Y����/��/�ڱ����x���;�d��������f��1���Pg��;'�,�P
JmOi6��4��i�}�I�+*��h�N۝�M5:��S�s}���� 2SN�Y�O�Ӏ��oϞ��>f�)���W����ړ�K�-�hX�ϸ�&�pi�hjjjL*/,c��j��9�U�8���)oϪ��Of���!�E�f�*�>Y�j�����{Ͻ���v�����Y	s%<��o����&o�c�E�1�"����&��g�gsܛ�A
".$.6��Rz�F��U���r��E]O#]�|u��5fO:��C>�*yJ�Sp׶P�Խ��W!��(�兒�|���UW�k���9#�j,N&V1����w�6%��M"J�h=E�%��EѢ8�.
��x��PЏ���pN	p6$B%�����h��$� ��s�������>���{'��MLsn��(R>U��w�f��1�dF�b�z?�M��:@��ޑ�z���2\R�����Q TEE��S�Y���KR�1��3KV�iv�Y�C�K��7J�NuY�:��KMg0�����H�����'ҘA�{�&&�����%S��$��
{�ہ�o���.'W�+|��J���
t�{�A��zXC����x���opo�����"��P��g�S�K���v��kS����#�/���o�kxN9Lz�u�������{1zX���G2���n��}��;ۇ����A�_v��v��O3x�[A�۳���_m��a۸�r�T���%���gϼ�v��W��@`�R8��J��(��Y lr�����l����-�4�s��-($kl��m�z�f��>n���¼���:O��w=��sY������a(���a�b�"���" �0X�@���{jW�k�@�3 -�{�E� ĺ>�7�e���`�J�?c�ca�T�~���Y���&eǨ��������� #��|�NA+\�j�9�h�sǺOy]t�P�<s ��84\B^V"
����?��� ���	�WN����ZZ���k�Z�>(k��9?���Ȩ��f1��S�ǳz��_�`���ՙN1
]�e/��4;Ią�����1�`���}���U[j��>Z���(���6ۚ���_a����C#nu:��V�I�����E��� ��w|��W�Ws
�=q��N[�ض��v�׾���
�t]�+"�i�БÏ����{�9w|��_����M7�b��~�ב`�T������/�����ٺ����M=����o�@�����8h�.wpjj�N��6�χ>�A�x�� A��sYQ�Q����	k���X�i%c�٢�z���b� ��Ҵ�e�e�k�7��2�x��0��sb���u��ӿ���֪Rf����Y����9?�!�U�L,{�9���_��s�4V5�� �ʔ��ō%����gs!D(�����a�X��<���]'X����y!��c�i����!��(&��uE�9�r�y�¶96�F��>����R��+HY7�(�aH�������7bJ��!�eaQ2�0Pe�}�e��:���a�k6����&\��;����2���dw���\�,y"��bAٙ�Ӫ�Փ^
���\;�|ݰ��s-��+�A��|{��[-��kT�chx�"kUƑ�Rd݋J�xz~$LM�8a�����o���p)��:�@��������W�x�����pҳ�%���i�w#�Y����T��˯��Ղ=���v�U��E�օM��Iϝ7?��u}:��e;����?�^���������\$d��ԉ��#�x�q�Aq�����¢��y�>z$w����}��[KV*EXyzZ1rxƍ���Ѕ3������rJGeQSEK�
x��d�ј�t��",��jD@#0�,BP]�Ԏ+�{�o6B��`�# �Q	�b)��S?�S���"WC!a�� Q��&���?ޘ�����X|�g̃2�k!��5���� ���>q� "`%�2c�\�ϱ��|��5A#d�p���)��Y��SS��+�eq�1�Tx:�JMv7/��%��En��o��1x�z�|�9I!�90g>#8�g�{|�S��g\����B���9e�Ⱥ��`<��G!YۋX=S�G���Z�زѱX���oY�V��`q#�wQ�ԝa���>��v������*������/��/�JC�!�x�x��`կ�fk¦�&���.yOP���<�^��o���*a��\����zљX���^����?4<�س;�s��:d�`={�CC1`Y���Z)z��MDe=��c�n8�?�s?�.?��B���~��XlJӫs:�?��n����O�KZ�d����U31y���3J�
�T%��$��9"�����H&����c(e���0 ���AEW|Ndp|����P 
�i��5`�r<��#�M-�2��=W�.�����w�����( )60J���#^�Uv�@H�(M�8�l�(�h="�Sȱz�S�[�4z�tXk�����=I�r/�)�9�p�0#J� �o��o��������yQ<�Ng��k����_��1GY�o{����\?�Hyf��{�r�5xq�K0���<	�`�s���y�y�]�(1=9�$
��cC�A@�O�G�@Φ�A9�xm@ ����܌�{NOO���
+Vm��q�dDF1#O�n+#v�gdU�&����1o���|��Wݐ�6�}�q�;d{v�
��B��jՠ���(�:k����{����r�3=^�^�:�}�b8Od����zc�1�]8��kqC� ��ix�O'X+v<ȄU_�2UySS'�����0p<��(����TH� p�����1�(-.�⧥�5�_D@O���ܢ'C���R�Y<cˣjV�> �P�i��;q���o橬���4�F�^}��2E8���%�l�3���6m�����íJQ-fq��`�����)}!��CmJa����b��+���ڎg�}q�W��ann&ǳ!��ξ[�J�;,L�x����q�V$�	]�=�ɿ�ï���9��������y�A���=�;�U�R�+k5-��9���y"��b�f�i�0w<�>���|�Z��
k��Z�
n�[����0��۰�yF#c'�@��ŋ뱩{��J 7�2���pY���`y _w�e����ed)u��g4X��@�4O�si��SB��g��r���}7<����~-v��n��
�X�[���!k7c~8<�Q`�S6��i�k�"��[��X�0KY�(�#p:0oa����h�BL@D��|���\�N��"���`���	�F��h6�R��4��[:��7�*V��)+9�#��kVPQx����̊"A
D�CA��V�Q�@�nZѫ�p\�V�'������[]��-*�Z̬�
`���ôЌ����֐�"�b)l^�󋋲Ty�Z~�P�������R�(�9?����MF��5�y��&���-�����P�����Z�x)�/J઒5-@C��$kIy���=�	����ow8�,1�jyF2���b(Z��w�M�ܵ���}�㠪�j�Ra��,8�?���G�v�X��Gl��N��iv3�:ˈ��N砤����l6x.@�p�?Yh��T��5�����+�jPp혵�=�v�Ѻ��1�Í��P��r�Ki�)�G/��y��!��y���d����A���j<�bL�D�V��)
5���c�P�	$�xpP
��	:;�!qq	b��>��M�⽲p�������c;�՜
�aN���i`�x;�zv���]xͲ&�=�(�S��`u;'��~	�Џ,e�H��yT ���:�\|5�Q��
�Dɠ@eJ��V�J���_/�%��*���)%�YB[��g�yu:?�PE����=�L�e��6���C�{!������ҌyaĚ�b�I����Q�T=�Y�7��ҕE�̓��	?��c����x�<��=R��A��ʘ�:ԁ}����K���"����}V��<�F�!�9� ��e��8Vu����X��O���m�v�� �n��w�\�Gcü���±�v���/5�W}�x��5���� ���(v+�2��ky�������v�8����������)���[zo�¿'m�,@��b��kæ>f�\|�ՃU276aa�jU�
�j��D����h�pW5��R�X,l򾱪�_���zVi�X��nq��M!���`��)=�}��F9�@m�f&OXi .��/D��Sh��螮�E��@#���|QG�k�*S�*�,��զ�q*�9����ɛ,e��m��;�D������"v���)��M+��{A*���'˞���NQ�oR����b���GE��x_�E�:X/BP�|GN�R'SG�S�'�R�j1NDy��!6J֯��xMp�FZI���EV����hR7�Eʇ���}5�)��ސ��Q
�7<%��p]��ĝ�_ۧ[���Y��X��	����7u��k)V���O>Go\�)�궜W+�Y���;_~��Q�"xU2��A�P��z����X�p�I�8yȦf��h<{otl�O�ѵ�[���=��9���h ���@����R���/��pn�G�n���%��+�28d;.}��~t��{�q�/�ff	tl,l�Ma��p�[�v�?��Nz[F���f�0�ʀß�?15i>������ٙ\�a�PQ.4��m"��o|�]WT�2�,�Y�p.Ulr�aA&��ȐMM#`��מ�b�i�}1�SV�E�()V'㪱{,,Zܩ[.8F�E��+�@l��(�=J3��L��������"}F�KiR�Bp�vJ��ІO��H	�t^��8H�C
�A�Y-R0e����|�@�E��\1�w�	
c�W�R���~��`������`�y���2�39硃G쑇w�.���*e{�?~�cSk���H�կD�Gw���"{��̯����mϣ��z���|�n?)��������>�1���
�5V������e�:�������O�/,:�w@>��OL7��)�mv�m��T-�{�1��I;r��a����t�^�5��K-���$7zPTp���C�R经��e�����=�����<[�9���m�}K_�re��d�uY�-7�Ɩ�&���m������&�����1[j�K9��˟�\$C�v�؃>ܫ�A��-��ԜW��߻/X���۾u�W���;qrʭ%pU Ua]���X�XTy�)���"J3:XLT�����qZi�܂�:2��`�dn}7X1mk461�p� ()�V\�7����J����к�BM��x�J�����R:x���/O3�FA��6+E(+���N{3��oY��W^�g_��)�df���*�:��C�Ǩb7e�1��
 ާr�c��CV��`-f<[ɕg�6�
�Յ���k��u?~�F�3�{ ���Η���V��}�/�ۺ�B�Fl��v�ȉȔ�U�
B\�v���b�����dT�Ѷz�ӥ�LƐ|����>�����F�e��I����^���UNi;kW<�Z_fG�ǵ�v���~�F���9�m�sX4XV�?�a����A��X_4W%��q�I{##hn&�2�����߽�A�������
��@���:	�em,�����^�:aِ���??��C^��7�´]tA��k�� �`�S�@l	�
�C��7��qA���H���(�B�ě���<(�{��R��|d8(� ؏��a���SRb>Jc�����?��n��\8�(�J�U,E����<�y�.���LA�³�÷�>���r*���&�0��۶^l/���Ju�9���q!��Zf#m�?�On�(���`�K�*V��T����v�R�g|��mlt�6l����똚8�{��ͷ\���ꫮ���"�C�'���͹3b�\j��¿k}�8*�&����{��?������k~��ʾ�m��w\7`��G����#I�t�����
���l��A,86A$gY,-|DiZ.k�J��yN�<<6��I���U���������d=kA	�J��XP�Ƿn��XZ�J��uKД�F ��k��De�G, /��18<�4&R��_�k��)�f1l��L 7͒b�Aq�7���]r��8��ķ����e�(��Q�U��K�}%�Pu 1!Ȩ�`�/:<K/��m[!^�f$�9d�ʒ�1��_���;�3]��& �Eߨ��}�?�Ǐ����g��Ipu)��`OWka�+3G�nt��k��=����l�5�7��-+�ݬ{.�<>OL��ۯ�{������Ïtء����=g;y������I�G�9�!;v�����ĭ(.鞠/��%C�u�����ұJ6��4��[�5�UF*x+/X�,�i��a(ȉ%��R
�-����*2�_�5kW�f&X)��
��9�aSԃ��n�*�����Tc7�蚗=��������4&� �A�PP��5(jkՙ`m�D��&댵�\�X�.��F��J�e}��N�=�¿�c���0K$�TZ#�t�K�{Zl��S\p^uv����d�n5�Q�r�@��g�'K�Y�1̼�pMk���.��r�`���Vm�ӵe�c����50�}�@'=/�����S��?�u.1>��G��j��P�4sQ��I��f� >���ڱ#��Ѓ��[c��68�6"�Yg������{����X���=����Y/��^��0{��ĉS���7�Nǃٺu�kjR�H�"O��*�͡^���ȌtNh�y��M#r~�|Xboy�[���H�� �U��1���
k��M�)<�x|��a�u��bFbN I��,�X�|~|���.@�X���0������ e@!$ș'��
�2߅v +{.��9>� ���M9\T_����W�@V�����C���J�5-�c@l((�c�߷϶���^�ĩ���^��AI�'�
H12*��^ĐY�V�����=�����͆�K�[τx=x�����F�!�c�p�����s��/X�6OTP]C��J�#����z��:�@���l٘�L����p�=�e���C�r�������l'�~E^1x��ȐkV�W�?��a�~���9�m�k9g?��MF&@ڶN�����]'+@�N,!�m���)�,k��+ћ8�ųe�6�eu(��G���7i����N�5�_*���`�Ȳmx����J/L�۰�y~�|e�Ɉm�u�Ќ�M��^N��6��5mө5�{� A^�q�7�<^���C�����\����<&�@��7�f� ��@)��0g�S�
���O�U��b���=�sq�*�3{�{1���"ݼ���k�>lr[��0s�T����g�Ůt1[�*�B�p�{�3���&v"��稩�~p���磔g�~�����>�E�r0�����h�2yj��aϊ|p`8��`?�8<��
�sS���Mr�dYɺa�@[1�փ���j���E�r�������1��Qx��%� iǔ�*��HpG�l��6���w�c{}�S0�cp�K�c;�J&L:9���4����k��a��!V�z�:�8���EN�ų�b��HM��5�����Kҁ��-9�T���lԱ����w��e�h�^_�җz���80�x�"���5��]�g
Ͳ�T�+Д���u�*�4�3����C���H�lWk��y�[�nS��P��b�K��xz�Vu��<n���*�p��u���T:��xN�� �r�ʼ�T���^�y�{�{�.�(��^�w�N�)^)|�Yz ���P'��[���%#�F�sb&-�/fe�N�fy�_�b(o�EΆ�J�5p~�a��}U*8'�PV���uc.|�+5��+�A[�b�M�<n3��
�����T��F����ٯ���K�D8 �`�KR����T ȿE�&����`����վ��3��,��CL@5(	������{�;�5���u�`�°��\`�:7�Tf�F��\�I�~+�o��H��b�9{�A�_�i��[���!�2�T�����#�S/GM
�R�c���m�2h'��AM�u�����}�7�tP��*�3��ꭺ����n�"M&sJɤ���(�L�������}V�>ޅ��� o��B�4�Rʷ��B�"��&�%�M��w�����:�H���q&&��Z
Mͳ�x���݂c��^��ѷ3�g�V�^^�Ƿr�/Y���
_�W�g��r��_�,�aQD �U�+�Y���`}i
�x�u���f�ȏ��.<Y2�87q+���y>G�&s��L�}Z����������x-�̤>~�K�8���ڧ��e���]�:Ԥ�R(+A��	�P
���v�N�H!�L��lN�c�O��{:7= D�!�������E�O���7��_8�D����WK6O��0����yZ}��7��]b8S��X@,l�XNlB�(cH�/�>�g�8�ڝ�X���d��˙k�ͨ4��Ջ�Ƿ|�x1��@(L��Z-�9.�X΂!����W��pf	
�S,��ǎ�m����>���ń��k�����W�5}z�}�Mp��H��~��6^A ��@U��b�]�X��&p>C!��Q'/)��A,�Ua�|�T�(/��N%bX7p;�X��r�t��WD*Z�V��ͨ�ݓ�#6T�g�gڍ�^,+R�g�z��ݷ�H���߽UZּ%�P����t�z�_xB����|"i�����v��t*	_̕�,
����S�8��#v�P,D#�'6���I2O<�y
�,��<��m=�U#��ֿX31��h� B@�����x"|�|��e�� %��Y�+_��(��k�@���Y�{<a��+6!��6�|��VsQ@$�b�s.���!
׈��us}�n�����Ҍs��-K;3��GOZ������И՛���NKy�q_f��ќ��p$U���PBJWr�C��!�o��}��3K|���z�U\Z����Xe����HcbStr��f@���g����]�}�6[�SCT�5��>u�U1����6�)n�~�Db=G�f����0����!�	��u�]��?��?��yV[f��8�)�|:r���g�������:��Fŋ�,9��S`]#�	�-N@��MQbc哵�<$������ �`�������z!c;B�Nk{���hp�?�����;.��1}����=�R�
̺1�윘f��+���b�ǐ�#��Wa1͢��su��q?g����ȫi{č�ajh�*�Gd`��Pڨ�r^�q�[/\3X�O�ɩ��lLY�B5�y&C'�T�f�K����dXv���v�����������3��e�,TQ!���:R� �bS*R���pLΑz��-b7Q���[�kJ{�w�J��G����`G��Ҥŭ��BOEe =~�u��.�0�V'B�@si6;�6u����e60X�L��R����S��~�=��RA�������k�57bY�w�l�'����	�?װ���,��h����قֆ]�*%��!KFCʡ�i�����ڀ9�s�C�Ϯ/^���<�Y]7?f�0�Ώo�L	Q`���N����4ax|�C#ܜ����E�	^��#G���NT��GP7�L9.1+�C1CF|_�\���W���wߝ[�@TdqM�3S9�������A�F�+H=Uj��STM�E��t%��Ub_��`FE^�j^��ʱ~Wῢ_o�K������HcnE'Xd.�ã63W咳��ߙ�H�j��ɫ����N>�؇� Lɍ�?U��-��ۨp��[��0SL^V:̅w��OG��H����O�)O�,����}Ѻk�x� �
�B���Y�D�um�`�5\Ѵ��ULS��� �v���S��Vp$�oz�0���9�$2|=�,�_���9�r*X�_�S����y��A>�&�K �}@�Z�~�&c���d��yۮGq�PO`�� HU%��'q��a���"�H��b��z� �S:���ؗ�={zF2rZ�R?|���޵?Ҡt#����%��2`'NM؇>�1�[+q�r)ҳ��xj70�HNq���8�����kg2�S�]�W�-�ʧOg�*F�`۳^�zV���ز����L�X���l�b�\�X��Y�~]�y&n��CG\H�2m�~�r�����Gg��I�+���f+V(f����>� �o�^8ǅ��Ӷ�SǬ7PX0��N=��<}�X-x�j^㪻���ȩr{�4�$��M�et]�0�|��G�A������w<'�Y��H���� 8��n�B�N˶|�����/��҃8�T��� hUg�⫵���	��ˮ
U�9E^E���[n����҅#��������Kw,踆��ګ���^��<�)pn?CŇ��87^FJO�2>�q�t#́��S�/�#|�68j�����ÐPQ��������V'�g�M��Zu`>�P�j+8w��}�R/8�\��G%�u�!���2��G<@�j�1[Y<�kE)׃bf���E6��l�+J��7��g��/�������lm�-8�7�!�O��v�~}�T(	��8(���]Ps��AҎR�"�Ry�ί�"�Bvn��e���v�ѱ����63q�]ڊpڠ�����v��1�7Z��o!.��OC�~��2t}*����L�I$����jCҴ]�wޙ	^X��)e�T�3p����%Av��AoX���sX�@5�a�"`��w�ݟ�����?T��^���G��H��X�R��<� U ��Dv��Ӵh-�����xq����+����Z9�^.e��ю�9/�(��p��XYO��� F�������U�G��������>+���Ӿ@�(�;�V���W\��Ä�����{<��޻��yH�����Ԟ��:��'�Q�S�*�p�c��\�dd�^������	њ��K����6�zԖ���۷�'?���O�J�E�+���,���jv&�h�������~�� F��ќsvy�x���#v|�DX(4np��J����-"aQ�pN8��eC�Ñ�/���,n�w~<�!.~�������� G=��D�),�!/(��5��Y���<DV���])"Y�b��wxM���f��*૶�i���֑��hX�Bܣ[�;y�n-�:�Pj�~�]s�e��m�;
�v���ܲek�˷#)�"B1#���6��R��ѭr�s��
��`+3Ii���]��ee�n��Y�������;^���	�j4Ȣ[�n�]{�u��ؾ��/�}��i���a�I���^�{D��۞�^�^Y\���ӮZ�?3;ִ=t؎�<�^��Uk���>P# �����0H��{���ܕ�7X��>��O{���:�&���`��Z��ێa,��R��������U�"�x'+Z���w� �W��I.�b"K-��z�<e�S���^N�x^��d�H����~��7k�կ~�c�<?�J��@a�b�s^�5�)PSz֥:�!�H�T�#�X ����Z���Utυ,.E@�F���9׀' ,�aD��9�3V��?�)�Mk�i�,CZ�Qw�(f����Ms���l�����٘v��z��s��@�o�{,��(OJ��w-S������x�N瀋��	o�>�Т�
^��V�U\�ƾ��_��_��m0����U�7sYr���z����.��U�9v�O�S'�z���������}�P 2<4jW^y��t�-62�<�Ղ=�Y��Ŋ++���@Ѝ�����@�
�Op�~}���h�z�С����o�ӥz�A�"��l�s��^���^@7���\�;��3�"DbKq?��lY{jB�TF��.E����xr��M��`�eRk{��g�D	M��q8���{�oe舁�2(�3����Ӆ;B
c��Y�<w�8�a�C���j_P�b�NF� �C���"@�F
�O<asF��c��I����7�r�l�!Q�_��p��o���N���Vl��Q+6P�ᆗU�
h��Uʶ�.{�*k�>�2��̝���E����a�L��=�;�p�a�^{������g�|����m;l����-ۂ2\m������c�֌�ٛg����Ӈ��z�_����ş?��˯�ʞq�Mv��^���G�O���/�q�gT�6�d'�����^��9��%�@)da��*'X�����������{(ɮ�\x�[�s����F3#�r@�H��g�c��f9��᷍��l�1^^��<�m9'EF9k�&O��t��|���s�ۧk���i�3u��=]U7�{Ύ��6�<����je���Mo���IY�Rs�̝�d͊3L�U��et�������?�	xu1Sis Kt����o���`�ca�} 3ȹBW�
�=?�%�aB_�(���H�Q�.J���C"B�j@��ר0� A�
���8����y��F
! ��~���8g2?���*��_+}q]8<R�EeP0`�1��4X�^�O�Z ��������Bޜ\���n��f�sޠB�O-�N#tC���4��L�RN8�@�2U7b8�f!N8-�\G�n�e���O�s�(;�C�w0�Z{ը&O=��<��C�k�.��^�z@
ټK#r�����]���x�,Y�'���Q�������cn<Щ/��z�����JcґO�����X���e|b�P4�5K�Y�bqT���?��O��x���C��&�Nc��R��8L��$�Fֱk��X��C�����=%�܀���C��<��~�;9�6�ɪ%G�`4�^,�-@lѕ�H�
g
v'�5���k������=7�	�P1���;`�d!a���I��*]��� ���� � X��
�TL��H����9�]<�&X�P$x���964�EL����E�Dx��H 7���Nd,�b�sa����f��`դ�W�y�j�G����Xo{:�^'}�+͍���l\�Z�5V����`�5,6�D5�>�A�HO�ׅ(����6��R�A��1��wE��j�T+#�����HWg�Tj�תқM�T�.G����?�o򋷾NV�� �V�4E�o߷�Y�/£�4������4�X2`M���әH|�ټI'z�2ٻ���.�0g� d�'&�TQDr�h�/49�%,X���〛qO,v4u�{���bs���l� �U�������\WW��s]R�M��A�KJ�c�D8�U�E
n��K�5
8�t� ���%*��%� �c��AE�nPldN`C7��P�q~���a�@���j@b�x6pg��W<8'�)�>1�sM�"�����H$*$|��̑����)�	�m�b�i�G^S��Ϫ�*�CU��Ra�,{x��}Kep`��������S*X��Bz#n����Z+Y̽\.�1\�=z�GO ����U��ɸn|�P�z�>���^�v�^GE&ը�zGw��G��d�X�cE�_��l���39s�F��{���q-�)/�-�6��BQ+�V�IOW�.��F��$��QT+n�Z����,��`��,-kzՄ!����P:q�:��Z�܍ՔH����w�i�6�&Zp�4'�[J�$"��jm*!��u����ez�hm�|,a��.X��Wb����,m5�^ ������sI�8�/x��$�&�V3>%�����B4�����}�vZ�Q�!��i���W,�����J�|�FXc^ ����������a(�C�^=6��v|� �C�^j��](��ߧ7�VZ��Ĥ|�d�����T��	|��޺�e+�������·�#�x1w0���IÍgxp�n��s�:�3���ۗx�&9
������y�]�s���M�����c�V�ϼ��Z�S_��3�< &���C����
�:�L6�`�@b�V�,Zj�<>�)��vx����}���l������©N[s��UX�P�\-
�x�FT�D0
x:���E��~*0�7��ix�e��!Y,~��7(YI�CқL�m�ϳ;��v p��b!+�ɷ��h,�:E��!Zm��S��}�����>R�gx\��a ���&�}( �����8��7�zQ��(�ώv��U%1X��~�a{���G 
��f�}	�j��`�խ�5�=��-�S�խiz�܂��
����rV��� k^@���?�cy�[�j�-6�G.�=(?��֮6��e8�
:�!
J.�1T!
��+�*Γ���Ge��{�
��x)����@��#)W���V���|.)�w�>��^�x`���QmG��.'����Q�X9ࡀ��ݿ�8���˧��8>��J"[�#��ȡ]r����EK��j��Er
��"RQ��"�T�z��p�� ��A����	D�A��ˎ�c���T���2�7x>��b<|�B����]�Uxn�,~"�$�'����r�}?Nx����Yx�n�v�f  �K����
}	��N!\#'z�8P>���:������nB����?C��D�W*��K��uOEe��2���C��t�%|����6�~$�VUϿZ	�=��S��;�}�{���pohbO����"e�'=8���f;���T���CϛM �$��>�1'�*�(F�FOθ�f1���9�S^��4s��ɴn�j��X��8��o&r\aUh��x�u]p��@�,����x��K�\p@䰘QJ�67-Y=����=\5i�8�o�^ߤdԺ��"g��8H�X}GӖ�v�K`���0g1�5v\�\�>�*?XC��;=dȇ������=IZ�P\|nx�a�@��eX��C�/��&(4d�� � ���%+������u�p�����Q�Qt�B�v֔�|w�}��
��q���ճ���o��8��)����Uu	t�E"jm�z_wv�˹[/�J��*�T���O��_�.)���@٤Ru?���½c�c[%naZ~���?�01o].�V��~	5��ať*R*oV�[#Se��Z/����i��~�m�w�AV7+~���~�*[�H���'�L�w�v�Ly)tvYy�Χ��2v��i�+҈��G������w�y���w��][����f� !� �a��tv�?2�o�BKf�4�Ua��EO��?��B\x8����Z����`����2QeT�~�C>�>�n��,ߘr�J�g���b�����Ig@4
�:�g�BKPX�;P�q����hL��a�T�����60M�F�9i�wS��EE �z&e�8�9���U'`1���H�m=2�����,�G  ȥ ��#���!�t�2Y�j��Ke5�ft�ܪ��7�vmM���5�\��A�H��}�z !^.��������X��v���-MUd��{e�sd|�\x����'d|�l�7����V������(H\��7�� ����E ��<������q`M����z�굌��ş�2z��1�4T�hp]�J.Hjűw�q�.o6\u�<|�zX�،p����I\��'6:��yv����ρ
�O��sD��B���0D����������v[�x�X,#�^*��|����W��(8*&�휺�p����w��@���>�)�V(BDØ�g�ٱږl��
���˩�V��=�#vC�����C���0%z(#B��q���l+a��6{`I�Ž!���G>��%�5p�}�c�R��m�](���P�ꀾ� �Ī�e�Y��[&�;�-�$j	�=���
��?�8����s���A6�K�bz?�C���iY�f����*��2tx���&&F�d,�.Hhn�z��u��$<?b�L�b��� ��͞������&]w, +��?�����~N]��y�.�$��8Ir��K�\i�yZCjX�ӷ1/�5�����p�c�(6g5j;����$.��a�ǯ�3���%a>O˟�B�,c�8�6"餱|��iE`�g
��(?���{���!A���Y?�����-�F/�`���U}�X=�%r�Tn�}p�O�Tq����L�#\w�QC�� �_��_J��0ҡ�$l֧� 4��u���Kj��a��AȝBΘ�׆36�5��h�ò����C�䓻��-���Fr�q���uq��>�e3/�FY��? _����u��U�rM]���iG<p׮r��ak�GͰ^��Ns)�q�C��p<��|�3�7�Ɋd �#�V�+^�
��W�l^+�i]�ӗO�v|R'��dCv=�CjU��֝��@>+�5���E-�T:�����Xp+�%��'(F�W�p�P���'��yQ��µ6����0"�Ճ9gXe����e2lCd�X��7C/[�Z�:��q|&*B;1��҇g�d-�E ���Bx#�okk�81i��By��l��R@�*Ž�F�#m\�į �݃Ec#�q���ڄd<�1�E:e׳~
4϶XQ��������A��0�BD(��Ї>��ϸ�gp�DZ]�{�!�6�����J]��d��@�����<8j�����l�v�z,��� %�m�}�d��5�i(x�q��V#p�bb�(����N)td�%/y��k9Ier�eW�Y��&IN6��*�U�����1w�?�c8tP����ֹ���k���H�R�����k������X��Q���]ۤ�_j�Ѓw�#�X*�:�gƅ��J@%�d�.�?�.�@�a�<����r���ܡ��pNl �5躓��վ�L����7��S����?���~׬Z]S�@y& Q�=6z̅�j�%䦳7ʅl3c�;`�j(�񊅐�� &�>rԎ�Y�0�rd�����{l=�
7(�8��EBki��a����V����P 𤡸 ��}�8�����Xƫ�Є�f��ի��[��FR>�����è��F�[^�R�3%5�r�K�������ռ�`<��/���y9�c�~�<����84��+��I.[-����\�(�~��!�c`rtJ>����C�<x\�x�(l���s�J���}�0�x0�L���p��T&�~��񉒹��t`�@�����pb�@� ɋ��x<,�~c��*!��.#,�|v&_���6���ŴI7hd! @��
S
�C���,,*�zc���D�c���  �ň\Y+`�!,�{D����m�/n�ه�an���<��>{H�;M�	�i�3��:,rҋ�w�e��_�m�ug�  q���7|���Hр�`]�<�'�>�{"�k�9(!��\ӣ���v`|8+W,�m�oAה��!�`�aF&U�wu�[���j7xwu0���$���ɸ�g쇛~��O~��	����J���M@�Q �	��,�[�J���$U,tv�cO<n��@A��!_0׋Aӝ��?��e؇}E��"��K�я~Ԅ?�
؜�dY��H� Ə���b3zǬ>,�?��?�ςW�f�|�4��bq�����gB��⛵:�B�T�'Tk	-��h�`Ψ�Q��m��CH���j���.�s/ ,0Z��� H�`�ạ�|b7Ɗ�����i|ZgZ�0&��� 7���7�O饢0	��[�����ǏkA��A��w�wm���_��	i6H��>��4��:X5�A�c���뿶�!��ϡ�PQ;T���&[�c���9���i�5b�sd^���p*�^�Z������\���s��z�"�^�|Y�|�]���S���j�Q����|����8��q����D����d��/����b��)/��d#$d.2�Ҙ`,>L>�U0�c��7,J��ȊȒo�ƳM#�}>�O��C�~��`�����;?��D]E��=$��b�r�@#�nD�"����C��Q5��mm9���h%B�����_h����{��d
d��j���XD^��/��`g)���>�|����h���a�\ ��{�]���a,����`������8'�C�<�������ll�C>�=7�R�,�FՅ�@��ϲ�{�T�޾���⹌�=��F	��� �R�*ܔz���?���9E�0����������=<G(W��^ �'�7�1�02�9������:��|�5~r��˰i�4�7��eec���Y���������0��I��k0�E�&�	�釞����EuH�<��s��0���Ca�L���U��2��m�ԋ��&|��ZG�o������m����Hos�~��o�+��aeb�A�����p,��/�.,�w��]	���!�������c���#$�Bˇz�ӦWɦG����i���<����M���Y=�U�@���7��ֿg���۴Y���K��[R���*�S���64�JK-UK���~��Y�HH�sG�������C���O����-���bIVi3�@�EzrW ��S^��7�Z�/Fg��������d�9��O���,6,�>�$P��d �Gr�%����o��L��:J�;��뒎�ZS�qݼ�p�k�}#���:�7��!��	��[�J ���Φ����>.��8�AC�\�X#C2n����7���a"EaϺV���%��3Ɍc5�c��B�'`�1@t�F�*����A�ǳR����'���w�Q��f?3�Dm�r��V�4�����m�:�+ӎ�>�0}d���������w[��Ph��½HXã�L���C��DC
���3f(��c���c��b�i/�1�L\{̰�9>���
�Ho��\�x�X�
��P ���U���[� V5?ϟ�l��l}���oTC)N�%�B��KnNʕI��fBG�4R�ؑ�ſӨ��F����n��D-�b!j��LaDWߧh�����rV���X}�(r�P �*��q\*,����J���P��	M�@������@1�G\��J��%��ҟ�]7Ce� <�??�R肇�ew��fA��y�汦,\j�9�_��P��q��=�1�"(?�opݸ�}�c���7�5��"�3�O���lY$��>�~=A+l�?N_��<��R�\Z�\d~۷Z���9c�<-��H�!��W.x,j|�)3�˦|�87,�Z�YS�	� ��e�?��q�wa'�L�l���j(�0� �AT!�,F�i9?l��>e,�n?&;�:k��(��!�?��}( h�0�DCk�	��6\��!b�T4P��nR�!1��3�l��ռG�Q��8��CD>�r����Hv�V���!��c�L�d��P8a���֫�7���q�?�9~��=����?��$J���L`ؓρ�<�$������<��fΆ������Nߘ�|�_�>'6�o��	�kCDxDJPX�'j  �a ���[@̵i�$�oq̮�&�՛����~�)�nE
9wO�c��6E��[D���,��FvōG+�����s��%�[t�3n���R{,l�����/���6��/0(�0����g���}�LBC�x��|H?��?�Z�~�����ѐ	F�/s]��ܵ.\�а��Z��n�\V�"0@�{F�����2�t�q�)��2K��h�^)ǐ�ؓͪ�E�\<Yw]4����	��g��)�i(����7&������':N{����;���VN�oՐۃ
�V�����	��l��e�p� I?"�=�S��Q� ��PO���ftb�^�D�T���F����9c���;�q2G�e��o�QPxFC̅w�1��\���;(MT�T��F���#�?$�HoϠ�^�A�U5�O(N��%��f��	z�T�����"bh�ъ��|N�"�@Z�E���IfB&9�,�ހ��i��!Z/P���s����T*�w�voeA7����r��n]��DTܗ���V��Cf�l����� �Q7��@7�Q6��+Z~�M{<W��kQ-q���ټL�F����K��ua�Fv���9cI^�74tHB$��h�3�O�"�3iT��4ʡ�-�8��a蘈?�C3ĕ��Ӝ�8��|��ӧn�`�#Q+��LK����f��|r�3yǇ��{<�}����ύ�$�,����T&[z�r�H9��(t��
c��b@Ӏ|�]}�cm��8�cv#��]����n���o88rW�Z:���V�e]]0ҜYŔ�4 %p�l���}�*x��"F߈�	^�b�:��̣�8i���"=�٨���4����  ޘ-.��Td8�w�h��°-v��|<.CA�|~a?��\�KK�_�R�ԪGb\+Y �b��Ѐ�Ti��LUʒ�,>ZE�_��u� �'���Ӷ���6f�I��v�t���)[S&4a�u>U�X�s���|Q[H��ܴ�vh��˷�����'8� �a�Ic�0�I �oȠtj�{��TP �L�_?Q�[��<O'2Ny�?''r<U���3���	.�����Xt�(�}aތv���Wr0���#�J�xD��k�f\%��
�TC,�+99U�kba������7Bc\�f��Ԙl&������h��5Z�HrhX�rprj�5H䆇G��Iވ���d�*Z.�^�W\_$v��'KR����d&�l͠��p�&�g�f�0����~Q��_X���F���?�8��f��%N�D
pChd�3�A�؊�������a�M<N
O�]��Dt��&u����bh)���D[��{��T,�F(�uߨ98_�~�]����I4��26Q�#G'��k��ϿVV�X�\/��M��'{�Ʊ1�T��w:�����ό�J��zcK]��K�O�I�Z3�P+�Z�
��:T�ҥY�'P�����U2Ĝ+:K��x���]�`}�^����V�Npq�fU��F�m˿����� T��1�6�\�p��er��73X��&�7M����y��կqpb��)Q�ҝcl��u�`Xv�6�Å!:ؔ��y����ʰD�8��1��;��T2k��U��C����%/�ŘH��5��7�~'�W�q<܁Mb���dE��>�d!�	��A�h��Ȯ��Lޗ��I1P�g�t�������6湟�;��u����毙�ol�56wMM�y�Ӵ���<���6&*����<�Y�ef/^����Le�4,z��Ҥ|���_��~/e��W�6?�/��[�o�Z1A福u?�@��1�f(�����8P��`�.�#�����d�gZ!�o�:����ϒ+.�\���oX%1��(�:����x�Є�iZ] ������U����'�z����1{9�r �=}�d`�Y��=�׼V�{�L	�(+��u�Ԫ�U���#�
�Ը�FG��L�wMi�Fdx��f#2%e���;W�V��b���d�X��K�����G��^3���
�f:���2��%�Gk@@4*��<���(x;���T��3�!�V�7{���ǧ�f3�ڨV�,�0��,��V�..�!"q>���n�.m>%g^Ohg�3FH�7�����$��$�%J�e�&��I��H�V^q򨤲*X¼Y��;0��E�S.H�����y�����y�E�P�J�)r�/Z���@��@?�D=Bz@�`/�3�Z�l\n&�c�PF?�FG9mI}�&�׆�J@�����u��<Fz��?�����"_E�������Ƌ��c J�JY3p��L��z,E��V�?,GF�4b��.3�4�'��(X����Z���L[��D������7��g2Xc�$��|�͇tC	ԬaRl��=i^X3���X�˰k!�]������(��aPV6tx�>�d�R��R��Ȧ�Ζ�k�[�� ��ߡ1�N�E��E^QԂ��r�
\;����*��ꄏZ��O���k�����I���/�X�ٲU��XeM���j�`e� �h�fO,�׽�u��YD���ˇM��D��d�"����0b�ȬE�o�,��}��45i:������czh>��kL�h�!�'%&TL(�@d�d:�_u�?2��@������4Bm���7��u��b�/�G7r���w�h/��y����HP��JkB�}&��#'\U���&�èG@��g2ܚm4 �.���\�}P3u`-��}���~?��*��ç�-���	BrhP
�j�|̏��X�7l��Q�h��dVn΄P�2���Ϫ������ร�_��-�E�Е+_M�=�x��GT���8~E�F�u0.�鄷	^���GS�h�X�O+Q*��8�c��T��p����}g�/���(�}�1t�1�U����T'z0'&N����ȇE�?�}��(䬝㱣#*�'�|\�������q�9r�ŗ��3j����?޾=!������u:7po阡�I� [��u�\�|��pJr�H���%w��=����K�汪�h�����^����L}@Xl7�|�qsӊ�5 �>r�B�;���<����_�z����[,c�� oj�+����Mق���"I�b¬h4��E����&������|�=��A��t#����ZY��U�(̙�`a3��1��V]qI�zL��n8P��YG��7h՗a�=4�?	��x�e���sq3�,��~���5,����F�	�Oڊ�,~��±��	Ⱖ�جi"OƦ/tmQ���҈��A6gE;
�nK����������R��G�� U�j���5m�tʅ$Cԩ��~=����P�t��$���g�W�<AJ�����v���,O^#�a���$�3��E�Y�<f��;N83��0%Qz����Y�C���k�5FS�����@oP���������߃�����7!{�<!�|ر�I+P��p�9,O��>����] ��Ke͚U�8��'w<������I�)/�[�}�[M��<O7�9��f�c�%���[�˭��"F8:<l�����_Z���{�g�a���2��6l��.���P�o����Qs�����o���a���d%8O���>� ��:�ıZ`Q�*�'�N�B�gI�,�����QF�$�Z��W��I��.����P�V���<��*��n�JY��B��9"ׂ̡�G+�!�{� �Z��j2�|H�S�:�[��j}DJ�q��(�5e���;oT��Vc�!��]X�8_Ը�(;u�"�%�!�jჷV�U��KO�R����E�*m��N��`mG�0�9*�ָ�U^�q�:�*@Gꗊ��Gus#�l�r΀���V%�����U3�d�ff
�|>Ãa��-�Vፐ_:t�j�ٺ9NVV��6���
��e�u��ީVc~��ǯWFr-�����Y��>��"��L�����`���"��_��������@��=����j܌���!��I]�����3��(�՛�*���-�7��笁;d���0W��
~�S^�����q�s&��͛�ڄ���ʷ��e�ֳ�uk����	�6fdl|B����	�y�u�]g� x�Gy$�h�F̎�V�h,�p��2f�����2�(�}S*�U�,D"�j�J�B4�=I�f�E+{���M��5 �j:���F�4�.<�r���g�/��Jy��+׮P!1�B<vC�p^�:@���ty�*���q����խ���C~�
��� E{��321Z6�epi���,Q-���+��v=.���p�K�8�B;+K���a�H��UUL��0p���T,)it˝j�g����#�^�#�s�'���/�;������REcޢ�wthJ���άtvAY�1<�I��g6�#E}��[��u�ͥ��)�� ϰ&��f&k��,��nTu9z����O�9<t����N��~,������cR���r>��I{,�1`U}cF�k_l����8b.�Ǽ�����n�[ �B���z�{�k�;�������=�\�T����񈮑��Y�D��)kh?Uv��K��������;�'+V���/���m�'���>�ih�e�<兿��� ���U�;�Q�������q:\(&�l-�p��B�S-�1k�v�-��%�Nm�����	�^ U��݋�/��/��@7%߭$wG3�ۉ�f:�f��E��I�m�ΕMg�։�������*�.�_7�V��@U��C�F�;������b�'��R#�.�ۈ�#uRy+V{��G��w���뮽J��ҮQ7�5��Z�D�#�������wn����u�Y�e�:U&�di����*��>V�o�^��(ʍ�]%}��t�۰�W#���kBqa�'Z&Ǝɒ%r��W�v^ ���\�>�HY�ꍤ��Bjt����#�ߴ������*.T���W���[=� �8�s5>V�o|�G��^p��?�i�/��!��IC�c�׳����m�,W^u���Y�9���	�F��R1���}Xʓr��[d��:?u����[�}ʱ��7��GF�^���K����<��E�����0���V��O2|�B�������~�+v.th����Д �������#r9C�航���xTe�r�?��q:R��2/}�K���蓣:Gw��r�%W�~h�ʕ�������f$���k1Ny�ߒ�'r�-Xh��Uj�8p�ڿ�P��֩��::T"n��*�qO
ZZ"����H%
��;�y�?��/ؿ	�d���\�6�
�|/c�O3���#maX)(�)�&�,*��zք�6>Si | lr����VQ��ch��k��"��Q�o���@Za������MB�%��e�S1���ʢ�	ز*�@/���`��-��p�f�︡�
�M)XE����q��B!{p���Y�5w��]C e@��oOA����Gz�s"��a�,C�j��u�A��~�
���B��Tծ6�BөF$��6�8!�Qu�"2�IxO�������Kh�fG��(���e3h2��zQY��	bNcsGx����p�0����@	�z���Hf��q��b�q3RH���kD������F$�eMJ6������L( �u���
�9��!t!C�^�7 �@����/����jҮbxl|D��R}�i[��a��	�$��󙔮�kk�DgGo���:�q����o;�����Y��h��8D���ߑ�!>��x8��@1��o�����P2l���|/����Ic4[K��ɒd�ŵk�yF9�؂��'"5WSV6m(���+"6mEh%�w ��<F�v�C@�@�{�X]��Z��[,��>+��Q$�1��	,$N+�)��ͨ�"1�#�آ�N@:�G�a��į��\�ؘ�rQ�6*��UХ$��}�*$�E*v�Z�b�]U,���M�EU�����nT$V 4K����ҁU7!�S��͍����`���K��T�~�
�|���ME�Y�Q�nM|`������*�lƞc��C��)�C�-}h�':ȕJS�iK�?_���3H�\�F�"�i�0��.Yh{*c���ײ�D�I�;K�B'��b�'
}�A`�{�{����ޒ��?��^�*���lﳾ�͎X=��Z2��^!��kA-i�$���&��,��`^\�:��n�2��3P�Tͪ&�R)���>�.�	F��	���v+�5	:eCnQb��+-g%=<�^z������7-.�������/}�K���`˾���}�9Z:���9�9Z)��,�kp/q�˨��E��*��:W�Ѕ�`� �Ě���3b��#��Аad �g"V["^\6��x,���5�Q�)�@b��0F��s�H��0��$���g�TW��6��nө72U���В�����d�D���x��A�ϪL��.�	(�sʚ�l?D筼���E�(��'	q�!Y=^�����2錛�c*劕j��	{�~Y�5m	_�S�u��z�����\C)�)���=8�qEP�_#w�$�[�<s-�~�O��a�Cj��:m�P�r�����Fw�>!�Hp߰�Br�gfM��c�Ν������oΫ����q���8�RdH�l��F�*U5�
�NWcr``�<f����=.'�E?����?�@U`GgA�����Kz�j���V�[�{���Y#���L��DE��V����6����^ ,�������K��+���|�#����\@$��U�ܠz�6}͌��۳5��������B�)uOIU���`�Y*X�CG�&�!���F"��F�j9v���\�g �[�`�a�NQ֡�fE̽��N����D�����>��g��ʆH*������g����1�u�������]����%a������5�Vv���W��UG��r�p��BcYU�cG�z�D/�`�����16Z���^��;t�����|%e-���hk�3��8����
Wmj�Gz�X��$�#g)�JU+�����̑#Cv{� B38�SQ������U��l~�z-׀�9S^z�\u�T&&;,��/��B������wK?��Sjh��W�hG�L�2#'��ǖ�+����q��gn=�Ċ�0�^��D w��;��p��� ��?k�~���uk7ȡ�g���V�����n���~����I)�|��[^���zpL'ͫX�8�$�%aN��54я�s�v��7�+�-W_�y��{���.��]�K,|�u�u�M[Wv�aX�F�W낯�ӟ����P7�t���o���0�~s�"7�$�o��o���E鉺-� p���b���˖���:Y�|�)��v>)�?-S��%E��EY+r��`�2Y�~��%�?�^FT��ԣ���c,�L�
�^������;e��5�v��1cC>�o�ZS%#��d:,�X�5 �*��'�fQ-[�Tϻ֊���{Z���%�)�\R9C� {_l7��8,��@��߰BV�Z/�� ���'ǆ����,T�kjD����������2A�D歹�T �-Y�v>*��~R�"ٲ%�%U�L>�)� B�%�ӻB֯9[ϻN��1����U>�T����K>�ڂ�)���\��Ⱥ���Ы����?�C�ј���p���R4�����}:��e�ʵ����d����Ԩ	�P�	sVL('t��Pa?�B�]+T���9����^��\6{MHDW��؈��4k�DӍ��j�}�8��1�.��ϱc�~��_��_���E�@����Rٹ�aٷ��Շt��V+��;��e��~y��'u�����,�F��@~ͼQim�EQx��}��#
m��bR�㮻�˥_&�j�#q�~�9rdhL���'�ʭ�1n�p�W˦�ےb�{��\>Ұ����`�����|�k_��Sf��1��s5��q�-�GN|D�C=!6�I�Z�Thde�곥�g�
�N�9��aCڬ��#G��sm�����L�����9c�f�����W�궚
c��Cf����X��D��2��@ϹV֮ۨ�YH�3Ղ�{߯
V��%��q�����w��sW��X-����JU��U9��rŹ�, ��^��N���M�.TA![P�Vz�d�؈^g�u���oZYU+W�wْ�r��3�"�ϓ�*��� @�*F��Qv�O*g�w����z7���*A���;/��R�Z������Wb�@1V��~�w�Z�)Y��G�?'?�~�
"�ʺ�v�zC׬�?��/���v�U��4 1ͫE�~c�����x<nq��-8�A� }Fh�۷\�:{�z =�,;{d�*���wD�1m��P�5Pn4�T��I����ǯ�hQ+Xf���]�z�z���~�����Χ���5�y�����}�3 ��[���!� $���սT���(���W	dr��Tv��~�U��s�7�h�Ȱ
�$\dJ��1:s�Q�Mҭ��#�������E/ԍ���^)W\q�Z~=�l���[�����.6K�/~�f���H�7��|�r�ԧ>eP:|�w~�w���a[��,�&�n!h.6���.���A�U�ꆯ��4fbq�n������.��YQV�ZŹ��~��4\��b��,��IIO�r�n�ֈɺ ��(O��c!�jC�Z�pܜ�TEܻ_��B-�^�2��M�b�UƻU��ˤ����T������Wk+��2���:u�;:���c&�sªY��l�*1�x����kM�@L��V]�� ����4mJ�����0�TC�W��֯�"#c���ڛD�4��F̀M���):O%��"�*�^�R\����H�`���z�=�dD�j�58�ӈg;Σ�s��J��Y��jYv�K�=�d�>��S%QO�1�U�T�w}E.o��z���Md�h�=�R�3�@�!��3:��~���X�L�
�Azy��y��F��Ac���%�F��<�P"�x��<�b�WR��q��Ss�2,tp}϶��ׂ�IՀC�����?���z��PBr�礝��<~Ȋ׼���[��,]��y���}�?�Ò����r�5�ɖsϓ��X���>�_�)����e�����?j%�<��U�� G�O"����)/��Fc�V���kn0aE�Sk'�ﰅ`t�z� �	d�X�@�� �9T��;��~�#y���-+W��!@iU,􁲦�O�2>Y_��X��<��,�zF^���e_'�ͤU�Bh�^��
��7�u����׾c������j��q�*���U2e�6�I�KRQ����m��yz�nٳg�\r�r����E��`�U`���{���&J�Id�����˱�1y�^��?_�EQ�mJ��
�@�W��MDQά�~���^��]�����ea�[o�U�٣Ϸd��(*������yq��n9g�6����S;���[/���&Y�r�Z��l��.[c��)��`�U��7�\6o�P��|�;ߖ��k����s6� �2B2��&�`EYl��h�֨�c�paC��?���ۥ�җ�D��id�t�B����*r5j��]{�z]c��#����9�\ 7��")輢�"�Ϲϫ�����R]��.ٲ�K�~�K_�b��oy�іXD�i��_��z��]��D�r	�^Bk�C?�ӞY��î}&@�R ,�\�
}�pѡ�:��S����ȵE��>X`����@fpO���� Q���A��k��P���s�̳Αo�9�������iN��d�$w�u��w�vɫq�~�1��g�o��=MNy�H+Ӡ�����y)����|�2Zg�;� �����N��z��g�����.��� ��g�/$w�	�C�ŀ�x�Ï>��lC�a,Z�-��8��%��	�@����Y#֟c��� �DW�j9��F������r>2<)˗ʹ[/�u�W� ,��ZX�g���Q��t�jA����19phH��v�
��,TS�ؽ
�2b��4�,H��D5�9����e�X��.�B�ظV��}��rV��87��0��eЩ2��Uo�wTWJ�l��X��b �ƘP:��0|Y��2}�y��'Գ�+�ܢ�|�����Vv=�A�!��"Jg����S�6WeAP6��@t��X�X(-g�EC(�]w�t� -�>�J����BY��K�QŠ�H2#4�0�Td��U�۷B��T{r���?d��\v��5�B���<G�0���e��Y�"/G����[^�U6��Y�*�.�Y�8�"��!��ݳD�Z�z+Crtx��vδyH�a�#w���q�.V�������9�p�ؓd�D�Ίeˍ��!_|�W0 �
�0��rYX���W\j�H��;�����s��##���ʑo盦T��;t�M�1WP˜^��K�<�pp������Mem~��ߕG}��;V�Yia��jo�;'���wВ�۷ߗ^r{�!0v��8>��Z%0*{�0�)|�S�4�Pr瓆�ս�	o��<���j���f�	*#n�r	N��']B�^u�!�9���㐁�$2N]-�RmqC�����@,�6�Ej�Ud�h+��JĪw+�X!mU�)K�A0cn�F;²�LNLY���c��ڋ�W����jgü�[��l�f��A�r��>���9���}��҃Ŗ
�"oČ��Ɋ	U��1cNZ�8�\6o���*5�r&x�:�]�H#�� �',i��@11��h��C�P!]��˲���c�5㺪��X>��Ƚ�T� }�g4:6ay�FX����n(��Q���x��F07C��y��F�,�B��R��ks�deGGg�9|�L~(R��=:iV�Ɛ�(YL������>"�"�P��8�~�Ϳjt ���� �9�����Y�c�+�
|�+_��M�e��.Dɶ�!Tv�ܽ��ͷ�q��ۿ�h��ET*1P�1�ZgA�����.�
���"&��V t��
�q��׿f�<�:� �U����x����ZR�0��i�� Uox������k֭�߻ݒ>��� �/��/m��B�G�����E<F��b�%����͊�@�WtE7i��8��u��L�"���$q²��nk�ё�!�mxR;G�GIP���0�՚��;��B](	�x�{n}"ǜ�U�?.	Cᙕ�QRp���¸f�Op^��
N��������g�{�.�7N�ȑU�K7�y+�r��(�M�TP�������I�0ra���Ūa]���)?\c*��Z��t�
�i�hV��P˭jJ7g�s�X�*�1Q��-����F��rE]��F��%��I$K5tךN�cZr��A �2����m�y_4��i����Z��>L�r?��e@=�?~ߟ�
X7d�>�Ʒ�������>A`㻀h�3�l��`�=�z]�o4��5BX00-�{�-	�#g\�l�m�>�[��X��c�R?RO,k��uu��B��[�(�B��׿�����`0"��'4>ڴ�9��2��2�4����a���&�1�npΨ� 4��̊h#$R��>.�g2nz��������n.X_��������/����!��^ ��@k�����2I�)�K$�`(���>��D">����2τ���["�P�g�OX��ݜ�*DQҎtnn)Zˁ	m�1 �,����"b6�~^㣅���ʙ�U�m��3�<S>������ߟ�� ���>�9�� ���D�^Ƴd�ܽ#�����T8'�|8h���s��6��aʹˎ!�3��Ȋ���ݴX	�B> E]�Ї�w����躄M'pY��\W���~�17]�t�O{ܪ�Y84�No|&:_���{Z��k��5$>����54�H�s��b�3���b�}2�{籉�'j�J���G�h���量>�-��AZp&�G�b�mmb�B�`O=�>��>�k����}�'��Z�v�F�욟04��W's�s�<�,��:�+rv�x ��>�,9�0|zOT4Xg8����|��8�k>�|�M��40��P���zh�aa�+`����O��L�=Sc�{&i-S�(Y��s�P8aP���rS(���>-5�"�{���M���~��;�w)l}�#T���y|AO��S���Ӓ'j������ p��2!Tدi~�|^�5�3�p[H�p<�ab��B��ÿ���.�G>������yoD�  b���-/ �
^��,����Ƃ� ��c����hNFs,�����ɤ7�'�m�i�yc�Vڇ?�a����}�����͍�>������7�s���P��L!�6�/�}�I���'��Mkʷ�\«��"6Z��5҂Ǳ���hnxc��y_�ӛ�s$�Wz$ �W����d(�a)���򇉀�����2���sH͖�o����}�~Z$H�4?,⯋VU긎�DyF~�g���-'k�f��u�w��N^��#��yDU?��y��ו�W�>���4p���q����O�
�h�%��Z9=c��
[�M<<�������>p�xA�#�e�^ ��6|Z�'{���!����+Z0��Z}��D�-�wz�x�gU�|�<���r��js�z|���|___b�3�G�L�B��p���A9Vw����������\�����4�3ŵ���yzE�Z����q�B�
�G����g���O:8�4p0'�(j��Q���ż�Y��+Þ�������9�=��Z�4<V��6�ۉ@�hٙ���Xsq/��/f��_d�6`% �	�I<
��M�\�}ف*e
!*1ߺa��0U4� �.9|d(&�j�X�͞�h���	�5�����c�3���5�y����=2|Ԅ�/����A�{�@b_���{�6L76�o��:g���Ő_�`}߁�"�s�u�b뉰�ߙ��@@�Ч���5%Z����>�(]�������-,��c226*ݽ=��:p�����87���8�x�~���:������>�~�]Ιڢ�c��:��,����Q"�S��[��g�dz���a��k��c��h�y��j��Kn$n�<^�uIRaa�c0AI4r���'�]��� �}�In��7�Ip�����l$b����L�����hY�@K���b��ap�O~�3�r4�f�Oa���.U�B��U���3ă�
!��.`�Y�CagB ���x0����܎�s��)�}t�����ߏ�7���00�Al߾݊S�5@1c#oT��n�5����2����s�d3��*w>_*zz����yP���<=��Ѝ�Ȍ��}���h�Od������ډ��L�Ml��+�u˗��Ń��H��p6)�
y�)q^�8�no��	&?]|�~8p�\�/?�����8�މz&�p�΃��_&�y���jm��9?��G��������ix��G�c���Ƿ���l(��0�
��6p�L��a���OC�
��Nǟ+*Z�;<��;���i�%Iq�A�`��V�)�4�4jq_+6#Qb�"�/�3hm>�� h�Rc��e�_�ͮ��<%]=�I�̚�x�]Za�d`�b�۱�ߌ~���Lt"j��h��76b�� 
����Ď,��~T*�d���;�8���<zܒMq��k1��s�a�#���?b��0����%T�I &�zg耉A?�K���R�;3|�����{)��x�����G��|�|��W�6س� �ņ�Oy�?Ο�/^̔_p�lݺU�����gYSr��!������S;-�%��'>���F�{��x��]���+
�V{��s{�'�g��3�G�{m !g�
D��oȽ�w�}VD�y�o���>Aˬ�ʳٔL��I�?/<���u����љ�Ze������p�g�s�>tD���;��"y���70�1�D�0��dCD����G{�������ʬ{1���g�^�k�J��_h�a�Zy���#i�a`":1��׹�|����i���J!!iֿ8��/|�M8NWwG�Ks! s����@ׯ_/o}�[�c��ii�~���Cdh��t�~���¥����h��h=f#h$z��믗[n���	�@0�g��-[�X��Aw�u�) �*,��Ny�ߘ��
`jr�������w�g�nk��{�N�x�K�ʦ�g�E�\f��(�B�6@�|�I+��
������_~����G�h_}�7�Bb�l��h��6RG4ú적~�K^�dFz{�L^ �������ADa��A��W��UV=��������F���
9�A����W_)��21>"#��r�]w�~U H����DL�<!�<|�zc�o��Tڈ�n��K����J�/}�|�ߴn^����jU�h�N���NȘ��o��h���O�3��W�C���GOW����ܿG����㏘G��R(�#����\x��&Pdx���lE��n�8b���Qs����s�\t�����)�V�etx�H�\����4���l-�j�>����ɫo�o���E\(w�q�'&�T���_ϻ�
��G��*��l;�<y�������޹K����h
 Z��H kBҎ��Vc���^'g�`�͓B}�g��^�23�ц!�B7t���o�Ċ��Rq�%�ʚU��V-�qZ�����cCOKg�*ݝ���RW����DE���w��񆛭��ٛ6�k�<��&�|���*�����o5l�!̢�}��_�ݲ՚z䳁<p�vY��G�ذR���ɤ�Z�i�6���P�~\?[S�������ꪫl1��G��6$�B^�}�{���7�2'�3���e�k��h�>�0靣;���Y�- r0������mo3��=��h�CV`�W+E��أ*+�j .�]�G%�	\߈L��O��ب�i����++V�1�Б����,>�:=Q�S^���a1�C���ի�J�^5�s�S�f������J��Svr������ݵk��t�M�;�Z��v[R��&ޯx�+l� ��\>(P=ca���( j��o��x��3�>��C�7�7I#R����W~�W����}��=],����<��òn�2�~���J:$�=-wv����49w�6k�y�g��e+�����/����-�g�
_8K��T0�)�I�VD[ɻ�O�oe�֤�!�0m�ᒱ*Z�����xa1@�Ӫ���+��������ϟ�V�!IZ{�G{���
\둃��;o������9~�������x����qR�<�{X����+�FJDVƋS�C�\iX��{�Tt�=?�W���Vk�T�K�Z��c!!�S^�A넯�42�M���{�|�;�J�h۵�C[?�'����/ ����/[|n����>=�y�<�$vj'|O�A�.l�9��G���>��gL��;�A�S�oذ��;�������-~~X�4�l�֟�0D���dJ��L8ցj��EǏ���	�5�Ԩ���,j�'lT+K��2����ٙ��֟4���0N�0H'�Ux��ĉ=8Y�����q�Xxn"�?2��]w��C�����0��h��;��Qx���ַ�%��ޝ���T�-oy�y�0����]�ش�'��P�̎�!'��Xod�4ʖOѤ�#�$�I�����r#�N�"�(j͞��4Y���ʥK,�a��R�Eƪ�J�%�q�1�ή��d�>�B�%~H�X����������\>򑏘�G�7�����Ѭ�����sj��>�0�[����~������G�O������˭��j{�`ޛ6m�O}�S�؊�M�H���/�5�֫LI����AQ��v�9I�p�(t��XY�_�m۶%b<f�"?�0[×V�/�a���
�y"�Zk׬R/��}�<�G��0�U��/.�JoO��-H�|P?7 �]v��e�>7
���`����"����=��K��?�qz��m��>(H��=컀����{v�o���MX�$y�������ꔳ��,�G��ɤ�,��υf�����6m��v�BG���	
F�X�q��iKu��R���]x�
�,[�R�ղ<��ӪaG�qG��!眳M.�����I\.6r��~`߁���|�8����wZ���ɇ��}�p�c�N�ʎ��q���W�'���ty��"��$V~GRg�d�YB�0�o�1[���,77)����8?�/�ɉ�K�������y�1�_�2�JƻX�J��5*  ��P�����Hދ����-$}��o �?&79�lbC�z2T2��gHzs�}!�
��_��s0��k�:�iP�����y�@��-��y�_����~��,��<4�1j�������?o�j�$+d�X��{:dO'��U���Y��(%K���_n�Q�����]O���s�}��������XИp<������=G^�����1Y�t�\z�UF�p���Y��T���˖�%����bIg���m�<t1$k':>������ :,AI����ÇfsQ�Q��h�gjpsb�#?q�����E�M�E��^@;�/k�B+�\�>ԕ��A�4�����m�=(x�~c�R}�/R��^�7=�`ǿ��կ���ߟ��=_1P]s�5r�7&�W���3���]���j�H��e/7K���&,2�DA��%�B�G�߉ޢ^7�F"�}#ȓ�o�9i��+<���$i$�U�A�1^�\_��WY���0#�a��?���������{����<�B��������0���<�ɟ���gC �y���׿���{��{6Ǆ{�a"$���"S�c�y��j�wȗ�����K�AC�=��/|�K���_�x��s�]�?\,��2��Φ��*��k}�s��z�^t�ҥ���yW��e�^���JZ5m���9�Q���6&������-��A�nX��n m�o��o�{����I�+���bwl�Mr7�W����!�[C52�%����䴾[?e�9���6L�h8f�7+}�
A:��Z���(�sB/D?\}�����/]�tV�����ph�ؘ���&�9ر> ��}�I���JdO?l7�kn��|A�>�LY�r��3O�^j��W�=��q?I]26���
E%9�u���S��ӛx"~��38z�b�	;�[�͈���k��<P��MG���,������gϊ�J?,��`�����C�����dQ���k��mF���d��+L�A��=��a�!��q�Fy׻ޕFrmq� �eq����TM���׾��\W�<e�RД��)�G~L����q�d��F�q�� ZP�<ɚ���7�pú��߿�v��B]f͆�=�Ѓ��s�w���L���zF�����#�=jud�%���~�*&
'Z|X���o!�b���UNE ���R�c����p�v�s-~��
����ϰJ���ߧ�dώ!!�W�ӨI�~��' �q8�^�{���`������8Y�ʕ��?/�m������}�[��l����=��a/���'�}eϵOO�k�ϖ덞�=Syvqs���uB@c�RI`��'�y*1�}0�_��,��y�fS~��{;�{ts�X)[A����g��/�����i�珌o������RR���f\!&Ъ��/+V�2W�O,���a�����zUd������M��0�?�iq�9n�W������l's����xa��%c�rȑ��^�|���� ^�������}sh�֧��I5X�xQ�Q��q�p��S�u����a�ؼ����xp����1i_����5���=�䥳Ё��f��rQXO�+9j9�T*�sCh3:o���뇑�^D�P�B���g�Y*.��(� �<BZ���%�^�'~�i�|�s��yŋ���/s�}��)=ey���>ԓ��~����7��]?>��}$b��Pq5+J�#��a�֭r�X请�[�T�ܷ�LV��l��~y����D��Z�I6?�C�NS���rv�:��\�!~%� ���?����d`�	',V$��.C01���OǌX���f��}�!x�,xp����7[�>� ��O@���͍͌P�� �i����`��%�������7==)��5��7�,T
LB#���~7���$)^V^��ot|,��)@1�D#1�!6�zBPњ�9���0mV���9iı��1{:{���B�����Iٹ{�k�L�/|*&��=P�C��8��g�|�)��1��c68'�p��s�����g���3`�����b`?`��0�9�,{V��y=I���مD�yqo����tp���կ�#����~�~G����)-?�Ž�^޵F�x��\j �B�^1�a�����G��R�Щ�:���N��F����?h�v4n�u�k.�6`E�Ʉ.�ѝ�j����|GN��,X�VD�`#�DՇ?�����w��xӛ����̈́�/�N�`;J�#64��f�Xf��惫⸰��=P��l����D���a�;=\6�e2ˍ�����I,��}D��+�(�yh�IbZ��Vz/��1�ZR�^�C�E��XQ��h>��r��C��,P��J��*(N�p�<��,p*�f��?Wț�ea�8yJ�M����� �`��s�;��|��dqds��� ��1���i��� ���F>�=L�����[z>Jέ��TPիr���A�,�$k0N�Cr�5����ú�0/b����"	,�=91e�	���U���I���p�$q�t�I4�ߍ���X�e�2 ��dŊ���Й78ق���k?��w1|8'��ߩ�����r|�()X��_h�j�Э���q+�D���q|��6�����0�ޜ�W����(`}��l��Ij^+Xb-Y7�0�C\�)���{�� �,H��_=���{�Ռ�3gB��������[�:����\�0�G|v\���p�?>>C�|���S�g7/��J��珠��:#E�%�ߢՇ�b-�o �d2j,�l����&��8�,e�dB��ϲ���{b#h��u��ۨ���?V	�^d}1�0m�� �;Xh�]�X�hcc="��x�ܳ��f�=��C�@�x�Y� a�pQ�R���̑l~q/��(nf��Ru�h?��j�q�)���KH��Й�}V���%��;@ZY�R7��������˾��i��L濓�ϴ9tJ&�vt a������)<�P�<5�����o?gp`�#Wt��Xx�� �\g&��D0֜����3	�3p�����Hl�ÿ*?�M���8����l:cs��17��ʦ�4�e
�,��!�Ű�M|���,�<�߮/�p�=��a�{°�	�<�.����u��3���	�`��&��ǉ\�9|�;�� TuA�Z]zR���w��m�W�@�$��� 7��o�/}�K�w�ð���c0��_���>��ǥ�ǩ=�}�C��
a[`�ִ�o�qӷ��~��k4b���t�7�ik×ʹ�?�8兿�C�0s2�sq������`��ۿ�[��9����p��C�dl�H��!������g{L�F�
lME���j�z�=~�G��>L�'w�3LO���A�������� �+fr�
�f����9�F��D�I�8����6��)0��1<?��G��虑	����d����(L�g}�b�q���sz;�<��6�����Cs���������W���y��<������V$�O�q�8�HY�|O�3 Ny��A}<�`6������b?�O4F3���P���ΰ6B�D�l5���������`��,n��(\�h�}�͖}̤S��1�n�3n<s^�1��;!���Oo��'�s{�c��ii`�u����`}m��Ux'#r�ۢ�+��)�g.|���'�����M�4��h	�0�w��k�w�l��~� 
��
^
@=�io��s`���"�t��|@{�,��Ѭ����_���?}���Ж�-�F�	|�ٺjSP�{|�%ףUT(�ݻ�����B�R=�P����B|�,��9}�d��s�܍ފO[܌��B��z����MFG�J'��Dn�|�x^=(V�2\f?��̦������|�����x�,��I�XC�b~�c6�?9JGR�T+�����������r����>�oQ��lI�l�7\�1L��I~ ���Jȟ�E YR+!�$� �)�1`\0`\�1��]�,ٖUn�w���g��9����;�;��+m��\͜9�-��gW5�?���U+���bZfO�*`A�Ey����.1�l����[)��a�;�l�5�GaY���H(���cQ��p<�-���k��7����Y��{�ޅǰ�����"�{��P�4�y{^[�w�1~�����W� Vڣ�#�}c�+m���?��UuN�W��ZE*e�|Qq�^�-�w��m
c̊;l �����+�u'j����2y��؊S��Y�ąN�*�����8
��Mt?!c��D*d%�ez`�<m��1X� e��8�}[������0Xm��%K�m�p�Z���,��D�sT�����sl�$���.F�<�
���3�56Z��(bKgRzL�Z� ���#�(1p����JX�F�A!Bs��.P�Z�� � ����Fh�ز�N�b�(qL�R�1�B���9f%lR�v����G��9�t�b,��7���x�	���8�}.��sj���ϙ3[Fǆ��zp���A�]~��q��ߢ|�VK��!�дg�A�WD۱�0Y���}�\v��N���Z.)�b	Mݻ
�Ig����uN  �1 @�l��
^�fc!��Z��GX�YL��Iu�����&��N�Q4�U`0��Lm��u,d��dT 2A�q`�)Y�KfNm�V���"��Mgb�:��Η��,��d��r�S��N�	��1��2��Z"���ñ}�5�Ԃ9~�'��ٓ�<�!S�q*
y
��5Pج¦���R����� ����պyO[0�}��h�A�ь� pOj��5HAa�/�OXw���7�Y�
>��,=�9�u.���Y��sf͒׾�5���\���^a���S~6��4I�Ƅ`�g��`yL֟z���Ȭ�3�f������=�ec1\��c����9�Md�6ky���._���b$E��� �a���B�Z�&��D�$�؁��K����d5C
4ݘn��Y'c�8�#0�!5yj�d�8?z�W)Y�O��M�sw��59���ٳba���иy��[�%
�;�.BQg�g��92�����b�3\PL ��X`�cQ� r� b�>�bT���xˠ^-�������G�f"K�L������L�������a��D���&������cl�P"�Nz_�����t����]�O�tQ9!��U���_�����%�8��ݷ�٧䷿�[��t캻���h�)9��c��7��u��k~$/�� �@z��ml�i��C	�z�8y̓/<_�͟-��N����~%[�>+%'�!e+���9&O<&3,ǝx�t��ҎPhG�~lR�?��]�SN9E���_�m�K퉌����$���"2C0	t.BĶ\�ϟ�-�;p΁e4ٽS_�j�\v�eu�t&��Ʉ�&��ǀ fs�A-���.���Q�̟Z�O~z�jRV3�1�
�L�-'ў�`iDs%�0 ��o�a��Dc�p�b}��K���.���C(�X4����C��U���M
e��s�9G�=(ȒZ?^�=p��z��x���S�Źѥ�!a�R8[��>>��kY��f�{B;�3�<ӯ�Tz�rD`3��%q�/c�A��ޤq.4�w���O��|`\<Hm ~���uD�� @;̕+�;!^t��O6��<������(� �z��k�rB����M���;������B��`��� ��YS�  �A�-���\9�%R���}���e��s�;����-�����'w�u�l~�Ey�;߫Z��@�>9�(�t�^{��7����_�z�h�� ��_�<�7�abc�'�	'�0�1�Uc5i=4<S�����8���<�+
�]n�yO��غ	B�q�ʬ���jo��0�?���4��P�h�y�\U�����f�02+�0&`Rt���E{>�#�9s��r��hL���)v�^�����}�m��*��i|=���cM���E;�ItS]�c>)�gŊq۴�������Bj7#��&�׮�S�y��C��82ִ�]?6 ͽO��Z����ZQ{��1f����G�޾��o�J	��P��k�S �,�?z�<��S��9�;��~��<������ʍwEN[�T���=�|y���Um�|L{�6���is���渍}�G�s��;n�#W-��;�ir�ed�_��7�G�B�� �<ޠR��6���>L:�p`� &�@7h�hm���7�u ��6֯����t�n�6H���b�H�9��[_2!0o��Q���vM�ic�Wۀ4�),,tv�����b_./]td�60=Q6�2dtn��|]O���0%�źk+_p>WPE��@ 
��1j���0F��gLJ��͞�-3�5�y�:����S+�A�ҹ���x�Y2ѵ�?�k�
,�Mco�8�vp�úB������WW0�� ���|򓟔[n�E;�q��~a=�=��?%�g��Z(7=	�(�+ȩ�Y����W;
._v�
�#�X#����[;�)W�N{��,ϟ�L��×����twed�K/ʑ+�Ȍޜ̘�U(]��LAd�Z��c�ve��21��܅	�f4�|���Lr��.��b5��XsP+AýMt=�O�m8������l���7HR�M4�z
�����Z��q]��O����y-�O�I��P�4ux�
f��x2Qjy4�q��lf��d��k``� ��x-��6�)�`��ٜf8"�}#�$÷)�d�xv4Ɂ&��r���B�)����^���Q�̙׎!���ϛ�}p�����Mg���|�l�5쫽�?x~�g� pK�.U��������Ö���B�p(��7��`�6�>"�g�d���2w�wÏ�X�hA�����-ȝ��[/\!�3g����e�aK���Ti�3�f�����F��;G%l��-۶=�-HA;F�v�;I���[yL�|�8�S�`�Ϛ�AƑꈺ
�����_�1����Њ��翐����̙77�Y??Lln��I4��t�������y�|��Ǖ�=&���s�E���q`�b����:'s�)�d��]�
�����X��6��f3ڋᩧ���$�;�L��ܺZ@����70(���������3 ��
w�r���)�C!±��êD��fy��6&���঺t�z���?�-/k�P3��q��d����a�ARY�.*úRk���M�m��b>���*��C��MoR�/�� ı  ��s���^{񅗜U��?�(�g���NȎ��q�"�q�Y��ky����.�M�����_|�y�Vp����h�3�Qbb�v�ʦs��Ckԁ��lJ��ɡ��c�5�ӒqǏ�n���Q�ƄM�F�^2w6��d��M�l�9��=a�a<�,��5*���V����O�qܬ`�}um:� �^��8��Ա���}c������cj���6va��Y"w,	0�fy�,X��F�<��gצe����%ƿ'"��®++���I����"�f�q��ʰnЫ�3���|�󟏳�p����ަ�~�/��8]'N��#w!Z6VkN�G6W&���J��`�qp��)�t2���5�6':b<��O��B
d�8�ȫ^v�
��g^�Їv��wҵK���ag��iSK��;�ͬ�X��p饗j�j��@0��{�y�7d�gf�X_��$n4�dL����J܂�%6�f7>c��L���[�i}��\N �1�c5P�l=)sh���8�3�+��
U��-�i�67����%%�k����c��4c�v�9�|>S2Pm����#�wؾ���xnd���_��j��v���������g?��c|i�0#��B����3*�rF{���ު��yi�Q�@]�iY��-�Ҡ����S"kHR�0Г������x���	�_��	�/=��=g�̞��i�nӧ
jrժ6 ��K���\�Grd�5�ό�{�G}��}�k��;�6rva~�+_����7�f�Y�n�6���Zs���u�-cO.�F�d5�fZ0�ϑ<�-@%���Lx�d�Q+4��B�g5|^�~�8s�h�Xo2��˞�ײ��^׎�i(�~3�k����K�}����J���L�eb���e@7yO��ܛ�k��`V���뿎�'�� Ա�Y���cb�
�×.��b5-�l |"B5��I�`����󥧷�E�>�E�B��[+��q���?&o��5_������3ϐ�;v9F}���}��9)�#�fuG�+9YԻ��Ԟ�.+V���-$9Z5R+����P� r�!>����>�1�җ��ھ�ٸ� h�l�7�'%�o�_��%��̈́�ua�sY��M��Y��t3q��2jF�1w���|�y�6Va��V�?��y�ɿ��������
�f�׎5��H��9��[?=�����co�CA`c1��j���]�E��MaGK ��9���{����p�����@	��dՑ�ep�%���B�L�vVB��U�Y9��3���k6�G�@�>�X���$޳�0L��P�����\Z�{��.7��{�L5ǰ��966$4fϤ��v��r��r9�����0�M�6�@N�h,��.�*`��?���p̒a�������,m'�!��Z�e ����2U�:HZ�>�L�j��Ѫ�Ԉ�l�E���&�߼n+���&yV��3
C+x,��cb�Jj�,���P�ot�V,��{.�Z�1Ѽ�m���B���(vC��;3߬0~�ޠAw�&p,���:J��,;���T�Y�R)�M�1�h2�ͻs�e�;�s�tǮRK ���[�QQ�k��:o�WUZ��r��r�mw�+/8_F�Z�d���"�������c
]r�I���^"s�-t����wOp���_���wj��~�� @̶m�����l}���bd���w�/�9��i�$����ؤ�8Y�����h�[ �%��O���ǤO�5b����`�2+k�7Ҿ[y������3��cac��ڠ�T�2�F�9?�ț�[]TlƘe�������v-���������KZ�M�EV,y$s�uI%�{��塇�SO^'��,9��N����]���������b�r�y���k��r1����]�=*]��b�Dn����?�?I~� �'��?��P��c�s_����\�������ŭn�f���9��8�U��� ����=�,���0�9|���*�׮Q낛�n �q�O"^�D���Í�{�I�}���=�s翭��U��H�p�m�)���p{��>R��粩�I����
~N렙�k�u[��<&7�s�T�Ɉ�g�xr�W���Z���fa �?��?W�>g��f�� H��;{��\�J
�9��3�UGɖ�7��� %��L֬^�, �SR9�%��#���?�ŝ5.��s��V��=�oF~��9L��\u��w�Z��	��9G�Ξ[߬nB�ق���u�}/�������?��?>G�=��ƍ��͛b�.d���.Y읤o�L���`l�2�F ɸ,�� �����>P#�ОR��Z�7I�����ͮm�C��7���jF��1�&��~��o����a�k�m��k� �}?p�Dw�2��ـ�����A��
O�������7�M?��gH�[����I'�.���xP�]#x�P��n����:+�?��� ���S|�����^�.`g#0s�q�)�6�}L$.��6l�GyL�=�0���l,�w��ݺP�@��8��?��'�.�={v�;5�v��� �8#i�X�8��QV�>D��`%�ka��}ٲe��|�f=��E]$?���!�ҽ����{?��b;�q��b�
�'2��/bk
(N���=���Nhx��g*�B�z�N@���u�W� S�7C�vI��}� ���u� (��[�@ ��>@j 4���|�Wj��Ƣ @�> �z�ߨ��XP� Y'���
�/Ns���Q0j �vb�:�S�a�#U�C��Z�@�E��x�`�Ŷ��a�Ê��������C? �;aR�g�2�*j�V��R�r�_����ө��N�N���G0�Aq�"Xa���&
�
�Dj*�7Z�����& x!ЋB.��~�a�馛tB�����f! �:�����Ad�eQH�F������Ƈ��Ob�������ܢf�+����˿T�
�u���� �l����3}'����ξ�}o��4SWÈ��aӞ�7���<`pA, �xV2ٌ]@�����t2Ku@+[}���h�$����=����;��&�M[#=��"3�=D��`%��2�M��1����������` ,	��{M�E+�?���� �֮�����[��gS�q�FA:OL�g��|�8�!���Zq���.��-�3+�S6�[ڝe�������XT>@�"�EĎJ6ۢĸ�f��%����{��E~���v��!���p�0����}�s d3�\�f��dVF*^ڗ��BOlex�>�k����PZٞm�g3�OGn'���R� oZ{�z�|��K�4���E��v���_�O�ӊ� ��XLHE��׾��* �o���ЮۅZ?�6����l6������=n�OX��`05||��O�~��/����f��|�+V|L�1`��
�y�@N�{��LZ����'���D�i�	���g�M�����]��N@*=��"�Whְ�̜Z�L>�����҂�}���"J���4PJ�$FK�f~�h��)��ŋ��� �������E�<���5�O�8hNcކ��ֻ�Ѻk��`������ҩП����/�l���m	2��=��f�Y�E�3�#�^����7[�kB�q��>��<]�A��{K=B��/��h�	�+�@�J=��~�z*�׺�ƶRZ�D�02��@<V��oP� 0bҷ�ܡ�$ѯ�ģ�3���(��^s��=C�;�X��e�M|*���y�X���cŇ���@d�X��Np�=�j��e�,�T}+?x>�r����z�����β��J���촞,Vp0E��^)'L��3��� ���ZM��N� �k�]�ijn��1����� ���[�)����U�xR���@�琡ں�d�� (�$Pf�AV�K֊���bƎu��,�m��?����[z��]��]�"~�N��sLg�S�����L��aJ�����[�!�hzІES�g	�,w��ò� N��G�x�z�"��Mz�p��DGc�^K��s�0��շ�yj�48'�o�vl�
ٜf̔��fh�K�k��cJ�RHd��E�ð���;GB'�*��ҹ,L7񚿿�={G+Č�`�Kѽ�:�e�J9�-��0�}G�����/�K�_���71H��t+�Aºd&W���@!�%P���s����O�Ly<{e`�����R3EN[�"#d�5~>�,j�_���ղ��T�h%���󟴁�����5�)*W�:I�5`/GЭ�jݯO���:�m��V�"s�����M�DR����A����YRp�*�����O#�F�;����>;%i����;�̌��B�t���<t�8�T�u�A�,��|���쳲t�ar�y��9�,����NP k
̿
�B�1�ZQ��[u���-U�W���H:�J_��|Ӎ
ّΠ�O&������q½w�*�8>��F�,5��}E�_0[Z�!�M��(`�x�����T�|�[8��dd-�F�t+�L ���5x�*nQ�O�[�,�EJh���i��C	�b$@���ה�����3#n��H��V5���v�I?i^'K��6ɓ�k~x�Ө�ҋ����n0f��i/�]�E�Z��eo�_J��ݲ`�|��;�i@�R-"���4�XK2�Ǚ��;�4�Tg������E(�� ~��3�����	*���䶕���fc�nӹ�̘�#��,�o��Kp;���@�FF��B��2P$0~:P\=�p���&�L L�%���SH4�R?�J�e���GX�z���zu�R�F��z�(�<nw�Z��k�!Ϳ!�}zٰ�1�rMq�1��C�n�u�.����(���}n���wO]���mTQLַc�{Β�YrQ�?�}�i��%g�h�Ϩti�W�� ��,�h��~{�/��Iw���Ԫ���^ɧ�B�He~xǂk���!��.�9&0�"NVkS����g�?W-�� ��T:$�ZY��9uE�
y	�Z��Q�����"�XM�ʽ8U���Gx�LCf=�Ex%fՁ^����
�6k���Z]�&C�X��w�8X�*��4Ѱ��������5p��A�=4|,("+
����n��w�1�Ë��M�����	[���b2�}���G�9F̐l�G��Uefź�5W��xn��3��*B�^Vj�蕙s�h���`���%�<:be�7���9���gܳ�z�%ǐSmdD��i���ԱgYcN<S�FS���	�J�397�9't2��S�b���|�ΠӚc��D���0�FOk���`�׶4���E~�Sr�'�1��؈,�?_+���fb\��B�W����6�ӰKQK�\1�������>�h��[�MY�l(�)��ŗ�RN?�tQ=0J���>�9�u���jr{ٮD�dU��Pۣ���Į5.�ae����$К��������1�*�����o4����vz���hmX�8m>���T��y��s�Nh�Kge�1�.�}%�I&�չ��v	�4CrZߝ���
��sK�{�.'�rRvB�\)�X��!˖.�MO?�kb;4I�4����9�:P�%d�̘�#�'.�Ŝ�3ئ�:5�3β>��3��sϓ�n]A1�
�`~u��ZIL�������}M{���3hJ�ޞ�����sΕ׿�5Z�U.�jZ$�%�"r!k� Z��|��_��6m�tO[���i�j���+9F��c����qV����U  �"�;E��ct%�}���p#�qi�PkN�h��H���tI՜�VH���G�2V��ʘT���v�;�0�B��˘ȔR=5[��-Q�eU�⳺$����L*�Wh�1��~֢� 1,�c�����u2 69gS�|�Q��ýv �Dֿ�72Yy��ީ�������ݏ������w) ��UGʯ�k��m��|��.���D_L{���(f��)��"W��M�Q:��M�T�n���"}�}�`��Ys��Xy��dg�q����ۿ�[\-�I�$����?��?��~���'�&�ැ�>L՛����3L�Q����n仫pH��X�� ���{ѣM�8�B������$,�J�����R�8�;�>K�J-3&Eg%Hۚ��}G_�'�jydB��H�+�Vk("s>@�T�9�WM��+O�������5P��n�U{y�`2c��݊{���P�t��u��l�e�{��J{'��I��� ��Ś�~���mJ�e K�{�ʕ-��P�9�����K��a�ڬ?޳���1�������6Y�z� ]�/tV�}�<�ݼ0.,�#�X��u؍UY���Μ��f�k�<2�n�3��ɾ��x��*K�,��^y�t�s2sV�lټQ~�>y����o��Du��'�g��Qǜ �ן����e�]����s�9��կ�a�� ~�t��o�]���oi�7��Y"֠��h�M�{J��:t�F�J��8���0�i��U�V�-�·��L@�&�]x���>�.�2��Z �4�`Yw���G�1��%���R��ߖi��Z����tYw�M��.ٚ3�L�%�J>�M�`�<S-z&]BG��Y+�b�St"���H�<@� �
{�9�����p��_�=�0 �/��r9�5Z̈ڢMO>��Z��9�:�v�nY�r��~�ٲ�5�,��;Y1�  l��Tb�Ӟ�7#g89�c�`h����Ҷg���[��#����h��Ӣ�����V����}�yH=��3�_ߩ�`,
hӐ�-^"7�|�B�b°@������=��3yV�/j+,m�7�Oj&)��\��(�pZc>�6t5#���K���s�������ˏW&���VI;��7橥*�ʨ� ����^��� ��J�$�6��d۞��m�62(��j{�&�M�&���70��ɸ�M���?�LP��ReS[=K8�N=C������rꩧꞇ���/��b�����=�ZE�ݬ8��ի���O�տ�rܼ�Qyⱇ����+�?,�-c�J�������ΖSן�	
�7>����r��^'t!�)��g�M*|�Y��*U��a��淿��yY�l������^ �<�B�ᑊ�x��r�jY�x�Jx4kA��>K,��[��Yg����������?_@<�І����tM��{*�aG�Qq��|v�P���@Z�5rbld؍u��AT�&��K�?��?A2�j�pM�R�Z��u��b����1�q�5W��ـ!u��+�Ȃ'2���2:��0%�{��G�s[�oߩ�C�c�ȯ�JH�H���%3��;:�&�e1ЦA����*~��R;�1J�C|�d��?^>��O��c���Au����~m����^}�,�x�*�]��2&�f܊*h��wUah���䦛n��K����T�@�`~[p���nA�?'���eK5�6�Ч�yR֟r��.[�̲�8������;�\�J���>���;��|�n:�k�qD��"��w���՗�n��F] X�X�����$�)n{N�l"��tE0�6N �̘׿�m��RM�-��*�28�]
��#�$��|4�ew*]S=� R1��B�3��0��V��!H��ޅ�S=}͇w�x! �P�RtLi�c#���ޤ$���j�I'��4A���?'�4�� �P����:��q~��~}>�ʗu[��x����b�Y1�2|@r���2]tP����	���к�u�E�{� ����/|�ʨ�	H���ʕ��yxý�d�Y�h�����;.М�+����s,�����j�W_�Z=Ǌ+���v��V�m�3�fD�����ӧ����s2:��&bT*U=e�\q&fyX���� }+����I��,6Ӯ]�T@@; ��{��^��0�&:����l�@�|e�@�t&u��$Ԕk1��~���'^>�rԴQN�<&)7���ՃYb��`��s�"��? ���PqO�ӵH��"�Зz`�0���T �� i�C��F.�0�Ɉ��9�8K4ɉ����,�KNͺZ?��.i��F)d� �8X�\�{ҵ���<7����ۥd�&�O���x(rK�.�7���կ~5{Z`���Ν?~�ȥ��m��='�4�n��lA^�a@�c:�1}��}�=���/����W;�0,���k�Z Ӟ�������g�%cVq�3jv��	(9T�l�riDjUg�� �3�j-@*��ɬ��^��T쟋��O�S�����MDs��K����[9t}�"���BA�cHtu��m"�����h���͂^
�ﯦ�W��UV<� 5����%��DA�v����Dh��T�sBp�v�g�����^@���MnR[	�,��-n<�%�y��$��[�&�̶K�G�;��y߼w
�����a,��If�gc}���+�}�ϡн�oTW.��ڵk����C'�w�Ճs ����~��R��}NX��Kh�@JQu5�ᾃ5��R��c��S��i���5sa.1����TN�xs���������� �����G�)Mgh�0����oD���h��Hjm�ק/�M�1�8��h?��f��>7_ǄC���Hۍr�c5���5��w�g.�CuL����!��(����
����gS#��S�o���#_��Pg)�4�S��8rt�(�ã
+h�M�L-�W�g���p5�����M��mj��NQ����Z6+Ǧ�RC��kƽ�p��a�C�>�ǴK6k�����L���%��O��
=���NS����}M� ��e�ݧf���W�������og+I�si�	�2:6,3zg9!��1Z��JM� O{�N���4��]2:R��+��KfΆy��4�R)#]��NW4ҷ��Ȁ/RM��/���1�!��W�*2!R:i���X�h�UW�}�&�d�%�.�OM�����2���̛�)դ�������	c�"恳��+ձ��s"�240���,p� ��F-�� �vL����W��uB�-���5�SH`��J��[T�@� X.元fi�����r26<�n������QAd���t��y�Mx0Ƥ4VԂ!
u��y���� ����|���V��H �:�<���$�BbO	���^�����تZ���x+��o�E�������[������;]W�����E�:�(�\a�޿��䆛n��R�6��4Ȏ];=�������e��Ŏo8K��B�L�o�ҘS��&�/�X�ם�>��%�Ok��j>{B��BӞ����cOl��O<N�֟z����K��]n8!���M�O�����)�y�n9��T���7���>�nL2���ju��
>Z�數Mls�4��B0��dұ�b��N�F�r�i,��1~�؛׮�;7�_�j3��+��(4m�<���������x�1�Z��,��9�|V�n�T��L!�'��Ouų(J(�Jj�D�%��1�����J��r���u�:DQi�Ϟ>|*rxG �>�|��?u���آ��B7���;S�=�x)�������~�2k�B�(��E�9�,��v�ˮ�a9��ӥ��[�d[�<-�7=%��yiFmߠi�bM��0�P�q������Wʖ�7��%-ꁦ72:��9�[4K�=cr����J\,��^zI6m��4�L���ze���C�c �yx�[���e��D�����[<���F͛+����is�7	�-��)t�E널�H�<���x���b���{��k��KP� �Xq�1Y'ra�Z�g'�Tݴ �\r��C.���X4FS��f,�mړw`Uſ����ܠL��-tfKe|��������b
^
�hjd��<�%Ō=ya@!���lJC��'?����}�,=l�<�н���!w��S��d��T�Ȃ�K�R�ʪU���/W�cht@�{�Y����'�i���������=�������'+^�����A��'?���~�+SJer�x���կ�E��Љ�tG�|�4�p�򗿬���1����?�o8G3��

ݲn�:y�Wz�(���3����w�� ��K;w�=�/�n�VՔ���)�zqc��-�1�7`�1e��%U ���6�H�1��z���l�dr�,��F�v�m�]�WoF{�jm�"z[�YhX5�a�k�E���;����d���3&�̝׿��qj7>g2�7��͚��{�Bb�ƍHϟ��.9��u�םr�-�r
�f�UK�\�]
/���s�=�Y�0Y3���Ɇh�QOWs�"���_�d���85nH��{�1NS^�����i�ٴy�j�k�>F�S�1{�cZN#t��-��"w�u�8�%,x��(?\<G}��@�lذA#�H�1V1��%����u�a�d8Y63�L��E����X^1���%$������w&�3�Vא
M=�ˠV���/�Ɯ��%��,��ze�PU������vR)�j�=R^�=�ŷ���yki���K p�iphX7�:��(7]�t&j���U�}�L?��u�?2�Ps��B���ه�d��{�ys溭�-��~��Y}�<�Ѓ�e���e4&�~�z'4f��pEQ�~�Q���~���.�ixƔ�M�;5i�D��	#��������G����n�3w�6MX�t��x���#%�Q��M7��Y���?��?V�����r饗*x2���
�Bї�a����k��ry>�b�����#��p�t��h���6�{ob%��묍�'}�04l�!��2&��(/>����%ya��̎T�U�3�xr���'��3�>�<';�������0S��rJJ��t���������MU*v/�C�&Y�$f ����Q�����5�X �:R������D�R��P�|���hm��×鱳fg�.��pX[8N��s�	���Oʏ�cy��-*l�u�����R=	�06R��z�t}�Qg;M��x≲b�2͂A:&�VKI�1�ǞxLn��V7)��0Y���DÒx�k^����|��؝��я~����.�H���!@��Ru���j�2�L./�<��|��߈����,��b)����3d=�:X5"NۥޞY280"w��^M�����ל�)���$�	��������f����K*�U��x
�?��<�V���w� + Up�A��|Je:�#a��Y6�-�h��m.c���R�h� w��m��;��"�}�yp��0�];�� �p���9��p���(bo�xޝ�~��/�����V�i�3�s���B��]�9�����a�͘5S-X(���v3�]��eǎ��s�7��n�219�D�Ϣ�|`��|,X��H�p�$�7p=Y�f��C�=��(\��	��)bQD��!M�+��^�i�t̠���z6ױ`����Yݕ�\
n����K*'�3��҇�/�dj2�/�
|�.oqQw�s�V�*�=�1�uTS
5S*Pl��gZ-y����>�O~��'��Q�뭷j���ɟ�7����"o�;�Lxf�32tː
�U�V�+�T�`�=�͛6�s��
��JeU��+|a_s~�������QGZ�x�	>$F�ˣ����;�駟�A=)����Ro���(s{Y�?�����%D�V���3�tG�ԑ�j:b����ݡ��s���q4{:=��u*�����4+Q�^��, �U!��u�⎫��X�`�)�RZ���L{��)���x�P-B_��Zw\{a�{\CP$�V�����i�v2-��
�\��tF`3n�v�&.�)�դ[ (��<?�W,�u�r�9x1�����~��T�����;��P�
�7�7
���}H���'u�m�7!]����e�6 ;�v(N���(�5֨�)�u��Ti�R�
��ct���2�[��3|b�KVPE���.0,>�>�я*C�������MM?�zDqd�"��Ͷ��m�����	���)��5�`�&�mj����}��
��_�����>���e�M@���C1W��+��̰V����;0+2D
������(�m�ʒhU�ձ�x�,f����$i2&N�TiV��Q����;�
|�����a��YP������K����BRp�"	�Z�/x��ʑ���u���ǫZ���p�=�oV����2e���#�1�1'��X���7n� �,lD,@��p��#$�+H�0գ��(��[�����ׯ��E0��[�'�֩E�X~c� Ўc�k��{*J�4g���Ƨ��Z�lJV�-?��#d��B������g��WŦ��*�����ݽ*[�`tP|��`��[�S3�ռ���4{@TX�v�=5��A�'�GsX���D� �{��+��)�Uů皏B�.���f#�i���u��g�惻�o<%M�o~���S߱���ޠ��WH�[|�����ˊT����R��~���?92a�����7��.�`7��CVӷ���$Qx�+ΕE��-*�?RG�"��K��G,j͚5��!��$ԠS�:g�&���I'�$K�,��<�ξ]z�]���F�3�=n��A������(�!g����y����{$v����kt�ӕf�(���\�!�P�nӑ���h؉�9�s2���qI~�1d�5TZ)�̮`�O�'h��8���K�����e�Ų�[c��/S&���b��[^����Jf��9\���1�w��}}����x���'1��Jd��] M����?�~Z����&�?iER��4U� ��?��UK%�&�'R}� �糀�����8���?1q��j9��3�x��`m�r����JVp�E�s" ���~V <|��u?P�������O����_��3И��5�-�	9��g���.����C��lAl���0�B,\ &���R��o�y��q�Zf�� ������1ל|��˞�:$���#�v�
���h��&/���od�=���2�aЗ!�HZ�E� ��v�*כ�[�xOt�C�h-
4SɁ��"d��פ�<Y���q�����cQG��e���n�p�?;��x�y�6���.� S�����/L�s&�SS�i�������:9�c�o���8��͟�b !(f���\b}pS��	;aj7�ĭ#Y�x���,�i#��=�8k���� f<@�bQ'��*���@{�>�V��z������RKK��o�
١�B����z\�`��7x4�kLW�:�dĠT��ֱ��!�ݟ|�ɒ&c��;��,$4�k�'
��-Ȅr���wr�;����O� �j�������>�A��7�U2��2a��%5������.K� QK�o!�9�,*�ֱ{O�ERs��x#�_�f��e��߇l��g�}���ek�a܆i�w�駱�t�A�̔?x3  ��IDAT�^b��YٴL2
�yR�d�N:;��e��K�Rq�!2ie��t��h;tY�	�;����e��{A��B�;��ĽMal����g�F��_��EAPW�gQ�2�%��w��V|��hL{�?��'��(%w���b��	Q.U�HWf�T��er��q���S�b���Q۲B�fh�o��-)�*���2��)u�XF=�9��ŜC1�=dD��itD�*�cΧ5O	�^����5�r
!�J���w-ܝ�m����):^�Y��Vp6Ef�6��rkѻ$�Sѻ��lΤ��9�c�y�f���oM*(��1?2,e2)_���	+�5��;\3͘';e1œ~ ���uL���je|FQ��3
N��P-���F�* ����;����K����ɂ�L���+�?,]C��	���e�<V���A)� ��|�7�r|A*���3~�<�fn���$b~���Iiyu�7�@g��bE+q��2����hS�#�[m��G�Ķ����ٱ�������?������}t��� 
�f,)�fY�(�R��|j�A�B�C
̠�3kQF�z.�&��B���|�)�L��g�5{����m=L&?66o\\{FO�2�z���H�g��}���̦Y@6�+LE�ء�Z�z��`�z�S�����l�;d�螱��{�8��Ne��:���;�7v��9IE-3٨[w</P6�b���B9T�#V�/m[.M�ާ=�o��s���DE�:��A#�#��/>L����64]wf]��m?�mMlLl�v&�mۙ�v&�m��}�u��9g��]�]]���[g�֨ ���p�Z�+(i���Tߖȥ G�M�qdM��2�0'��^:x7-��R�af$eS�[���"*D_٢U����	�&uj9ad-Gv%N(BJ�J����
�ǎ��B�wh[��zZ'.u	3��c$��6:qd�l��&�%�#^��V�z��˚93�ٷ���g��Sq|ܥ	���ʦ�&�8Iz-/@<2��TG���<�߬[��X�j�jZ��U�������q~y�J4C��h��"]�j����R{rU�R��4ǣ����T��9��w�Ļ��<q�;�F^���.������LT�"� =����<4ƙ��+�����"�+1�>��T��$-�*��y�D5Vr�{�l�:�r�Ԋ±�Ey&�����1��d� u���b>�ѐ�N/�7AaU��R��o�tY1�7㻇X���pNcf�Ov>6��þ�p��wH�\��lI�`��I4�+�=�J��!p���s��ɰ�F��X8E�8�SԞ0o3Ĳ;(�w$�J�0�'�%v���
������ 9�:Lf�Wew���c)����p�"Ϟ�Ê����Xag�5&A�H�� !O=,��{�s�Лπ��.�ga#6�J�	���������-�%qH>Z���ϗ0_rP���R��٣�!��H�֛�P�E���7>�ic�����v��:w�:�I$W�kj�o�*w�[vq{��ͼDM(��ʗy(�S�}.�AO�?�p�����i2 X��MB`<���P9:�1o�}0h����6wp �4�\t]Q��@
&uUS:F��f�fD�*��y��Q�y�kSnq_�W$p�^�����Q��R����^�_�<q_�e�}�B	���N�o[3��!#b��V��.�e���	�Ȋ����~��e.�a$�j�\k�����l:�a�K�8���d�X��y��e���s���	$X��D����Y��S���p�?��B�i�)��F���Y�*
P`:RQh���e>��!�mN8�Ev��q��B6�~#����3�-F��������2�������ҟ� �R��U^��~�+�^?p�������濑B�����ݗ��o˂Y�Ws.a�J�b�Q�hT��'�]��M36�U��4C�'G���{wj��r��F���!`u����y��)U���>�a;����f#���UԚ�H6�뎛*S%�;ڼ<��3�Y<K�6��������C򬷟���d�=w͌�c����b��e��q�(_��1'@'>+�>�]�@���m2�ΜY���c*�x�z��T�S嘎���Me���Od��3ǔ���˭:h�l��1O�k%��S�:��쬧��SZ�ݾ�]?����S�ܽ�E�/�	�\4�M1��6_y���d�j���Ue1���ѐ��Z���,�j+b�4W��d�aɞ���D�����qAL\K��_@�q���s��Zn02��k�4�\�k��<6̵���[+&�$� �>���k�������� wf�:�V��>\�e���x�����*�;�M����F��g��K��;Lyk�����Fe+� 5iQ��.����4�������/1����Yj�4n*�����u*�֐��P�ɿ����w{�����ϒiF�7?=�h��.�bW:��Z��.�� ��U���ˬ1�x����Y���Ԣ
�W�ߤzB=Y�B�^_{��9|vڤ���%LuyU�e �-r��Jڷ���n����(�8��rk6��q�Aec�\�L���o�*��DP�m&O{y۹�o����8�3���Bi�H�~��P9�������/�*����3�%�#nR��ViӞ^0g�>D��,e�T�}�:�9�i,&y2��^�8x�d���4U�pQ�0��8a}�K��``������F[�2c�K�QW�n?���9�>�~?��nkw��-��������}_��}�8>�i���J�� +��L�=c
�+�X �kdw�4-�
ʘ��9I�b?F&�s��ל��本�">�IoL检�*Q�[|�ɖ����c����8�&,G��d�}wJ5
	;�#���q��t�� ��{�P��w�-a澜U�� ��@	���?z�˸KN�|�}���͜VK_�Q���?����ZE��~��}�6[���f�f��ߟ��U��0Wv���c��Ev��Q�	�YH�"�W&�W�B�xc�����RkV5�-��x���������z͊9[w�<����e�|Pi���R�<��q*�,p��*6�n������&��R��q�
�v�s�z�q��=�Uv��u��\�'�������i�H@7���I����ӱR�V�֋���q�$�+�Sw98H�t"�y���ݳ�|�@�ٴ�p�+Ŗ���P���u�m������Xzl���Jp�� ��B�m���=%����:��"������&k,4�}c��I KW���Y1�dx�O�ϓ��zM�>�zUn�Hv��/x�6�XE��S9�	O,�����PP"��i���(BZH�]l�n�"�Pnr0�i���b�o��$�Ѡ�j�Q���T��.��Ѵm�~�1>E��浱se�2^��$��w1��P�h2�Dt�oh6y��:ltL�3}P��<2����t�	�/��N�(��#x�bL�����Q��?0RI~U��?&[g�3A�� �M_F�I}7F���}a�A[m�/���ؠ�p��o�qD6-"'�_��t�_O�ze��sT�妅�t[ބ���؂v��~`��Pq�)�)��&�鄲�~�2-5ڐ�# ߫�D[��QH0�P��e~�Vy�I��C-�L��Lnk�6�a��s�7��}օX3o���b>UY�3}ف�u��ߟ�V� ްU{���@w���C�t��t^��w�*�gH���Y{iǑ0�\��~X��6�:��!�_6[�Օ3<'lߌ��>���'X�&Yy�4xOʕ�5�M�iDc���`���k�`�0qA	�7 ����I0@��w@@���'3��: �D��q6Ap��uX��R,�7qş� �N�����9{	#v$)�8���Z*��s� �������=�[�9�[yK/]���ZI����.D�܂K6�M3��,��r��G�X@lv]��.˹]f�S��T��,E�pQxོ͕K�m�'o�;7��\�1!2z_w�lN��������� ��&����v[�a����Ƀ��
�d��-J�����,�vUP�?�Av'���/-S0d�����l�2K�A�ړ���u�N�咕���N(����j]���O+"٧6�<�O�7��$ޝ���L���,^!=60��E�9��}���agM��%�O�4���b�ˁ�^b�H�{
P눻�#����v>iX3��#W�^3�_I��r���I�6�lc�����p��n�2��v�����4(i�n�d�N�ˢ�3ރ��+���Ӏ��řp.p���c3�]�b��]�5\'0���ۦ3�C.CS�k�[Ҋ(>{O�&1t�/��ȹ��f�{5'���Ϛ&h&���o�^[,.g�t4���?�cbm�P�%����X��'��ۧ�)z��
��7^��?�{�S?w�)LК�;Q:�3�z:,�13،J�toI�J���{7&1Y?���=�����%1�ޡ���V�p��Vè��M@����8��_����A�V�F)�ĸ�ު^�WՑ���*�.ܙ��h��c��|���DlJ�S}Π��ӊ����?m��,���T�&�%����������{�N�m���#_@Gc�ΙA%x�����6ɸ2���
�e�;���,��u�2庫���������~a�/x�IMyHvVb9�6�^��̨(\��O|�*���t'�l��U���=Y��?��P8g����^i?�o�Xy��3�"aZƟ;XGT-Z}����wy�f�o�侓-��Mq��lL0�R6d	�_�V��1$���i�c�OB�0a��� @b���2 ���i~*1���/�/I�M{�����O��_�y<?�xJ-DP�����qrb�G�ǂ�������:0��D6�:($�#���%X=�il	q��%���}U=�MG*/�~?�.�WQ���^w=��,��$*(?���.�����!Dq�*��NI�<��]�ǥ�T�8�7,F�i�����\�W��x^���+7{&����<�`��;@#��Ϯ�,h�/�s���K@��e���I�6U]E-�pj��a�58^$[-�3��.��e�$�������!ѫ�l�hO��91[=պ���\l�&@�u�2� %?�DX�s���bYow�����H��i��l�">V����B
�+0�[�GAKI8	�m�[�@�Q�̈́�X:Z�X#�O|B�@X�^���xwh��!M���E�q�QAsJo�e/гInv�{�������a�(Wi�5�>ig����}M:��=��b���W>�����Є�De����+TǇ�	t>;6�y��l9�F��v�6�������W$J^7K�W���`!r�Q}��%��ƶA�� �q[���� �A���M)�]�j�v���C�ڂ����ې�oS���bg7���C��|�خJ��}�h�=u?�.�E����Sr��T�ݸ*{�ݿ�%<:j�ܹ�o1i�y~5�Uq�d�D��kf���_�rAc�����śᅟT���I�}�a&|0e����?�6WN�t_Flr����1�y���?��(��f6�����7�[l�Gr#
��I+7� �Vk2~����L)��z�EG���x��W�Ӡ�~l ?�-ؕ(����Η����2"�2���ԩ��a�������(�Q�ffe�A1,�f��yj�a���5F�j=���^�ŃS�_����{|��ҎOj/ ���=�p�6�4ͫ�B�+ͬ�`��[q�MR�Z���S��gt}u�|X��2šT�W���#>� I�C�v�-�r��l'O��__q6V���N����Gw��1��x�����y���pP�Ӝ�鞐��ogiVģ�A`ZڻJ7�8��z^���H`�L74|������6E�P���GJ>DJ/\~6�]M|]`2P���q8T���lF}>�g�����6ZlFe��M�2�´�뿁�g��c�����Tڽ�z^�������s,�����|2��/
 >0�����mp��D��V���#4������ G��4�	�iC��Ԓ��tR�L������P�"�
S���ڷ�ڕ�&��<'�����{�c���t��ð.���Y2C��+r%̇�f�<�0/c����k����և���� E/-F&Pɫ�{:G�ifm�T]/����$_#��s�lBi�[��^���R�Eb$ZiF�(�#�TD�4x��F*�$�����p}��R��k�X���n��E�Gs�w҆�<���=��͚��;����e}Z���#̾�!4���)���	p<�v�0K&��\�M"G]Z���gf��?����%���7`h��.�P����m�ҵ�}v~���B�4�����Wg5���g��|6<�f_�=�i�;Ё�t`W8`}�� ����Y�۝���^f xsL�=��Y:��W�/�2햌nr�r�w���R�A�[���T�b6N�m�X>�6�.}|q�Εf��MPl�O�+�Y���R�oQ�l�U�.�H�����!8�'Fͼ"�EC����)@K֓��lY���q��H���;�^�r?+��/<տ	>Oěb ���i`�n @����`�!X�~�AFepB�04<7H���Fh�ܼ�iC���$�o��0*B`��oScU�<�K�*��8�B��Gi��'{�"��ί�+&B���V�`�j�����& Ͻi��*+�|���4e9��4a|�����������93D��;s�*-9Uܳ���$P�O�����*ίv���!��?V-:Dq�y�0�O�G�<@_>�nyo�X��D`;\L�9����xQۂ}�;T~��V@�(��4�ܰk�>��T)��1��?8kMi��Z8?A����y�D�!8�M푕�4����s�2��29�3L{>��q��3}z����8�-��L�Y=��@>�d�Eq=�BZA\\�s�;2�Zqbc�\�N�^ՃC�.�r�X��&\��ό��Q��@Eg�����DW���+!$1��P�O��9��ʟ���	����q7yi�u"���53Сz�����bs��U�:�sb,���˘\��W����!�{?5��c���Sc��y�:[>��4��Jg)�l��
�M�r���(�����&��b�@2�33�͠Q�Y���!��U����e/�\3@z[�5��4�+��MUnw/>��J�\IY�׃��z6E9<�F}ŭ���2K
��?
_��������#�lfE� #�k�^�7�&u�-�A�{5�{�ߞ�**��rI�$;=;�V�,��Z� F��/Pd@��<��6T����w��p� ���=���)�h�����'�3ٴNr�d��8=}�����Ue����?����k��t������G~�@�`;}a��){พ2ki.�R|[-,z�0�V���ex��/�2{��.D`�6��t�G�.��?ו����&$$�(2���M��l���O��2%<y~�,�s�I�i��;:d쫮C���[(�O9��KW����@�Ԛ�ݫy3nd\`��@�!V��>�XT~p�uá}sam���!*��F�� �B��2.���l��,��ȋ ��§[�7�~�YD���yj��Xn��Q��Z��ct
U׈��.�^S�g?/E����}%�	F��z������z�:���8�A7�Wg��2ݗ�E������d1z���T��(e4�#���\��a��쬧�<�~�Rٞ0e;6>�cO�8	����f ��:�y5X�R9��[ۜ?�%P�}�/�ҋ�	�Ve��]�t��!Xգ�[c�����k���!�th��c\m��	�EE�f��v��2G�R���5�1�π�vR
KJV�&2115K�T]Ϭ#I�������O��PRel1�&�On��N@c�ZcI�)���J�6��e���)��l��"�H�T�Q�V6�`ɼ&����A#��e6�!���<����Q�&;g��X��X�P*�+��˳"FOX�+��b�!L���Րd����(������p�G�.3�Uƌ�0T#f�/v�9�թ��0��|�����^+
���ud�]�,�)z�BOG���^��%y�=��'����i��u߅�*�:���1�i�ŝ�J�Tń����6 D���@�Y����&����+��(������� ����3�������L��DO�%+�½d�W�}R3;c�=2V�|��[���
�c�.�yf�B�BK-�X�А�s��s�+����MF��P����!NK�B������x�T�aӠ�Zbsݞ��:��e�%�;4�p_�v�0��ÍH�X�U���{�pa�jbi#_��	RԩybN����N�H�߼�y���"2��V���ui_�����k�X�]j8��w������F��~j{і����5��Ԅylze�S�{�P�P�9q��x�ۦ��Ɉ��ᶉ�ځhP����8\���j3g�K�c.G��h3�*W�a-W�&˦��/a-�Ȃqm~��CBZ��f�k�⦩E�5�A��10��h��&��!S��q|���t:5Lh�<8���P!�vxӻ��U]{�y�7����ЩyI��k+�&u��o�f݀��,���41�����;U����˴)9�q�1g���?��R��8a1C]����^?a�˶�� 6����WMDA؂�֟Ɲ�-�E"�W������������Ǿ�8�:��=���i�o���������|ʩ��'��,�vz�`s�(�J|lG)��џ�|u\�S��2����l������r���#.[�m9�<��%&(f���]�"#<R��o��X��1�ϥ8}�_'Mf�7��G�M�ƌ��j����*s�PR"3��	r��S��m���X����7��+���3SbV�	{ ��+
�fN��v���/�����/ΐ��Wl����SOP��_��|�)�ف���+t ��'m;�W����Ԕ'[Z���ο��h������)g�,Or�}}����~�]D?��+�fu�'���R������t���lን���< P��k"��i����jND�����$8oњ��ǐ��a��{r���r=�r�!��N���� ��Z��=�'�	��7À�x��vs&u,�Ѓ@��w����VʀS���N�)���V�h��d�C"�ĭ���m����y�7�@�N;��G����(�P�*Ćh�L��6�������;$����ʢ$�;�K�2g~�D�\�qUu�p|�*Q�]�5��8�	D����o�Yf?=gD_S�o�	΋ꮇؘ���O3&2Vi(��:+u$3��&�ځi������h���"vA'�}~,���sݏ�3�!��0����l���Eٌ����]&�9Xq�$f�]���h9`rM3�1��l6Ĉ� Pʔy����(PW[ n����u���m:6;f�q���7�0 ���B���F#�e_L#-����414.�sZ���0֙�`������VWd����kc��N�vӜ�x���
���z{Ðn�R�ya�qE%��r��q�}�,���L�j�"W<(�U��~�]�giդ4*�Wo<k�~��E+NР�g�>b�f,O������c� <�X���� į[�ѭ���1#~	ڞC��x&����{�M��	
&�d�|%�@'���^̞���"�!�|5 �	����V��y�z<�(kN�jj��p��>��`\ g�r��%�A ���y+nM�F���|.���{�I�L�-S�l�%z2a�d�f<��ǋ�<�QxY�	�%�'dn�K�-�P����֏j3�q�g�2ܿ��Y���1ط�Ƈ����#��ʻ���C:f�+ڶ�5+��C�H�ge��������}Vai���j�@ݤ�|Aw�q��K��Ҝ54&�ɣ�����)N5������{����4m�g��(`X�~r�H�H�\�����S��+P�4��ЉhM@��N�*&��o`��L�YB�����b���M5���"��׶�Ҝ��":�� u�'��[U`�_^��>_f�U���\�,V��������}Yu[
�g����a[?7��n������n�r#������F��ϣٮ[D-�O4�'j����9�^�E�O���:mwHeKB:�J�']#��e�	-yGK���I���yg�dm�9z�K'�x�����,<�t����1G�؆OE����2�:�Tj"99bDE�w������m�f��m˳���_m��1�1��Z���G<�@{kK�
.Ԩ�Eۼw�d�ctɾ��%pƃ�b�~Y�WTk��-c��
ED󰘆ou�2��]צ#*�QVK0����b-��*I1Ê	�r�+�i��1M�
9rU�hL8;�;٫�����c�^��ȴ��������a���(�}�FEiAE��h�3k�����faF���M7��Y����|�,B���)>�^�E�sU0�1_�	qrݴC�!�o��Z�2�%GRs]5/�X�]F�&>�����AX�M���g��P����[��:?3YLt���:vH{��R �C�b=%VQ��sa�^X�<U!��a�o�c������9��3��6w8v�"�Q(�\�B*�V6�\y:�ߗ�#M�o��4�>���ګ> �څf��� �����k��^����MW���p�N߸��n����A��Z#����8���ԨbFFn��mR�y�W�ǵGA� �}`���N�q�R*���L'5U,�ċW�L�ZiM��wծ#N�|���f��*�j8���ru���g�����ɚ��T>n�\��;u����q	��Ǆ[���_0FZm0��K���	���:EH�Y�G@�O����]=_���T���m�r2Z(zz�(E����>��ִ�o쨈�U�*���B ��[�lk��r4�-?��t��8�o��+'z�C_<�3�� ~@t����eveP��Ui؊#�;��B몀�^�-��Y7�:~<_G�E�*+�j4�G������s�~}r5�A� sq��z�������[��I�c�!�vhJ�����R�B�4��@G�c"�f.l�����jUbA��ݱM�����hz��ǧz�t�E��醧�N8p�!���ud��s4*�}"��b�Y<�6�S��`�����$C�(�JV�#�QD��e�TG=���W}P��tڼ�����&q���u��>�&��ڞ��dY+�|�)����&�D�_�4�L�Ԇ��9{��k��'D�	+ۼ��4����0�~��hd�u���g�{����xD�w���`j���0�(��~�޴y�Cˡ�ތ�#�w8B��!q�>X,ލ�Vz��������O�V�P���v����5�x�ٔo�rY ��&%d��X�qm/4#�PԤ[�����������K�~�V���a ��%��f��f�l�y���g��Σ��TR�gE�.�m��-�)���M�u�w��Ix�+�*��l�+�iSD>{=f�X�
/f���V����#���Ql�>���6��j0��5h��E�~��a�����z�W�����M�f{ݪ�JL�tqp+wK��]��觰�:m����2p�H1�q!s�3!9�����u�y�k�/��XZ,s_���|��Jʋ�k]5!�8�`�e�Ì����b:��~'��Nu����ʍ�ڻ�(D�
�8�x��܏�G����U��J�Fa	4j�i�`����1�L�f�P�Z�YOxĘ�B'�?���,��S�D2HR-�_���0�����a�F����jn;�r��~ʊ�Y?�Pފ��#�J�&����pe�� I8oo4MkRp�;�4��,��S���ͪ���l�����Ѭ\ ���Tc�H̦9+�R'շ7�����8���Ź��A����A�2(���F�\�;��!�4��ܯ�܋q�O�%VR�i&��!1D���~+��z�9���i���j9��_����V��0K�<�3[�9[����� L0���q�r(ڷ�m<t�φ5�=�!P��(gN�^*F����d�GN6ĺ演�Q����w˧�ޏ�j�Ӷ�Q���4�ph�L ��	��w��1����ݝ��"��.Y���$UL�R����O6߸@�=����X�˖F��@���R�!u��v�+� ��x2���(���g�͸ �qZ��P��8�	ru���-�#���~�#>��3�jC&2�@ӟGv�C��lV�w>����5UM,��+�4�M�`�h��R���4���..�I0f�?�,nT�ϖ�>4�[�<x?��}G�%U���0�D��0=馒����Y�4��t�lF������ ��k2R�Ԥ�^����GV�~���O�'�Ŗȁ{`������?=4�RzخAI����\ZCEj�ϔKϡ���_�sUX�$=�]�>;nfQoP���({��܀�l�H��՛�w���o�&��_�Aq�[�н�Iݟ��kxG����wi����F�B��KIh�o�S�Fo�����q�7xz[r�{k�˻N���@wN˂�+{q���Oui&��*ٸt#�LpŬ/���L�5���W��xبN;�W�n�'��*̗���֞�����1�*�ZnUt�h�ZӰ/ǳ
��/R� ������P$Ɋ���d�f��,K��Hj��Ll�rQp��:69������gi�c/̷�Z��K4*S�uוp	�땮qY�}kϛ���:���dD	l@g���#��E�fq��Tύq�s����KU'(���Q$��t�zws�"oh׉��F(V�MC��x��j����+Ȗ���5�j����?s����hu�,�0���=��\}=��d�
�c)>�&�����d�칤�]mҐxc^��V/tE��}t���aT�gn��~���kͪ��`����X����h��|��QGb�{9����E���cE�Z=�U�����Ø�C�C�e���K���k�0"6�d�}hʱ�}��5u��TǕ��G��\��A��K]��=��h�]�l�E�[_1+��Re�Z�ݢ�]ã�m=�]�,���
��]|l�coyiJl��	ǖ�1�VN+E����;�7$��٣#�&��`J�!bh�^���`�����IlW�0���W�3�ƺ/��q�b햢��ũ:<�MS�I��os���L����qFv��~���aDmlp:�Sۊ�pU�0���U���W�NC�d�t>I,�ě�����j��usi�O3a�1�j��gc�Z�Y�y�9c�U��mh�!�7 R�e��v��W*��<���滻J��\FrR���b/U�����*d]g��M�B(�K���L������s��'�(�A��&��=�����G��_ys���S��rW5�]+���e�J>��vI��.��MJ͒JM���F*R���[���f��+d,|Qee�B/��=kx�]���`Ѫ���9��uCX߅��k1���-y~�%k}�=�@�x�!p9�g��=��́���!��`�����'瓮�_�x^�o��@��'ұ;�u�D�oxS�rY�k�0%�g�^��>�h��=�#.U��_ay4�}��R��F?�J���}��rq�D3�BN�:���[��$���o�E�����&��d ���s�z.�7,"��������Ie�9��J2�fqLR��ņ�&�:�E��{���3ב�*���ĭJC/]��fd;��,J���\���
�5����{O�H�%>�O5���ҁA+�m�mB�8$�4�e�*}�j+�)����{��s����g�y���7��r=�z�S���pl�rϭy�z�#�׻F���[/�/f���R��m9[s-&�1��/R�%��l9�D���%
h��e۰#�u�kB��t�reM}[x5)q� '���sGӵo��R�n�|��"��)�{��;$Ӷq�m�c�Y_A���F������k��v���O�nxLg�m����"�3�*1�Z a:���I{�L��Y���kX�5���-�b	�	܃44�R�<R�׻�4؞�G_������#��͉�a�;̘���l4�ݩs$��kͮɾ�o\��� KR����v��3T8D�m꫏�Akc��TE�n�u�}�@Y?��}�� y��Z�4��c�)MG�ї:���=\�c��J��eV�� Q�	r�뢞��UʥOs��꿼���.Еo���z����t&���9/G!GJE���$�cfb�t㻗��b�(���Nɧ{�L�²��$ط2\{��	X���<�8��C��1 ����J Q�L7u�_�n�3 d���C���ݻ6�:��:���0����<�K�x9��7����w�jZTn��&�9踰a��0����ǋ�T1�����@|���8ːy�[M�Y����g:V8ݿ�f��F��[��r[�G���p��軨�y��˷����QP�ˆ���mu�3&Bf���o��d���0\A�΄V�@Ƨ�����Ӓ̋>Hg(h���Xg2�ix���}DO�4m�x%�̌H�����]-�?�Idր:NPTP�\����5�l��ѠC�YC�?:����~ޠ����u��y�y�8�$�;�+D�8����c�a�(I�h�c�;��r(Gcs@�ĵ]�+���%�`�'�>�#��4ٮ��G=��h�W��Ψ���~�~kW$	�q��x��.��� �m
Q;�V4}��,Ű�;��j�*�*��K�I�����������?�X<s��(�v����ʻ�sBA|���1��oY��}�'m۷2��f�V7�43��X�m������R��y�{�tbh>�CG/DvP�C�M#��O�at��dy�N<�ȋ� "}���L}�0�)f�� ),��0:��6C�Ҵ�N�!i����Q���d-�ؒ��x&~..]R-��/��e.����b�[�E&+�{;۾s?	I7���#P�ߡp��'�{��;�~,`x������6&Vpg�F�����\Ы|f��3W��؀��n�il��Aư��b� �j���f��k��92F��.v���ya�#I�g��m��_�*�����P�ߕ��a�^<�89"�A~*��J_��bf�Qҧ)[�i�V�+3*�z��*O���2�r��y��m�i�<,��%�྿7�Po�`�1(��O-S/�X��v{�M�]sC�zw5���Yt+7*Hb�㾤2�À�O~ZЃ����m�>%/�ZyZTw)k������K������j6��~�~>��b�@'��35��hGAB���ß�r�k� ����N�h_D�~m�g�"�$\��\�/�A�I=���\Da+���������Z�W��%�ʕ^:�I9����ȷ3eE��6�lRҹH�@16�L$�P��Gn�?�W���kh2A�^�g��$x^7!�&�������� B�LjA<��"R{^y�<��<N�U2�z�Ê����ɚ[���V�~:+��}|w�1���_ݻlߜ�XY�B�#A�,�1���'?�I4�S֝��3#���}�ヶ��k��ֹ�E! �T��?Th�'�/b�]�����R�*Vx��T��uXB0o~ ¦q�"5M�ɫ��os������%�(�Y����FU�����/��y�r��DѢ�J~ �t�{=�^��$�	��#�_�� ��E�ơ7����ҽ��#�EFn�ɸ	z:RU�oxx��X�?�06�oZ,4p��XY��~���	
�Ӈy9�%HkĄϑk�O���79� ������eK	��!Reo��a�'[l�]"��%��$�(�)A:�%����9qRl�{l^,��<r�-_v%�R3�J��2�╌'U�Oבb[�G���8�
���7+�fء68�ɅĠ#)�B��2L�6e�R��}�>Q��"�V��g1G�3I0f߶�qݱ�Cς�c�7VOS���ŬM����cy��Y����!B���ɀ�1�1�����v�����ro�Tۧ�����\�4�Ut���֣�g?��?�����\#�>�9� {���K?����s�A�����`�r��u��� h8U���)n�Y�N����R�]h�*��*�L�+�m}5���+�_��%��*u���E��9F���y��a����L.z�Yu|2fͮ�A��&D4�Z#�)�<"��䌦����'�&�A��xX����oӑ���I�FB���������5��|��0zw	t��7�N�m�{�仐Z0Z���h_����;��w��`�G��T8�O��������rZ����c"i!X�����Du~�he|�T��d�E�3\������eۏ�K⫻i�g_���ޅ|�c���mqY���Ѵ�>�*8�qX�ȠZ�f�|*Ԁ����O1��Э��O&��qᅬ!�^f8 �b���]����00�xՈz&S�HmXkU��~���w0>%qP�U8Q�.��[�*<ބN�v�Y0���xdg�����4��#L�kh��.�4����#^=Q��6�
9 ��o��L,�ߙ	k[ͳ�Z���l�CIK��]��=�zN�V3L��<# �6����/}!�(�QN�R�Gj�4ǟ��n@��w2��
�,cջM� �cRxB�ݫ�,R#)��W�m�����}bu��s��(V���?	r̴%�=�1�n�&6K�_��ˆ�=�6��Q� ��0�����%XĒ`0!W�b����[��G�Ə��=�5=&��
���pL��}��a/���!�b���H���/(�('�,d<��hϏ8�0�b�2�ڶ&dݧޛ�s@T�H+�$,t��2K��G�X�^EMcFv��d&2ۂ�eYM�8ZI7=In�D���7,�'\KXŐ��qa�6�^���V���.s�Z���t˜S}�����@��#�b ߖ���it?�ca�cp�_�D��"Q0�Ӏ�*�DE˴���qA g��@��a��Z��Jd`�d�X
����bP�W�4�����2�!H������c(��hS��+Z3q�U����� w@��n����\OY�LADٔ[��fQ �L�Q���OU�2->�ӅvvW����4�T�X�Ey�۵�F�  �Z�v��V^���Y{����Wsº�����
��xd~CP����_��o��%�y�J��E���s��t�Iv�'z͍���f7����,A,��/���Dd(�AA��Z߂~�<&�D�%5��<��|&a�����`��]۠�2޲�y�t~j<�9~��G�?��!�9�Aa����@(�L	�~���g��:7L�/�����u
<
R���
$x3���y��Vt22���KVy}j���-[��p�p�1�Ⱥ�{X��֮;2��<�kj�nU��=�=ϩ]�O�m`�f[�n�]#��Eg��������wXc*�����!������#E���	���z�B�&�C`-!gT<R1 ��5��>���;�$�9x�+^a�������L�=�8�ą�llv���\�M��#�o��j]�!2�r��R�����G�M��N�`3#��f��M���|��ށ怍MYo}�rJ(�E� �α��T3L8��K_�R�`�6�5���aY�z���\*[<o5ptʔ�n8,�V<�%���_�<��4��7�:�vf����>�-�3r� �+{��m��͙�O���3[�G�-�G��jj���P���d{hƼ�E�r�adF8�9�}���۷��-74y_���}�Z�t{_Z�u�Mo�2	��]`�Lf���X��h�Vv�5��cc��z��|�� Z���B�O1AM��!�������P��[�/n��-�#��=�	N�t��!�ʱXt�1���!!�b�ϳ��*��k-Oc�m@$��!$��eW �to���ޏv��ɺs��/��pZoI�4�lr|4}w�W����񬍏��/����DBXR��{3�\����,��莴Ӈ�w�Y}")��	� ���Ζ'��{��~�j�P'��C��/��,Yk|���kr���it$��);�3=�り��[�¿��7��u:N��{���`/������$O��g�����=��cNGcA���:�l��5���Kq��|��ڱ���Vڐ�)�zc��}��!��s
�}AG��-��`�}�L���y>b��#.�����0"�0B.������9��KC��]��{P��W�rn?�!��7�e�gX'S�j�6h͵����*�{+c�����~���dm*��]����G��~��Ie̜Y���=z\���G��O"�/��iC1�\��U�����{p�~Z�>zZ�s戮�?fc�۝�99Ѱ�;��W������^ ���[y�,S�L�{���66���$ͫ��t/ɣL
��(�t\#��N^��K�FQ��=���	.���l'	��K;(6����l�F�;�jW�ȚfRV�&�~����g0�>�\;㌳|--_���~�/�Z��[=�����z�pݢ���Kie������<+=��/�'�x��=i�֘�x��~���i�G���k��u{�K/�3�8�'��LJ0^%6q�#�8>�h��y��z �\&kQ��9F���0�s�(x/�|��f�tfs�����+�'E�8�<		љD�0d��#�,�ى���Dƙ���	2}�����"h.�c]����'�*g�9����SXO\O�qRP�!�JO��ݺ�lw$���k֬����:A�48ɡL�v�u_K�`�v��Q+�j�Z�CIy�%,�q�fV�U�
��u�s��DY!���R�>b~���M�/��j�aOm|����$�������Z��{vϝ��ӛ��W��5�`�,�+���6=����;�\�4�^�[�'ּ"�g�y��Y��v��e�n�d�c�����Aa��Z���i�sɲ۽{�v<7f�z�o��N;ͅ<�:mv�8)��đ�O�=c��G}����SP��^h��bzc��a(��"E6&�D�+:^��oi^��
�J(K��<���{��X4�!�ň��D4}�<���P�U����,&������,�邔�o��	�$^5���=��g���V�В�[�K�,K�g��O�ã�+	҉�,ڪ������d�����7����[*��wK�Sʼ�bm{�(��L#sK�Z#����#���_�`4�~ޒ����lI�'á���NL5l|l�x����/��b�y�a�=>əg���9`�����F=��Sltt��4��v;��c�ϱIP?bc��aU|a�	�vW���^���y�l�&y�{��]�轉r �o��o�k�q%��_~���D)�S�_����z�������S �K�ySB�	�L�
D^�ޏ�:#�^�}��)&��K�Y��)DhH�9����~
$G��5�ZP����5�,}��r����j(�e�A���-]���E�7�9� `hi��p�+4iY�4���\�w��6>9���@s�.���|{����o[���M�Y�E�N�sK'.�c�ȹ^}�7/c��/��7��G{ ]�|�z{����y1��Fmْ��s�6Wp?���SN����8RJ���;��x��"��^��zp	E��&�k����㫛6=n'��Q�  Iԝ?6e��
o��+��	�V� ��!������+^��g�@�cA��Dt��3ͭd��1��s��`},IA�����;���nd53g��&�R�c<� :�,���{#<����^S���XF� ��^��cnH���J�f�zbI���z����FV§�,ٵI�Z�ɾ2'Tp�����xF�M{?aɲ�~��oM�=̓�H��MP4��BL��t�������[�P\�Z����˿��EO)O��}��=��ԭ�uĞ���C���ڱǮ��kץgٲ�RSHG��/������?��O�|9�c�Gy��]s�=����L{K�]�¿Y��I��o��>�����b=�١���1�oƴq�&���O�p�|�^m^�
����GP\w�u�pp�	��A��c�wdg7�e���)��i�,Y�9FPJ����`+�+�N�U�Gʇ��U%�c^�6wL ����v�9��>�����=|c��{��v�c>�l���";e�J���,�Z���w��$�̂�N.�'y%����+��!��'��K���=�c�-s��R�J�����h�t\XK�����+�}��;�<��_�U���߁��xd�>�{�;����Xc�'Ň	�Ï�pX:��k}�<���#�<˕����ֻ��kiM4m��U��bMD�g�߳k�E/�{�RK��N�/��/fN�&βɫU��M��L<15Tw#�*���~�!*7��]�C?��ُ������U�)������o~�uW6�V|x	��M�yC�K(F�����G e�g�}U��0�!�!(F8�KxpN>ˉs����j� ��x&h15��"ry-}R|�+X�E]P��-���پ!�)}���\��,K�VYe`iV��<@\*W���=͖F��e{���k���L^t0��̋�5�I���l`pvڵM��Gg<%2�.��b�l��̅�#HX��G�I[X�R�j�����x.�:�H�7�CN�����d-M�-}O�^�ٞeH�B�]�¿ԍ��*����X�: ����g7�p'����崨�_ZN�C�)�Sw�Kբ��Ұ�y�L=�gV��63������{��`�j�� ��m���C�6�K6Y���ñ��?��O��uϐU-Z]�dp�^�7��ω�zXj��y�!�����*՟s�z,�qy��g	l��ܛ�N�.���k�\�"8�S2��jȒ�a�wZ}����R^A���t:o١���cɫ~����d�[�:hO<��Tyi�HR,��Z�]���\�YO$܋�U��F�9w{�x���퓶eێ,�ײd��h�;7Hs)��%�!N<�g�<���c����ەQ���	JY���+�{/�rqT�Ȓe��z��}�6[�r�mٱ����X��?MvO�<�Mأ�<��Q�O�Y}hZ��41#Vo���I�Q�vȊ[�{ܶl��欳�*�Rzy*�Y,,=6���h�(h�U��%�����C�YA�K/����R�S~A�?C�y��emɲV�%����0�����<G)��ȸ��T4N�:k
1���m�g!l����E0Od�Ha�}����׾6S@�v{S���ط��9$3U���-��cTbw����{�/�R��ozf��6����$,���t/O��q��$�К�q����K�+��4�7���j'�u*���i%H�^�mS3�k_��~����!��!�0(š����S	���^����d��x\�5�j������������gmbr�ο�,[vH2PmԞ���m����M�:)�4�?����W�>�,b��|�N8~��%����`��w�m~v�'bd1�J	����$�e�~�!�iXlR�{UeѼ���׼�5E/-"ea�qם�����w�/���b���nk�^�\�1cFA�Nn~dIȃY�A�J��>:���]*��f�!Ų!�.�Z�*8'�qxZS|E �q~��
���.���u��攋��4#�gF�TBV�ٰFS �j*F�ߔ���>�{d���`�Y�9��\��_~V�� u�/��H��V 1�+��d�`(�����v�/���7���������=H&�u�]^:f�-v���m�s������� O�֬]jûFl鲕����;�زQ{�)'y�J�����{�"ٞ�w�V�|`
���/�������ڹ��V�X�A��?�v�x��ȳ��5�竖���O{�����t����n!)���f�����G�f�����ۋE<:8vHX��M�9<2���Z�I��Z����I�߼�< ,��2�ʊ%H1��t}X���Y7���i���~,�s�<M���m
�CP�9�
�P6 K���R!���� �(2V�q��hgҔ؞`��d�QnA0L��GP6��J���������B��[@!R:3ɽr� �m\ż�H���Y��{��
 ���y��fB��Տ��Gp�q��e�t�HoH�߿�6=�ɦ&F��Y5�Om�dK�bkWeW\v^:~m�%{��-�u�D��c��V���0�)�΃�~�;��;���68�o�#%;��b��m�=�̟&�1�S;����/��ի�M07�ζ�~���{��%�\�A ��x�^np�7���H��3�����CPV0�1�X*���rW�f;�uZ���`I#�# �sqNA>���'��Pք���
^T^�M�`
�F�c|�-�׃����HB�\^zd�]�Cu��$�"b4��HT5U��,����e��T:�j�2ku�Y�	b��
���\��_��@��h͕ 17����+#����}
멼6�!�Q̳�#5d�w��;~�*k��ǜh��%v����Ș=��öb�!�b�Jמ�^t�u�zOv���w�{]R��ҵ``�|X��?���ߦ�\���j؏�3_�o|��m�в���^}�v�k^�Y�XC�w+gk�0, ������X�:��l@(�#��f0-66�~i�}pt�hl`6�\|��W�R�� ���H��Њx�b%|q.� C���C�V�`����Q�]���cbd��^QQ1B���׃�y{H1Q�2��}��z�R�S
��5������x��&-�
�ߖ��
�>]h7m�׳�Sn��f��?�{�
Q��r� �4�����9�������x�}~��󁒅�)
hdW)��*����y���=j+Vn������7$I']���G���F���/����v�=^�F��}�.~��*���MF�ʕ�=SʉA�����ܶ���.��O~I�*��<0�ԅ���pM�5��޻��	"�N�j2�l(�?�я��� Y���{.��U�����V7�F��o}�L��_�Ln�R0@��ɳֹ�{�O��;b���� ,tq��W�0G(`�5BT� %֮����`ۇ�r�b&�cP\��(^��W�ҹ�%%a�V?�60���<R�5@���D����Kmf0�C@y=�v\K���;�tx)�������f}�|�H�-r �=���Tn�09<(]�9�F~^$L);/�9^��o;���]l�Y�k�C������u#6�d��عծ��Z��G7gl�ь-V��3�X�¿�h:elddgf���&�s��o?��v{��G�\
�أ�v�N�e$�fvo��6{���{,�F�SD�����?�C��h������KH0x������_��p�YXjxp,�P�U��SO=5#t����'�E#�폘?CBRyZ��Ǆ)�}h�cP] �t>����G���,�I�F�JHIgA������>Q,JTV��;:��l�{�<���e ;���ؙ?�Y��Z���]�ᡒ��l��{��b|y�f?.|N�X�>�6bM$����I�p>���"���gV�����x��<w��7��	���o�=���u��?~��vc�ݲ�5��!�n����o۾��ȕ(��G���4�����7�X�¿U�N�ECg���W+W������2͎����h��@ڠ�b�U�z@ic0�X]*��q��;������)AE`"(������2 8�`a������M&�Q���+P+H�y��3��$P	�ך`�F0 x���q|��W0v�S+�22��Jb�7V������J̍TO�Ž3��4�P�PD=�{�k��_�F���t�l<��P*,��&� �C� g��A��R#h9{�����,���m�pD~�1��1xy��{���+	�������A����	ni�3��k_��?+�Eo՘nb��ݶcǮ�HH߅g�{x��T�̳Ƣ��GZ�Su���H��#ɵ���0=�:����i4������d�Q.��=���ܥF��D��44�����C��O��Ii0�0��#���M��N�'V��KL@��|�`�`�tB[X�k�軕���=�ǜ	A&*��?����x\k�vQ/���:��(�I�3ޟ(��B&+�*�C,��;dH �r�:����J9w
�%�Z>
�b����l���P�]�>?��`l���<���i6
%��(XS�\�6��9y/���l�|9+�9W2W��Ox6q9�}��H�s�4ʘ+Z"��K1���z`�(N
7�����=�����q��栘�A���G����"T��0XC��Qʆ�c+}e9S=�S��J��l�����d�Q|�+��E���z��ڸ����"b��lŅ"�7�\��K�D���E����BK�Pcq2Q�|sV�s:�>�wxE
^
�%h�������l��#��m(kz	d+�h���E�b09���e�k>�<�%)��ȥ㣱 ����ܷ�T�,�u�NA���	���me4�y_��tEPˍ�z1z���3V#.�>/�@7�̸�*<s*�:-�ޚv]{;b�yUڧĀ����@�����1��`��=�{�̣R����{��E/�{|go=���:Ӛ��6��?�y���aU��� �������>p�c[m4-�H-�9��mp�Z��d��ǾЖ�(��k�z�k#d�=�Ȣ�A���	�U�G-9x�U�E�by���Cשu��v�ɳ�x�X-�	%Pe���B��!ڦbU�������*��"�\D�z2��s9�`�}�&���aȋ�E�m�Iq�kjgHO�=���sYM����ڰg)�c�՜^uS�o��ٵ�bn�*Y���y���g3��s���]3g�*F�gV���_��{4g��sE�\Q��C@������r6�,G~�{�.J^l�.�@�p�v��mp>��N(`(��B`b�r���c"�Y�);ݫ��7�����b��u������0�O|�^�G���m.���:�_��`4����r�3zF������3|�*��8A8�Y�4AN�֕
�EA$�&!��w�N~9,�}ҋ�O<+hܫ��")
	J�U�b�n�2%1��IyZ���htXx����{�}�D͌*]��_aD�b��wQ?�)�U`����^������(�p�	�qi�,��YQ��ͭ@��T6%���*�Å`.�bC��Ҩ'X����õ��׮T�,��χ�/Z�P���8��hY*Q}%��g(�B0	�/���S���΋*M�0�CL��9kPP�2�uY������Py�����0�C�`�x�:��T`�)I{gEC��P�Vre�r$�cs)<�K���>JvblԿ��#��ƾ�[�x��5��PW�\�}�'�۾랻3je���3��"�.���yD�;����l��!o�y���G/�f�8��6�bD���m�շSC�J�Q�`�K	6Zp��TS�H6�m����h������X��}uǠ����Z����9����{#���|
�	�ݟ�{�C�A@$zqR"�^),	�s�~�o5fU�k@h��#HBВbGz�N��ۇ���w_	y1�$�4���nCumtm�l��~V�.�1R#���l�[]���%̹�Q���L+y�*q+�F2���^�c����X�¿���L?�g�5�.�Y��̔�� WPM�{��e9�/�_~Yb����f=��n�%��X�,/p�a�~-��u���L��r�|׎�UU�.s��9O�%Bϟ �,8��g�u�c�	�^��ye5*CT8�����$o	+��V6��:�X&b�ț��8ߍU�^��"�7]�O�S�A��P�N���X�VJ���,"�:���n�R�i/��k428�k5g�Y�	���3�� �C����V��a|1�C���ǿ�س��L	�1��o�/{�m[3=���L��5���Fĕf�`�j�ֺ,5Yڰlq�%P}��zo�XbX�.��r�^
v�M�0�F�L���k�cD�������� Ās'�R����}|��T�-*{�C�,oi#{GX3��n��_�ñ�,)�5)%� Vf0�ٯ��
Q��x��̫n�W�)�:8/�'�*,~h��>�=�r�6���a���O#�Ә��i�hOkϪ+\�w]�n�gX��sؓs�\ا��nf��T(ɐM�H�|�g`��|�X��h�S��j�K�F�/��P.qt�5�����V[xE����,#]�R� ��\ӔM��H@ĎO�4v��=]C'��=Yt�0�|C|�j�p����eD;��g��֊���1�1� n�Ź8V5���9��5[��,~,v?�FLYE ��T�?*w5v���X�3i���"���nR�P �:c�X������in����U��e�4��_�1�O�gQ.�Oĩ��L��֥�2
}]���u龳}���~n�Cy>�d���6�!��"_ �����@E�^���}(�P�fV�X����f�)�x�q'dV�Ĥ�G�mٚg�V����%�!+�����Z�F
c''��-vX�q�j�+`k�hQw~N���3a�^�NX�ҧ�PbP�G���GB!2g����PB�y��+K�90����a%_͵ܶ�έ��3W醨�Y#@�
��<�	U�Gx2��O��ד>��se�F>�=q�W\qEf�4��`�S������z) )�+�9w�~�扌d 73A��׭�ViZޅ�����K���~R�=8_�z���'��1���^�-҃Y'�p�y��g��@V�i��K�����
`��V�'C�4��7N5	��1�:'/y�K���3���)�:�&��d�y���'K^�	.&.��O>�j��~{��fcSD
!�[����`Y1�Ŭͤ���)dU����GL#Y��F���QK�G&	#*3)C	����!O#&��߅V 
�I�<"�F�Ne�
��^P"�G�\
E]��1>7�^BZ��V�̺&���:G������JT��!��2�״6���:�����9���z
ȫ%�Kq�n�[�Qݓ�Kk�כ-���u�s��j�+�"3$�5�2���G��^��N8�=ϥK�����n_?��Ńv������lyY�9�t>p3|���U�gVOQOG����|�7\��H�HL��f��V��&k��u�i��op��L:�~��~�7��_���\i\{���]Dlu&�Lc�4{�N7d�kX��%������Ɋ��YC����Z�Ŏ����N��ڬ�.��(����u-<�d������,AS���z��u%���6��/(2zCR���o��0^BK]���u�μ�V�iD���T�UDl����Dh'Z�b��we�f���lC��O����~ �uZ��W��(���!&���d`R���3�p�oȕv53��9�l����䦧�_�G7 �U"�P	t_Ǣ�y	�YI!�Ed�j|/��"��񤝫e\�qۼ#�j�e98X�ɴAN9�$[�f�O�����ª�P��K�����|�7ۿ��������^�Sة�	Pa�sI�P	C_MA�� ���1K! ^��C�G�j)���'�
�ٯ�r�3v��,x���_��(���Θ��/
�s�]�ys�L��zI ꘨e`Ȼ�=d#D�s�L*Qu�����y]�	����n/?�ZPRН���Q�1`�ƺ֩F����Y�KAc=��&
\x5Z����4��a��⾋Ɣ<���Ø@���կ����J¨lN��(�8͂$���ڵӖ,�����>�[�/|�Kɀ�ϖ-Yj��#��q_Ǣ������˽�����^��+��9�H���n���Y�W�\�=8O?�,��<X)Z+^�	D)<��#>���_����|�#^��f,���� ?�5��׆CyQ%/C�v(�'�9��~�(9~t/j΢���5����lV,,e��������Q�Œ��$ "�����qi.��z�h�Ȑ0��=�/Z�<�JR�1�'��R*�������R��bs�H�t��Z�E%�EZ�s��'[U+E�YJ^�+���q�6"�罠���@m�7%�̟����c�~�^ӱm<\0��z��ב��нy	���0������R���7�>	~��~��6nz�n�����;}n���=�<[��P'�,Y:h�~���_����^��A��v[�¿Ճ�59Q�`��]#v�1G����d}�U�?�arٶ�q��Yv
��/�ݞ|�q;�e�Y��RW_|�G5jg!bI���p!I����ۇ?�a{����3ZGmj�|�6��(l�}"@X�����k\�h�	o]�g��9Z�q=>��X�jT@�8�\	&Q��[B^TG0N~7z�Xx��6*�X/E����xu�*1���u�־p`�S�]T�A�-���y=Blj���C�3&�˜0W�a���=�X�ū 2ǣ�E!U��FC�q�Z�_/��@�+��(
���e�����'wq-Y���;�1��3'W"(��<m۶=�s�C�����h��=�y�k�A%��g��w���2I {n�3v˭?���m鐕�%{��_�5�����^w���V��UW������vNI��Ƣ����dc��\ȍ��N��m|�Qk�ǒ��O�t�UrL��o�޴�׶l��w��}�ݑ D�M(�#��F�W4<�dY�
|F7�׈L�N�!��M��T�b�Y���М�sa��@8F��x��
�,S�	�X$���*!#Ꟛ���D�I�="^�Z�RFX��	<:���l7�' K[ޒ���.��_�3w�F���������q��3��U0a���jq]��՝{���7�!�-4�5�>��Ϻ��� �8���q��<��Ig������ܙ�+�?�
�zQE�������o�o�q���\��1��?�>�[�y=��Rԭ�1{v�S�s�6[���zkmbr��Z��}�����ˮx��AA�u�v��?rJ�/�K�3&��Y�kIz��^nL$��u߽ގ>v��o8̞����L�?ɽ��)�oO�J��Э?�Ņ��ظ��8{j㦢 ����)�.���B�_����n�tz	8Q��^GFE�5�G�g)XJ��\��,>5���*����BB%$T�����e&�@4Eᘂn�#��`�ApR�k��vX��/4癝3ǡ����i�iw&�u+w���Y�\�փ:o���v*�^�J=(ʔ�����&R�������|�yWp;��el(�4>9QԧaD�c�F��@�ր��+Z���״�bn���]�J��v:xql�O!�F�<CFRr����oذ�~�#u���o*�;��Uo}�-Zb_��W=��o
k�b�z�+���+�mz�qk��؉돰'7>��~��F&_���-�����V;�S�_���Jo��hvx��@�������;��;�V�\�&��I_���u�G���6�`�)X�� [��1�,(K���kXO?���@*��𖷼�q>�,����?m?���E@/�ᴐz�N�Yt�8{W���B� ��,�����o˞��>�@R���^�Ғ��+!
S�uH�I���|�>�];-���k�gAO,�p�^Z�zL�L�Z�+��|�[���gd�Ǻ2���	B�������&6̹+�r�5��	2�ٹƤf*lV.5�&�������A��KVt	k_�����s�X�b)
����?���Z+���~��N㦮����<�����{ϝ��C�@J@�S@E�����T� ƭ�2h��� qd�	':DM< ��g6�A��+Ib��v�����R�d�?��S��-�m�&3�Y�T�R���L��h7�@X
Fbc��	�b�}�;�q� |�w�w��?�)��Ul ыJ7pd��������H�0J���	�$�)��<�J����ıD#J���P��I��@4��D.��1"�U�
���+���������;Q���>fbGVH�̙�ye�:� �ǅ�G9K�k��(
�v>g����g�W+X'*9-�W���fce־_���ݳ�{+�L�]O��:��ÿć~x��n��!��e�ā~YGxyt��|k�����m���y�!i�ҟ���N��O�s��=���o��VK�x]�\Ǣ��L_���0D��rˊ��Ov�����I�*-��!��X�C8��t�y�{�:��ƥ�'-ߨ�N]{�L��@Y�)��ׁ���
03x��4���V=�$P�(�)I	+}w��kr���B�\��b�;RW�rHiʒ�	Uz��+��>���6��ˡ5֔<��{���k� �
d���?� /�Y�����%����,�)gP� a�
���Q.�z9Nީ�J�=�L[6� �`���c��BI,��3�bє�u�O>n�F,@�%�� �D���-PE��O�S��4��i}Y����<:�ÿ������OL+s�)�ۈ����i�>����l��z�ȏ9f��t#�+K"�L���db}9������H�Q�H���l �"�;�3N����Z�!��|���ǚ�lv�HmhY�F��1�����Y��7R�$@�����R�n�SѱN��G^�8�ԘG!J�1����������6S�������P�q�ְU���yMA^�Q�C8��"��d2�R�z�/(���oֺ�ː�I�����?��X�)L)��-TF�c���$���O�q���-�׫^~�S�K��p��ۿ�A�w���M��w�y������>�o�!���[Cs��_s!�m՛S6���Z��rr �ג���2���Ĩ�5�!f��9�E/�ͺ�wgg3`~�a�j�a�;�OѶZ�VV����Ln��'m�ݾ!�p�$&M�*�t~YbJ�<� �"ZR���lC�����`���q 1��6	l,D-N����q�����=���c�^��V]A��y��"�^����%mJ1pH���+Ȅ��f������^�g.�_�M=7��
ݕ��uQ2���Aq��0ψ��=A2~e�j]�X��o8Ya{�F#�k����xĠ�����i�=͵�Ѿ�Rkv�L���mHc��{�s���W�ʧ���8X~�m���<;�XO��������X�3C�������,����lt��ɦ�|��>gcim�Tdh�
�&E2�\�¿٣����l���^y�����s^�lOۮ��l�����F�(��Z�R[����a[w�R��#I�[�8�2�#�KO,�E1(
�ن,���`U�W�_�;���}T���X���r��bPL�t�$KV�
���A��C�Kx�*����v�������n�M*�D�LP������υ�h��f=��1��
��2�A�1j )���`p>QL���QS�L�Ab�b���s����]��cnj��r�v�ry�z��0�-�=�N�n1�00�{���!}�!;�%��3���۞�F�φ��:��4�v�I�أ�lLϻ�pF_2F�3��w�O�&����;��9�i��g.8��$�WZ�@5�W#���:�t�?�g�Ɇsp)�v��.*0m&���l0�?��?م^XP�b���G{���ͯ`�\��%p�0�YE���>��f�9����H��s(���C�0F֢��V\��͓!�\�AyX/�>�5<��"��h���6?���$%X��P�e�� �,ƙ���A����H!w
"�Oтǻ�F��Z;����C���ľ�,��̚��o��33��o�s��&�^�9��3��潔@l���-oՍ��z�a)~�'��7���>��[�;e0�&Ӽ�\u��ܽ+}~�m����J�犲�f�d�Ye�^v�{�z�<{�F�����/�Z����'�BIf�;��~�n��&��5�Nx��:f�/͝���'7�3<n�rՎ8�(;��uv�y'���MǺb�p��^z�M7��"�gS1�K��B8W���Eb)0���lB9&����|�7C��K��{D����uQ�-o"R�Ua�XH1��x��l�wO O-��cEHE�L	��6��Y�M���3R��m	r��P�;��g�a�8����D&�����W1�"~��dp>�����`�2�*�9���i���b^�_s=)�Z����z^ܭ4͢oN���\���zT��*ʹ���
쿈�NRӿ�����\�h�����/
�ꫯ����ﴖ�<;��+��,	�I[��4۹}�y�i72��ɲ">s\20/����~�	�������n�G~�ȍ�t�N���*�¿�G�Y0Z��ot,���K�y�?�X{��׻u����/�ڵ�rNu�l�L�S����X�r�� ���o���_��c�4��;X߸���o��"�3\�cb�	A+,D0bY��,�IٿwW����/���<#a؂��6�%Z$�*�~�И����?
��Y�<�'��7T3ch�ƫ��x��3mB�<X���_u��.R�,e�
�g�x�j��8֥�-1+���3��^�?�x�.�����Ox�bŚFsabE���B��B�%��J���L�dk[sR}�ݾG�K��BŖF+�q�Y){���m���Sݽ�^^����~eE�&`�}�_�ߏS�eyƬk%H*7C�c�Ĺ�/�ܾ��>�ev�y/�����)o��x����������lȊ�ױ�/�>�wı��Ѧ��g>�Y����� �v�����8*���6:Fᬺm߾���o�օ��ZL�����x���������.� ѧ>�)_���]��ψPL��Ŧ������ fHH��8� A�(PX��s��糲U�AHΏb�R���
���:�%���M���D�,T�AX�|��2�D%�
�1)�z��_��_�k/%ſ*PƘ�k-v��Ǫu�kS��
�	$�.a�3D)�9X�Ϫ�C�T�����JaP���_��`!�i��>A�F�!���"��`��H��9�%T�NtL�@5��`�:�t�&.������d��Y�ֱ��ã��̳ٺ�r���2�;STޑ�zŹx�=O����\��x�rX �7q�o��^%��K.��Q�s�)g�`�LN��̵>�����{F��j�k��V��_Gg@�QY����W�CP_p�Ey�⩂~���?�1woQ�E4K9Y0X����Q�෾�-�.��B/�@�@��
D�E��3,y0,BY�
؉��*E	E�D�Q�/����|��F��.=��r�=�C�"����@
�r��'b�,4��7j̑� L@����ΪT�EtI��Z�ipN�s�)���2�J��9�[��*!+[qU�d�c+P��c��cL`�!E�ʶܻ����c���x/�"&҈�(�]p~��'ltx�=���6�kGz�n�[��R�"@#W�<�,�Q돷#�8�cqO'��^zzs�-͗,�93�=�,�'��X����Po��@�-�l1��s�v�w��x��_�m���a�g񙆓���k�X��sN��?�Yͥ��q��/u���d��M�\饎�e�Ъm|j�mݶݾ���x���k4�%0>�Sݙ�����
�J(�E#�x��21�*( b��JP0*-�6�'˓E�LD%)H(]TQ����'�������#��Y"A�� )$��n���V(�eM�_�X�!���w�k�Ϝ��{|���3a�#`e�G�q���C�Q"�N����wz%��x��ށ��4Шp����5�Dzyg�\u}�A�ɱQ+7�WI�F_��+�Y�MU�-�D���X�]J
#c�4�mE��h�s)�/+�s~��l��r�AG�^�L���y��
2�JwH���o�F�G���xR����p���y*s��N�j#���x����e��RT�^�+YU$`d�{˃+�mg�wʭd�!�x��;�g�UC�e�C�^u�U�(O;�4�H���T���&�5r���| )��X�vK�ɢs#���d��'���|*=��Q�?�ѹ7�AX��? �]V��V�zY��k�J�Z�~��`���)� L^������)oa��TyS��UDN�[q<[�?XW*/�h�9��b�sC(���'��@&�kdl���wHA�
*l���E���~4�C�.���%i�٤��[�}W�fΓ���̠R��M���ʜ���{ �v����6��=���J@g>�|�W�*&�{docpѷ� �bzzf�ڱ?y��2�3Y�6=�%�S�!����݋�S{h�sT���g.̸R�t`Z��m�ˈuWD�t�%�_�k�� ���`���`�F<�k`�I������E���'?�Iߔ�A�p��?~-W,�����W�v&�)���,PY���c��|4�N� ת�c���`�^\R�����p�E�YpLE�8�0Q#m�K s�Yo�f��|.�iމw���L#�de%�u��iK��ol�+v�0�N\~=o�yQ�D�7oRק����T�X��x����p�u�0o��$�T�GU,X�s�%�e��X7F��l ��{s[�)7�j�	�d�I�yyh��@溪bB�AmdD�����y}��_�}N�7���������̟�nȐf��J_�&��V�Oϴ�ɣ��~�ûlp(y����ʔ 6��F�$���&K���6Z�"�~�E���f��d��m�z���K�1���R&,����� e! (���O���-n�IH�d��h�h}Ja��#��%oɲT0W�Q�'z�+�:f�"�x�AB���E� �K����0R�N�
��F0�@�R�Q)1
Aל�ZKi)�b&���<������H�a0�7��%�5=	 ֔�y�����l#�1⻕�a�r���I!���g#�-r���X\�ۂ�Ӝ�f�Y�i�%%�%~a�;%t2p}U��t~�Ԫ��!*�8�W^��ɑ<!ŋX׼Ϗg�潒�HX@`��dՍ��'m`{��J�V�Z���I(Zg2L���Қ�� ��}5�x���du��Cm�ܵ,{i��H��Rő4��0�O����[9_p�^��w�>������M�{d�S�c�,�����˳keMŠ��T HG�B��x��rs�Yd[%�D�dh�r܇(�x*׀`'\�d�q�QF��D��7�hΫz4�.bYDG*cy��[FgPS��C}�f�u3�ۿ��΍����s����<+�*q� ����ׯ/�S�]�j��bs
&� �G��<)��R"XΚq6K~OJ��[�E\ks�,b,"Χ��2�ߨ߇ ���N�C�VL��<MQm�3�۩�1���<��|��6F��~��Y�H}���+�$x�PQ��<��QfK���0�־A��\��G^�d��3{�g���y������_,�i*��^|��2�a����^_0L',"�}ڵ�r������z,��c�,LYw�?`���>���x�*� �BP����[��#�&��,J���Hu�`�}�m�y�G�x�l��1"J�P̭�%�n���@���8V����͛zK��,TxO��I�L��Qָ�4t����Cl.�A�~���$�8�g*�=�f#)����ߏP�{E�¸)&#o&��ϕ���܇��R�ϲ���D�p~]��}���o~ӫ���?�q��C?���eĐ��׬C�劯!�F�}��1z����ح�0�j@��EL9��큪�k���/��/�ܲC��h���;d9��Դ���zt�&�F<9v������mL�(j�oh��Q�H���΋�#.f�
��&P�Y׫�$�#g_�X�F�'���{���s&�G���*X-���P�^��+Y[H��!K�&^��Y�xK(�X�ZZ��-?x(O�q*)A^S�G,I0SPV����-Ԑ��<f�S4�͖�"���ͽ���*�`����-'k�Y�y��5���%zp{��kDa��%(��vT�Z�>�`1����6<�*��Zӕ���j�i,k��f2�H���HY��}/�r`F��e){������Y<\�@PDw�!�u^4%ܦg��R�����9GW<ZȲ��Q��b���$���~���K(�]�ML:k��_���;��$�:�[c�}_�sӼ�p��7�SA���@y�E���yw>/A"��WF�^cJTQi���s�j:�֞����4�߹���ӳ�wLcy%�G�n=�z#=���*"��6K�P�-*W�,�w�`�����<:��)���Bs~���x��PL��D�P��zS��s�[ƙ���dzɍ�"�n�1�:iN��|��¿���5���6y�	(հ�ZY<�'�]�/��z����fV�g�D	�J�m1���[�i"�:V,�SP�S��'���}ˊτW5�κ?1o�㗒yH�JTN��,��Y�m����ڟ�=�OV���b���)�d1���O|��1�S<��D�%�y���He��;��G'$ة����^�������b�u�T��'w`b�&Y��$k�{�f]�X_{&y1��z#�1�ǲ� � ��ڂ�<�k��;h>y�R��baC`��@�xn������9�Cc/0�����F/2����,��=���X�¿�m�6��$,�k?:U��m¶թ��6Fw�7c\0b�t
�ο�ń�4�C����F^�������5�f�ĲuQ�IE���_�F+��F�ә{=�,�Ҷ�ע��:b#��<���&�'���a�#�FU�-�!VL�W��(/NTP�(����� ����wu
���9у/L� d��Ne;�!ť� \1��S6����,߱d=[s2��	�	/�W�Z�!�\[�j�-]�̃��t<����.�O��ؒ�����Plѧ�*%�h�id�Ǖ8D��g0t��)���d�������`�9`���E�pl������/{���DV�m鲥>�Ln?cc�6�d���Es���
�B6�Ц-0�N�W>.Ta�L	�t���(�'�vۣIVP�s�⎐N���Y�A�N��Xݓ����+u!GTz��Fe�n��4���M"B�����.��~XX�w8�o�D��9����w���{^ÇzD�b�������\���y]kGA�R��	r�	�ס:R
x�� 
 S���p����jVճ����o��=�P�m�>b�G��i�
��*�G������|Kqʛ�BVv;����$����iLi������u�o$'��%�<1��o��\����y��'-+����ױ�k�n���vZ��	(}�}�km��徙֮]�Ʀ���f��[�~��<-	�G6&�@�տqkK�D���f�p����v�
���`m���i���xq(����"�9"]0ޓ���y�qn�:���v��y�}����O�J�"�M�﨣��F��w�^��~�Cr��,?������sX��\s��7��M��W����_��_�b@���}��zPԮ!�Tɂ�����*�G������5RD��5�C�9+�	��O@�G]޴v��p��,�JF��9y�q���=mKl�r[Z���J��)����$���MO�j=�G=��b?�'Avj�Ɉ,��
�F�q�Y���>���m��?X��%Mf�_�'�hc��?Psh��j7��ױ�?��f7�VGI���s��n^��Wم���d�(�sءk�g��)�'�z�]w�u�%�41��o����o61�෽�mnݱX���/yIg5[S@uY�>_��~�~7!*7�xV��18�4|-v�K���������{ /�	9�����VR�o,�D�����:2	d����C� k-��ɉiMTp�D�Ku�ԴE��=^\$ŦGy�8< 	Ш���5����E����iT��?���(�����n�����.U2�%�Ջ��:5s��U���k�:L�\y�u���-�\��ǾZ��w�@~����,bE|�w��C=���_b�]�^�EJ�ܛo�E��=���v]�����l��n[~��=�ȝ�>�~ g�v��=`䙝Y��$�)u�[�f�x�Ŷ|�R�ԎO��&=�ӯ[Ln��I8�����#�����޸%R����]�S���?���`_��ל��~�Wx!1<	Tc1<R+ƓO>�/�>�����3���ҏ
����	��Q����+�O�����;����R��I ���תe���Tc6���j,��CQ����Vj/����}vֲ���l���:)q<��K(&��}}.*o)J�n���uia=�n��s��݉-��-�J:n~l�^_�)k�WD��9�6�VS���8i����������#��j����'�3��ח��d8��H���E��e�'�,Kط<�E/�K=`�r��V�q71:n�sn�'}�L=�ܳ������m��<kU:yy��zꙶ����C׮�+��F�=��;��IF���>�9��N��3N;���^{��Ǽ\0�T�+����\d*�L��)���,J��~�}��fk6�Q)���
�"I��Ijg�3Z��<�x�#6.n~6�m4Y�p�I�X,�o|cZ���
.��`��Nq�9)g%�}�"svr<���z�Q�����VI����}���I�ޣ3���l\��{t,�4~?�WJ�)�K�)��g�3������͘k�ǈ��ێ��Ȭs�w��y�������q��z������V��hbZ�d�o�fO<�m۲�1�ի��I'��%����)��d���a���g��c�G@{��V���\�d�Vl��ەW��IcjĞM����~b?�$ؓ�54�'|��m����9�BW e,e5ؖŀ�Ǌ�aA�z�E ��&j��I��5im�[^�="_XV�g�Q��6�P;:�Pu2p4�	ୈ�a��4��HG���y�+/A�wI��r(Ы2\ץ��=<)���p_L��1�O�ڪ���;h�e��[bj����b��mt���^�!Gk�!��������M�~��ݓ���^
ts�>^�k^�;��#lb|��Fw�/��~�������l	r&I����y�A;����QGW���w������.��|��>ϑκ�c�+u����Sq���g����u62�ê��my��$䟱�]f}G��� ��:"�w�����9�W��J������g�E��br�>��F����{�x���}���*���;�Y����k�+�$'a��6T�+6c���덂Q���*9��-��_��L�+����P�G���"��9aD�"���1^2�2���|�
�1��n���(���X]���2�w�����GM}�za�0x�r���w��&���3s���gG)q�?�"Y�q._����*▍���g�d)_�k�8��f N�y�+_�kO_y����?�coV�o�Ϳ�?��?񹈙����?:6l����Ϟ��H��#���Y�i�9�A�뮿�N=�,;�����Î�N8�6w��	!���;ow�!����j'�t����X5�?��F[�jȎ?�����4�c��J�W�1۾c��%�Ɗ�k�a"�ُ% ������C�1���C#0\�ˢo�34]��t�c�AZm']��Ϊ����<*���������Z�^fA�H����6��"]K�������X�y	��>/ap����e0ڨ�
}�=�s�;���E��k@��;�����;�)ԧ e��4's����#C�f�3	o�S�����\�����^c��#���:�,�����!u�t�MN � 6��u~�9�V�f?l�=ro�)[�n��?��F�G}O��Q����ϭ6<2a?���X�'�֭q"
��=�Yi�y�^��X��d��v�y��iR[^5���n�7��r[��{k���"ob�N�ɢ�8E�Jε���<xKa-�9����*ңW�EQ,7���p8a�ެ��Xp���ٽ�����}s�M0:��3����R@ΌH���Y݆�U��N�������)�/�P���ΊMlP�*��y��*�8��ň���ǡ��ӈ5�E��#�TВ�'�C��b{	�={�uf
 �N9[ڿ�S$�u�?�;�:����)��X�|'xM`�[�pσܗd�2[�z�M���FQ�u/�����a�Q�u�s���`��w�{lx���v���E�����w!\��g�ޘ��ݝ}�����NZ���`j4�=Ѣ\��-O=h#o��/��{׻��X�� Y X}�����z�j�k�GKMp��ǋ�'��%�c�_���V6�h�6#ŲS�+�+�!�XL���*�|����U�}a����0��RL���k�+Ll�Q�C
4�q%�s!.
���	�+r�9��I	h�u����B�뭲[�e{aÜ�q��}W_}�{��f���|�����ݣړ!�9�{��s�l������MM&�0>�{a��¬zg9���z��f��
�x¿xT{�����{��ղK�V��*�_�����¤���P�ȳ--���
�����eu���{�m_�e��K� "mADE�b�h���-&Q�����"��b�-�`��BD�FT�" ҋtv�������|��~�9��{������ܳ\�ַ>�yN���]�AY�x��%/	��������,���k��qՒQ�>N-��U.���f��Y�x-C�(N��9>�#_%��lk���bm�m��R�f}e=�l��g]D�)t��8�����|�]���g��X���/�:�|�Qh))JUH���<ήJz�ĸ�X��u v�׫�<某��c`YW��؅�[#��i�9~:xp�VdG�.}� �>�>ѧh>*l�e�;4`sk��q8�}����Ͻ�֮���2d���� ���zu)^���oV�':0X�n�`X�|��$�H1�É- �r����� �F-6��A�bn�\~�_X��$6�`}��Q֐�?Gǘ�^i�öYub[�2�═��Aơ8h 9.�Hʿ��|�X� (�FP�V��H|��{�j"��~А~���x���V����7|ܾ�8tͲB.tL�`g<LQ5�L��;5�,���h#[�<�s��ʿ���a��Yk�=eH���\�(��?�nr�c�Q�hw��.ŕyvg�5�7l�Du�n$���Y�/�"�����X��<�Jޑ�nl���۲�J�2�eO��)���wo���w�)ny6]�W�8�)���1�0��+R�ʩ�|�{ʽ)�#���I��O���]�7{�����E�Ѣ^5R7�L2X��e�s��$�|�IV���Qԋ�o�L{�4��e�����ްt�n�)8���kV?֬Ò�W�9�^����%�Cm�3<��6������������@ ^�e�h�Ǡ���/FȂV�2mi�T�b�J���bT�H@_!�H�Gh��RӾ&J|XM�Q�y�b�",�u���.�-PW�����`R����V=�Hx�I���Q9/���JX�t����[n�3t��y�Q�T��r�%��:�[�떱��X�^�[���7|���8&�tW�.�v�����~�oX*ЬZ��/n����Ï�vTN����7��Ƴ8w�q9}��3Xy�ќ�MqKK�e	ζ�egY��|$P���լ<��I��S��OsǗ�����>'*��������|�0��.�̌=��>��]tQd�6�o��݌qu���¦�=Hݑ��m Ϙ����;<�ȣ����]����"�2�z�O�4 |7��J�և��7G��~�3�mrg��w���M�{�N��`�5{n8ꨧ���=.,^�gN?@?OY���s����Y��E�j����7�y��=�4)ShK[���p����(#�Q�=��l�Դ--,�5����WD�8�a����m�<(�����%��P;$��u�3CT/a�=��fox������j�8��#�	+��:�ظ�u����?����R��"��dfZ��&an
��/*�+���85�}��ap�?�ߡa���	kW�
�7�7��yX򥳣'�^Eϓ*K�����0��2@��Q�*���}p{P�L�|M��a��2��4�k�TO��C�7����a�\���e3�o�6jz��Z���`�	ƭ�>V?�"���+W�Pm>�⇹_���I"�s�!����懧���s@��Ca�ڧ,��v�,�=�[�(���Y�B�7�䧡�ws�M�Im�����vا(��	�	��VC�˾���j�S��SN��˼��¬��aϐ��VK�x��|�;V��V���e��x��h�nv�@�ɏ~�c��a��Z�CP(�n��۲������M-��q}�-ʈ�K�N{�*�s�����{J��n��p�Yg����}�d��#�/E_@��
B'�+�/�z
�^t�������9+,�u�%�}�'�,�������_�첼��r$�-���E^�&���/̒QI5m���L����ζm蝑Z-�6eE_�r�e�a�k�+,_��W��>��O�M��T+�_��B��@��mT+����g>q�rN����ծ[���%�r���4�<��wɋhDR+	kO�,KO	6_il�`����%?��U�V@�?0ʒ�_.�x�ڟ���U��:0����y�v���(9��Q��Ch����E����?/��� ~��*DЧ0�{(���;�x���g��Hݠ}P��_�����|.�J�'�]ͳnf �:�R9>~�!�ED�o�`�P��}����eM��R��c}�N��4���~�㟲���^�|O��Ю���#��!%)k��MB��e,K��O�h\�"b��7�#̂��0�ꈕ�+6=d+
�}��TV�k�b-�����yN�f��G��U����
A���3���n+�&������O����?G_d�Ϫ�):��/���i2E�U��v�IR����i���f� �{O-"cf"�r�?�A]�=B�_��W�k����eFY�E�<?��,3\{�V�s��#?��T����f,�_�Ѷ����0��=���n��PTG���R��&��o��P7�6����yG��޻�W��+��s��i�Q��C�AT�°H	8 7S��$�E� ��J���ۙ%�dmx�6��-B@=�M~OG��X4"
�RĈ&����j�,OO�e�����h'���.ޞ"[���5LjI�GA����������&MGƃ����i���2N��E�k3kV�Q�Jɐ+i�r�r����W��($�y��mA96%w5�՜E0l��/�B�&�\��%�7���1�ph��~sK�H�:���>k�H>Č��j3�ᶞ��?U��9�����P����z:�j)q[�,�tp*$ �k�z�ue�{��&Fb�t��(�d7���<�y ��+�q�WGY�ry}�F��� =7�?��s��t��X��u�v�U#j
�� F�LDj���m�r����H,
o(t�SnO���UDcK�Y�'B҈:z2E���;�1����KII���@eT�o�q$�~�9�OCh5Q�0�<�@��H��QJ�s�/H�[� ���/�c�h/U�(s����z���������>���)���
���>M8;\Q�&WR�,��lT϶�,�� �b���k!�|�;��c-fċ��ѷ����',E��1���[�Z�|!J���X�s.B�t=4h�Y�:&Ÿ5���h��=T�������Gu�X�;���Sr���)���=S�xD�!�U�Y�IcE`_M>٢1�á$;���б+��ΈC��ԒQ�D��'��W�u�Um��)<�n~1��8 y�˅�Ȱ5��f�%BX%#�K�~���=X�J
�n��M��Dj��V�K�����?KWm�MT6��ь��U]����\��)�	�w�+m͗)�Q4ΙE^�p˾� �$at�W�}*iE�h{���qkI=e"��m&
/�2%�\��EMqT�Y+�;�[�PQ�Mݴ��L�z(sQR+�9ޘ��-诮k�/�m1f+�w���dS6{oᘸ�,TB� >�篙Oו,�&o��y�	�Q(��s��)�Сs�O�_����2gNOn�#D4��Bm7k#y4XN�Q�/��C�1�a�V�6h��e_�J=�7��Zr1�0)%P+��>?���)�jV�7W7��7V�Z�u����4T���|����{�M��=��1��n6�=)"OC�WT�Ÿ���0��l-�E*/�,�re�v�0٬ �os��$����>,�d<��Aw����U�E/�!�@��C��X ���/}I�m��ro��]}��Vs���dJ=��Ʈ���/�xw�dd�"R� �'bl���$2BX��x��DSH/��-�7.�o{z�,�P�s�m�W�(�]�R��!:�d�y%M�p�J�J0d��\�aK�A�����~�s��y=���<�տ�Y����@۰c��3���Ot	B<Ǹ$�c��p��Q����b�����n��-��1�T4��șlM�k�B8�evi�x|�+��T��RMR�w���B�#d��q�$�uHť�b}�"�h���Ȫ'�@� cJ�ʾA���d��>~��*̼�9����5�8���d+���IG�*�5�&���Ƣ΅��k1�$�ܟGQ|��������x�5؂8,�Kc0����馪[ �a�m
LʉU�1G;;���\(��P�\�|LZ���u�!�ƿ���Q)���l
AC��\JW쁡T)��;�)r�W.���(&��A��H�=�C���{p4����h������g<>��̍�&��8Z� P��j��eU�I�s
x9��;��H���9)t)r>�&�硲*���#
=�O���X�"ߏ���T�E&[��ĸ�CD��*��h�Z��
z��-T�̪/%#�Gڽ� 3J5����ǩ=V	��~��&��[����\�W�Q�y������5)Z��������aJ�T����E8��Uμkiv���~���7�@�����J��9�ƴ;�o+2��x�::+Yf�ìl� pߌ�;k� 7Tqq���F��7B?�Z#񿑞�ږb�����|%<^��5�h �M*���B�c�R��������H��EM��\�{�"�7����;�;O���;�֌R:;���x�o��!����iҎ����g�C���Pv�Vݛ��g���c��E�wnM�y0�chA�}�g&�����3W�N���ם����`�ީea+Bf�yXI5A}}t��2�s<a�i�����z�IM�3���L)[��m�H�T�)e0�5��"@
E�SL�m�_�BXF%�)�k�c��L��SD~x��d'���O�z�a���m"��V�7c�X�_罴����}K��z'��|��exoK�TA��[�mlb�ް��'=J�x�޷���ֽ�tY�=5��\�3�֊�(?'u���|�ӣ������ȡ�S��Q��T�F������Z�q�CU�$��y�Y3iy�!����o��Ψ����)nx޼���a�:KΤ��(aҹ����M��h�7JVB,������ ��/Z�>f_T�� ��%哽�8�9mmry[$O��J9W�G��U�x��=�x��<9-�x
1�Z��S�L�xX�{=�Z��S��)q�v��&)�V�I����"Aj�a���[�$)%�v��a���c�h1U�I�� 2\��&��h�VO�q�Q����PV璵��r��y����s-,M(��`s�V����:`�A�����,�ߕ�����p�QG��sS8]�\J�}~}˯��<��Us"J@M�y��3��{��lq Aʊ��_n0Pߔ��58<���@�b_֢�W96S`�|����~���� te�q}szYt�WŅu��3���
!�d���������d���־��V�1�R��� �c?��f�7���crkI��b���?����j�	��� �[��ih�/������B�Y/*����ہh��K)�)��;��}�1F�ĢE�æMBGg�l�y����52+J�X�K��a��/^b<�rw�m�d�v�a�����y�T�9�~��������o;��W�J��q���w���ۢ�"��|ޚ�R����)Z��f��Dy���yL�"�u�$W�����.Y��&�S<~"��H�z�/U���@D?,�e����{P��M��D����8/�4�y`��+�YN�o-��A��-��Uua7�l���x}QS�1T�e���3�����~�Zu+�
�y���c�1Ѐ�)��y�q����~��[r��$U/'�iXq�I3��Be�%K��A� ���AR��eɀ%{W�^c݆@[tvw�=�\�X�$�_0�������������{��^'�/pMn��_�j���Q"�R���/���(���b���=yWq���B�ޢ-�#��믿>�
����B0���U���+o#���xg��Gl�	��ҡb\�;�L��E��Uա��>g�y�s��1�W���>�_g�>���=��¶���q��?�����=蛡t J�����'>�<Q�y�E(���;#r���[��H�QI�D�澰ے]ü�¢Ż�����ʹw���R��k��^������J�ț^��4gx�s�-�y�TNK�~�âӢ��O{z�k�ea���V���f��C�A��.}<�ce��DV���6@��XZE_T~>\����mg�Z����?�c�¾Ta-*
�;-@=	r�P���*>?��#I4&fb��6�B�\���?F=lUU�f[%��,a τ���%����w-(|?��s�T�2?-����u��`h�m?~_%�Ѝ�������*��g?ks�¿׾���P�P?|򓟴�#T�ƴy<���#?�@'��=em��֭��"�i���Jٶɼ��l�΄�ǳ�O{��L�ɝ�g\�l�p�����&�|�/¯o��ݐY�������=�����p��Ǆ�p��X �|�t�bWEA�k���lٲ|" �JV�౎���'��mU�H�6����,l!���F��b�ɡ��呕�a��}�"=��������~-�o��|��0ط9��prȰ��Hj!-yL!��rHߏvr�c���g�����և/~����LY11��ΒmC���ů;���SO��:8���^���/��b[���7m;�9A�������@�>��G�7�����'���=��~����"�(�:!�C����|{z�V�a3^�w���`�شV���n��e(*�êU����-���a��e��]�f]�ߟ�8�\�.�}�����'[G/�w`аYYY����c� c(yؖ�+R��OwԶ�jR�*#�oB��;�p��z*�4�)������p%+�V�U#�z)q��0̖����]��C��ې0�1E8������'yY\~�������ֳ#�0.ޠ8���z�E
LCu0��ۻ�=��*�a�����Ɯ���S�ׇ˿�p�	��7d�'�n���p�]wY$b[��i���&E^p�E݃��|�����/¼��a߽w���#a��}��b��֮[���p�?	���ߔ; �fbrr� u#�+ĀO�]A�����}�(i+�)-�e���"�C�������~7S�s�N�<GOs`CV��5� �~��hd%��Y��?I�Y�U[J�Bt�kr/��HG;�C�����cm���߹"�wιa����&Z�ᔓ�̛֬~*=�x�4*UxҊ������Q�$�a��Y��:�?@+�p��>�W?�fU�я�.�=��2�p���L{�J�#~��K��i�{`s_�;�ۚ*<�όx~ظ�'fq�rW6[l���u�6G��Gm�?�\A|��Y�SLX�
��'b5!�|�H[��-�l��hY�SY��y� ��X�a�0�ը���8��Ba%��b)U�fϙ�'�ߓ~/.���^EV�x�V@�/�
�^w�u����N���뫮���,���^>���Q � @��#�S.U��o�i�c�°�^KB��ު1 ���\w��`X�p~����-w�{����@B�ΪUOm�M{�_
�M��;��sٞH�C�#��0��qY�������\�a[X�<'	,�/��~�����;��=��!1��f1`��җ�d��3�I�D�ôe��p�J��h��^1׎DB5�bHJJ9�laӭtf�
��BZJ-yC1Z�n� �؜ΰ��Ѝ�T��I� ã�?���B<��Wq!�hFZ���O��-���7�l�n�Wy�w2�V�ZV=�xX�����t��l������T�2n�Zm�E@����L/�0����c�3Ꙕ��p�7K����ņu�CgY��MiqqʤV�6��$q�2B����� |F#x��|�.����t5e����
�Lm�W}�#CuYM�=�C<��"�r�`dl4./�åa�XH͈ޔ�5\F\ �� �M
?QØ�@�P�ƅa|��;�y^�2��z����s�����/��'�c��) Taz�CwO�u�d΍%�nI�4�
�Sփv�k�L���o&)?�4������Z���S���:-�M���v�OWGw�<0��ss�ӀQӖ����4/ݼ�+�s�9���~`�_����芧��֖����K�no�<�4�b����Q��r<�h�1��D�G?6[�5*�ٶ��u;O2�>)e��Z�	`��::��M�_砤����@;���Ë��E���/�x��q$��k���4�+c �Q��e �}�O<�.�E�ڊ�Aӿ�=��Pn�R����`G+{����ʺ6̟7� Vs,�?��tǬ8@;�������M�;��I� �"�Í�"O��$�2 (���#�?���?��?�/|����W��/(���-����S��{�.���6<)Z�C����V��k�eo��������'�������2ۢ�j��;j/(+%��E��*tQ�y���z.�����WCw>#�G���X?ߡ0�a�
ݺ��tu϶�J�fx�����5{j����ua�^;�6�gI���%�R���C女p���+��nV)u�q�psX�vSXs�TI����6�n��=b7�?�b�<n��ִR����t���Ȩ�;�n�.��_�o�}�C��N+\$���e�cnˎ�ɄZ'�TQ���(i��0	�t'�P����ڐ%q��*Y��?�i��xF���O	��`t!�d@���.� Ý$Y�_=Ҝ��-�fT�:�֦�����a}X�~]� \�g����x��C��Y��N4 ���MF�F����	�6�
�V�����{-�#���;�7���W�5�����Īա��k���ƀ�����B[�]K�i��s��VD���p�aO��zsX�a��*����[騄����~����ͻ��s�N$ox�����jx �@l����g�"�EEBB���Ԗ����5/یs�_u���������uM��RW��U�P5mi���j�����\��_���Z�v���-�V�%�<1�j�ق�!v�����I�U��9�<]�O�����{�Wx�oSX�iM6�g���U�[I�ݬ�粽�I���Z>�߰1�u�=F):���d�S�eȚ>몃�?�C³�����Ǎ��'J����3kd8����Z��QO;&�Ǟ����k�F����mA�g=�n����j� H�PZ~���t����-h�Xpmi˶�o���� ��w������y}���z���ʯ���Q;{�_�|��&(o�=*��>�ݴ�8��_g��W(��ܠR��\H��/|���^�2��R�c]�$1��0�|�~��������t���/<����xU2~��v[N{�s��
s�.�c�����]w�6�t��;c��5���T��!�w�WZL~Y\�I�{���|�>�Ʀ��G2g��ea>���ub ��e�p�~���VOa��
�ָ}(�W���:5ߞ�(�����J_O�M7�d�1ա����(��� ���O�H� Ҿ���U��J�����i��R�导� ��9�=�г�q�f�!`���A�0���9>u���W_}u�m�Ea�ys��y���f͞V�z2��m�r���|�5����7��^{ì�9���U���o&iB'����������a�����a��9T�����oF��~�j��FTra@��+v��;��U�<h-�do[vv���
w�[U���o����r����zܨ��0~r�?U��ߛ]�z3�f����z�*�J[7��,���
�b���׿��]�O����(~y@ZL��^~��-�=k^\ ������@�ي�2cq���QGt�u��{��U+-<T�3��m���q���Zޘ�%��/~�?����7�����q��W��6���ׄ��+�巈���������fx���;�>������28���w;�Iy[ڲ�ģ{<���jCi�ݼӮ����m�$���y��6��gaTY\
`Ͱ��l;�W!��"�c~����I'�d�Y��	�b�Q�N��������O<eq'|�;��:t�;(b�i����On��y����S��*�^�7+�R���m��fϝg�W^n�����u���LY6i��?��n�:(-'��!]$�����>����f�q �/\`!{�ψ~�c3,0a _�5=`۲}e���L(��̘������@�u�E��8\�`��vBj�S�UΊW;�ݲc2�Y��r�c�D2t-~��`��>I���_���l���MA'9�o|�F��^Q徘z�B����|�*�n8萃��˖[�?�G'<��#�E`4��\�6ܗ�3�B 0s;y5asey�jg�ǒ������X7��?�x6,2���B�=����W�j�\F�O����
�����G\�mi��*��0��ϕ���	[�V����%�����{.F���O�f��Y�[��A�VT��OA�5x.�³4jBA���O�~�к�{�F� �
���Y���Z����O�G{4k��:+{h�����z���xB�X��}��]�5�`-tf�a�q�ש�Q�d
��J�!i�!�Ց���^X��/�� $9������e��V��(`[L�V�}�X�FZ��w~K�@�������	g!�<��/�	���5�暩�����:�*�B*���{�"X`% ���~};P��HH�}�mn{J����3�Z�V���Xv���ζR��Ŏ�ي%tS��
QV�(�T�b�'�ݡLq��ϊ���H�ߏ�C�{�Ï~�#�ü'����J~r�$����c�CF]�і��7��V�e��vU�F_�P��J�⌝�ʟ�݄m�TMNu�g�k�E�Ɓj^,}�9��L>�z�<H� ���FZ����7�).&c	�X�WyAS]�#XQ"Ucb�
y�y����C��Ct���#�+.�;)�c�>����[�o�_�}*Y�R�o���']F���X�ԓRP� ��^��͏J�¼s�k&�jod �����_�����Ð�}��`��<PO~+䞌�����1�כ�(���?.���Qyc��^ײ�6�^:9�܅b�@�(�z�[�j. �[�����e kLx`�f���N-uo(k/5nbK-�$�G�=��A�K��N�Q��{:�f�Ų�EQߓ�>
j½p�[XB��Z�@-�gX���u����MI���/�B��g����D�@��(} �]�V��9
�3���[���;��1���p4t�J6�E��E#��5��(es"d��>q�_#��j_�̜a�R���w�{T�W�͇?�a3�t}8jd���Y]-;���%���]u��M���p��W�(� ��|��A�í�x}(��hpȂm������0�({�Ϛ*�r�?�V�T/2S�FEp(D�b��𚸈��=^�Π��E��<(zAh�e�6F)�d|�����I����ڱ�A�����D�_�GJʟ��$eP��@%>(�8I��WD��͵���ͱO��fVO��V�Ŗ�R�fd�o�3�<7]SY����~�%�Y#�Zy`<��m��fc�^��k�u� MhgFf��yK��rke�+�Z��/^�r�/p��`<��ۥp�&D�%$&?�#�`��R@^���5�e�*l#��lb���>�*�U�Vc��-�֥ב��B�d��R<\JQ������^�F~�����Pl&/y##0�P��țsF�)l%Ũb*?~�@d���K�Y�v���&��l��ª����Q�@�t�t�b��+Ua������Gख़��gˀVV��f4��6���暊��z���sm��3����tq��W����V�~������R����uq6?��=��?�IG�&-����($��m6)E'%���>�z�>�.Z1�k��&G&�X�:�֑Gi
��@��>���}�/�]�\�ue1s��7�Z>���H����
e"�N�FU���0$����jH�Q��������1L��������<\�7m���I+��c�!/Y��pH�o���?��&a;o4H�3��a~�9�;ƒ�����FyzJ��#-*�Qa��s�O2q�~��W�IǺ�z/r~c�(H�,�}�))�)��G!yإ�<gx+�_�c�X0��؄��,�~eD��M�䔬���I�s\�dI�O�gAn��Ip>'�A�)�t=��gk������,�f��ZȔpTX��%�s���t�:�9'�!#�EC��z�#�����M�K?#�~�;JF�2589�]���,5lJY���Y�w���04�.�T��0����tTlQiz�uBz���jg�j���9���t�VR�Q��ku��ʴW���8�}�Qc}�V�����z)g%"�KO�UB���C�DV"x��+7����?
DI-����1��krj�q�b3-R��z�rC��5cA=K�ԑ͔��x:&ŏ9V�[H$��PD
1�D6��;j(�筧�{�~GAWh��=��A#��b]K���Q��(�;�<�&���`S�V�J�S�HcEH1�-���܄�Ac��W3=�~kԱ��fe�Q{���к�J3�߬·R�j8�a��ڪZ�IȔ��:-'O-B�db�zG�k�'��/�������ڷ��5����J $q$pa3��w��h��0)�=��::Owg���j�����5l�^i������2���#-*����^�h�q_�&���r�0���=e�g�CǪ�i���PЊ�9��E��YH�63^�o�;
����N��!;ϸpu���?d�,�t)�Q����@H�{�+]'��3؊95��0VA&Ǖ�sOZxձ/�0�E�;�.�nʍCc
�:�s�OǤ�u4�Oc��i���a�&�c��]w5*VU�z��Q�d78M�=Q�����h&��w���o�a��e��
ӣo�(�&�b�<� դUa����)�YY8R�,��$��ީ�gx,�����'/O�s&�
�
!�R&��QQ�����ߔ���(�z����^�+��<�Ƃ��p��<U�1�h|)�%e��������RE�'#�X��?�C���?olճ�uZ���e�]L���	՟�Z�9�:�����PP�'�Y{�4��	a�Y�������?�䨄>Jm�:ʝ��m7?���OJ��P�E���_V�x�]`�KC(�j۷y �}Κ+� �u)b �� �_~y>0&�:�.�&.�L���g6Pe�kA�v���,]���j�l����W������=TL�
�M�ܟJ�'�T�7�wW3"��b�0c�q�x� Y�Eԙ�c�#)�E~"D	LY���9yT�Dqr���sնx�׻���TG)�V��/��\�Ej�:�K.&x՛�!5M<G
�)�$���+�cW��y�ᤓV�=��==�J�7�m��Px�Ǭ����z�Ø�[XX�ɴW����]mC��3�8I����n����M�q5N3�==i,��U�BϬ��Y0���B~<�I�l 3�T ��&���Am1L\���Kp�f	[m_1��!��������O����b�^� �$��$/�Rca*����(�K�$����Q���E�(�F���R�0�S߂r�a(D! ~ON��2d���z�������﫝sJ�Y��XT���t����W�e1���{x�P��T���q���q$I��!r%[�jIX�d���z�<��p��ׇ+���NW7׫�<i���6��M���I$��N%��o�J]�d
��|����c��@�%�l�ޡo0~?��B�pË��v����D�&�?� Y%*�A��'� ��K���	ca���<|t��欣����u��ӻ�
oy�xkE@�[T� �(j��7����t|��b"EJU�A��X���D�U9	��(��Έ3�3�󂹧0k��TU,�w�qǍ���ʯ+4+��T��74&tnԃ��cn��؇�FOPV�+����ܳ�	'�8!�KI�˥Z��;�d|��q� �6�<�0�<��ʧV�cc[e(�ZCӗ��l	��>��/�ma��w�yG���_��}40�
;����V���?�~'R'7����&�,f�;�!�� 4lrtt�A�i�X"�e�w�.U�
��f�2�����lU�����
1�z
��(>�������M��SY�:&�z�F��>Wa+�����1I�,��_���S&�x!�B�SS�õ������4��&�����3��R��������[��ݏ?.|>��`���o��d�bU��v�iv�4����(s�'�|bڏ ����3���w�֬[�ſ|��ê'�O{�3�ҥ�����-^�]���Ӱnh��e�Z�%cc[�|�֝^�����љ��
+W=���DK�?t�l�bQG�7�p����Uk�QO?6��*�R����N-�<
Y�~Mz�bXF`�{sT���#耱EO�J�AU����G;,|�<����ĳ��8��"R��{x��d�VP�����E���d��ZBQk��W��ZBaފU�x�V�.��'�=m��&�E�|\��Y�F��ys�KKR/�m�������4W��|������}O���Ҽ	����V\��`Q�oi�R����/�{��a]T��w���9,�M}����~���p֙���S�@����([�ʴW��	@1���Ι3;U{�o��M��H�Kw�����?�)~��.�����}���?��!y��7c���z�^hȋO�y6YXF>��cͶ���#4�X4X��,⛅��
p�F�E*O�;ؤ�*\�7��d�Bl���a��yy��M+�UQ�D���J�
�H����"b!-g̞�{�y�Ɵ �����֬��p�C�5��r�~<�Z>^}������o��C�f_��O��p��[N�s�?�lI����
룞Y����_�bx�E�	wYl��#;2<�Уa<-�g���	tW��K���m
s�v�[n�U8���򽉟�5k��;	����as���zVX�nc�����z4�<� m!�x�	<4yx�^`�#{�'�MdYy���������O����C 5Ƚ2���h�d����^���tN�!:��]�"_Q1Vު�ڑ�$�����mC�WJ�U�L3�7�"2�\|ިH���0��[woC�	��d[9~�ܥ�{�dk���И���?�"�EO��^t���1�c98�F�0�U�m֪᷿�9��	a���>4d���ӈ���V�z<>�V>��z�r곭Q�A~�ӛ��F��Z�.ȴW�I#��RͲ�W���3<�أ)�H�ue-�Y��G��ąN�E �o����`g�y���TSx�'���/�5�җ�4��_�e���'ێ�j)�V�r�-,N��aq��M=�d[�SY|�{�e��D��?��Qdx����˛$L���ӱN� y���i�B����~���r�O<�8��
�%��@�+W��{�p��ˣ�9/.��3�� J�[�TaRl�J��<��,���.��#�?��p+���W���PO�B�ء,�����!+��������>��+Z!�ërχ|'�/I,P
,x~G�׿��f	(^���b���M�����+c���V8g\e�QԬF��9��'ק��L�թ��D�PR
��o�C���y
)��~����/.J��0�"O�WI+<Hn���%��+����}���Q�j�ĸ�GT��
�R�3�W:�EtpB�8�fu�����A�E���<�#�^����jQV�j�u��7����՟X�]�ܙ%]C�����qM�:�8�,wA=>a���ĘZ���7B�8U*�jB�4�!w+�˒Ŝ#�gC6�ERS=��E
��'baf,���~�|�m��62
�Qb#�0��&Y���IǦ� ���檼`<\B?��Q���+�'�=x-�a����\\l���e���`^w�Q���OL�uk���W��ು�ƥ����[ݳ���`�YJ%�!�^*u�M*UR^n"�{!atS�^���O��2�L�>�{���y��U�F�8�BGE�f�E���L�\�ĥ3�K^���O~Ұ� '�˼=e�A߶�GDʟP�^O���Cё����~fFA��B񵒱�C@�`
���G�&��	'�`s[ʜE�ӷ�������T�������ƅ�V6�r�_�V`��j�~{��.:�3�#
�&���L�z&}�tRp�kf�ww͊�¡��Fk}m�Y��h�f�QBgX�;�Ǯ�W���?�'}�Ї>d�>&(�?x j�۫ց�(�y*%�&+b4T!�K�[U�;j�E�����F��-*��)  �G90U$���J�W�J�z��b�Ó��]:v��!� ����Kx�0F�(:'e����9�ȧ���k��5���:u�9���u����-�bŊlA������UO�L3���	�j��O��]ʉ�3���{Pxr�C��G�aH��*�P����[������ ���Zgq�f�q��)��(8٧>��N)@�>	5��2��l'%(�O�xK��
�R[;�0QhB2�^�>�-��4��c,����\�\�o��2�h�񊮗�E4J���Q�V�}��P��u��4�p��>���'<��á .��]�E	�gO���ݢ�K�,��E��v0b^H��<M9"�T�_ٴW����#��}�s^�={��5�+,�.�~���~���Ҙyq�8���1ǝ:����V�V���
_��YU	"ڽa񫠊���<jH��2A�Of�_��2�t�bX�8����w�(�;��d�c�|��4变r���ɂ��fAP������@�I�&���������������}����k3 i;��cC�^{Z���ݖ��_���0ؿٸ�6m���ts�qǞ�v�3��p��	�@J��3*�g.�O�2��:+�B��������0{ޢ��!G�E��m�;V\n�.w5���h�@�I%7���d ��ӟ��n�����  ~� Ą(E�KJ����SF䕨���b�0����D������־�4�CV�����lq��
������A�|�q��L���D�w���	>=���¼{e��KϷ@�v���s��>Av��n
#z�~���1��%���·{ "��>!���Q�0>��������]w�i�Ϳ��?��N�,�T�` 1�1��$�İ/`�%M���G��M�
!�k�C�3�f|݊���wb��Sqt�d��zvO�O�����X��w��k�i�j�A%��aNT��.�?�x��E�=w���:��|�!)d��6n�W�ϕ�_c��]��{+3��O����K�f4��=[��Z3����h�����E�ȨU5��j�0�:���M�!\pAx��^��o�&\q��k_��YLLmW1Q�&k�S�>b�����K�"��k&n9^xb�hdbiۂ��կ!��j���I�ce��NQ��s£)�*�@�d#��+�b��c���$�}G�yOD��"+��'���WwM�P�B��E�+��B�B/�h��_�<�����@B8��������E�r�,
R�x�į/�����;�1�c����)��H�D�9�1����s���crO�f��o��`*����d�׊sa?P��M����4��/_ȋQ�󊗽܎o�Ż�9s���?$<s�)mC��>�9�P� І�%���)4�zjB)#�O�z֩,J�:_է�7��$(�!_@�]Y)bGT�NJ�6��`�Il����@r���>` ��\��p�r����0Y�-�˕U�;߃�.J��	Cų��H������{r�RZ:�S�B�Hd=QX��/R�οނQ�.�G�����ENVe=���}�zh��q0V�@*���+�}��Z�@,[�0�}�7�*c���£�������LfOx�P|��zECq�T�KIm�k�����~��_<�@;g#|G�~�Be��wA{H���CW�f�q.ox��E�C,<���/�\�1(P� ��K�~��~z8ꨣ�;Jx~)^3���/䞆�Ȍ%v�����WX��z�M7�
#i<ł��Z!��TYV�D����o?+�Fi��]v�e�\�w���h'E�+\�5�Ӕ2�I�q�9�+_��m˔t�:�!0�Aqބ��;����;L���t0�\�Rǣ�g�{˓�c����(���̹�]����X���z0Cmϓ�),e�C2��T u���gE��!U\ �u(�(�;�qSj-����3�Q��\s���/Xؾ�	�
�"�f������?�+Xy8@�Qp֭���	�O���Y �sl?ߕ{�x�o����g���O�$�'bM�}��,,X�Z��6�	p��싱��x���x򋱮�t��w,:��X���g�5C�Z��`�q=�y��F��Ɍ�zZ�Dq�
kEn�o�"�M��h���{��)��b|>
�N�@�L�`Q��m-��@�M���w�-&���x�O~�܂`���/�{�7V>��$

YҜ��d�� N��eeyŞW �}Ja).�܃����X����+9=�2Tx̋�ڢR��)T��o��d�_�t>~�-��Ň�t>�影Qצ�IP¬�Q��΢ �C]W�	{0�x-CB�E�Oޯ���<y}�7�a#o��Ʊ�m��x��[����2�ѥ������m�$�6ʱ��x ��?����{��^{�:�	�1�(��A�����9�ЖI����3~�G��c�'���C�EI=]\YA
mx������c4W	J���X�X*��b�a��O֤� S[;3�G�_)|3�'��%��%7ٷ{�y��XM����x��5X��GǨ��rqY[���4pM��G�z���U�P�6R�XO�c��ݓ+(�O��ׄ�qY�+�~�H<��,:)1�g���|2��̞~z,eQ�#��Z�-�~z����w��[�K
VcH��C�}���3�SCH��@ʠ�exCL9,>c�1t�����Ka�H}��G�t���9/�/0w��_��WٱC�v����X5�}N�/�X�bDe[\C�O��P�)%��6�><���ذO�q���|#����nAt�"�|q�@#%��.��P��J�MF�Y�?ɋ�d�MB���)��OhY%rk-ќQ:�[ ��z�%�BԾ��P-Z]�da!����?�SM���J����$X9f�l�� ���D0� ��x+�uU��{����Qܗ����a����l�+FΟI�dS�h��'Q�,��(/ΗEoO�J�EPJSR/���ל}���kxl��d趾��ay�׍k�}��5��uQ�����cD6�[J����!$��'�M
�Ѥh�țf�a5��߶��·	������K1yY�7�ٟ���;�7\3§�w>������w�Q��uև�Y�Q�Ωt�s�y7{�\�� �cp6�z��a�&��\`o�!B�ԋ��X�B<�#�G��� D���`>~�d�,���QP�E
PP7<�I>a+/AJD������}�Rg�qFn��!��J�Q���cb`��!�K����-������^JL��(Y�LL��e>���d��Zם�1�u�@��mOׁk&��~�m���|�3��/6����d
�Ca��C�0Iz^{@?�|���X
�#�|e�)<H�k�H8��
s� ���J����'��SO=�ƙ��
E�K��s���k���4�4�=�*���xd�(SZ�8O�����d�)��v�NT��%ijOpj��a�>8G��]�앰ւ�ךk���n@縵R��8�������U6�����2R�>��x���b� �()[M\�A9�*B2%KE�X�P���ؒU?9�ө���R*��� U3���ۿ5�Id�*�^�W���T��hC	̕���Q����(��4[�t<��|�+��ҹj��9�""h2E��#�J�^0J��9�z�ߏMY��������gD^'���'>a'��v�(k�G��vAa�X\r�%f�{�[�iy��7���"��BCR��X�}D<�Ya%b�,:��\�����{!EM��d29��H$�-��_�a'?������Y����Lsр&~��镧���y<dybrJ��5p������Ʊ�� ���#���N����{�]w�n�_ F�m�]n�$��R��`��*(~Vᕼ�}�3dぞ�J�+�Ȃ�� ��N*�=�n���9:�f��q~��"�?�S�I���V:V-��/�5�����%��-�j^���,s�÷��"� ��R�4%�j[v�裏��|��W�DM�g'�t���p�KɃ� D �������*�$i+�F2�y%wQt,v����{����o�KȊW�/��bJ� ϕx4��%����Dj#�6��^"�<���#EĘ�e�����'j��v)��\�;�5�\����CM�Da�Md��Z݊댧���
eP��"IG|]�p��y�"l�U)�c[�7ҙ�������X�BQ���R	b[�����A
�)�%�4��fA:6���Ci�UO��	��|�BB�7�Rj�����
�u�%n694h}�M�6�+��F������*�qP�O�KK�3�U-�_�1S�L��>mIe[c�8v�R%����ڗ{�g(
�~*[A�YӢJy���C@��e��Q6�3l,��k��������ߓ��WS��Nŏ$�����Ҵ7�(V-1H�C��U�XWL\�4)���~�����b�m����ZX�@�����(�w��?�m�Qm��(Y�L���,��s�U�3�����a@���E��1���Çu�:>�x�0�_,����\xα���y����D=T�T�i���{�_� T�3������^n�{_4�s�Ө}���Ry0�<N;�ܪ�ّE���J㷼�-�}�z�8�[��m�6Q�{"�` ����+_�J��!�O|߃�(���/�+����R����B-�����q��m`xlM/�F�P�^��TV�ȴW��=�o�!g�D�z�*��!FK�"b����CDV��T2�Α�,�?������\�h<��x-cS[ƖV8{Z:�H�׼�5�ȧ��<�*h՗ZL�(�������s��/��3Qt��G�ÃT�f�*�Y��yHo#)r yU������/	Q��2�?@'�����d�Ax�5��0�ô�s	���	5�:���B{��G!(�6؟&ߨ������6�,��a���>=����d�����o_�p͵�U�O�tWg�q������MZr ����+?&D�i��&؃���[[W�R����B��b4<h|M~������X2�Ǌ_(���
K�"����`�\��j[������(�ָ}Cx�����k�r�=N��y b�_08Ny�~�C'|~�G��A�!Z T9��=��XX�,>$�	E��R����G���������Sjܔ��Tf��/%;�寄����!zx%!b��Jx�b?ȥT��e���-�&�`z��9���"���B�!o����G����.E1���6a�f���bbX���)���R��<Q��W%F��4O��b&���������o��
ay"E_��{,���C*�!���������X����u�[��Vر�xE�%�N+�B�o�<�?F`؉E�@�T��^
����ʁ+�䘚ë+������9dWPȂb����rDC��[c�f��I��}c�q�>o��V;z��H�n7�0��m$�ے���3x. H��o�h�IE�+���}�E�����ٶZ�"���V�%�g�D���E��_�%j\� 
���k^͇<���rQ����+�s�8�����M\vV�ǟ���ʿh��l7Ӈh'[!,!^snX_|���'�{<N�X���˲?��g���|vu�\G�F�o�zƭSA�=�xA6Fs��E���7��DSma�;�!h&r�Ց�S;p}��s�?�g[R�u��1(G�X��ͮ� �,�,�(Y�� �4��<+�((*�����18 ��,�Z %�C~�Lh��&d�3���2ɇ)?��T���(�ڷ���ۙ%���TM{��lugV���n�s)��9_Q�X'
Z�Lաk�I
���iʚm͝=ǬtQ8�j:=�����r�-��ũ�dR<ZU���X�g�u�uR"�� ~x��!�Z�#+�,Ă*ب�rK�E`��/Xo�Ḋ���U�3ް�?��O�7�����_��_�؅�����YX�4Ua|���4�-�U^$h1�Gq4)���2��1I:�!��7F�ƫX8U�"�-Q��z�m≰�����_)猻;��k�TJ����������Q|��^���M_��}�K�o\V\]�$s�`�z��>���d��
b)
��@Lo��f��O,�F�����!V��a7�/y[=g�IQ�y=�>��R�x��IֻN��#Dm�X��(.:tѪ%���7�$���XM�W�1n̂��@�?1��lC�Xǀ�[�2�+'����u��	H&���DH�?IGwG��ŴW�q�k��������I%����'��-Z�>���dՖ��N%ٔ�U��1}�6D��Ќ�5�W��U�Țc1�dl$�0<��9�Q��W�V�~݄�����L�o$j��ppO�N�?��8��҇�9�I��C��#���F�TM�Xt�z̿��=�� lKy.O�k�&C�J�<Ť�3��.�b�?�fo�K�B.�X�r�5i4@}`O���C���)���7�֢��M����ĵ���\CV�g�(�3AU��X�R^����D�阽���,E˾���S�Һb2k��ux�8�h���W�D�"P�9�43 CUOy �k�Lݷ<�ƷBA2<|����YO���VD��+#�-wf�T��==s���ٴW��Ty�[�^	*�3�E3$#�gE.M�9����D�)�llk�%!�����xeQ��E֥�s��e�Y~!Cl���6��˛%�&�/
�
����+<!k��J����\C*TI(*	�1#��S��s~?���י�&	UOR���:��"f�b=�>�\�:O�_a��G��O+���U;Ey�y&zD����n ���$��Z��K#�?U��E4n��"���_{?G4�$;��/gƛBV�����{.YR� �ښod�����7͟?��M�Ԓdf��+��H�Q���׾6\t�E�$D��r~��sP <�LEbp���z��$�'��T����b"���7��h9u@Sӟ��!�g�#��8F���Y��9%�E�,�&�4�t}�U�:MT��<:mp�����\�׽�u6>�؅n^���ã�?6�8i�։<o�5����ق�n�=������O��{�d�ƍ��w�&�T���D�&%���Lpoa1�9a���Ț���@�(!rI��	���g��_�z����R)ԉTVń�Be`�9,y.$79~�!�bƱ�:Y!���3Q�L�+��W��ն/q�����h� ����7j���˾�e�m�ehK#Q"]p�Y�O~��+��v�+���-��Z�7^�C�"k˶��1`���y�ؼ����b��C��v)U�i17�p���k� CNm�JHM,A'�'�^��c�'�������
˱ `q�|W��^��(�a����J"��K/5���������}�5�� ��7����>6�����!�EcY9�ٳf�{��'�-Ӟ�����O��v�i���\��5ض�'f[FD�F5�'!t��=R�R������ʿ��  �IDATK|<_}x��Ǫ�E����C$F[BO�ࡒ%EZc�&�΢0�^Z�|�J�m�d	��ZQ��9��0|��9F��.��2k���9v ���+̪�C߄�[{N�.�gK�-���u�p��ϸ�W}��o���GN?���]u��/]�p��(+� �k˶��v�!t���A��4)N�EL��_Oi��P%�s�,F*�����{,dB�����o�=��_,�B�������*����.�U���eL	j) <�n\S��e�b�E��G޺�0��x[K���CG<�w���������W+N:��xa�V����.�BJ8*$E]J�����x$�^���#Z8>
�(tCD1�r����%�&%E̽M%��P�6���
�����VHj,%:Q��J|q�GSi��?���jKt���el�H7�`�{/[��?��?�g����~��߽�_?;��T�����˷'[�dbЩ��j�	��LLe�'��)&�z�h�Dr��5�����)�9L�xxa���'^W��ؿ�f��F�Χ�5�����ب�=��S�s�i��q�����ZX5�5DiKs��F�E���U�|�W�n�(�s^�������>��p��܍��L�3�҇z���r���1�})
D� ̻�cҲ�FB#F���g�T�����"��p���#<�J�[����2�$�
u���CY�r�J�������dm�߱@;}���>8g!l��6������p.)�^�~_�s@	�j����}{�"�Aq�~#�c��)�(rA0��]�a}8��s�Yg��~[.��,�_����}g	ܡ�P��W�@��ZĔ+R�]�FW�.uƶƱ�PZ���:-ORM��S�ҟ�\������ ����贿��~�zvϬ[�;�[�v�(���E�\x�_������y!����3n���������Y)�XNr�Q�ziԓC���'V>�+ioU�m�(�,w~���z֞��K!�G0V�/v��C\K���?��k���J��x�a��^���:�!X���ndyRؾ�I!�祰�/L���J��gG������Gы�Mֺ�N�C��Їrg%�=lјѽd~�}������^DcQ�V
�=�P�M��>����<~�,�>G��Fk�#�2e�{ Bu��2��5����.�����6� 9�S���{^o�y�Oc��^��d��j5�h��"��ui��a`���:�+�f��"~�_�x /�1���+W�H1�>Q�)7�S�� �}ݚ����Ś���G�Ņ�,��x��\��r�0-
Z@����/�rjF�_�=�_�I��2�����A�؁x-z_:N]#]��H����s?���=#&"h,�џA���C��gh|	��חmiAW1"�)�HV�Կރ��G��M7ݔ�85o���}��;�h�^1��8���/~�w>��4�݌R�тz��o~�7�x�aq@h�0=��Y1�~D�O�q���R��)��&�,:Y>�z�]�c*���v�R�2(�B2J&2�e]�-��yJB��Q�C�аV=V˵�-�~~�P���Y�=�s`�{�+^a�y0�:�΅B4�g�������0��̈́��,jfy��q�������*�H�PD4��Aޙ@��}���c�,7VaZh�D�x�Ɍ�Y���&|}�T塘�5���C��3�<���og��G.���?��ˢ����'Ƈo�T�鞙����Wq�vu��1֎�&U��\<�rɬ�v��L�<=l��ΏG��~���&�b�b5�����6����{�"�_�I�&��5���-=����
���h��G<��o�鷃�Z������J$��B4�Z0u���4v���Tϓ.BZ=��b�ڎ?�/�k�,�d���l�"_F�����4ߢ�A{�0٩*Zp�O�Hظ�{|����[��S�q���?�㣟�������%Qyv�϶�?O� �#7��S��DO���\T�|�Ᏺ��p��h��Q���G��w�����xp��U�+�h�vw��C��Z-�,�Ks�RZ�aÆ���^��D��v*�k%���TW0^��r�|}��DI���¥~(~y���=%c=ݶ����B.�7n���v�/Nd%�Y���Z.��̍����0v ��xF_��+dO��Yq�Iy�B4iq��i�>�����@Ź,c�'�=/�S]��ո@��q���.�<��ȌS���_���~������V�`�EG�B��ʯ��OZjB�
�sd��z���'�����)��p���|�q�-#):�����̙��W��e�~����c��c)'=IG)�UX����k�w*)���&�Ox*<!�89!!W`�$�O')�<�W�zo�����!�c�9��9�~�Y�
�(ɫs�sy ���/��/_~�G?��w�m���<^��ZT��4 ���X��.��ҷ$õ?�;{�"����:�dF�g-zr�XK}�L�^cYqx�'�����1���Nr�_����h�X1�1�O,�����/|w��[��T���_�����߿��7\s��M�o�T��RXr�YU��M$}֊����2�a�714�O<?�(������q=��������o�г���Uc���]PH�k��{�`m�+$,W�IAR�bŊ�ɷ��,h%=�7�=ďC�p������V�C笐�^�|��7��y�I'���&��骫�z�%�\�!n�q���1d^h�����},_�(�䓻S�D����g��[^��x����/�QP`-�B�y0����P�ђ|���{sl�og��G����7��w�m��6�n:;��]
�zqmo����+�O) ?�䎓��i�mb,��b�԰�jõQ
�Oબ�q��5�dg�GY�x�_�����G�R��0~/#������>��Ǉzd�J���RH�ڄ��zƆ���?��?�Qu�x��Op���;��7\{������x^�c���șI�
e�=���O����ւVTƾ���-��Iw�������]-J��9}�y{���j���6Z��L�D�B���*����y�����[�����~�����-oy�O��M��^T��R����
�Qp�V���sl�뮻.�p��H{����I��W��"���o�#��څ�כ����x�O4���81���>�+���L��^#����Tq��vi��9�3�_y啗���kg<����4+U��\A�+��зU<�����pǈ�{�ޒ�I�W3Δ��h�f�;�!��� FyGq����֊�W\������n˾g��G�K�ȥ��M���OƋ��Ύ��!�Rф:T���PK�\&Kd�kr0@�!x���p�
	��Ysf��j��;n��N�O�&Չ�+tuu�[�[���w�p�	<�y��{��8P�[a�}��YR��r���a���	����7��E[s,�{���/������*q��׻��X�2�a�l�h;��*�v����z��oG����9.���줮'��kL����d��'-��������u�kf �)m�ɛ_��W\q�;���/���G~�O��d~��#'d)7��<���x|AS�2�
u�}&.5��"��Xg���)/�XY'��/���:�c�)~N��؞����}r\q�f��tW�^+�-Z��YO|wQj�$�?��u�\s�����q^����W�σ�+���(K��m(�������#$R����d��z��>
�f������M�q�^�]y�Ag���l+'�w�����y�{����\saT!�tw/����Cx�f�{{����ng�q�s�����y��Y�U1�r#�6�Y4;�fʩ�ҁ%�v�����+_�J�c���8;�.��{�0fY��9�����<�Fֲ���!ت��n�������:{������+�,����#������^�|���H!-e$��x�\&���*e�|R�I����h�<�`���8a�G��w����}n��n+�:��������ݯy�k�sϽ��q(ύ7�8��;Z�'���|��P��^\����M����m�������ۗ/����u�Y���ٽ��.�&�&s��=��me��]<��O?�l�n���mrmN?��M�������O��O�|����&"i�p���P:R���h㦈������1�&������=��1������ӎ���ۿ���+���}�����?+ޭ�{�����7���#������{��7g�x�:';��	�T��	���|�é%�QU�B�H�5I��3�C#�+_��׿+Z�+C��z��Z�kD����+��s)�����a!FY�8�c��ړa,�����>���;����x��ZI��"���7�a��o=����-�&W4�8&<�x�6Ɨ���g�]��O������{����	�w[�� o{���>���~��{�%��y�Q����dxy\v���0]���WI$CV~R*���L.8����YSa��JI�aҷysR��`F��,,g�rV
S.�=���R*ل��;R�YRuk�4�`pB��RP��;E%b�����y�m���@���x�?�;g�G�F�#��wߓO<��/�.]J�w��Y�f͉(�6'������q(��bի�#Wz���z��Fp�Xyka��%�F����x��h�sSk���^o�F�go����9ȧz�Wuu^�ˮq��R�G�X;���@�}��J�8G������m'ʽUʕ�;*b���Qf����8�x惵�����rg�(���R�RI�zŗꎇ�}����'�\J[ܛ�{T����j_<��{�������C:�8����7��(m�������W]uUwTB��гf͚Yq0΍�DԡS8�y\��%j%dcJ�n��f+��w������7�3N�2Ǥ��5Ǥ��/����&�4��1��uR��'������~v,���qL|���K�������x�~W�Egէ>���ƒ�x≏���?�hT������R��n^�#�e�m��3>*<w�7�d��g�W��H���Low<^����.���,����w	r]�d�Prz�K��^Jo���&��4����@��@�����uB3�;�Z�T��{���;z�I��ܶ�1�W�XfPƱ�~�u����gOs�1�V.��~z�;����y��ٳg/�ے���.u-;^�A5~n��{:���������k6��㸩e�|>_�h��yvM�l��`���K�=*�����54��M�D�%��&��9r<�cw .��K�,�׭wٲek�9���7�%m�?9�l˶�
m��r�i�Q�{O�d�&�(o*������k��Z�%�z׻n�nm٩����ҖqH�M�J�������[�Җ��@i+����-m���V�miK[�2����Җ��eJ[���-mi����oK[�Җ(m�ߖ���-3P�ʿ-miK[f����^��2�R    IEND�B`�PK   vOX��n�% �, /   images/c1d4a215-2c3d-48ac-b15d-f6239b4c4b94.pngĻW[]5Z��/��w
/�xq+���^,8(R�)R���w��������;F�8$#cﵗ�9�	�J
R�(�(o޼A�������&��EB�~�=�.��"%��b�d��LT^�͛߱�����vҚ�o�`t�^0}� c臔Nߜ�L�,lm( �&o���9����ٸ(���?q�s��*_˿y��&�E�w���Gҗ��Qj������DB��i�Q�|8\�VU7���IW�Kj�o� F�VOL�� E>����0����a<l����6-�g����)H���(���/D�tY�d@��� 
$���������~��2�]�4)L�ׂI��������� ƒÿ�`oBo]v}�]y����C@�7�����u�aM�gz&»o�^5��s��G�i��%���bQ�@�A{�&��P!k�p]T6��a��V����k_3���2?�T/9�������Tu�X[��I�H�4��-X��\­�����Y �dO_#V��;\�|�)S���-b�\tQ�g�%�{���UQ.<�-FSq��#=��Q���M2���ʇ�����.�	�`���6;M�t�{V	��E��Y܂=`�$����vO���8h�Q�s�����7���� �Y�ǬL����1$�q�aw�L��T���@��_s�k���5����u�B���j�ً��mcs�%�"'@ջl1����������cQP�WSGX�������|�7������n�d�dtW�cJ��kh5�E���Fp�nwY�><����`������7��a8�9�TjjhBj��!����d�^n;�Xgvu?��`s��8�I�Yg�R�6{Ր���9w���}S8WR����M4�j1���+U�o�0r��k����O�y�6V�5�FXfׁ���zcH��9��mh�"T�	'��[DP),Z*� �T���(�ni��tt&�{�w��(U�{��P�6��mWx����`iX�Pp�� D3n#�O�}sGn�3!��WN}��B�=!Ǌ������"k�\�N�'��	�"�z�>Q�qYǍյ�ҟ��r�֝�8�����t,��#VS���e�9S����1��}�"	bX��!�,ѷI��{������4 ����8���������V��`p�|�l�D����ٷ�ldZ�*a�d�Md^��5�,=al��Q�/
Bл�oYT�6r!�?�罵{�+�nQZ�`�Ze�P�\�u�m//�~ Y(����C���bm~�tA�/a�i<�@&%��j��JK�l���rf��A������\��T����jmڊn�2�b�`���a)�:��v�	�!�K��ζ�*�� ���_c��ABίP� ���z�ߒ�L��t)�?�h�����{�<C������)��@�3l+��U�Dcؤ����=�� Jq�X�L�n'��av�I�b�ATܳ���bl�Xh	�}#���^��Es1p��^�v��j8��IG����I�9� �d�dMč�.�ފ���~�L	��Tׯ$�Y�ޓ{iS�1�������t�
9W�x��Cx�x��s���>�_� \������8�)�H2�����剗�kY?���L��˪Y�W���{`�VQ���l�F��:pGQ��c+%�\��r(枖?��T�<����:���eϰ���B,^&Ki� �ʚm�	!��%����uX�.[�T![��As�vD+�Z��V�����¤83��6p�B��
ˌ7@�-�;-�.>�����F�ޅ_;�'��0�i3ナ�KZ�ʅ�/��������*���C�����ֽ��@�>����C��qA�|Zwh[���Q�3�Mv��%R�ߟ�Ҷz�g�N6���}� Υ��߀k�z�u6�����\�1n?�qd6x��w�)p�k�G��\BZ�ì�γ)ЏQ����5K7BJ��p������ �Sy�%j[�2�x���>;ѱ+W����m,lb�M��SnY��!ǎxyP<zK���kn�M�@��R�Lֻ!�����	��BE˔�9���Q�t*K��>�j�˚jwVw�}�~�$��(��������|����c�i�	T��(��W�G:$]�J�"��Ц`�6�[[]��QV'���eWԗ;9��ذf�XVٲ�/�^���a����$�҆i\��Pi��H�A��[��7Fw���^bV�P���݉���m����q;FK�|F�5G��vW |�c��4g�^�c��"�H�s�=U�Q�y�tǜ
_�S�zr���+�u|,�フ����kPE�`Q��� �>c[��$�Q�C,m�����㘔���y��_��Ʊ�s���ɳ��{��k*nVg2�u��1�k��<�q�go^Z���m}g �f��د�&�ab��	,u�iv&�����O���L���P2�V'��P5���2��ύ81q�3ZV��̗$*m��c{p��A<�q��e>w"�I���(�.�@�L��t�sϿ�W�p'Ki+��p�of{�ӻ=��R�������P�Ly�8�'̊�-����/����N�R�Cy��e�r~Һ�m��-�60�������<�|~*D3��x��bF:&9��PM�����r�d�OV0��d���e��-p���C�jq�� ���Ȏ��� ^�ī0�"  ^��!ݘN�II��n�Q�|'WQz��Lr��>r=`�_��������Z �������.~�zσvX<��Mޯ��.�IP�GL�n-N��ia�	�9��6�I&�K�N������0�O�()�g���\��0�P��j�Z�K��q$ǭs� ��2�7dK{Ֆ���u����3 ��;��r�b{� �$RiӜ0]��p��- �M��������}6�*wl|��_C4m|y��s	*�����/u5�f��{W丟ge���0�#�I��S���P�CR���w�g���"œط@5�M"e�ڷ��i7��ȳ�U'��&)H�,>�%�� 㤃I�R}7�i�@��|V�""��\	��G쓂�內$��r��di
x�X��Uo��B��I���b!�A�C�&��H�������+��h�� ��qmwR&x%��2�gzl-:L$Tʾ�Z!t:�{��!�tr`�������`��b��2��9�q:}v���f{=�=uHy�+و��t��rΐ����W}Q'��z5~@ʺ�/;�d���¶�.����v�=]�Ҍg�r^���}_C����B�� ��;�@{�źO�O������<"_�nYȊ��o�+E�@�(���g(�.e�^��8��.�B�dG3]��DZ#��ѳj7̞�c��;�h܅��|T������8�nai�ߝ�����gO��1�r���̾KY�@-�K���矚D��%�1U���;���>C:�_��:�Cſ�Aѓ�6���(�}s؛������^��Q�t�ͨJ!ѼX,���	;w�5�ۈ�2||��=+��;3��I�T����|{K�����E��b���m�$+����w�7$�?n@����.1�����FQ�iX����G����e3���d>�mc�m�H���w� '�<�q�%^� 1#6���[r�v�E�Qo��V����^{ǩ]ҫ���9ۇi_G�Ȏ����򨳝��v[���/*��o4�㰧�y��;^�a���6B��F�x#�lf�x9�D��ws'L��R���u�-+��\>���J��\��֬��c��<zk�`��sa�!�-M�/w@0o�w�[
�=�{{"���=����33�4����8�"s+r�K�h��B!�����k���P�Ǔ�І��`�����b��?<;	~�Ũ��H�f �����F�?{"*i9���P1�.�Y�N�,3 DSՀԖ��9����N����e"�j해��Q�HA7��z�>�q���Sj�� Q��2' �*DN�/d^�[�X0h?���t��Y7ouf�I,��Ƅ#l�Ϟ�A�b��Փ��1�\��������υ�>_�fL�?Z�Q7I�`��ﶯj��z}�r���\����zV�T�������5v$�}e-q2�H�R�R��'s~Ķ-$?������ց��2�M����UV��fg��	;��­F��F��s�]W�G����d�W"�\�1��ʝzp�*�5��I%��%�f}�v�ҵ��?L�lGM#I�Ez
ا�1��&K-�$9�k��i��-M7I5�*�ђ����;f��|�z/���N���?@c�<��������/������})�$�-P���{E!�Š
"�^g��茤�+g������Ձ��I,���Los��'B�d���G�#8p�BVƸ�����3�ȯ#wiz��nB8����
l<<ּx���m�u����H���t۷B�hQg���({��s4=B�� ��
	�P���= ˸O���n��uw�b�v����<A�#�uo� ��"��:�$q4!���8���Sv\�S-Wץ<�,�uJ��(m~�c��p�$�"�_ �w@f�)Z&��ๆ��qE�2�Ϣ捁:m�
�����,�����1$��V��-	u�c�?=�vR��뽖��~�&�j��JQ ������h͹P2�;�H�Wb
��_$�갡I-�eL%�u�i#�ߛ����k�t-�M�Ȣ�ܣ����%B�>ZqH�-������r��" jt\u{��$N����ѝ��٢�ʴ�B��S�W�`[���d�%�6�(��r"��F`A\a#���������JH���F3�56�L��1β�\+���0���1�X�}�Z���#mJ҄*���w:h?��ɺ��et)#CMJl�b����9��AR�XUn��q�Xewkd�umL@y��E)��I+�7�̇v���p^�ӇR�T(̼!u��ȝ���_r��-r�
��@��v[�*춯t�nk�$%HD�_�_0*�b��%��\�)=Y~
�
�f>z�f��DҜ�[%��+7�±��;W	Gm��F=�Pȵ�${�6�F:��E��;�j�4�KR�7a��SI'�2�I"�	�)�r�F�ct��a�<��<�(;q�UfȌ�}���Ȫw��@K�䄀o�������s�H�Q��k��u���t{'Pwm�JƎ	ƚ����V�s�p�99�_��q0��0{5�+8�����y�d��,�B���R5uZ�B{l�ل��T��K�$�o��%">>��Y|��M����>�����Ȑm�C�U,���S�Dq<x�*�
$1Ԙ�^�4GE�P�ц��m�ǈ<"��:)�E&�^P�87�^Fw̱s-�)�o�?שS�����`�����g����ȧм���8���j:�O.�*��@+�� 3{���N��}3N�@��w\G����Q:/�����=�Y~�uo��Hr��Yc�q��Y;s�wb�UB7U��+L�5��b��o�����˹���|�F�J��:����P��C,kP@r����[�D��`�cj,eȆ6�#�Ͷ,�a!���qfB�fs�E��\P�G��[�S��T�m?�K��V��傢�u �*��ޤf^�hW�l4ä�1���U��
eǵ�ʋiw~GAT��9@��� ݜ�����s��Lq�!?���2�T���$C+�p�3�m���.�s��]�IM�;��Y�NtWDj��ty��h}o��[�@q���4����/����G ���wu��^U3�i6�ٲzO��R���M�J9�hx����P��~���?:���"�6ۻ�p���g~��d�G�(�S�>E3���Մn"��4k��������LU��.z�
���,�1aL���(B��Ne��-�؊�c�@��m���Ǽ�9%d=�S��vV�����ى��f�r���;w�L�����0̷hW�1'&�۳����6h�\<˗��ُ�!&e�=�*t��Y�1_t��}��v����V�ߒ&_���a~c߉���}��=^��5Ar�]IN��Mh���PpI�Me�^�MS�{�v�C#,-�ա=m߬�6:�6޵�y�<Ip=����uH�cG����J�n/�؂I�F?l�?���� �xK<������u�b��ngD8̪��}��Q�x����ǃ������������UP4(�^�q��{wH�oF�?m�80�eA��Xj�zw'��O'�kM�v����s[��Ў���	Y��o~�%�X�����\xh�sz_XFI_K�����9��g�`�o�g3��:g�)t�i2�6�M����I)�N��}�����ďo�^1'��g�ƞ���O����7>۞7\����}v=�R,H]q�L_�f�o�����d��M�(�W~�/޵7
��莗O-BSd��E�:61�YR>F��As"N�;j	�Kb9<j�����BI;f�t5���_����-�3X�?Bo��U}�k������?��|��t;ρ; T�E���Kb�H��Fshߘ//h�<=H�|�-҅,�^��Z�����\l��i����!����,!���Ji�����#�+E?�#3��%W9*��j 2B�UO(�;��/����>99��]�:��|$G�m�^��&�x�J �<��^:�%^}���t���%f���[��3Q2T�D���r$^[�8�I���V�H#�e����ڒ;�s��ǹ��+^ylP�P�JE��3�(��,iŉ�����~�q���7:�%x�@EZ�N�괪{3]�m�Yv��Dq������_kd�f5Y'�ߔ@�7�N�9�;QAU?O��	ݢH��1���w�s��Q}{
�l~m6���ה�a
4�;g��k�́Y��R�2���-k�`�5�&5�&l�%�:wh5Q��_��L��,���I���T�ƫȵ��9�!�,���ͯ����v=0���X��0�'���͂{���.�(d���-[��X���#�������ēh���Ah�i4$�S������xVd�K���w��iu���*�(����u�Nؖ��T[z���Nܴ?�L�z��!3�y�C
Y�Ҙ��l����O�
~�9`��7%�9(�v�!���.ZU�<Yĕ�)���Wb�2��++�^��ϧ�$�����T,P?���m�8;r�9{�~�=��WC���&tWl�~hβ�Uo�@Ic�(oD3"��:�~��O���й�6����5�%iQ�m�@�:�v}�\�f'W��:|�<�i��yH�lψV0y��|D|�Lߠ�V��B�H�+v*v��/1V���'F �th/�.xzf�K3E�*6����J|�r�)�ME��p��4>e���q1� y{{s��9��k$�� I4�	��^*�#z�|�5E��o��4=<T�]���N`]z�2�3�4���i�z��e�d���q��!�9�\��+Ӵ�����w�1"ޠ��d�|قB<���'�2P��;�A:UZ�+Yy@tO���Q
_���Nl�0�e�E�J@Hc3�E)f�_-�� _�(�t�~�ֺ�u��m��ɘ�3�����Y�!5`�6JNNn�b��/��dP��0��X��5۩��OQ���NH�_��l%���:�|������M�[�X#]���(����L�PB�&��|�a���۞����E/�O~�]D4�9a}�I2�ꪑ|E����eǘf=
$��OL��x���rTn�ޱ������M]�m{��;�C5�,V��v/	����W��s�R�'u?9~_q��H`�P$�e^�;=���]k�s>�.F��j�8~+��^T�<б��Y$@�w�i�����ekڬP����G�_E�4F�\l�{�m��'CI]�sQ1м}M�m��_Jʚ�/&�C�Q��׆	K�U ����ٖ9��S��ߐ1X,~�ǫ�������8�ʨ(V�B�`9��@w��W�`8V��j`7�w�.�9�[-3��C5����_x����oS�H�iI�Q��~PǲH���)	M~d��%��k�'�8q~�N�/o��$��k^�X�Ɬd���y÷��Q I���o@�q�1<��|iV��1��8�2��Z
�ҥ�O\j�z����+o�K�;��0�'C�<(7�(���﨡�T��d�8:�ߒ�>���~�d̈́8�ܼٍ��u��{~�h�Q ��H>cB!e�P3~c�֋��*4�n��Q������mWg�j"�1Õ�JP2��nb�2���$:�}�����!�`OՍRHJbޡ��α�?A,�8�%��I�j}Ƭ\
A9\���f�(�`W����<��@y�<n�CA�$+Ǘ����і���Oo���hF�c+q�����*�r�ԗ�J��� Eq1z�/�B׾Sr7k-e垊ڠ���\��u�l�m�&�*��C�Y�2ҡ
���g^�nփ�k��MLFN�f	iFY�!9��J-�ź�Ͼ�����E��X�,�GU�]�t�h��oe).K�_c%���4��:�_�;��vUޤ�ݑ��9��w���D�N��t������+i��~?�
M!8TTW�}��ӯ�Ν�ts������n֘�mrq���Z�#�f:��CVMG�z��>��策Qᗨ�k>F�߀�A��ϼ�hH���b�04�]�U������fX�`m��΁�<!\�����ǝo5���e��M2�6� ��}���=��|���W�7�<QG�,c�u��Ӵ�I�G�ߡ�BZ{h�I!�EG��u�_-2��z��xl��A<�$�ޢj<߯M�me�쇪`ٞ |���N�nB���J��g[������獃>�5KR�z��0��&��lv���"�hW�Hz���/M�(!Tj�Ճ�3��6��ܒ�og{ĥ��� �N ���~%4�jB��8<�z��}/��� ���Nִ���*���S��
,m1B^hi+A��&_Y���X�LB_nF�(V�T���0��ʠ��8���B��bS5�rHb���"Jɘ^>�:����:��y�Ϙ����b��O�.0�uf I��3g"�zM�!��&�� 6%�zld{�YZ4�Ҝ�X�)�pR��>T��$�Y�|Z�_>V/�8p����$r�{�{\a-�Oz��Uu?�*YK�����g$ݶV�����ȼ�q -.�׍.b�� �{ܻ����/��6����-W���t�
6$6Ie҂բyML��i�&5���(��nӊ�#�-��}l���W~i@�W:�uG&fȋ'�$�YE	)���G��s���f��&h7���
U��~�Ķ��ؚ �0�O:��<��p$der����^�������b���q^������0�n��B��'��уRd�_���E�j\���}��ө�}�C�Q�ʛZ_�P'b0xf�o�g��o&�N:�W\e��^�
Sz����Rîʎ{IܦVˢCcC��A���TG��M��S?+H}M:�d-�͑�[E�"d��z0\�y�L��4�/GIu�]-��(�8*�,����~�CbD<2���f��,�.nӄd��*CG�^ke�h�$ ���5f!w�IDو9��U�{w<��e��|�V���Iv�����Y_���?������̓'F̦]S�Fj���_K���E����,n����%��4�p�n��A���o��-5) 7�)���c:�v�X]<�˒'ӂPV� T�2B��&6A�Q�z��fJ�bY���-�5y��mﾱtN�������t'����^���b����I��3��������)ڶ����^����n[�S�+\�uX$��9�G��F�#��C�1z,PL8ϩ4��O�V�������Z5>�&�!d�������]XRL?D	��2v�u��O}/?��M3_]�0H�I��8�4d��I�H5��>�I�6觪اƳ�'���Y�o'�+^�\�.��b��*Trm�1C�����Mi��ny͊H��'�ď*@�v5����ӠXp���U����a_,�Mi�Y�i�h�*Q�����NU�jX���Q9�0�f��8<h��
C'W��ufצ@�"����G����X����=�|<���Wu�Gf��l�y�����s/�6T_�B�Vש�F'��������Q^�XM�P��tS�J�9gҠ,�&)��wy���ʡ�p~�C�X�N �����G�u���Z;�Z���e�����V�(�A[������OA�y<�����^�r���U+�����g��{ޠ�	_��Ũj���/
�^���w�����d��޸��)p�k�2�OK�C(�?]�e�ҖUյ�����k=bd?$�J�`n�ږ2�]v]�2��=Ycz
(n�ټ��.���?��[�������K�M��_3E�{��k�J�<-E���n$YO%ځ����$���x�`-����yQ���G�	���X�\IEj/%R 	���~���e�y�b�2S���ҩ��3���d((�mZ�Z�?E�������5��iI�|]sܝn
=j���)�����f���L�f���<Y���l����D©Y��Q��*����u?Vʨ��� �6f�`������q���y���٥鎮�{��b���j<E�����
CZf�F8�Z��p����<[��!^V�cd�H%'��⑟�xO�Ϩ��[��"�p-`�-v�N%��A�	�]�b��L�f�5�_��lk�����JW�%��(��{��:�&4�[�B[;�����9��g�k�c�w�ʱ���D�U�
�!,���Q�b@3���C~���0_�I�w�]�,�m5<e��ln�u�����g��I��������N��P�H�pZ���u
<F��x���D� *���e��ɈL���t�����y����	ٖ� h#����q�e'�QL83Ӹ��4�<�"ק�9.�!QL*d��Xw�X��=e�:]�@���*�-RIT~��{=�A�J>�	�葛�B��e͟s&��i�*���:Հ�F.�1�!��D�A����/�oI_	4�f�4݈W5���/)�ԟV�B����ic X�(Ť^�yD�����=K��ͨH$Q�ϯ���Z��(�Ң��!t�a���`~X�/�fS��$����6�(� ��t�L�uex>�x�]X�]n�@I=�t��ҕ	�(HA��F��{[3�Z|ݢ�5�O�]^?o��x�q.��o���[�B��ԃ�ٶlM�����؉�3����&l���m*[g7Iŧ>RǏ���3�c�l�*Ɣ>&���~���I<��>�2�-e4	�J=���1A� �������%R�m��y[,�E7����
�!��
���d޴H�{�N�(������nӱ��앢c�n�%���}���ӹe��'�m�f��]}Q�]o:��)��iD1�/^�؞�3GV_�uf�|h�����q���p�V6sO��ao�����pM,�����[���7��x�b�%��i�]b��ҍ9�.��&(,��x��P�[�=�ݓ�#!�Vs��Ng��9M�����v6�h3�k���)��S�A2�SAq�����A�ĺڐ��R�?��M���u��E[�{�&�;	�g�a�~�k����n��R�K<Eڳz��*� �.w��z������cև�C��w�&s�;ye,���Y�3��#a��Hp��M6V���	�� ��o��<u8{f!*j*c#�F��v��I�a��Z�����:���I+]X�an3�&� W3.�LLZ��f�����;�ײϜ��������H"Ukp�L�Ja���OGX^�O)L��qA�۞;���si)���>wi��í�k)���<@1#��43�\Y��.8w1A^�2n��ɣy���b���X�(�2�r�d${���?'n/edx[�{m^t4>��*j �]���VxA+�� �m|�.�?�k��3�1��,]�h1\�'�z���$�󀛳"�`ecD�|�+����=�O]+Ɏ
�M9p Ța���9?%�J�w�#��\�=^/�����^I�f߸U�2�΂�K1�ʄ�t5���x0h±�������}T)e�	'��L]�z5��8ȟ�C3>TB�.���\)�ʸu���3��p`�[G90�-$����D��p�[S��,���ٙvX�ci�Gi�6ex�Ү��,!�$JH��z���2ѩ;�/[�!6�� ��_�hq2�,*ћK���MGԥ��X��i�h7{��@sFB��K9�s��-�p�._��ʰ;���H8Tw.�;s0Q�ry��n�b��s�5V�&�Ϙ�H�V�d]9k�"��Nl��s/�g����}&C��r�x�18����X��������RA1��Pb�t�Pr�D��}��"�wv��E�~�����{�Pd�1���@Qy`@qI��jn����"G}7D鲜���닽=����i$�P�IHZ *F�X��x#w��8�$~��x8�$�U�N#��B�\sk���Z!���i���dj�N@��ݩ�����m�q}����o�-ML*��5C�uh��2�	q֦1TpNI����yS#�Jw�Ut?�	��x�����g��&�_a$N:q�g�R+oW|�
�� ����xQ��WԂ���{�a�~�� �Sv%\Y:vP�خ��:���yW�c�:�O�&��Ny���V�-�p!��~�s3����;dH+���[�%T���sf��s"�^�į�TU#O�<u(Id\���(J��w�6��C�wF�la�d�������.H[��2��vi��K�7'���'k�}� i:�'�(��*Ͻ��:���B1�W#���˸�φ������[�VAT�P��C�N&���%r`-r������~8�a���5!��<�$�f�@6��#��AA �t���h�eM�'x��V]i���_5&)��|Ǖ\�L�efܢ�[�i�u��`.�mg%��
���!dOc�>:%���u�xO���-����8�N������U�քE�3G]�C���l�/gF����o'ȕ������އ9�i�6�f�"Q�NhZ��ʴ.��)T)y��MƐUE�D��nd��h!��g*㷁����q�nRw����lAb9���P&Q 빃IB0�4{)?2��L*A��w�D�E\���Ŭ�Md��uKG����t���V̲B�
���u���IJ�������}����-&K1�6-�%�+�ػIGT�le�VH@Ihۍ<��Bwƺ8~$�T�L�@�I{�U�5���^&,u��w1�8�f�}����kvpy X�݇(S&��?���$@�jN��@+*�4����-�,!^s�,�}���	?��gO������Z�	��0��s��'�,��8�#k��Z�9*����+�r$ن�z<ab�$A�T"�p�k���X�Q��j쪖=%��[�
�����S��{�-�?���3g�xD��|TB�/�E61�ck��v�#��i3Үb�8�9�!�_�z��Yq��?PgM1��~֣g���l2To$����ʺ�-)���~�7 
��R7ۼ�����%W���O�����Y�7�p0����+r���wa#C������#��?��C��A��zw
Sh���%�J��l��JxW4��d�{M�p�LI���ߢ�Ut��W^�߿�1�>־�)�����v����a��K�X����R@�;�Ee�TX�z�y��鶱�;��:刱������>�g1�R��|��z���X��CM��������ZFf���U��m8�d��ک�	&���U0.�?9�`1VmY��Uz,�/�����2�7������:�#��?��x����S�"��.M%��z���f��p�9��p+�_ք*õX(L�=#�y�jJe�ONp(��`��p�_�s�"�$���*�i�Ae��,��C���8��vc�u��ug�;,R�D�U
#j�e��/;�P�]��܎pa&{�A%�f���4Eg���sR ����y��@�&�sE[gs�r9�K��,�"�\Bf�T��=�;)})���~�F��1W�W+Pҳ�@��:T�N b�o[�����a���z�Dm0�q|�΃*C��R��������2RWM���"q�^0�r��Y����qX�)����a��]����qlr�j�93R�;��^;���Odo�Z��̢���{ѝ\������4���l����#?1�/)YTR�p��Hr�j�܏��������V���UG������.�W�(�SJV�V��ೱ��m!��QP*-�,��R���� ��AO>/DѲ\.޼`Qj`�-�=ZEZ?�g�R�r�!*�o��R���IV��}ƌ$�&!���؃��v�2����J�*ڔ�C(JS��w���|���.gr7?~v��(>��w��Ug�R���m���x#�>��G,6��h��9F���p�*r�W����[�Xǡk�fT���C�2n��	��6xy�U��Y��p.���X�����'EW�[����Ӻ�J�f�n��쮍:0Y_��I�]�̠D��2V��6�81�"����SVF7^�6���,}O޼cE�{���E�\�M���� �蟵��9?��k6�m�`9(���h���'�6�|�F7Z�Hd�dF��E�kM$�%��&� J2G䌚�I�D
���/�ңmVϿ�xU����z��_%�PZ��D`;��%gw�y1�e��.�bQ�X�_��/iaϩ������~	�����F|����L�D;�9fZ�~P<��쫊$�jk�:
qq��)oL����Kێ֟�K�N?�dp�^���􆣐�R�y�Wrt����OTO��yTcro��B����ߕ�v��"�������#J�w����<o�뛭��T���􆷢҈N�ɼ����0��f�������t�f~��2)�2���Q������Q�3�@|��'N�`;�x��T�[��R.6N-e�HH۵F�Z;#V*@�t��]J����8��q�]�Z�����+�����7���}��~���&`�%ݽ�vR�8��l�ak(�4OǗWU�����}�3�?�@�K����&�\d��+yv;*��3A���F2���<�=c���
�@�0���v��Y�Q�Ul"}����a@ߺU2�����{�+,A���#��!<@6�!���C���Ê�2#��sh����Q�]�u�r�a ���x��;M(�T�ˑנ�ݟ��v�>��������}
�,�V�oH�L��Ş,���/D�$@�0E�V�<�>�{x�h$��uJ���+휚�͢��Y��̅iƪ<)F��0��d<d�X�����I���	�Lߥ�������	cP\
(U٨:i�˰}�&�V-����� ���E��w���4�"f��r����1���Qŷz�� �{�ڍˍ��9����Bn���?("܂3�Spi�>�/�{��eJ��V��.����	?6��tZbJ`�)Z�$�?���0,.�S�cߒ�E>�p'������uG���
�K�T7P6�cHFI��w$	X޵��?X9���=L �&�<�+���}�x�d��󮘴��U�B�}]ӄ̮G��!�&�'��\O��$�NMܠ�p��z�eF_��G����1�?_E٫��G�n���5`�r8����l�<+X8��2WA,A�(>]��Il�i� ^��I�����[F���T�~?=�`a���������1�_-�L&�@�~����ڵ ��7ܥ�.��M�XͣD��ԧ_����d~W��1�ט&Bw�Q|H���BD��RD��|�xy�U��N��_��l�&m+��" ���q$���N(T�w_V[�7.N��9zl�A�>��vĻ-��p�S�/>��h����sf�����U�鶙|��UE����.��uz�?i�(r���j?����~�gkn1��yr�1��7�|e��$��z�H�����f�w\��BM�Oc�Ղ�-�����h�ܲy�a�DM�]X��登�z��#L�ơY`�SZ3�=�6>��ܔ���8�J��J�iw��r	y�Y�%��nG�����Gl����鰤L��"����O�l�N��&600�Dc��C6�\�DB�>� ����I{ʈ�R8$n��el���)�ϒ�Qړc~�O�~G�^��r�YDʣ6�kc�u��న���i�[�q�� �Qo╲����h�P��	W�dg�)J���ǭ�k�5�P`�8�BN�l�� ߢx]i�Eն�}o�}_�׍����+9=h���z^,��!R�ϡ�w���Y�ٍx�Z ���h�V?��$�!qvZ�|d��d��_CJ�j�v�.�y�j�9﷉��sx*�O46���p�2U2�E	e�By�|91����7S�$}qG'�)��Ub	��F�Ұi���6& -�\�R��2�g�Q�����_�u��5��?l>X���m�ʷ���t�!�z4��Ӳi��L��GJ��doP�m�XMzz�A�z�vT`v�-��xr����#ci&*5�;��Z�d�,���Х062�c5��Έ���08�B_����96�p�rt�굵碷��?4]c\$���l�f۵����6�f�&�6k��Ͷ���d7qr���|�w���չg���J�A�:��[�;�n�!	�W�l��f�3awԸ�W|v:�u��$�(�zV�
T��CK�ۚ;:?�@���C|"�a�2q�2nf���8��,r��P�,q����J��O��5S�o���_M�����,�/I{y�� ��_�Ƙ4��Ȫ.����o[ZU����)d��V�|���ͶG�︙j���K=�),��Zʉ��U(�!/W�3U���qF�FT)�#��a9g����Pi���&���jh�!4(�M�qnGB@&+��'{V����ɶ3����5�p�yJ��KK�yڔi�t*����%�d���uƯ�C����zE��jY$T�')���H�2>?��`����`���I� ^$�P����ڽ���]�aV=c��y|@����󄶓�'4�h)2�#
@�Tݢ�X*��B35����O�7:*в�]� Jk�m5@2T'mH��d?�M�ܿ�/ p��[�{������9I
g��~��\¼a�V�4�Bc��5��X�b\Q;�.���6�+Q�	3,�4�F�zD�<[��3�k_u���t˿��9&�=�=�_�0�g+u}��&�U�3��Q���L��j�i����� �9"���/���0��P7A�9JG�)pU��~���z#�XS�$�>`*��(�FŹ��0B��6���a�Ͽ���tQ	�k��D6"�����Mu���H�%J=a�\&�h����p��1X�g�4���Q:� ���(�����0 R�A�h�i��O˳/���_3��L2�O��5Y����+�����9���T�C����:�"��B�_s�n'�^����o�����ϕ�SO�����K���������5��B�����e$���qp&�W���x%����Жp����S�ha3�?j������T���C��P�6I�~�G�� M�
z(k��/�'{9��[�i!�݊Bqή�,�P
�t�u���%\[/�~����}��D$�l����u����������a;�� �G�}u��_�%���:&)�@�B�L��'{}�c��ܯ�����s�j�v�+��P�X�d�z�Ʈ�c+������$�BR=���;H0)��JayOQ�;i̷T⛮�.�)U�ˮK��r/���|�V�v�w�U@�1�������i�mw�K����ә����M$��m�hp���t��q��0�,�~V*|^IY�}ԅ�T�L�r�+*��#o�,Hӊ��$p��S-�NiC4��|�~ny}[�r�R�xΎ"K��1��25,��6!�ҀS��
���ތ�G�K�UI�Åy'~:���Q�q^�V6o�� R������f�_:�$��F���ӿ��Q�%��j��� q例��Jp��M�H�8��U�o�R��3�Cmq>|�\\�^�x�i''�����"�om���8��qU-�0��|
�r�	���B�F�UD�{<as@Y��</�� �J'H�-Np�7�/Ť8\f髡�n�s�Pi`}>2�s���]zO�ԗ��%6
�C7j�Cʕ�'@)�O���y�MYeϖ.����y�FVg&��e���}a�����f�-' �|��Ma.�"��7��%$�k�=L��"�~_���2}w�x^zZ�!!��*��)��&հ�w(EH�xK��l�ÈH�RO�Va!����>;��렉�������b$*d}T�}a�.'���Y�q�{c*�t�ע�R6������.�d��2���Z�sz�ʋIvǫ�˛k�*;��6¾�+?:�{?d�ڱ6%�,]PXy�>��
������������jdt�Y��IG�zS�h�7���=j)]��/��}w�R�J?U媝���S�L>�������ih�w�0sR�N{SCCUV{�:����JP%~\)/c�����|�䓉*X	�%xELg�Q�.0uQP��<���ٽSaʹQ_�5b�Ω��sw�9v�B�
ǎS�:��I;�$��֑!	u*֓����;O�����q��B�(B��K�_�<
=�r+f�*"�26i�X�M�ľ��`��3\q�՜�2���)��x�:ǟ�6�X�:���"�52��!��;H̽�K4���� ,̓��>{\A�D�g�$� �<���"��lh[qc�.'N.[�*�aa�w9�����\��6�����[~�v>��P|��c/ +,W��i�3���(2��&�:���]^���X�����u#X�>q,�����	�ڽ����4�r>�-J�u�A�]BpKR�-0�s�-{B�֤���Ϳ�s �������Å�;w����1���49�8�x:W��ɡ�/0M��:�L��)��z;O��"�r�8
wƙ�r�"["�6/����q�g^��n��}O��P�����.ƪ��Mc��.z���T�	�,��3�[����V�,D���_q3y�~:�}���ڛ�X.�x��C�3'�;S��ڲ�};YP	�ƉB�lJ���� �p~�U0�ڬ!q]�1%� �:��I��vB�ؓ�"���	�#��Pu�t�*\=mg>�H��(Ӕ �:������Z�7ZE�?�&��I��X[�n������G�	Q~��D��}$�%�漯��f��$�ήO?��ć[����fΈ�L�m����fm�����;C��.��*�9�:��`\��G���Ӑ�Zy�ƴtJK�Sz<`B3rwX�8�p�R�m$�����KM+�%�%	�.Y' tu�늶���!��/#����K������G_|˴od8�����T^:�C%wq�Wke\�o��o�=�,0d�Yk�B�Uб��	�i��˗=D�Z[V�W����֧LY��;7#tSH�����6抱k*~�F���g,�#[_�t�&��y����	����P/�*��Z��6>���}ih��B�(�L`�9U��1Z'��8��$�t0�ϼq�Uϊ�v�6���=���n(�7R�����x�#�͏mk�/G�[��.Bu��x���۹6��`���y���PZO���K!۬Rnc�(��y�y�H:��͠a�-y|	ɤz�Y���rm���s���^�n��!��]������)��U�ހ�p�s����+�h���{�W�V\����l�v���l�r_����^��?����͛wGn�G�\�0F�f�q�W�>K���
��"�%I��}^4�p�z���"��_ܻx�ɥ�b�YaE�1��T0S�a�V?�k���M�b�$凒?�ᾄ���g{{"L��s�!������9���^�g>���"Q��n��$�EFh�hB��(�L�+���Ֆ�K&JX�DV]���DIk��缃��k� ���5���}��8W��,@�xT�[�c��fB��%A�w�{?��{ծZ�AU�?�����R�J辝�x�w��s�,�[v�h����&���bNf�)So�D|L �#+��eҵ:5(�"�������0��D��N�.B���T�l�#H?�h�Ă����L�|�tqG�@�&~b�N?o�F���P_�F4�KK+Y,�B���uo�=������[���ҍi+�i���w!0�Jkg��9ŋ/�I,�%�@T�
�K�[�����G��-��3�U�~��SoG�7k�Gu������g����{`�
窠1'G�*	�=���b�lsg8���F��*;�#n����nd�
:�͠m�h�|D�����P��#�r�2��_��yK�j)QJ����n<��vJ7��̲	�7q�~�@����@�������WO���f�m������{m��2�ݩ��"�. Ioc;�L�I��fR_o]��@��$�'=DLs�Ʊ���DD3:���i�&�)9	V�E9��)���m���"o��׸�w�;u\���(����]7*u��.��b���sڷ��Pq�ҋ��hm��x��`��A���R{����n=\T�64ƿf�^����`�9*��2����w]�s�+W>H-[T/����q�Q�"��R�u�סWɧ����LnMFl7�bU`�$I;��Q[zc9����gYA���%�A��!��zb�G���B�TD�ILP��zZ��eFC݊����I�xɢ��
�H��n��[�U�!m�]��D%���Cb������ЏK�K�^��s'2��AܵY���<�����LtԠ]��X���{�����/.Ӷ���DP;pi��F��N!c$�I��X�3��N; �w��1l>}���doGv?ld�m��Xr�a�
E��.�'ߋ�s�k����8r��8=�oW|�5-P��H�k��h(���T/ma3�0"��y<����D�?�n{':�}nkK�7�eOK���y~�GA�L=�VZ�(�����}>[�
��-Ls�t^'�S�@���{@���kE���*������C"p����&sb:����!��(����O]�υM���^'�S�w-2����nrh���E^D!-�G�J8�� ��b)�Q��ؗV����F)���v#�D<�3���!TcHK1�ۑ]/@%�j���T#nf���锼��T�N��a��2[��C��S0���ܿ
1F��52��gO��5��d3a_�}/�PT3DN�F�X!�j��'Hk�93��ru�\秮�B�F�-[�a��)����o�q��,s���p$0��M����gv5������YQ9�i��ҨUI���&���mb�e����Uu��p�B�=�_2L��&v��4�w��mI2��PsJ7�uɕ�O��RIƛ�=L�^Ld�M�?��q6Icݍ���Q�FW�q
��}�@L;8M�f�N�f6L��3N\�ΐ3�g1&���P�[��q��
�p<� (�D�iǦ6;�	�A�Vl_}�]�� ������1u����6&�1^��
��'��ʓ��AlhH�S�=�fm�P��=�I�k���0���W��`�
aI\�5j&�b��'w��l��<�X6dg��qQ��I巏c��p��^2�7_{Q��)"���/���[{�m��C5�Z������C��W�A�������W<]G�w�I��.f������%�^ǌ.�ۓ*d�ĳ�K�԰�3gtдȣ6�
yy�cUM�����EE�DDb9ɉaK�"+I��;�:y�ƴ��r�m�)�d����c�S����]Ϋ���;L3V��6 �U��GH�A�"D���e�/û���=b�Dfiw���p�-{}H`"+.�-ǐ��+�[8F����sE�1��dndˬ[r}u�bF�Ȋ��ȞqF��OU!Yae�s��������/��oP�T&ľ���\����^��θfK��筣�>��[c���G=I�!g�g�)�6b!q´]1�L<��!);,l�_ �`�N�����K{�T���
��:� 0|T[��jeh�d�H�/�yԚӂv�̂��ċ�lJ��r3��5Q��<�W1��^.K�Jg��������O(�`��[��u�j7ӵ'!��)c4�G�����D>��4�>ơ��@;��u�"�����wse���P��FԔ�����e���<��ek����YX��u)�b�
h�M~�7 3d��$�=d��I��a��05�K�up��"̕�r7o4օ�8|����&��,Al~o�r�CB����P������8H��qw���u��������g{���·�1g=��ɫř��C�.8o�?�~ gi#��`���@7=3�,~�'vۋ�����ɦG�
�׍��9��"$ݹD������.�����TKK�k ���{��yZ��oM��k�s�L�^�ώLM�}ɱ���M��҅�������,�a�|o#3�r��O�n���2	g��z~x5X4���j@l�^�^69��_E�1hg��/�:w͘w<;�O��H#�ã�z��q�F)M���*lq�,sG"J�!�R�o�s�	M�l�J�:Y'�F*Ȓ�O��NtĈ<&D��r�ɴ27r�(+J'+�p�El���4,85i������&�!�qk6����V�$�nC�	Yg�Nu5��.�ͬaf03L�'A1��H~��F�2�}h*��lG�]��3k�l�$D��By�M�~�1|��LD�UT��r�2p�5����r�mՅ�
w@�`Bp�1���%7?�+�y�����4sG�����]�pTK-q�}��a��J���I��AJ���< .`B9��^��sqz�=#�6�&6����h�R�5�%���&�1O���V����*y����)^
N�e�X�M0�řE� P�G0S�
��8�]�VǦ���[=�?�ʭ�i�,�R�[Sy2���j��T����&\�����(<��V./��B���D�s�嵿����+�!W�v�\J�l�*# ;�xr�Z<=�X�Ļ���-C��¦7��eE��f��Ϙ�2�uOi{}������9�7���t��h]����n�d�W,�:�մ�
 ;�:\DJ&caZ�!�򢋰,u�`!/������Jc��w��%1�;|>z��k�0n���#�O��d�qH�Zu�o"TM�r�`|��o&v� »>I�<֘�y�
oʱ k���4����j=|_n~����^f�/"B�X��X��>�%��:�a�֗��i%�X�J�����3���c��^d��7K�EcT�A(]"���%��eh�+��!}"!�����1H+y�j����{�+r�ҋb�iȨ���P�y2�;�K�q� �Mru��l�&ҿ��za���j��s��{g�	�|\rs��{[>����??�s���tzi��~�#�%��< �ٍ�pmha��B�l,��+�<|:�>w���v�D��Vס8�Q��n�њ��t�؍�9-Ćb,䣏��?�����_J������sH��R?N�9S��h��^�#S:iI���oy�R"dz��!M�1h�R��`6����3�f�N�9�F�a��?W.�$�&��H�)�F�*�0���MB�K]��5;�w~�� ��7>���ƒ"�@??�j�n_��'����N/�S���&]��#M�x���|2�������7V-|�l�łȸQZ��j^�2���_4���֐��6�J���j�ԕ<���Q<{.:�D	tW�R:,�L��1{����g�1z�Ǩ�&O����B#�%7O��WLu4�+P�g*O<�7Pӄ�u)�q*��	�7�-?�4]&^SktZBq�BÑ��y��7�g�-7[M�����3�fޫ߬h��b�J� )�� ��#GU�8J���m�yk@>ۯ�ɉ�ܠ>tG�������h�K��K���u���hy*~v�x��ȟ�tEݷ�*�"�!�xB^����&�q��p�~xE�do#P�F×�1�����:Ċ3�g�t�/�}j��d���ƎiWe)���<g;�h&�#^��\��ߟɅ�$�?��o������\]�{2au��6] ¹���R�V�c��ϗ���RtXZ26���_�Q��k�����<6�^��1���_}���@��un��u��i6�w�z�L�;��d?�Ǩ�o�ϐ ɶ�'*v���#�/��ؘxl��"�@�(T�,j�&D4�4R�Arj��g7��J�^S�0��.�ȣ�5�^�X�>�Bൕ�>"A��90eߢp��Ͻ���쥈��N�W�r�O/�#a��ʢK}4����%���Md^+�{�a��u=�P�ͅ��x�`e����l���\Mc^��oǮ�n!z6��Go~�K�$^ψ
��&L�P�K#(w�YS(��z�*,ը��	X��.�u������SЄ��~�b�1�Y�Fjr�A��+�A���~d38���#;);�k����ʕ�X8�>��t�60}Ta�BY=�O�ٯ	��HXf=�ک��2x�hBKeEg�Ygf��부�^̩�Ѷ�e��1� wE�$�_T����`�Z�^Sͭ0%�+�}A,��țñ8��U*3ҐKs��������P�J��3�4��)�y:��M{6�*��b�9u��lcձo&,�y��rd$Y["��T�A#�J�po���}�zkݴ��Ĳ�޻(I,����Z��f�귱��>uE���8�4��\�>�Wl� �{��V���tt���!mW�)(.������\��tb[h@��u�[V�^��Ŭ+��Yp��ą-�V�x6xkb}��X�Vbc�E�Gl�۷5f�<�"���{�#��im_�hѤzvE֋13G%�'��[�AV�!t�����R��G�`�z��GZ���!g�XY�Ѥ�p��}v�C�?ͧ����oM�����5����"�*�
�}����k��f�4�u���9��)�#����b���6��ݼ&�cN��$�	(�]O�3E����o�$P�߇�H�Ԝt02���oY��ja �I�t�z_yi���o8�H=�Ww�
���@�q��qiu��iA��d:Okx���)]��1���A<�Λj���F".kꑞO����ŉ�)�?��W�~h��OP��l�?�»����[���}j.�A��%)N�I�Q��6����ӎ��ʩ\�\��m����Z�)��ݑ�p���_�n��<o��E�D*�f�u��ǁEo#�I/ ��d�k�ݡ"��l5�WY�{2n��h=������[�4?��:��%O���p!��9߲$�� u���c�zU�pQF�Q@�N���������������H>�P�G�׏6F�b�꫉V�җ���o���}=@u��s��޺���%��Y��%.�}N��Rk{������>�#h ڿb}c�"���>��<P�2햰�74��=��T:�ҡ���*0�+E<���Xz���
=f����/.
7[�10p�}�KIY��%�P���Wp.=Ӫ3�n:9F�� L7*�KWv�(=��[m�o���W������H��_���9����l�/�'��u8���&�� ��a:7EO�s:.���� /���|;!(��]��6F`���S	�L�Ea@��n����-�`k{�;��FJl!#��#�Ö���خ��'����VP���-j�}icrA��@o�&��7��pӒ�e6��M��CG����{g���w "�
�vk64f�Kl�{��\:*J���O���J��U-̐Q8?����
:���Q���Ҝ\F���Ε�Ƙ
�B)�6VQ�A��Y��,Q#b	�Ŀ��َ��+�m�t�D>��]Kf����MOŴٛu��W�-d���J�T��R��P��)o��Iހ0:��5)3��K1 �0��w�ã!�9��.&Pㄳy��?�F�_4Q9�"�tq&���سL|�K�!f��yZ1=`��A�z��� �4��1�J�%���5?����D�j.?t�a�U�u��⠁���|׫�zG�-Qu���)��BV���l�m��� r�0[P&Z5�v��z(���A����R��A��?�h3�s:�+A@�������J��U"C�S>�4��dh���y�=&�zBB%����N����.�����;���݅�C5f����\	kTm(�ۥ��g	v؝f`L��+Ώ+B���7����~4����x�ڨ�z���jOM�8�	���>��$�CQI�w���o?#�y�Q+4?,���]�k��t��7j���R28���\�<������O�ZXz%�=7F�(�?A��׾�ƪ�]�Z{*��ȫ�ы�����a���?za]�FZ��FBԂ~5"�ѩB�?Q�"�K�-ZheD���մ�#YJ�D���]_/�����!Y1)���
#�T��nҳ��o*8÷�������Z�с�s�t�	>Ф��%��a�[�͠�K�����?��i�$�`�u?L6'�>Fa#3�aP�	ă�B(�a�Ǝ7`���PE��P���"�z��4��}������S�b �XԴM�!0����V<��<R�fv����r����a0��_8ޯjy��F��˙�v���ա�u"�ć@�����xL�{�讹��>yiZ�������ii�Se�?��>��o�ܭy3�5�*!Z�瘏h�M�Q����hw��Sr���"�TA{����U3��|Z� �z���I�?a3�9��d|�P	f)�`� _���NwYb� �Uւ��W�K��U2�IE�6�鳂���ȱJ�!� V�S�Gp��8��N�0~7�e����Y�h�OK�^L]��2 7�Ӕ��2BD��op��m���R����W�*=)���6��<W�@�k���{�$q=CϤ6�!^u�G����=W���a���B-2D�6ꁛq
���&7���V������Z�e��>�ǞVN�ᐃ��R�FD{r�@�3���6'�F"��62�B.�0R���gdVW*����5\�����{{{bI�YH)�����Ǜ�s�l8�B�	�D��"U��RJ*���]Q?�el#���-�v�"ˠ����P4)]��Jڞ�[�6��9��>���xm�,~1����!�ɨ�TNGN�O�Q6��wp��v�\��� �;O�.+�d�!4�%��6�P^�)�F(������lc6�U�|6��mGϷC�:�&)J�����|mVX�� ~��(ģdm��~w��C���8�d`��[��"b1��1\x�@��*Wl�x�]{�義׸���c�H���O��!�p�]��)[oule�� +�l�0�,!A4,���j+���_� ̦Pa����Q��Y4�"{���絾�����GwB;9|?��bB�R6�Ã����|� j���0�=��v�zz��� C'�!��7��h�.#iF�ݰ�i���Se����VP�XR�w
��ߖi�L,h�|X�L�ƫ��O���L�J��y�/V4��f�Yż�8�C���Pӳ��Q�\?��+[��k����G�ۜ���ׯ�n����0�%�Fe�!�0}L���nP�:�{��վ�.��CU�u&%�Я����$��q=�0��xQå��XҊЏ���飀	�ؙ���+s��m�s#-�D�������|�"=����*뽿s:`�9���$�GF�,�љf{D��̿�� .��W�|Y��>�a��e�Z�<�e����&�'�O�V���RԗG6�D��S��5��ӵ�����(R}�����w�̤�	A[\�mۑwOsE<_*xt���~�����UK¶L�tz^����IGU�Lb���T��t�y�m�`^?{�k���d�,|[�B�����1`�/ F��DV�{Je�mۗW��ZM�R1�-yx�v�a2��]����u-n�L!꽇���Z�%��:�5ǔ�O�5*��ޒG@�1D���1L�ͥ~u�=�xU���yD�XM�Y��M,�N�|���]��-d�j41��e�L�H1���ۜ�?�+uEN<et�	(0��G��kK֒	=凵 ΡH��P)��x(�.̑������sIC]Ͱ�T��ό��U]p�\�E9�_��k�fx�@E<�ӯ8��[΅�·�W�5�:{¾ߦ�DZ[���̦�8qn�ZL��N�0N~ﳍ$y$�Cʮ�m�N���BHo;����z�Qs�r�z��N����t�#;���,S5��'`/h�Z^�ҹ�=1�y�V�ӊ���2�j��I�l��0��ft1�L��5{���Y*6r�Wd�%/��+�}����z;^F5��XPL����-�%|	ļ����Dw�ʋ��k)t���i~���R�2eq�`�$��BBB�̔h��b$�z�T�CP�C|�a�x��ވl�j��Xo����ɱ��T�nJ�F ��4�:,�3Kf�� 6ҁ|�9�:X�LJ=g�*9�H]U��&I+����=���:M�u&m�۴���ʢ��c���,� ������Goi�4�I��u�ywg���-����m[*>�*�ݛ�!�-z�eq�Y[�Jb�$��K���E����i�Z��p8eӋ=�)jt:�#��˄<M����:#\��=7��I�d�]9+7�$�#P��nW�����bP],�8�-�	QK�˩f�xd"sc�����_��y���b������� �����q��w.��Ίn�*55�A@?Ñ��2%��#1W^�%8;�-�_�\��K�bA�$�?���s�`>@�bb1M#�(��H�z��b�l��G�k������� �-��Q;N���K�ٓ�~j��J<���8Y�V���]��ޮ��6�l��X���݄�,�%;c.�A؍���	3��`�
�H��=fg��b*���8 ܰ�Q�]K-R"
�޺��4�oR�}S�l�[N}�iu��S�"m�1o�n��-�����ڀ�����i���w��&��=v%���n�4|I�l��BNx6��aaP:�.ƥ�E��ƻ؛U^���?���4��6�yTJJz*���r�G�CC���p^)��۰���2�Tŝ��F�A���W��`	�ٟ��a/cxC�%�xB��\#�������LN��D���^\�m#���8�K:�G��9�J%*-�0N�/�4�^�Gk�9���-KA>��$������>K��a�q?D9����PE|n+�����u!�v3ZE�e�a�۔��1��J��6з!�UOM'�X�����4�e"���.ޕ7U2����3�S�R��w�~�,sx������=��~X��0���|��.�Y���S����sA��m�i<ŉ�,M�x���9� �E�)��F�_�S�k��}�&`�xb�슓�'�(�����J�y�1�}���F�Q�c+�_��а>�&��e��e�^v
����k{��	��J�k�B�떦Dڥ��;����M�a�Y?��M�ql:�����i%ix��|�
��@��d��}s�5��T�HV�5�Sf��:p�ȃ.����&�d�K�:!I�/:�@h迸O��O$��E�ը�.,�,T����W'�I<�ಟM�aS/�N���$�ӂ7���?���b���U���0�!��2��C�Mܲo�w-Eܐ�i������.�v|�t"4֡U���m�aP^s����a�������$�cƕ\Y�����A���������S5W���K&U��L���e\�9�H:^��`�����A3�¤4��D�z$/���כ��vM�Q0����K��5��]�o�(��/4�庌�K�C�!@Xa�:��5=
�h�gf�6a��7�&۟d(_�P��.���i����jh��&mw�0'nh#�ޡ�4�������h�,o=	����	)$&<���C�H�fդU�&����wzX�Q��o'�W�< D�p�W�Ȳ	C��L����
m�pw7�C2��fҲ��N�p{���"�J��9.t�W}��D��(�L�kr��S��}�+rs
��/�K�U�*1�K �Z3Y�H֮2b��^�n���nNb
�Ɯ��j����PB�8N3fz�����4����~��ѧ�I���w�ӥ���2T!e��㉺TC�[��ޛR�����O�BsOһ4||_'��t#(UZ�H�u��:y.y��揞U�e7�l���ޚ:W�m���'�*u�w)c�u2�AS��Sx;��"�]'�bB�o7�Lюvj�H��c�Z��/"E�����k%�Okf�;� YNW��%�o����n(��D�r��t�z��C��C�g*��Pd!l?���?;�F��n>�}^*n��PM)켎ZBɩ��O5���8򭉞�� (���fݙ��%�HHX�du.��0��xP�M!=�b�<�I�oln
��}k��������D��\�u�0aJ�Zڸ7<��
>�'!}?'5�)�rS{]p�X��p.�C�jE���ҹ�����,m�'���
+ء���H��@Y�oȌ� �x�&�'�X_�%��Aӗ�Y�T�m�/�;��Á�"�(*�FW�4g���>%�R9c��|���']a��q�#_96go�g�wˠ�^�����eґ$�mG^� �ۛffd�Uh���&�ϝҦ��K��[74GSb�_�]����R�>��%�7�IkvAʴi"G�b1�:�$�d�#n���ǭN�8�������ԶTV�C��Ֆp���J�V`�ʃ��D���N��q;��7�P쩨���H�}���b;�1=$������Gk�e6yqVn�p-pAA�k�����-��{c�ô��e^/Ny
C�+�?�t�rɮ�9#�*iU�b�b��N��*g}��ڞ���j�gz�ފ̏����5��n�Wa��I�)@k�T7�T:�U/�=hSk�"�&H�i�tC�U������`S��U@���Ę�!XC똉S*�q��T]�Z�96&�������yO��䉊���-BL��Y֖��>Oz ����U~��l�Ҙ¼�5�d�萌iG��q��X���#�=�LՋ>n���נG_���s�)���W!��\�A�h�j��'��O�d�¥u���1f�P����.��H?�<-obi'+�����2h��&%[.e���;�c��(9ndt$ׇ/>�MjB�x$��z[/��]�rL���߼>�n��b�yӱq
�q��i�@[r�aF����ݮ�V%�^�V2$|�4����N�|A�8b���(����w�k��3��2][�&ΊB|����3���F֏F;k��� �P�<R�zR���S��HhMM7��Hh��8^T��	���w0	��U����w<"��1<�*��&�57눺;|�l��m8���;¿'"N���)��y����� �v��"��|7s�Su�(�7�ʉ��q�����$W�ʜ��9���&��8e��W�X�O���d*#	�7\�|;�Z�Iو��J�A�����/�}nw\'3?��!��I�>�$	�	����wX�h�Y�H1ڽ/\��ݤ������$�e��2V�U�dG����<w����ح��UУO=!��YY3߈�7O��t�Cn��h�ҏcXU�KuqP����g�y?#aD2]�ZB����(`��Up՞�;N���N�ߓQ�W���F�C���z�9�>Z�v�,��I?��8�`37jWGW���R�^e$�!�C�{徳a�!�LV�Ni�X���'d���"n�ճ���	`��F}ҁ.�>���`Ze��gr[��Pc@6���ሓ+����K�9�~�T&�Qq��n�]⩸8�+������x�L_cV�U^K���l��"ߔ?�������+s��1����^�L[�ˋX�e��k���w�9�N���	��P� *�{s��T���O�ZQ���p��<�*���&�.���0՞�)0@ޫW�ni@"<$Uf],e�߂Tw��~4���'
�R� 6�O9�Z�3��ޫ}/�[�����1�wT�)L�!��}y��CH�A�Qrۄՙ;���z���F�B<5�H'(Q:tT#[�aa.����s�����}�ļ��.����o��B��3�֊��/XpE�j���-�~|�qM^L�S�b0`ē�.�n�wR&���볰�19?�VY9T���D>������v���J0Ȣ�闫$����͗�,QPk����Y� ���<�\�O�<�N})�Y�	FR�s����e�2�UR`��x��!ΰސZ�ܡy�c���#���u�!R�s��v����y^��"F�)"�:>�В��|�Ա�H }��>��s4�^���޷R���g_ʦ�H{+-�: �%�OtO>�b�}d�Ȑ���9_,q��5��%�X�h�@ˑ��u�<�u�n%�������<�5SV2��\Q���/�H�qU�mz�%x�4$�(��j�N�x�ú�bm/Jf������ޯ��g;	I�9K(���q�0ۿ{r({�[f�@�xe.+߶�Ee_+X	��!=�n��ި�6�+�4U��V�.��vE�5����_3#��d*K){L�����@P�r��vY����X�k7̇�7����.uMv�V�Q3��ܢ�=C��5rծd���V�i�#��	�g
�dV�?�r��������%�����L������	9���o/쓳�-��X�ca�r��J�r�X,���<��|&�rz���D0⊥T]�+��&Ӛ�vHa����A��� �j��3g�wt'���s#=�=��ڗ�Cv�;k#0H�KNy���O���+��W*�7L;b������F�T
�j1L�htT�͹v�Z�5e�afB�ת?k����Tv'}[p�~w9�G1Yϕ�u��&;j���%����z��r�]�������;�?��kv��pL�Q���"�UN�5,n�F�Bd.�LuZ�&����_�
��.@ѿ�Ʒ�K�}����طw���\�=�o�����F��4"�EAw#�8=���Y�y��PUG�:j,ե���XG]p�ɛn��7_���_��8��P���
�QU��q�1�z���0I6�p�64"���op��$O��q�;��Sx���ȸ�x���p�7��{��#EÉ�W���8��%H��C�w+3��@�e��g��4���
�.^~h^x�����x��=�Ŗ�:~���}�e�X*A��=T� g��?�,��koz�<U�)\]��^��S�(r�|B��("2ʩo q��.�=^�ӆ�XP�@u��8���k�/_��m�k}�ndݖ^���w���K�A���Zԁf����D�p;����s�}��(Tj>�w~��CB\O�~�����m��k�D6ׯj�ZN�+:Op�s?��Nr^��r��_���勮���!pͦ^��қ�x�X0o.��z��V�o�6�c��<���g�+�8[��R��",�=7��ࠟ�rt_.�v}�a�P�)�)��:F�'��ӊ�"��8�dkߝ���4Qa`�fL�0��ok��S[�3%��E���n�q�Y�n3���*UIj��{~���<��Q���d|�!�Dc�=�o~�Ee.ӑ�S�\fi�/}��x͋���v2��:8M�(˜�y�0����X4��;����#*�yee��]ﳛ`��H�CJ���Uw��4R�Q/�<Ƥ��~�b������b)��A�he�W����np����aQ�d5�`5$\eH��L{d�vl�+�O��!n_���42�p��+p�!KKWtn#�� �p.,����Ԇ�}��N�Y�1~L�\������t|�gc��n:�����_���Y|s�3�f"q��N����х��x�?�~j����-X�=�>`)�� �ڰi�L%�VJ���4�U� ��9���P?0y�X�	�X�Ԧ��6x���~w�b�9�o���qH�-���x�?�*�[����l�(W�,It�hɢy�~z��k�>p��f�*a(!B|x0�n����_���>ƫV��)�;M��t��ID�.��kjNf)n����E'ϔo����>�ݝ� X�{�>��;OC{��;vs�V4�]ȩ���	�nU�sd�;ǹYI>��j�.��ۮ�w=����y����1-��4�H�g�V����Rh8�����q�a��m-w
�߀]���Ɠ�de>���w���ZA�ԑQ����Da��p���������}��R���wb��Q�0�:g�DP�����gv��{: )�`¤q�����F�_�?{"�=uD�F�шI��7��I��4{�qL�}�ët���ߋ���g�gy��>��w�����F��M��G�ځ^j�a{���2�ʱMB�[y���s��n����Xx��s�vӘ�C���Ҁ�YY�W�nٍ\�[�)�C4�-�WXԎ;f��K��g=��m"Ƈ"ć>U*K>��S^8{|�i��������Q���x�u��/d)���jx�ًNNu���
�4���\Tz�:ё��>r�{�r/}���ð�eh ��Ƈ�$�yw�,��5�Z��?vS��vKT���]�ܻR���Ʈ��W��@"���{�z�j`�v��p�id`ut�e����Ne��Ͻ��F{5�:R��U!C�q�AE!��}=����VW��+���s堬S�;�tǣh��c�h���[�­6�j���[E����b9�����K.�Cڊ�W�^�?>v�T�����Okҕk]�����Q�̎P~X�5!����q�%�w������ɣ0y�xp��z�����5�<qU�A��ԩ���8�}��v~�,\v����}�C���~ �7���6�74NҸ���cMx�1��̩��ö�m�rъ�֊�{̘��|�#��*m������P@���g�+N��ԣ��s�dR�:��ip�7\^�!ޟp�ȮC��K���4GX���w~�{#�(��q����7bt��C	�R g�r=�G�R��Fߝ"��r�t��O�<��������Gί[{	[�,��}.|h+��2���󽲋�*���G�%c�����$�{�Ф;Bh4;�3g�ǒ=�᚛W��{)�u���]�=s'�ѫ
���l�7`�
(��d�6D@��#C�m��٥�ỿ�eP�%���Y�4<j�fL@�D�����Nc�9�4�j�F�ڍ���'ᦻn}� ���g?�RtE5����MW/���q,�[�������1
�z���U��u�}�{�]�cܘ.L�9~DO�Lo�� �1�pI�-�+(�������\���A߃ˮ_�}��A[̓)8^����)�����Vs�K?�͉w8�5��yN�<y��Y߃+�>Mw�Ÿ0D�.B��c�g��8�sL"51�#e��11����B=m��9���?�f����H�F���.~����Ë�±����&�튌����B�Đ�)}W����CvG�'IX�G������OExL�{��ض}=���ۻ��u�b�8g#�o%`�G���~�(����vx�E����jh2���s�|��+�6A(�ƽ�ދ`�7��yT��3�Oר�Q_�S�a[����o��=�E�.�w��/���7܁��^��ә�r���R�B�xz	j�輁�Mou��ghL�0
�C���")ǅ<mm{hթV?�)E��/���ߊ��v�wd/�[�{���Ω
��'{;�o�����s�A�m�md��|ґ��*���O�k�����֛B���$�=�{�]�䎧���}�ӝ��$%�q'��:����?"�ޏN����A�ˡ	߷� �����}u��u(�n�v*���`2N�k&	=z(~�"7�I&BU��R�ix|M���[�0��9������-�7%Y���2�8\p�W����G���E[TAڤ�A��9��"�u��X�q;�X�w=�zbW~e���?�b�cqؾ{`�E���Qž{�+W]x�#1�e	��GZ�֊���x6��3�����W- H�hb�� ǎ4�+��!!���D��|�t(ȸ���Ku��[Y�ՖL'T�C�:��\�O}��!HP|��Sp��	��
L�LP[��!�4����/͑�qZ�k7�q�?�PډP½�7?���d�1E5��8�eHhL��XӋ�V8{=]P�����xu����~�C/ì)�9�b���b���RH5uT��PO�P�xr]��|ꧭɭ!�����.���4��v�*�whܤq5��V���ސ�$�e���ш7�}�4��Tn~����M�뿠�I}�mIzT����w������}$�������O�Jk��1��D���SIddR����A���O6��O�hD�|ܙ����q�1{C�w�"��4�C�#�#m�����R*�4H��S��΋@�&��Oo��O��׾}������^Y��|����#c����#��1O
E����{����пϓ�~Gg=d6G5$��)$�U	�?7$Vi��@��p��Ko@��e�27�Ou=�9�w�y�����>l���c�+SExp��G�Ô1P@�8��O�Y����-P�ik��������U��(X��|�=/��v�g��:�NYI�����B\���;JQ�Ȫm4�^�w���	n/���k0���p��k��J��&�َ�P��D}��y�����!�^��������S�"0	TQEn�*5��@��`�����b/vdΏ:6�xt�u�����y��U�m��}��fSI!!��[���&6�
����(v�w�V� �P�* �{o� u�����ϙ9a�黛�Μ~73s��{�=�}�y�{��9|�l&x�0��y����ö�޻o�oZ�'�mk2<O��PN�E�������O�Q�������8����x�#j/x���?h;dI���/F����������U�Xb�קK���m�Xo1�)���<��r������fKZ�&�W{p�O��k�Bfg=��Ǝj)
���֐:�?�#�R1��I*d�TRk*۹�F�<�o>|\�O��=���o��b���B�%�^����J>�ʾP��T���?}Έᄗ~���a��D��z~�8����4�%e(�JH�^�w9�*��}w�%Wqy[C;ö��_~\�B-�]Tb��|p9軾r��� ]es�W�ᯎ��*�����ǰ�>; q��4py�:��uRo��_b�=���;n�	���A��ȹs^�57?���1]�PpC��Q�"�]t�炭k����z�O,�ʂ��N)P�L!�W?�0\��0�,�Reo8x�Ãԛ�9��>�0`Xg�KMW�����^1$2$bhgn?փӿ���(i�5<��ǈG�_-E�["f-6u��"r���.$q,)�1ևJ��,Hp�#�����_���xi^��#�p��1W���t�8�K�O�/��S�!C���礦*y���Af��$��=@V��;(v�$���?Ė4�|ܒ3��-b4���.�ĸ��l�\6��P�z��Kn���E���-K�I9O� �㙔+%�mz��".tv ���ݱ�ޤ2�F��G�P���P��(�H�$�t�R熈� ��&��F2Y�ㅹ}����U����.��{v,*�$F1"v�u'�u��Yq����W<�����R���3�b����C
����G��0���g�[��pj9eL�L�pŌ��,���yg����ٙ��6\50��*v��Gġ��ŀkR����Hq��'���Ϝq�<����Ҷ�N�'O9�E/��c��
�V.Լ��
��)����_�bI��I�]X��ʙ��+n_�&����e�܏�c;0e�TQ)J�������"�RI�ޗ��>$r�Y,�K��R�Î�l��oz�iκ����T�Χ�A�^�#�j��<d�UQ�%���s-�0������[�#�������u�}�N��8S��"��ö#)F���dv�v+����`hG~��wI�{T�Z(y���~�ӻ�Әr���8�o7�� w��4���l����Q���#\�IX��{�C*��v#LYg<n��i��Ȫ/x����l��DL;q���)#�vެ3>������L�*:J\�?u��:tߝ���۟�ӸƸ��?L1#�#�]���c��{=�[V�VK�dZ���9��Z�T`�&���S/,�'d�qn�aI:|��ÐF!�:ƣ��k�&*�Y�*y3��c�;[e?�<�&H� 7��(N�ܯ��������������w�;����O�
��5���J��.O�*/+�	yN��y�b�Otq�;4]am�z�(F!p
p1~$�u�>����Õ��ǿ����֪��:�b)Ár�|_�#���R���s�1�c1m�hcd�1���� ���`���J*~GǙ�(NY^�B���ōo�R6�|��R&F)�Mw�,��#�"���^�Hq}��fn;mĖ�r���%x������ܩ�3�4����YpľZH{��r��=�3����u�4M�l��)��9lt�.[������/�^L�_�^�q�0TxE_�à+bd��v�xy^��}���""��<���q[c<��'�V扱�Z�p.�X"F��*ݻ1�rGo_?����o�P��چ�u����7���g��G�N=���(���XV������aY�{;p�8x���3�4{�0~ �u�*w^���8�(����Zq���G���[oy��^��-��Fd�`qjNF��2f
�\��m���9!��y��7��g�<lW�	=�,#�k"/X�H򅫄(fy���&W��P�K-;{���I<>�E)#,iW�A��=�Ql�I�#���z�F�x��7��9=U��631qG��A�J�WD�ܡ��-�
V���v��;�ݴ=�����07�t˃��=��X�m+�kRys��0l��k"Q�s�Q�q�/�ڃ���a!$�'�֟օ�/�k��=�D��{�CXv�4�F!�E��C%��9/�ݧ����3�:0�,�u�?񇋮C��)���t>*���u�`�bX�!�Ȱb<�E��<$չx�;���|aC�b�w���PB y��\ZՓZ��,���p�����.o|���~8����	:%��#�\���%0l)
��h\�;�`ch�!�L�p�*h!;�Ø��l�5Jy�p4�yő�c����*%\[�ҥW�W�LjG��TG.�h��G��RV|�?\���夑k��~O����FZ$"��	j��x�_S�1���E�[�~�q�ē��nr*��(�%ð´���>���9i?��f���܁��s����8Ͱ�$#��� ���Ĩf@1�.�Io/J��P��c��e.E4rˁ�y�������H�1�����N���W��4�#FG�ZR�q��\�epb�>��?_~~tޕ��1HE/QK���!���~���h��^�NI��<|��#F��dX���rA�u���s:+�_�x��"2`��>���<�諘3�u���j?x�	T�q-�ZR�-�s�]d��Zv����1�)Jl�m���Ei!�ꣾ�m���V���t���\�
w��XK�p͍w=�y��X��káM!7����$�
<���SF��9�)_�=������,u�:�z����H��GF������=IX�D��n�ZY
�#��+��{���Z����1U��o8Ķ�I������Ν�8�HwH�Q��f��c�+E�˫�ᠷB�K~��e����U�TR|�����-���~�/}�bL�"��6x}D�ђ]il-I�4�B��rFO!�;q�i?1)v�M��s/���T��9C�Z�^]��K�<�-y�X��7\�Y�-ǆ�'�|M�`{������4S#~�Y"��_���>P�Rs���I:���G8*���WufJ%�D6Z�:��>l�Ն�K��Bՙ�����u�]�:�p�-��}�K�[�|\�&z�T�U
�h�zy�B�G�^d\7��Ȇwr��?Ƽ��L��e�d�P�͘�EO�K���0�����_���N:n�#e�$��|�a�QqÛQ�O��s�Y���:麎c{mHE|���蚎�õLi@ƹ�""I�ѣG��TV��J����9�jx�g~�zۙ�gn��6�%�Z�e������1�j����z�hT�[��c?�C5>R����'�ǋ��.�gx1":��j��Z��M�]�t����^i�R�ަRmQ;`G�mm���ļ���<lW*�Z-B1(�ed,�_sw�[�˥�݇�J�TShQ|��.���}}��m8poy����Б���n�h���)n�����9�/7�a��Ă�5<\�Cr���T�M*m�/B}�ݶi|kd�v�O�}qEݳ������W�ݱ!������!#qb)x��i[���u�C֛Ե��6.��c3_����Ϟx��D�%�~��M��?,��?j�ZÀ(��8S�\�*t;���`�¹(�<�E��� �?�Ƕ�?�����$��O#��QC�C�TB���dP���8��K��<��/��6<��˪s��,\8�ʣQ,t�9~���v*qV�#���Pjh%(��r�r��,)y���U+(����V#�7��Ј��J,��^n�rfJ`�M�+E�۬������16���iSǩr�JICt�yDf>��'ۢUe���O� :����y�H�xp[y^)w2I�}v���-�{>z.z�*b�˅"���${Y2GW��P�X���*�0��v0�[_8�c�{'�L�L�8<�e���Ͼ�ȢS���¢cgV.b1I�+k6hl���[E�؁Z%D����9G��U�g�zx�'~�VXx���VXo������r?�ջ��r�+��$�F���x�|k��Q>�/��Wu/�#�/��H�=)�Q���*�8V��ް�N�bm1F�����vȈ ��c��$GWg�-X �����~��m!,�cO�P�����i��Ҡy����]�4�,�kH�������;it~�w�����ٍo�:6�����$��R�EזF%�Ԫ,L��ga�ѣ
�3�U`�p�G~���OlE�Cvz�$�Gc�P�#͖h׷b��`%����w�E}K��*������}g�Ŵ�ן:z�8�vf�e�ל�7b��ni�y��G��P��2ĸNDY���UƢJ�w��iH�Ŵ^6t�=d�-��#�SD7�3��C��ۜ*�:��+��_�p΅��sF2�F��7�E����7�\�i8�����\Q�+i"���G�����]BG���<�:C��@j�
J���n��uN�Ô�Q�P�ШC9�I�N劜ۈ�P���m�׉�6>�=&���gg�u�"Do��=F�iC<��K�|Ɩ1���;���"�m�T�!iZEw����2�����CZSAo��<CK��/�|Y��v�7\�{ϙ�M�[�%͆F�?ƌ����Io�/�©tE���Dj1}]ӥ��zc&Ū�5��!E��E۹�Ki�^B5vq��~Q�sۙ-6���pl��(-�c�F7�ƪ�!+C,�l��>���I�g^����<��^�ϼ_�8ׁ��M��mi�|T�I�c�m72�k���n�b�9RH��d�<F���F�!���9=j_;��k(e�P�SXթ)���k{j��u���Z��&H�_�a>�hk���ys��Ѷ ��w>�l7ǵP*w�Z�A*�V�<�:� tLw�yK��>z.���QnfZɡ���e�*@��{Oym�'N9r�1%{9�T�kS
�t��{_|�!E�f`��\��9�GŨ�Y��("����f�a`d�HmIyKҳ*BJ�B$���>|fCH.r��3��A�h�"8���q���Q�m[V�X�吏}��R�?_/b�/H�[I��$Q�:�3bv��}�7���v�.�2����uFI>A��JX���KĶᨸ�H�}P,�g�m|�M��=畹jJ����M��JM�44�S��E u%c�0��4�v�yA��EFx����h�&V*"����T�s��4W�u�
�(����,/��y�������{CW��#v�䫸!q��໖����C䔙��yCk#ć��ް�u��[��]FN�O*e�=ᣪ06ln��Q�2�eV�5,�D`�H-P��-�Q`��$D���+�.�Z.�G�:��%�mиbl0u��OqH�9�SC\�(��mɫ���.��g^���V�&���t5�4���A�ƒ�Rx��*!-�R.3K���æ�6���l��""��$뇛QT��z\K��F&�HO=_m|�M���ĳ���;�f5i�$5D�q�
#@+�t�,����&4�dhu��>�d����g$p�**a�q՗Z���ymV^�Gg�"�]�HŘȼ��G�Tl�W,ODy�aƴ��7Z�V�|�\�sց� u�%�,{ņ�Ħȃ���'u�a`��Z��*���""i������Q{�#���r�ٌ_K!><�Y����Gwԁ�x�;���\J
B5�GGGI�q��9�؆�s�_�TA>g�Ub�"���Ǚ?�s�7�m`�<⠙p84���2���D��;4|�K��{�������}P�K�6HV����E|�	
^A�����jSHRZ��Qj����G�4z�����>T��j�����Fz��Rs��^�e�����\E�Q���dqrcm��}U^x��u	_9�@|=����*�����_�����/�����(�ed�"iW���Y?�0�z��z�>�6X������c,����ÃNi����g�vLZ}y�<I��(�9p���{f#�b�lK6��@$�F����S�d�E��7��.Q\W�v�e1��$�X��>eJ$-}��W9p�hA���p�/���֊0���~XA�փ�{2��s~l��W2`��$IP*���M�[�m�CI��)ZϤِ��X�o'x���bK���̠vL�1��o���ϼ���i]�i.��ۯ�Z��Ϊ���;��>lc��n���߻�����&$���
�9��iXan)�0�����io}�h��䳩��F��}�|��G�zP��ێ.���8����ܑ
)�G�5�>GQ$b�)��G�4v��'�X.��ˈ�n��I����2hXIL�P����C��vj*���::��^�PD�ީ�h�r΅7�� oR1&�z ".�C#�K8���T^{��.�o\��aDS*���G{	�f�����X_s�����4 �Z��|p+w��gC��|�H}���A��r㔱v#I^_G�4���N�r�=V��q�-� b��"ì�+��ԧN�q�ah��$���.�[�x���/�(�f)�5��k��w�l�n���Ac;���eS�dy$"絆˰�� `@1�T� t\1d��}�%U8%�<1g�{�r�6�������/�g}MX�k�Z�ei�$��rI۟��ϖO���(KJxs�U���i,�*�}&�Ma@R��F:NCd6�	-45�s[>j����*
uC{М��/���گ��zci��}����:�˃w��s�l���jR�V�8k?�5��{v�����!3�����([{d�a�i�.��`珼��z66���f3b7G1�)r���a`p�N6pt�uP��Z12�Q�+�~�|���޼�vj��Q��Zp,&�W9O���q�"�<{�C�5:�Ry�E7I:�;�W�Yr4��gҲ!e�"�GwgMS%#�Z5R�X�l0=�g3Dt���bY� L7n�j��~�3�#^/�y�K����l7liGy�:Mө���q�Q���/�u	�y�C-��KÙ��١��5k��.�Ѧ��x؛$�w��fN��񵈘u;�x���m�$��r��J9�����D`�s�bÀ�E8����^E"m���x�����W�bD�r�1u4���$�!�Bձ!f�q1�(:�|?�vC{�c������Ҁk�3�#��l�F����r���}vݴ�=�H����)(�u����x�����$������	���5�Zz
�|�U5���S�->�7U�2�am3���TQ�!o���>IiS{{��-���'����@ZU�G��5�CK�Y���Nұ%g懎���bܰ�0B|��j�������4�J�n�v�(QC/�E}=5 ��������<^i�1�����N̛ۇ�|��Y�e��	������\��#��u�3ye@�~���'��3Mx^�F~�m��mL�P�狁i�k!�߆˘F2�z���\��1k�!�ڀ�� h?!�\I��V�0����J��F������uT鼠�_m���X^ʥ�*/�>����]vjYX(uN;r��砧';��DĸahadL*z8�=�]���̝����2.�k#������'�iw���cZ�V_�� )!NĸSKi��5:Q�����O�f�ˊ��g��g���5�3,���p��T�@�!�+�Dd� <b4pPΛ��77���x�?�F��`D�YŵO}F�ϸ��l��n?4yl��ԜW�sf�$��Q��������#�@�1R����2i| sM�z��Q��p�D��UG��O����C���+��]p��D'( �j�l�� �\�B;0�̲�^�e��>�D���8�( �=�R�g���N�Pyvμ�7��NJ[��_���^I��ޡ�jb'ӆ���R�@jṵ��Y(%�G,�TtP�L;��rD��a�$1>�!��aƞ���xx�M�����݆�"�
Ȣe1�I���yW���z�V0iy�l��DTh_��^3��y�c"0V��e-z��̳s����,�N����R_v��s�t�����d5z�z�z0=8Ң�s���>?W�7�>O=�<�W�`~�#�z�Nm�=S�pЭ���qc�փ|:��!�:�rvL����I���W���m��_X�_�w9��W��`�.�,@*�<aG�-y�5f���Z��s5p�$YgGGa��}�Arx�lf��cr�g�N�L���]�ܿ���B��a(�m�viR�88�/7�ƻf�l2cB���	k�Y�mA��ot�z任ʍw���/�Wr�Sr�\W��2�S^,w��Mb��)�>��S�Fu��?�������]]Ć΃}����kW�|f�<v^c��K��;h�I%��a��4��L�ХV�P���Y�I����z
�y�{��v$���ƻ���.�i������F{�<9'�$lZ�ްZГ���Bgp|O@2v��w�k�� ���ft�b����=K�t���L���	��X+rm��k���%\q����G+b�i+'��&#�]x�ig�lyt����EUd���Q>ƛ�c�N�4���BDW��U�9s�X-�o��w�~�8Q#|��j�Si��QX(&���5�ۅW�.�˖�!��>Z{Jpc�V*�*(��h����ڀ�fn��E}(uWj�9���O�*�%��\6/�pQ����ݙ��\~�}(u��z�&y�TL	F��,i���CE�0VC �+�;M�\��Q��ǽy���)�fFŇ#��L�-O}�>��l&5��XKy6�;�����G_��Ͽ��װ"�5'�[��\�~�h01����ܺ�a�2waK�T�C��r�OD�|�h0���Gѷ��f��7hF�>�n.B�1��y�b7���x�=��`y���¢�xy^���b/��x7@D;qv�v�khax�3��CP(��w!����M�%�e�^R91������ԥ��?ތy���x�H-k����\ջ���r��JH5����P,����1��>�����Ӷ��2C��k�ɛ�?v��w�nw'KI�۹�!��0���bQo_��_��<<ʥ/��v��U����s #�T���U$b8�'��%b-�uۄ�	�sml��$�7Z��6�M_<�IA^_Mᵥ��<S���W{7�Z��1c+�|��a$���
�X�2d�R�Rl��m�o��Ö���]�'���b0;�>wJo�H��?��s��h������:����`�,���tVە�L�v(���i��}��gKW|�A���bƘ=�T)�����5CA̵mO=��=����`�'���	�o:���޸��>���'êఛt%Pk��rύy~˥;)Z>�+��S=�,��h.�>v���G"��J.�|"6�2^��v���n7�usj]�S%�(Ƶ��M�#����ݣ����[n{@��k#��v��'��-7��Cm{��łܳ��	�	K��b�Xv�<�z���\q��F�7�����z�}�K�R�T�6���Î 8�s���\��M�q����g��w�����<�!���5Ô����3&u�,���\�$�"�Ւ8����g]ܼ|�a�㕜�ݦbs�� cR�7��>%�8�mq����ut�VBC�ˊp�~\���9|��Ŋ�;>G���z^8G�)��>�6�?�?\���m���ې��d�����q�n8�2Ճ�1�j��]o�K��v#=k�mԽ�9�%�������rP5*>�\��a1����?�<de5�.1+��Q��'RF�߶JO�ϥ(��Jv��Zy�i�=�}v��S�ɆA��M����9sQT�d{9"��v
�c�8ɜ�P�:�N�A"���_��?�J���S��ӗ�tĤ�]a�͑0�Թ���J��(2K9V���bl��`A�<k'A�v!��O�tG�Y�-Z�k��;���u��n��,�����I���)>\��Σ� g$^��U���z07C����"0��d��1�i,yD�K�{v���]v\�!Z��.�O�˵���� i e&
a�%��Q����9��CE���a3�������QPRuMYl�T�s)%mS؞|�����}���IZ1-�Tjn������g�SY�Ӎ��7���7�Ur���J�������l������f�q�<���a������z�5� �p�É=A���a���n������Յ2⥗�J:��Y�p�clYi+�Ӻj��MڍL�z�Ĳ�".q��`��y�;�~V�y,9���#�z��,u�s�bn#�|�뭜V׊X8��3Ւ���4��4R��,�c�Fρ0�q���ܺ�������#���]��
ަF¥�R~<��4�:�`�Y3�_lAN=�`�jU�q��/H�����rD�d>�Z*Y��؆�;ʶ�*$+˭�>����.�N'B�Oy�"	U=��QB�{�Fq�Ɨ�O&yԍm/����9�hٳ�l+dXiL6:hzw��-߱�F�gV*FK�ce"��٪1��fF
J5�!������|�W�G�~���vc��'%mW�����خ� �Dx���u{���NCr��Ѣ�~��(�s�}�
ܖe�`�c���eh���K~���euv�y+5��jp���������qA����-�GE|�����wWi�dCA�ֳ~s	l�C�Z��g�lGyN0o��&�����2���-i��rS�v�R�EF�v]q!�R5j�Z%���B�.�oW����ai�*9�������z@G���Y��=T�̘5��d�78�c#�3+��Q�����}�9Fvw�f��A���{���uP�L�(�^'�s���@���F��\�M:��w!������,�z~�2�qD��d[%�١���1�ڭV���&ʘ\ш��ް�aa�="�J�b�4a�9{X�J��h�f�>��Q���]W�?FR��w��B�Z/1�Y!p�
;%TzH;��N��=���m��/,��!j�a�t\���✗JQ�N�����*6���<hs��Z�����?<;���/�E����S�f!%�2ߏ�=��l��t�a*}�?��P���X͖J%���>�U�<5�>I�Ai�}���:Ǽa��d�N�Q�#ć֤S�u��-[�����E���Rk(�\8���NԢȜT����$�EC.j*U����ŧ9���9X�T�m��i���b@-?�"Ө3u� �>~z�?Q�:˗|_�x\z(Qe��S�������Y/D-��v�=kc�<i���T���2��������p��͟��[Ȇ��9���n�t�0J���;sٱ���MD��8������ߴ��c��c;�w�m�=*�#�;"lyÁ[ꍢ�#���c�8��MÊ`.9����[�jj��}5�U�5W���fCm~�V� O:�;^���6���G*����0���Q��b���==��<�zzzs��G���h��H�y��'���;:;�����._V��J�K�:D��MD�6�5�M��<�[١��v@��Q%F�v;��Q!pD��*���'�u��8B1`��ֶ%�����Q��	8�3Ǫ�����7>}���� I��[�V�C�y׳���Q�nZ��u��a�`���_oC�I��0X��>�wؖp�$֟��!~��,��F������_bx?���[8���"��{�hm�X�$M�" k���r�)/+K-��?�3����Wj��5�U(I�F.y׵��� ,d=ކ��[4��rx�l�м�U�|���g~��ǹY��42�rC�F�/�A�E5zB�����a xV�0��?\�W��kD,�,��q�\o����sC-;�<�曭�Oj_�CG���P�5F���餷��~����
Pd_r�=�Ľ(�<�r�&��yv�Z�?���p�(�|�>���G$����6�1Q�#BM͕�l.%T?��$�^a�۸�[UZ�恻�y^PW��P�R擀��99V�"���a��q���G.,/�=��I��B	��*�'J��{�� 5Gn]yMC|��˷�_Uh������:�T,KZ��C��""��ρ�W�I=�8@)2�兩څ���G_9�]��\wЈ�b�����y�~����YI��nf��Ӷ|T�k�8+�
R�f"�#3G|�"(O?;W��hc�a����+�����NJr��\7�21.Zac%�{?x��xbb���2�n���V�O��&9>Dh�5��yA����9�h�6
N{�-�e_���2���ܔ+m��(���}&���5���v�%�m|���|���Z��c��&��%r�V��&�9V�U�;t��ς;�{������|=t��ܳ��>���%UGp5���m��`�����_h|۰*�����G��SϣV��Cҙ��@�SÀ(G!L�[\��4��]w��\��;�	�I�.����%�����{���?�ꩮ��5���}��ʦ�cj��������V�ep�z��/ج���\�K�r�J����;U��}�R�AUO˲�Xn}����$J)�39�[W�R��D�mzVL����ڶ��:HtU�o��!���"�WO���G~m���+�)¢w�Ѻ�3�t��B@�H��Iu�z"~��9T�z��y��,~Y�r��؈L?�OK��k��R�נ�ϤqmG9�x������j�6��rL��lֻ�+�Vպ</O��5�a��Jqc�rȴ#��2B��q���͛�3m��4��/�Nӱ(�F~�l3��~$}�ѫ�|Q���ᤅȺ��v�,"q��~&B8�7@.��Zҍ1�)��d�w��mC7ag�Ԭ����\eXv,�U��2Ĵk�3mocUy�hnG9!L�Q���\���l���Q��"f�������&��y~&��b>ƺ���l�E�+����5L�:Ň�R{1����Jx��P�aѦT��"���ߔ����AM
ٳ�b����m�n�8�F
�>gY�f���7�Y]_/ۃ��ŏ��� S�r�ax��H{��n����Q#&��8��>����T`��0�'Em��bH���Z�Z�mB����ؽ�
i�I�Q̛3w����~���~*J^B+
`��r��4�󇽭���<X���J^�W*����;WSi��15e6:f��L0+��{�Hr��qV~r�I`���CI�TǅIO܆!"�kl���4�D�	0�N�d�N.6I�5�	�xF�)�Ԅ�)�������h~�ۄ_|C��ѹ����3�����e�*V�>_�~*E���3#��f��J�Z�"�}+�R#>����q
�Fe��������P��PF�'|sQ��:\���������0��-M��!܉��Y		��`3�i����Q����
d��V�'� ����H�9�����~��0�c�!��x\��/�X����\��
f��1��t<�v8�㵻lh3��'� �.zv�&zC؋����~!����W�?2��%l� d�_�{�ⰸ�yh=W-SG���#�xjU����]�Q�+U��>�^��{�Rk&[���9��YZ(!5���˃j����M����s��&���&Z��τ��b�ϲf���ޱ��
�D��$��ݡY�zq.�Vf�ZߐT��R 5~�&�� =V1��\u rq��|�U�m4���{Ujj�]�R�w��c��Y� �/�ux?q8��q�`�Zu��IGZ�j� ?��U�l���w.m�q�`f���d�E���y�Ԓ0^�yA`��	FK��z;<SȮ��9��* ;�n{�<��h}D�'�w�7q��?gb$��3��Ǒ�/��>@��R�а�j��/`e/�v��0����h��)GoQ�F�f�|<���)+�de�T����.amM�fPS�M���~������H.� �6<�4�/�	�F��H�+���as�
��][H�y�X�;_S�y5�ȿ.'*_~`~���V?9���o�t��p'�!�K����$�}}ۀ<g
x��3�Q���Èq&ls=0��+?6��b����D?���uY��y�Ű�R�1u��3#�����ߖɀo?|�J�j��ױ$�:�>��_N�o����e@�`��ͯh"��+=�����3��+T`tW�y���J��|�����9,S/��S�9��M
�*;�1*_D�G�����q��u���&@p+�<3���;�]\���P�[p�1�Y�U�������AI�å[7��J����v���9U��G/`�ZI��Võ�y�Kţ}�j����ǩ�E�2הR�U����*҈@������M��9�p������b	HN�D.?�>�u����Vٹ�K�	��!y���M��#]7�i�ߞ1T�>R��6�h׿L��uJ�H��/�2�
�,]vM��6��$2���g��z��P!������f(�y-DE���#�}#*83A�=-���%��)z�π��8���p �D�P\-[U�i�&���͏�%�����ac"�H`��[�wP�W���<~B1�6c|�.ń��-�=o��7UmСZ�	~�rld����9��L+��_�Nmq�%���x�U���<��h#�Q�9����U2��K'K�]��-�x�	�w�]]��8�o��6a����0�[� ����X�ҮQ�a� +�#?�-�H/Uz:��T�c;�W�!v>0���RZ�0z_$V��]�$��c9�t�\��:��UbV� '��-���%M�8njy��^ZG��lS^���*�y��&9�?�^����(�P�"�LϨU]s%o�}����ɔ 1S���Ѣ����L����
r�rf��W^����L��&��i�	f����2ii��T�g��[2��Q��������~�ϭ�0��p؆�߳�q�?u��������5��]�=�.���������C�Hv�螮	V���A)R��y�N�+d���G�}�;��4k���͌s���rP7�|��� K�	')_<lʁ�*�X�:[JI"ڻ�a 2_�����q��C�_G�po�0\�`��@���Mbt�I ��>���y�J�f=��>
�����2��*h�}��&��7R"oXv���`D��� �DBiK�IB.��Jr��"s�q�-��
ѹ�d4���Z��a���<vSM�n�RQ�)�6j'4LI;)��䤐.
|�S)�̚�>2ք���
�K�����z��E-z�N[�S(��n�J��hh��o У��M��T�4���2I�5�u���'�� ��K[��U��&V���~�b�j�L�W���|p����Q�� �}��5��z�P�|�6����$r���-��A����B��x�P��/�����~Dt�{9�j%Z'[*o��ϢX T�PZAɴ �.<��鑇�1m,�ǹ��ͷ�Y�6`.��O���M}�|�)���y�F�
:���@�m只L߉eE��W4.}h=o�����9���	���˞w�m�W�qqw���3�:�9SH�U�ԬɇK�#�tÉ������-�=Uq��Vz<r�_Z��F�H֤~��ѕ�)�>�K�ƞ��	W�c�G����&�s��U綈��~�~5N�{T7s��j泵�9�K�3��0�����QY0*�%Ә�e�0(�WwFN,R���-�om�����5;�C�;�Fd�7�a/0��̇��3e?��<��J�TQatZ�gR�Oa��fA�(�3!�y�Gm�hL#�|�>2��5�#���jՅ��f��o�Άu�M&��|�3V�{�qa��^szJ �{�-�2������3tL�jѯ��Ǔ�q���*�h��yޛq����ݡ	u#���7Ɯ|���3/��q�A1�T��֋+�2�ۘ�,Wٕ�����i�x(zd���������l��K=�8�I��*�8Ѕ���⪍Ӈ����2`���;X�<���j�oJ���4z���/��^��n�7��BcM�թ]Z~-;U�����Gw+�)�S}"mp 8�����l���w�{f���h4_��W��:�b�w��$�0C�	����h~��6e���c=S$�2H��]�By�Oy7.h-E����3'PB�6�Z7��I��-��Uh�NR�zF���m􌩋�"�F�$-��S�a�?t�{���߬���QH؞G0��9����~`q%���W��y�-���Gř������|y�sK��\	��Hի�u�V���brs_j'f�e��.�5�~,���c�n�ӽ�5\��l�c��<���(��Ia�0��u��h>�F]nF�!b�E�q��:��o���JҴ倞֗�C��|Y3�
f���XYX�z��|(j�q�=��P��zB�G�%J��v��^x��U��&�}d�W��+�!e�-jL�j5w������I�Xը�b}�%ض����W�UT%��ҧ�9 ����/�{�A�c�p����	}��;�
�$��T���9�ɴj�@���X�q�fJ2:�8��ߴ�~��	z�t��d֣�O��G|-��bRsO�H��1��As�w��З0� ��]��O�\�"��pլ��!NtTg_�k��2�M�6�B�;}�۞�_�w�sՍ�>#j�U�X�YФ3z!��ą�F|H����8Q� ��~茪�.XHW�g�Ny��@8k���Ϙ���\\��X(�AՋ F"/�'c��K����2��z�Jilq��I't�戥% �?���Њ��o��m��'Ғ�o8�?�(w� �__{
�A�Y�F���߾���G��*�UE)ey�ھ�y�'B��eX��CۅD;�����;��/��i���I�g�1�)��(i�V�@��,��9d{nr�q�\#����'B�WM�<�77b�Σ��XB�N�}L����_�����x�2{�b�^��])f@J�d��}���,�~
|zcu�����3c��:�?8`6��0V�f�'Wa��Sm�]�"����皃�N�^ٟ�8�ي�Dm�WW�b�DFo��R�?����GVo����9�>��z�}�X2p���ʡ��Z����ә6~\��x +}E�1r+Vd����i�w����pFo>p�c��c�Y�hCW/�	�G==U��gz���m���vP�tz�]�͂niM�f!����Ѳ�������c����czS+r6�?�9���Wr�w�x�IxO���N�<I�_��^���k6�jC�O�o�q'�.F�X�.濈 Z������b\䎜�E��]z��������U7r0kg�k��$X-R/F���g�חq=Po�+�h�x�2�!o������gw�x)pۻ��AFYr���3{��%ԡ��BpRdBe v�UۑRx��~W��,���Մ��u���ׁ���%Dʼ|�33���+ٵ"��]�i��(��;_�v�`�����r4���B��w����v����?����{��/��_�N���a)�C�$׈��t=��ޠ�Ve؊�W`Fư�g��~�Q ��d��9�����͸�#QO1�.�t�������#�!_�gb3����RF�V��뮔�T�������
�l���s�^zт\���k�@��65��������Ᏸ��Z�\b��T�` ��P��x�q�&�z� ���N���kC�{*绞���u�>؞���6+��s]|��F��&Im1�iW��"�#G��ht��s9�t����<�����3�#�nw�`�,y�C�
ɸ�$�녩WV&�S55l���O�?�O��A�Q0PdgF���q�2�6H�(�0f���a86R�X��%�&���˜[>nJ��{���I��=�z��'MR-ؖM�����bUC��mQ�šY�$�䱟2��>����E����~��(V1&�)�y#<�����m��쾧�I�5w�?��5���Nޱ�M����<W}��*$n")��"�rٶIl�L�n@��0U2���h��PIv��0�O�JE���0�<�N�];��$[)5�V
MU��NH��OH�Sz3h�@H�u�,����v� 8�<�;L���'�;%Z���&2%��V5�wĹy�W��e��W�ds�S9����22�C˩=�:2/5~�@@bH�������H���yLt��9:��9�H��5��{Q���I���l�L��r�䁳���_>V�To�������o��'0���+Iw�V�N�f˽P���*ֶ�N�@q1:���'��NqW��� ��ٚ��˳�~��'�u�4	M��~PC�������@��ýe�&���n�>����	,�����{�o\4�h	���T��u
�I�Ս-Q}jqR�Ɏ��g�f*�8d���qXB�zJ�=��i}�}F�_t���1l��rz\������^��а������*u{�H�?ݝ�`���Sƶס���5Z��Vo��y�5��Iɾ�Z�A�sS2zZ�:Ֆ�^��^��B@x ���cלѫ~�tl�͗8�7��z������L��p۫ek�"G�qY+����p�w~�p�N�;��tb����ζ�!��af���J�`��쾺�z�{��l�^�#6~)��M	�����8�):1O�ӥ����\�;D/r
�n���C�����a�u�Q��m�-�)a�Ce�Z`�s+f><YQ)��P�p�됗d��I�ܴ��Lr��I�M8��G�?q���+dn:0ۣ~�Ӹ~�*���Y|�=�C��f䍱�1��Q��I@�X�R��(L9#1F�n������r��3	\�V��$^Edf����Nβ���]��rK��X"�(�b�1��R\���;y�{����3^� �"@i�f��$��l������LE8�#�'�+Қ� � ��n5�v���ɋ���cn��Fe�/�d�Ա7$����"�C�Q���I�#��*ʎ��,�b�荔�C@HD�%�?�NճG6�R"*��֋9�xȊ�˹"�����`;4L=��m�&�c�.�K U��"z<�/Q��$dЕ��x�Mn���[�qŒ̛�Mڧ]C��âZ������=,N�(/���D��
ʻ��T�����;c��鼰��C����Yu��� �\U��Z{o$�{��7/����!{�x*��'�ۭz�����j�[�a�QŚ�P1�_��LM�������}f@�H�L�-�Y=��y/q��������y�:\�L����D��:�rކdh��@�+dKv� �S��%�ng���^�R���r�Kf0%,oS0�q�ѿab�M�A_5$��l�$D��fZ�Ly$K3Txsf�}"��M$	�}T ����:F��-�����=��+�l�WԷY<�,\�ݯ���B�ޘFQ�����{��p�,?�8�)Rg2����� ��9��4��D����bp�%U�"�}{��nD-�^]ݠ8C.q͠�t�W�*��	�q��螟��q��Tf%��)���H2I�e<X�.�%@2
�V�ȉZ���A=����K��J�p�}oy�B�*D܅��ʶ4�-�z�_������"�%d�7nkf��*��/��-�D�����JӮ~�:�XP�[�H�滎b��+_�H�a��~�%�B�O�Y�S?�2�I��K+r����U�_yە�0�&�##���� �� �w��*�z�s
f,uDPࣰ>�8�9n��m;��~p��������F�wEc'�\�Z-���7��H�!�G�w�gNmQ>=�#h�7�a��o�ɰj�Wp���sf�ܯ[����΃�#�����b4��J%�D���A=�K�<�����%.��}?��z�P*����T�R
@b���trD�s�Dpfj+�$�U����(��L,�Y�&){���.RZA�v��%rѯ�����!�%��%�s��OsD�e� ��`?<�UV�gwW'�x�5mD
V��	f�q�;��J_1�|g�g��Г�� ��n4�hDZ"�S�!2��k/~��ƔUR��@�홿�(CM.�:`�]�<��9���j�K[MP�+2�C�,r-��8�]��[�W�xNմQ�\�Pn�B)�fQ���4��g<�{��]U�s&�{��윬������<����a��c���q�s�8��	�
y��FP]� 
P�0i�jc�<(�|���^�������bM�a5��&��t��eWHe�Ll�6���W���_v���74-�α���d|�N����ٲ��Dz~(ۄ��ڵ�Ӡ��[x��6��z7e�����q����
+��^}1-�w����mm &-G���DAPb��˃�˽��W~�c���0R�C�f���F�����k��E�	N�<'�l�"��6�,���}���N��Vr_�hMy��k;���F;owk�*�l�Ng%���ח�'
�Y,�a�1���pZ|"A�x�aб��Ef��a�Pq�xm���ۃJz��t���ۿ��7Y�@�^�eJ+�4%�@ȥ�bǲ��>�K������O��9;I{AoLB���z,A.�^����C��[~o��T�&�ާ)�������!��J�`o	U+^'���k��o���qidtr<%:���d�.�EΈ��5gV��Ʉ���r�]���NZ���+�f~J��&����3���d��2!?\��}�8��j�q�?h���Z&���:�mT�F*ߞ A��A���R�.�A��>Ok:���4L�'�௅���)�h��'��+O�+�Mw�J�UZ��D ���k�{ӷC��ۧ�<�	�1f��D�A^[8"�Q�[�#�&���n�Vp���_������*�o�]w�!��38����~�:W򈤵����gfQ/H�c��E�ʑb�[M�2F�h���=m�'�k|`�Y*��=�Ywn��o��l��̓y"��Y��>(W{4�h���QE�d�������x����;n�8�!�;�*_y�l����Ze�*�;_þ4t�����_�zC6-#�#�>��B�-Xғ1J]�U�F�i����O�E���ׄ�<�J�y*���-2XT|���i��D����bL4�^"FÑ/	�YQ����
��i]����9�B�Z˕O>��i�� ����>tm�	��η=o�[N~eo0'�����,��,ZW-�V�$��%ZM�~��I�^�����˸ǌx�6���mO��G.�f�����LU�_�!�@��H϶Z/D�Z�F�r_~������}/���N��ɣu debW�V���L�k<=Z(��7��xn��T��/�bA��xa��7e5�6$X���s
*(�RI`W�B��\����w�H��rp���e�ds# ���x	�1gHC/�`g�i<�p��Yh����ϕ�2��_��E�|�S�։�8�	M7Y���Ӯ�{p�s���2u�ܖ*?�$R��}�aؼ��vI��L k"H�@W�3�Q���H��XMu���G�s�D��G�8����g�	Kx�6t��/rHP�('\����D���]�m���ٓ
��6V�mI��ݺ��d��a>&�$���,�̜6��L�����=�IBL�ט^W�wі��m�����"�[�?��گ���q�3o0�Q���lh�H�)�h~QĞ�pc���*���C�����$�QT�>�B����"��#8L�"'��b�Zai\D��s��_���;Ԡm9��(�y��K���T� ���`��V�=�E"���� dM8O���<�����|ZCӰ��I_��Ɔ\��"d.�9v����:�
����fTz��N�Z!ۮci/��}�ߐ��΃t���_���7�H������y�����J��]���K���E&-�C;��L7����2g؋g�~���~Ӹ��&J��p�ۅ���^�$�z����.C�0���X��4�)L���c�G����6�c��y��{��K�S���*	�\�m* �-�Ƕ���Dǵ�|.��5�GlJ��:&�3���t>ysp2$1�9�(�����v(5�k�1��x�b��E�u|M�ݕ����"^��8�e�|^����A���>5�W�$�p����=�X���X�����cw��}��=q7��~:Ķ��\���'jS~��l;�W���	��w���k�0Б%��soU��E�;���Ԯϱ
i� Eh��# R�ۼ\,'��4|
��ș�ZΛ��7���N�41q���l#u ��MW3n�����Y�����Gt�s�\~��b�Ό��b�$�%9E�������R#���Tk�N�2�˩M��dt�BFcEc���]�ЄYqSw�It|��G^�s�Y�m��z��,��~5l��+I�SP��7�3�x���OW mTc���ʚw�&�5}�WÒ5�bˍ��=�g��">�$G	cѦ�R_XA���.�ֽ6 �jt�{�ifX���	����Q�I�#���n�;�����Z,�P���+M��E���h+�m�*�3�;������6|�G��VԑŅ�<ȗ��;�g.��̍�7?�E���rDa=�O�c.qM]�DLE%��XY}?��H�LR���&aI%���la?l�c����Ez���
 ��=@�������G�T�y��N�ʄ"L�<Si��[��g���0�l�i>Orj"���@v:t���Q�����f1�r�b4�� =��Ec)���aj��1]u�_L�p@��`n�����y7ˈ��&I�\��j-t��h�����Q�:�L-��/���0�	m8�_U�u���l�2��E�1��v��D�Vl�sR^�K,ⷩ�A������(���Z��bc縳����Y���;_��� ���Ɣu�����~w|���i����$��FDS��5/�&AY ��m����0aֆQٙ�A.q�Z;���Io�K%+��.���:�_�t��þ������ﴻgԬ�<��(�5��~�6��u՘R�$
qi�4��Y��u��n�
�5���g�5��z+�����]� ��2(�y�Hd���Ș!_�{4~�R}�!�a_2�;-�Y�S��8YSp�F����C:@�c�����		��Ȧ�]mƢ�{{�J*I��\��K�O�q�=��+��e~���;��/iˉnt���%8ű~�w��f�cÕ�a�D���:DV���2�)�;�S@���b&��J'tY���N���̢1ߍ�d�W;��֎������	)E>��@��tbuA�_v��l��O/���^T܋D�{���@��;�V��|�q2"�XŅF�������j�_6��/(+�>l��S�_N)+!�M'��N�ߓZ�M�ܝ:��-im�5���gmx O�>��.��U�I�7�ˊ��q�������zڿ�!�G��'�b-�}
�K�D�G[o7��P�]{�kf8M�ٱʟ���#��B��e�q�n�х��u	(�:��}yE��ݸБ� �ŵ)4��]�7UR��q��_�G�z�d\�?��B=�}�$�l��"�r0s@4��Ԅ������HU".�L�/M��������ʨ7���8͜h�t��)���_����T���v�����HWq�7z+I��1J�o�����'7��F����ʥgO�"Oh#�A[cg��w�I�]A��ȘnϲP���T�Vy~ts�R<M������|�kTJ�_b'%��9�^n��	�~��#�!�)r-�h�\��z� "��v/7�'��Jr�?,�{��-zdP��¯����dXz� s��K����hF�h�`�ja#�T����ǽ�ӞM��$_�ƹf���ؗX�h���4>E$%a.r��}҇��*L��D���m�5��Q�Eߢ1v���D�mo�Ġ�b�u/�9Pp����	ђi�%���AM_�~��r�kQt����+���|CޖTxg&�������J�T?@c���+L��OjH� S�ʁ!U�Yo���S��)��OXo~}�����᮴�]w����|��D�#9�s�b���?1�nOcz���dӺZ���/(��G	�֖d�a�e|/s�� *|���3'챵Ԝ�f�~�ƍ/AwK�������H�nE_�A��.��@��3��̸�i����vkS��Ob���5��CfҮ�P�:�;0\��>��pJUN<R���t�ǧ29��	���C.y0�c	P��p�܋�t����R&G;H�������j�}N����5)E+6�Y�&h� g�ˑO��4����G��E���5��;��	%mS-�I^�c�w䇪.���t$�.	e%�M�Q&KM�q�'v��H� ���H�:;7W�E��rk�XÖU�)�^u��nC���_�;�������ƷJ�cU@�	�|�lۯ�'�4'����N�6�sG�Y�N\Ͼ�3���c�cc����|���=�:w��T�SE��1P�L�߰���vqb��,`l"ݖ�D��j�C��	_]7��]�9^[�
�IR��W]w8o������Q�o�W'��)�㣏����u�"[���
J)1���2QY	h���YB�����`&Mf˼�o�%�6�4��a�;2�?"��ھ�4yi�U+�J�8M�nG����&/�����%ȩ\o����U�2�/n�E�C�,jV�ڠ��E��B�w��p��\�_�nv��ӧ8�s�J��R�#� -�<X�W��^/S��*"n��n6洓�~�w�̷�Y7�D ��lc��?��7��&�􀳖Q�X�)�N�(VY���%�sQ��zYCMeq��h��4����>m�>�ID�Ӵ��/#S� ��kԷ���6Af����9���j�	F����0�T�YfcԬ/U���w"m9^�/To�E���
9�a.{�Y���mP�m����!�o�Z�vG��ث���Y3}�}Ы���#٭�`ö+bH�����,km�/�٪%J�23ڽ�.��ϩ&���Z�����	�����H���u_���`��,�L4W�����P���y�x��(z��9��A,du��乛L�x�T��0��#�
��LZOr�1��|}P�b�ˣ�ط�%�W�0���TD9Ł �.��{���������u��Ї�3��DX�$�4k�6��|,�׬�,f!�X`�g(��P���[Y쏹�a�2����jM�fu�D�·Uѿ��OB�/lK�/���5���\`C8
��P����?ˣ
��v�K���gƛ�����̌BV��]m�]mk�CsW��zM�Wn�*��'��5�r6Z�5����mߞe�Q����Rb��G�7wF2޶?o)�ҳ�"�{*�:�䧦hޭ�����0���a[�&E�~�r3u��,VDS���_�=�*D/�^6�����ĮoEQ����,���핞F&`�%��j�9?�'Nh��U��Go�bY����~t<��?��}�֧�;ś��������~,�^E���h`�|"��wj}=j6�.~mL���P�,a�M�o�$E��Ԧ������Q*e{>�-�&Vo�B4�b|�3>��e�0�	���^�������~��l�#�|���-������ؐp�3]8t7�[i��xB��]ť��9%��m?�M<gy�-v]�ޙΗ�1���-��j����(�����`��TG]���I7'-�:��/9Tq�L��K
%���K<E~�� 﨟�Y���9}T�d�@t��+gl�7�k ��`�\���v��]ǹ��9[Q���u�<X,�rҊ���՛B�N���y��e�a�7j�m�9��翬�l�q�}�F��u��r�ꙵH��9�Qlإ�ΥE�aM�M�.x紞3�ӓg3������,,y	�Z������y���Ϗ������`�N�lQ�����yq��Z��v�\^.��������6��jr�U3y-n��˗�3xK��l���+����c�1d�]���k�q��1&�=B���f������,)�8[����RJ��1��F�0��Z�u�G�끛�c�|�E���ȩ��f9�k�a<�v��,9���"���@N�:��B�?(�m����E���Tc@璩pտ	2����0c��LԢZ�(�jQ7��t��1`�Y�K34˳V��DaZ)Ǌ>�)~I���� k�D��x�kJ0I7&0�F̣Ƿ�ER��\9�A�T_����t�_���3�8b�HU���mƹ�(
u�y~�w�q�d��	r>[��ep:B�u�Cv�(/5f��-;s��zJ��s�<ℝ�|�A��.o�G��J'~���|�������؊��N��c����F�ab�X��p#�)z����EB��"-�i����e	x-�F���>^E�57GNj��qa���̇L*�|RF!+���HQ��rŶ���oأ(lf��9��Ĉ)�?�X@�0`���|��\A���sI�=��x|�!zV�5Y6W�?�Sl%���e�ݯ��0J������
X�
���MǛ�DV���4��!Gg9!���<��μ ��M^��3�nL6��֍r�ܚ�ڢ��V���s�������Ϡ?���f�=�v5��1�@Yp������zk���ד��/fF�T6����'E�v?`��E.@���=Y[��n�_��7WJ0?:�*��ZoG��C�8`�۱<19U��:"�`D�D�b?�;�&[�M�9���_gM��m��{�}�L�>���|�_X�IB�{���qf�
���jk<���kci�����{��]ko^BWsfh?��ǡ�-�.���V$��_��W�7O�?wx��`��(���ȋ���_.6���v.���q��G��[P�眕8�L�l�?��r��t4�L�|δ��m2铐�[@���i�L����K��ݸ)c��^d��\���?�Q�v"�뙖�z^��hǲ=�2,�F�ط:�kK�.�0��\4�fQB���P\RZ���)�nH���TUg��I-�
p��{�B�v���X}*Ÿu������y�@//G��D��o-�]x�x�T_��㖺��r�`���y���yFSg�4uT�r���z��,�F_}��߃c��.���ܯ�+H΀���k!9��[�Y�f�TA��|�=�����ÊRdƩX�!u����7�V�-�I�\eZe�BO��<����H��hO�֊�<ڿ�K�
c�+5�2�B����ǈ�E�ȕ�<:�m�������u��8���%z	����d�k,���pam}o�G�eL�kI���ફG�&l�'���3V^Ͽm�+V�����v�PY��O9f��7\#������@Ԛ�ԧ�#?�.�<��v/�o�x+�{��9]���a�U����/\�23y$xX���+�'�C����;�h�7�D�_:N�ؤ�q����p,.`P 2/>'R�@������l5��%��R�r���5'����E��eG����&��pP��^�e��V��5J�l{[�m�6�VW��ϡ���Ʈ�d�H��Y(U0V���^���$�ٵ&e����&ȗ!A`,I|�O�ΏJ�S�b�C5r<��qcݷ��&�M��[�YC��{�3�H�1ع��/�䇹
Z�1NnS`�\�w�nC�ʙ� e�]�c�C��p�\�C��@*ߥ�U�9���RlB��'��Iu��4q�͠���^C�x��RIZ��b�B�����q!	ֲ�քi���� /
;ɗG; �2�K���C*wq��B��2���9m;0uRsH<��pRVB��6�x�e#����EnL���w2T3�\����<���8tn��VFZ��QG��;��N�G����5/Y����1%�a��ƒ,aNk�q���أ����4:����ߖ������s��߇p5�v�;�G��*m3���D�i�y+K����vu���=vc#f�� ��������k�q�΂LJ�:`܏J����C-z<7-�,�ձ�B�N���"�җA#�&={9:�����{�kMk�V�� �e@��[����oS�ç��hv]�p�f��D�R�0h�UR�vЌ<i�v��؟�ˀZ�#���2o�h7�{�����N�+�i�m����2i f�&<f��:ޥY|4z�L#y�M�V0��@�<�X�o��.3`/!���j�rf�����ɠ���1w�H�L=m��>��|h��}�4n%I/ �OJ{
';+�ZT���@>R�XC�8NR�<E�b�
��SV�dA8�*���n��r�x�:ex����WwO_�+�2�
������w?~UV�Y���d�P���K�����]��ȸ&�2�/�i��^ϕ�v�Ձ�+�z�̽ց�g�%�R�O������F��Azg[��� bG�x��z�x�Bn3��1�4�"AQ�<9�/$���r��g��O)�W��&�"�h ���O��J9��||(���`�ٸ���������{>jL�V����7�G3��_�}ZI�r��;:F&'>�'D��N�bm8p�^ϣj��H�#�j	Q̱;0K�c��L�.�p:�LYޖ�CiO�U��������#�f��n����' R�SnW��	M0vt!,��@s�́+b<�ڕ�ާm��_SV����e��N�C���*_;���w�tM��c���I ��F]t�����bS�oeQx1e��c����ګ��kW�������H�������iF�'Ku��ݴ�~b��UF�q�}+���U�	u�������u2l:�ޛÙ����,�8�7P�ߓ��������c�g���xUKkV����jk�ޣ�����V{�M��ZU�w�{b�رS� "B?��y����<�|�����''��Հ�L�Y����l��M�a���k�^�����o�fl���W����bF0値az3�t	ظ+��x.�3�u'��d,I��~'�L_͑S�u����;�Oh%P�+�r� 
��x�Z}��@+@ �� �B*���������n�KP|v�����s#Y��S2��uRS�A`�f�K�s[Y����U�F������� ���c���� ���9��%XW�hU� �͹bǮ��'�n�����=ӌ�j����8����C&G�>���T��g9Ѝ����I���!�<�-����(�\�j���C�5E#f���w�C�C c`~�ۃ���0��8�AB�u�m������W@?"x'?�b�׫r5Ki�cr=r/�쓈Hj\Nw�Z0�u�z�L`t��9 �u�<����k�1<�/�lJmB�H��]\L`�?�_�����3�90ֺ��Yҭ ���ӓT�c6�t8�O�eTM8�������c��LWsP��cI�y�}�J"]F�&��3�����A��0c�NaP�`�b�����m�M�����
�!�J������x�#�rs	O~�l�/�� c�so�a�:���-Î��f�*~��fff�+�un?(�Q*��4@O����q�m�� �%7�ް�b�%���K3C�$�~���Μ������&�(��	M��#Moz{�Y;z�^�M�O�|����s�Twn�Hj��]I��c��3�d��"�LMH�GE�F�Iz�(l'*�|:�+bbB=9d1�r�҃��L�`�"�#�W�O��X�0x���h��q-u�x��OJ[J���p+Ώ3+��1h)�bW�0c���$�����i9țgq~2�si���!7z�+z9
o�_be.�+>ѓ�+@F��� �1�p���K�/�2��� �x���y�<��!n�m�̳��v�]�s8�������.F��f����5���dG>2�#�ՙ����^=a��#m�0"I6?�$5х۫8��\��3�XmTHG�y�(yd����B��9r�P^ѝ��'zf뽑�k�iʍx*����(�|�f{39�����@�o�H?�U[��<3<==-�K����G���0f���?0�!��m?lsp3��L�|��J�w��/��.G䢷���9�#lh>��?|ٔD���zO��@��BU�k����B�zgJ�\��vO���$�\'D7�tdZ97�e`
���W�����>��P��]M�*���G��c���$_�9
b��ę�밍[�g� e8�4�8���O����
=�q-B�@ ���95������E���zU�sac踞�[��~�T���[S�q���T���a���a�	��Y�C�}[_�
�c�c�@��ʸ��z�����O\ൔ�*�]�ũ��i}�b`�d�&M�ؒt�W ԉ�?�M��(�͵r��ߦ/p�ど���H6�g�g*|��p����t�O�~'vM����9��l,L,����h=�;�kߕ����*��`gN�>Ya����Zz��xS'}�f�k���BÓ��%�'�m9]����z�LRyl��<�z��I�����n���q�����H�~�E��E��Ս�v��/䳊��_O�3� >t>��H-���0�� ��Z7��<�@�l��[n6��2��K��}%����Y��[�mv	��l;y7	�S����&�K���y��O]�����[=(.?gt�&��CO�.��>W茂\�(�V�����,��H���&$mj3�Q��>wj^�t���x��,X_�֙�̄c,��n�Iɗ�I�z~'�vEL �G.!�������6%gnC�2o������GX�&&n��\6+&����]jF�>�~n�3� V��o6�X%@��d(��vy�mTo-�i�-4���%|�赑�4�8߈��X]��ڊ������"]��Y|a���l,�c��aÇ�y�a�\���~�����f�и@��'M~x��\	��^�w�n��F��1i,��2Gׇ1�@�S>���#�`�����&�#������囨�\�O+`#�pol�H��c��S�\��A ���m]�:�Q�YZ���a_'�	��5�.3sgݶ���g�v�o��Kj����f�R���O1h�U�i��قe�@�W���t�H[��2A��*��:�Ù��q�{�����ÒT�V�|�2X7����>�\t�龕�W.�Q1����]Ԧc�].�	`X�w�Ѭ��+TBrkp�h��7	L�F.]�:�26�.�)!�>�^P����u}2�=���Eƣ�{AD�_>��0��L;*���!�Q�Y����wL?��/S\��]l��}W�YC�ԃ]��%?��A�=���I����4mF�| �	��C� �N�Xr����L�'o��Y��n�V�����j��N�b�CNG�����D��$���C'��F�F
��O'J��E�
d����gv�WZ_�:
�;	�� �	�Ӥ�����MJj�(��ǈLC�#l�U6o�뵲���@��l4� �:�x1�^p�=�\x\�^��^@9
3�+
��^���S�}���$��oɪ5�{CY|\;��/Mך9^/�C3<��>����E��	�l���$]�Y��jL �RD��&��vߠE�*e��NM��ib��;`�������Sss�<_b+�h��G��c���������B�d�7֑��Fyj.���S�ܣO�1��w(xrSf爏c<��B�cBC�R�r&�q�'b���^���4�Tb0����o�4�N0��_��l��t.z �08��[�w�B��Ĳ���헰^�(ڗ����^��U��rTЯ��EFo$Xy�?�~P.e��:�kr>�Ǵ�Ȩ��m1y���S��i����E�$Zs_�Fs:E�U�t��dn�Û�}��\����,X
�;�����"e�eT�WM��%X��܊�� 
��;d�D�^����X�Ǉ����[�{��j�jxh��g3��
T��Y0#�t]�g�	��?�V�^��ˤ�!^)r���p&/�}k��.�yr$7D7��k!�,݇���qػ��N�=@�����V1����C�m�X�>�oMk����
���(��gV���{$Ǌ�A�^�#q�6�]8+�jJ�z�A.���M��͜�7w(������]|ÿT�&_�:�Q��d��š�r��xxlp��5ؒW~�~���������byL"k`����*B4�F�Cj90;�k����+1�o^�ƌ�kte�L�.Q�Υ�6��Ont�A�����(.@N������P)��%�O���-�Sm8�qxO�j|W	��~� 6�*�=1t��7Sv�֖u������+@�>�Y�<���7�|	Ϲc3�U��y��*laR�*���e˺ Z�}�ZJ�J�>?%�~�����/imߢ�D����I�ȜYޱ��ה�HJ����Ӂ�#���w�K�V_عR�	_��p��#�.t6�t��*������� �X�9�:���A}]*��j�@^T��h��$��sN��Rǁ���U��[���wfp%�#+D`�����Qt�z���l.�#���J��{A[4� �'u��(7�ƈ���_�ʋφ�<s1[�3�ק^��Ǝ�aר���q���Ih��i#�Q�����y0�=�1uo�s��h>�&����I�b��bF	g���Ľ|�DGZ�y(E�u�g��ؒ5�bm�cf�RnOhc��WQ&ᓼ�Q.��Xu�,�a�/���UT��Ѩ��B�k�apܛ�0�7�;-��UmA;؈d���������6�/&��Po׽�?����	�R����L�
O+��v��{y1���ӱɼw�%�:���/�1&���k��Ȅ�fVkN3cx��ʑ���e�0=�\/��g(|ɕ��mڢp���|oki>a2P<~�̀�N6$蓕�s�Z�s���(-��хb�H!�q+�t!����v�ٔKT��h�=�L������r������H�m�Y�o����O��@�[�*� �	)�
,Ydۧ7`c`N<#`HW[|v1u���o� >M~ی�t��ZM����|V�W��!ޒ/�T&���We�>�%=�?��Fҷ�Ѩ�7�r�:YI��}y(������jsۼP�5?D�:�HB��yq`] *Y_�sdK�'���Y:���T��SZ���ǎu	�l�#F ���RQ"���!�O)��.��w���*6͹�(x[A�V��u$�E�U]p&�J!����{%�f�1D�ߡ��^����,N��dl��{���_���z�^��z��.ul��-��^�v��2spɨL��{�ʐs��=���@��y�p��p4c9'�:�5H��Jx�S��|����Pg+�oy�̕�Y��
���AwsVsI�����4j�	;��¾�sJI�a63��ĭr��4޿`n��Y0Y���[:�Ss��j�n�h��]�_��a�LC��u6`�e�FN�����WrӘɪ�R����ߩ�m��O��U��L��[�U��f�`�e/�Q�C/���4�Ʉ]��ָ"�����VӇs/_�-[bA��w�����t��F�.��-49k���X�[����2�������;���ў������ّ�	�Y�/c���h���%;����e��r��y�?�?��Z���Dw�^h��V�.uc;�U��3j":�2��sS��Ԉ"���s*�I�bn�9�����Bjz�#l�)�Ns�)����j���|,iŽל�����ԍ1�����֡i��%��no�'�a�@>�2^���Z�0���{���*d����FS���3��R{��"'�uO�y�Ɓ���`z�0�})��8bƷ��%���9P��ķ|�Sb��&��<��x�R����e{���C��@�vT�%Ij�=�³�QR�Z�>{�?�NA�.Z#�䘁Ƽ�ko�"�;��у��MGޡ�K�.�k)cb�uƔ���U�m�&�6s���x���Wu�}����(�ae��OMξT�� ��5�W��q{:v��[�	�0"+0����s��A���KH/3@�d��1�
ҧ|g�h����VEi�Ds�M\�K�f�!	�~��?����U_by��IYȡ[I�Y���P��%������#�@y�MFl�bq��Z����)Ȗη��w�./��qf�t������q�ʼ��j?�:�Ո�ӊ����h]ۋ��C�,�������7����R��V,�菘��*�4:#מ��u3~�����LÛ.�,��~���0�P!���؜U�`	��(��v���wA5ݒr���e��*��,���m&�����~�t�߱œ��ɴz蜼Y~m…�#�������ն��y|��q9�+�,�3]�z�@'�q��"��?)?)����'����2=�	��n�g�0�6�C~���S�o� d�y�sS-�aoA�'��oY��(�6
���0�2��o}P�=:��CJ��u��\R�4�e��hy��2��0|JA�(պ�b;�.d^�,'^�ï�ԤC��k��xh����u�X���L�F�8�5�W� �E���d�vO�n#]�����h}?�JqYH@~3Y�ލ0*q��硢&����ǵ����N�Z q���ɧ�j�Pw�OF��n�Y�ߠ�%H=��?���]h���4l����ϸ�G�a�zon�V�#d�)nw�΋�n/�-������1���ي�<9(]w%��1�K5�u�9Ԟ���PߚU�����f��b˾�����㖄g��iL��g��?�-m1��5B@۹D<X�o��BY�;�Q�ߴdω��D���D�8�}��4������h5^�Nnc�����0NÁ��<�r�S�8=xL 'e@�F����*ne:�J}�Ѷa�����6�̔�=u��A�	�qv��Fb,���m�\�GV��`<?X(�+qd���Fԙ~� �쐇�o,��٤�iy�JG���j�i��Š�`��*Ens[��H!�?�kab5y�-���v���-+�1���Z�|�i"� �A�#���� A�z����m?���j��B����J�fL��6���x�>�n�����l����-rnhtu>(���9��yŽ�m�)/x�C�y���p�L����a�hN/i��G��指M���!�=Vq:��+��X�Ǔ�lᖏ�¤�2W�1�����+��_J�r�sLW��O�w���}r���.ik��#1^����/S^R�.�
B�+~�ݒ���3�뛌��jC����#^�a)F �i��S!��T8�}V�G��"���G�T���>)�4������3�'>�T�q�X���E�W["R���D+{�Tmפ]K�U=��d8�;o0�,��F<��mtJ����Go�����m��$�C����f���#{�,\��ݤ���_�b��b6+]5����Ql����s�BZ��>��'��r&�|2nR|����yU'�:���ѷ׶o�i/���D���`�X�d���n�c[���(����?��^k�S�`�+�V�;Ƴ��М�%�"�ߗc!ƥ� ֠�=�FqD�}��_�)r���?H�9~�L?�d� E�VkޫL}Y�X��{��3<x���Ђ�z�Q�SW(�A�$�<�u$��;[�J��\\���C�^n�F1*ᰯ�Ĵ N��_�iS��Rz��)�|#f�����iq���9�6Y�������W��ιkt�T�]F�s�����G�Y� ͱm��Iض���n?���h�A4�z��"��@,��-N������f�����9#�����W��٢����v�K|�Ț~'�B��%QI~ OA��<7zV"����9�Q(���H@���*�)��i�D�V�=�s��%�C><�@::meom��~�}$(�z��u_��IBxmN�n<@9a��c�/�*\*;�G7&+�S����M0;��#vw:��\�$֎)�E��U��U1�����t m�#�>��+�u�e'{���M��~�7��W>�%"�j��דR� r�U.v<��cW4��->u��A��:���g��Y�W������@
u)�l?]��^�yp���"�F@�@6##�2-��7^Y���/e��4jh#ٔl\��#�����[p<���Y���Q���S����lqLPٺ�ESȷmt���qJ���R�0I�cQjԝ�N_�����Bێ]��;N��ܗ��]�R�$���lmS�59�9�M;&�d\�2]:�8K�߲�����i�a#�3�x�Eƿ\��m�lu�����Ic��l���H%�`ː�=u9j�o3?(��{���|�u��&D�bI���2�<G �����.u��GD.�$#��h.���/8G'�}|�)O����}ق�ѺA��Uv�p����s>��x�e�XUd��׫�)��˱+=��^��>8���:��;�������Sao�y�˃f�Uu��'��Ҟ��A�Y�D� �ES3�����^
�ב�ZZ$�	8�>_uo ��9�-%�}ؑ&���ϛ8��y�pUe �^2�F.���x������~G�w5'nL�?�/M�*� ��X��ݰEm�������:>�
��j
�+ۅ�(Y�Do���}��sw)�og�V��:�千�@��2SQE��y�?�
u�I�)\}we�������ot� s+ᘫڱ9ĕv�¼u�i-�����(K���Ty���[��a2��:D���]ԛ���)ձ�b��e�7o��
O��N?$�]9<s��\����Ɋ�<[f���J�R��>�Q{r��� 6�~<#�S��o�T���sx�[3UI-H}If�v����usg{t����⤽�WnW�����<��#so�-�㦛Xz��F�� ��a��t��Mu�6����yi����sZ'�՟T��=���ю�_�~w� ݥ��^����/�'����x5�V%��ڱYzzU�Y��ݨ(n�Y�ZM*T���׭��|Y6�w7�\�/о��{*=�
��Wk�"�����
|����WN����̧/Si��o�B'��PHDAM�k�{�]w�(.�[ w�a��&�s�*73�{,$	��ĪY�� ��d�]�:��
͕1�r�>��9H�!��-ɍ8����\�:0��DXSҒ�Q����M=�=�Ab~Z,"4�KO�P�(tgn�D�KC���.�X���Xj�/�z�W����[ݐ��?��t�L��rO���
�1��jn J4#L��K)�cJ\��v?�6��GxB�R�V�'{?!�|k<�Qg���9��@ɞ-�/H��W@o:}Ģ|
��:��(*+�I�di�r`g�N�5df֌�	��I2m�k�ڤo����'y"����1�a1DV���=�O�}:�k��������D��gK�`�\�v��+��v�5�zK��=tau��T[ɃM?�9r��8�@9fz�T�k�7���_U��c蛧�lX���?���8�g�2�E��X���R
R>i����6�}n���Z�f}R"m` ��5���1��������skq��T�Tz�lt����"#��_�ج[��+��_,W�)��~j��D���G�do���6Wo��]˚emlln/z�6t�B	lC�Gi�I�kL͞�<�l�3�+��2y�Z��x����5�Z��a����b<��4~��o��[*�,����rȔu��O��ɱ�~�Cos�-_���;��wΟH��ϒ��p�w鿾����m�'�c]g��7�Q��0�s�Wt6�|Y������ݜ�ᢑs����?�2�dZ7��t���W8�]�~~�W�X��ۓ�y_Bɩ�(� s}��WwAF�o�0��;0 �UF�2��2W��~��h�r�<��� d��<��k����$�z�F��R�^�S��� 
�ZLhٮҏpd?��W.t>�u]s�JcQ���.�]��ݨ#�eB"�-��*�K����V簐=��o���g�)іl�Rv2��_��ː�9O���=�UX�e;�Z� Ț_V\S���%_V�	Y�bk��_��k}�펶�f�,;��ӎ��g%�����+��rr�x����G�kl9.?b*��-�)���5aM�GX��6�fujTw�v�j��9Jb�YPEz9ѓut�B����!�j����\.��g3.Pd6K惔�v�M�r/��}�Q��`z��A��v���<�L��T���Îg����5��y�]��A�'tt�) ��.(ȑ�A�RX7���~�%����[�_W���������1R��Q����vk�ONY�D�K�.�N�U@�����&�{ ��!����R�)���%
��F�j�?�����];,$�����!7Ws�Yl��ĥO%	Wo)$A�z�����}�
.�ƺ��9��g�j��Ag�=Zn�Y_,.�Y�k��&�H�6���b[L5n�7~�2 ������f�`�DĞn>g[�J'��M��`*ff��T�+T�-����n�Ǜ�ݸҰ^�7�U�m��\�Tݿ�ݓ�Y3}�1����&�ɫ�ޡ�4��%��7Ÿ�R��hj)"��G�Hq�*��Of���}񘓌���I�?Uw��G^�9Z�iW<���u� ��&Ul��ަ	����5�iUYQ�4Y�,�����?p��E����>)4���&ON��֞��*���y��uM�"���l^�Gm�a�:F�R�b�nE�}V�Q�q��HC�z���1���"�<Y�Ť3��3��8H�~Д9�L3��!6������2�k�.~`#��6��,�C�Թ��p3��7���C'4n�D��ޗ��1��e�	��-C�����4@>~s�c�|�,��M8.3о; 
� ��$�:ZHT[m��~�������D��s��:��>����"��{�*+���z�kp�`hP������Ёp�4��r���=���_ڣ�\��dk�+�!?�q�Fwq\Uv�~O0���g�u�6b�����L2W� �;V�r�x�"m+<nQe�|3A�cۀ�m�[��M0!��8�z�����]��.�An�� }iDɤ��L�m����ۭ�>�bu�����d�wßzd�WR�����FzvQ�H'��m� �R��$�zg\������7�c�$Ga�7��cn��u�|d��DD�2�;'@�"�i�Ƙ%�cɑ9ǎI��J�C����9��x������$h����6���S+�c�#��[�P��fGB"�"��Gv1�ے����5���<s�yN���S�$�c1��;{��ʎ<�^�����`������ݤbL �7�g�)Z��Q����`
�B��^v<�E^br��/�ei�M�ika�;�пҗF������)�G݌�kCQ�k�d"��������./�:���Ͽx���B+b��W���a/����¬�]��خ�{D�y@��I�}\��Og<�$$�{iCF�=�G�*�Z���;{��46Ica�NJ|>���Al.NV���a��M�}��T�;/	�:�gmq�~��(F�'�C
�!���;$�`�-
�i������w�%�4Q���ŏ�ng�ο/�Ή�)f5B�8of�1jHJP���1f�9Ϟ�1��0��(Y��7%�%*�-���iG&Rs�g?����5�L��ͻq�˧�6���Wj�Y"f��/��B/����I�J�2�b�����x(DR0XE��}�F9����^��$S�D� ��h��T��Ld���(x���Q58����Iv���iRM�s��֡�uk�F�=���4�����*
�����d�x�mz̒Q�CԮ�)n����VĬX��U�'��^���iE��;�d��af�7�ZŹ�{Z��F��dSvW��e"!�\Ŝ��[M��-{�;� ��Q����{ۻ���=���5�7|�¼�Bs�;����k͇�d$K
8-s�8�J�mR�l���b�q*�W<�O��=?��cx&M�>�ӖE�Q��UCl�'J�2�\x��o�9���.L��p�2����B1���p�]3�'l���A�C}H7o���lݝm_nBب�&SMݯ00��*��:�s�`Λ�}�&�֠�����&�l>6p[7p#G��j���*k�-J�mvYI˽(���qf c��9�l�L5�0�<�^N-����^�&����Y����m���s������9Kчn����ԃ>j�y����?�%�� ���{�uT=g	9a�yK����Q�m�����c���ܺ�����ʘ��C;&��w!���^����f���oB��O�0;�eͯ�'�t��Z�E��������Z�\��������@I"a*��Vz0���3h�u�������L��Z �Jp[��'W�k��[��Uo�A�c�x����35��JӚ?r�%|]����ʹl7w�;�7�����^��6�&��%k�U'|%6��R;��H��8�����a��%G6�7G��a��q��ַ�D�����ހ�����,/�U^|޳r�9��w%�� ���5z2�z§k�\[$���R?.������q��^�tR����x�b�%�tj���v��9[��)��R82+���^rU�o%���x$ �Qa��\�����X=vc�ʬ����V����.���ﴺ�vK*��=�XhO�I�o<��9�����nx���Y}��fnq)<�֬
�N����of����ֈ��x(��y��ԫ;�
����|�e-��&$%��x���>�ͦ*iʳ�Uo��O
ގ��v��Ļ����#Yb�;��TF��6y�������2���l��%�o@SW����%��	�|j�Z"�%)2��4���'�n��>��ʷ��m/�����b:r�կT���?���#���Y.�}y��(�cq���X��]����V/����-�6띺�� ����rګ�Wt��H���fʓHT/|��དƮx�u���K���a{8���kw|��L��Hs����J�����=��V��Bj&!�U�"�����`�G%�4C;F��2X���j{o�7@���7�D���VV%Qg���PP���lA��Na0�a�*��&Eb������1�̔.1mK`⻥�}�JI��%�/l�߿4��tvv��O�K��xe�YF(�4#�۝kk{-1$�9��-�W�3{�+��q�.jɏA&IY�#�j���°���VÉ_zE�l��@	�i�e�wJ��j�Y9#v%�M��QV�W\D3,Tx Wf�6�������㠿���V	�b1�nM~z�������C��F��jt�	N-d��J��£�ڏ�a#��+��h>�v���nR�"���!V����]h5��l�R������_���^W�͓>ޞ��Wuͥ>����9m����k���3
��O�&!D���=��׻!m����Y��n� y���w���Z�$�x^��C�����j�ջ7����Cg�9L�8VN<[e_f �)~�O?�Cu�P�@)$�@v��q�̦u�i�����bT~��E)����+U�.��;�A~ٿ'mS�,���{?���ΦG���F�R}�tT�l�+TIad�qϓ �&���W#G��jf8u�=$	��QO�OQ�������7����`�[V�����不:�|�^t���iW50F3QIvHZB��Θ�j���^�%�Z��edI�v��D���$r�D,�@\�q�U��m=�����$�D�o������osh��F��u����(9���b�Q���b���!I`x8��R�+��7#����>O�8<YH��Vq����`�[qpKT2���R}���Y~��{>����]�ZR^C��ylmV�n��-�jt�53��Ӭ�0�J�#c|&$�������/�X�����'����|֖�n���ߐL'�p.�DW_D�bhh���V�Q����t�I�K�5����"=�%&MIaW�Ĕpi����	�~���� Us���/cG�b�i�4��/h/�	�]�Rд�#�� ��o_ �
��q��m�8?֓A45��>S�,N��)^��At�� J���ɡ��Ag��֯|cA���{/�������t<���|���Ib��j[\�VP}#-@�IBRJO��Ƭj��􇊿�a�x.D����Z ��5	u/A��t���l��[ɦ�\_mO�RJjv�T2Я��x���ͧ+2���xR�����ӆ���kG7Ė��`�@ ܄O�&L?�Ȓ�n϶���j6뵤� �_˶�_��gX?)d%k.u��$��Ծf�_���]�'|��;���J� � J3�7FQ�����<� �:�}���HԷ���@
6��|�bΦj�4].J|�:��=�.�铴y�%�s ^�
���@#(���Y219&�8�Q�/���Ʃ����y,^�/�S:�o�t��k�����2�h&�Z{��)ڣ�&
�u�|GLn��Y�����^��>�&���sS
�;�3puiqL/e|]EvC�`E�'� 8��[v~� �[�P'�5�gK�(��y�����95���pS��	�M � '-�'��|��G�D�p6�:M�����0V�b^]�*�/0F�l�����X���~%p�I���-oG|)��V��N��J^l�8 ��G�K��C��	 ��������1��QMa��t2�5 k⫞�{�t"�7�!�a��"�d�.;SR�����	�4׮��!V��A{����4�ً��y&������'��z��U��,�o��:�PHxl�z]��Dl�9�[��fr���������=�G�b3&2�&�)Q$$2�G�=ҷ4 �r��G&�������b�c|l�4�w�z������vi���N읆3`x<"+�1���3]mm6k�'|U$-���yg��C��"F�~�������<��_�B󴾱O�ATP�y���V��{�׵T^Q�WּǍ�LQ��ˑh1�`_Y�hn���O�_>k�ɶ��{��<��+d��g�̥�~�z���R�/ֳ�z���:��G���6�(d���J��*����R�8���L�|N9c��(���*�i��w�*���}�&n�i���k�4Ã�eg��O����l�����:���'�}r���N$��@��{\�/_���	�,�Z��c<Cm��ƥ��0H��m2�w�;B"�(u����w�P���f+7���I�nƙյMO��<f�Պ9���̂��n6�Ȭ9t��j��J�9H]J�8�� ��nBC]v.�!]9f��~����>Lҟ�$`��{�\eS-D�G��˶���xTc�8"�]�!�	�`�ޙ�4T���um�Qa�p2�����I;�L�űW�8�X]�v���\׌��z�;�|V�h�<m����J�i�ç2ό��X��%f�/��l7�������%"[�w�<���������T���-j�8d�.n��ӉeGΣ��ˋ7��������Y�{���"��:�����H��.���~��E��hgХ�@y|ܓ1j㊹��� ���Uwce�>�7cW��ϗҕ�jF`��n���>�䂪�M�ɬ?��̭Z<e6O'ビT������]���Y?1w�\v���j:�cg ����Z{I㼱+U�K�y�|9nS6뭉��b�0�_$��ay)Q� ����N7���ͳ��܎��%��|Mi&���fZ���=�ɽ����(��ö����e������	�ts�p��$�}3@Fw��>v�T�R�hY��>�1^�@Vrc��6V�3y���qԋ6����i}<�}֘�W5i���!���b����:5=�y;3zw�,s��L�K�hS���.9�{���\��U�'M�R�����A���G�OP�vR�����W���|��?{�A�f�We����W���\^�~߃�m��06��_ ������iV>��j���;3jW�3��ޒ%��zk���'9d�Q��XR����C��&W��B/���B��|8B�����KG_j�'l����ͻN\p�m8����V�����5����[�����Q�̢&���陮�p�}s+|��Yi��^���I��T�

JfO�*4�v���<�� �Ŷo������л������{QYU����`1k /sc��p�VX]�{�We�F�_�('�O��s��vF#�ȹ.����
\�T�i��垟�Hz��3����#�nۍQ�D��	���}�I"��vv/��o�g�K��6���i��$�Òf��f��:O�� �,��R��uށ���y<^��v�@��"~ƿ��%���C��t����L�*#��}�� ��[0�z����3},)L��_��F��5@m�-lW��1"�E;�_�H���uPK� �K��8]��U��� a�Yi%[�:��z���^%�$ڎ;x�S����w�y��uJL��l�O��)ƞ�L,Oj���c7�Ze)~q`H�޹�)>����e�G��7뾜�a��\�S}]�4*)�x��0�^�����4u0�D-l��W煼(�y�5����a�����*@"x�&��P�+���<gg�H�٬�O�WY�ͷɕ�������V�����d2>�β
�p�9IR�^����� I�i�'Dw5�P�P%4У�[)�2�}�:��'�%~�׀fOm���]*��'��Ӆ��S�Y5s���#�X.��R������=v%�͟�2�e�vQ'��{�
�Yq��-�_�C��qNGW�\��f(�3b�/��������s��B;���?�P6;��V��V�c�׫<�+Y/��δ	)�!8->IR�c� �e���D�T�� Խ]oX��/��a�t��:�J�j�p�6������nN ����e&(�g'? [�8g��w��B��R�r�4�)4��W�m
�1~���f����U���?M�ɔ}���N�RU���}����4�H�)���������:+ŏ�����ծ��Q<�Mv����8,��B���r�)B{}���������9Z����^eU�����Y�M�g��������ᗱכ2��b���oX��Q�S�X�A���}�������aT��ď�p��
�
��N�/�x��6��48'$ܫ�Q<4��B�0t�tg9�-`�ځK� ;�W?;�2^��"��GdF�f��B�I��J���T�*+}���1�Q>���H�t�,%�� Hww-!Jw,%�� ݝ��)��twו��Ͻ��9�<s�}ϙڳꔶ�[>���V�<j]tJ4�>����4��w=�%0z��;�B�Sd�5h�|e�sd�������U���gh���pVkCn{��2~�|<��,�Te-��$9�b��gXa�"CVW�����*���:f�$n�S�FI��+�3O1M�ڂi��4|�ƅ'�ur>(k B4��9�qP�;_�48)��Sxt�[�9-�T
/�����W%�M1�������[@�Rױ�C���L��S4�[�w��Ѧ�& �}��!0ԴbYM�k�9���}��^�,��7�_%�]��"�"�q�^�����9�S+)u��d�����o�޺�h�vm�G� �㫿E�~����	�K��o\��B��'����L1�� ��o��{o�(ހ�;Hm�!~�&bd�٧��`�׻���t��v�i��W6��H��(1����yn�xd�mK�=~���uk�X1.�S���I���E^�Q��㐖^6xW�8T�v�qq��\��u�C�����n@{Ϋ/pw���X�vg�'q W҆g��0T���3������ٞ2�MR����#��)�N�O=�C,z��Gl6���g":�;�x1�������]ܼ���pk'�]�|�.��\�w��
���FFF;�G'�Oڢ����=#�XI�ׅ�j5���j�mx�j�fDT%Z9Q~�(���Y�����g�`0��p�Atm%���x�y�u���I��ʟ�򶵿���d/���'3���V�����y$�?8ͅ4��[�A���V��9ZE��6S-��1���`t[*�9x�\zqp��{��d}��bʣ?�Q�R^�B*B뺕�1t�B�`�ޗfI}���o�X]֠m�v�����	�8�\��M!���^�\��u�",�J~�E3�Uiԋ�+mkQ~�^�<��_���� �/�۟�J�35�|��e�\�9�:�����hne�=��(|BBd�%��`\��H�s�ؤ'�̧.��M��k@�V��f�A9ǴC�]xY���'RL�i�mM3 ���tt�˯��F��L|4%c�=�����Y�ͪ���~/Bi���&?�]�Z�]!g��El��6	-�Nf~�w{��������,�@">mO�^����.md�B��N� � �r�X�QS#`(����.�|��	$��=t,�e�p�#��j� E�}g���Blx��y�3����׽�h�������(��sd}(��L@u���T"����O��_��̌�}��#��5���Gmb��"ћ�մ�Ӵ%`4�d�d����G1���JQ=��d�=֠����x�,`��_H����>tߡ�c*�|+vF<�)pR	{y
~u$*2�q�Pp��!_����#ݪ2)�H���ڏ��)�D�)�	q�|h�uBK�Ss/�z�pRH.�C�F����B%uM�F��U�x�]��K���`9dJj�Bk,W�¦�����oz�/�8c�-/�暋g��5!�a���pb��q�?�yW˱���(�M�!�>c�����Y�S�udܨ��1���;�~W���Vٲ�
�벥��e�B��%F CLE"S�ZT!t��D� �r ��zHg�9h�B�z�`�,�<2��Ģ�����8��b��0�~2�L�B�����Ot�me�e�+-%v��r�jkP�iA�eNa��������HO�ɖ��]W?i��/��������d�~�l/�j��y%|̜yR������+�gyM(�'xP��w���>oZ\^�.��,��If1�KE6n�q.�iS����̫D���/����x����<}e�߻Rp��8����$I	�����O��	�����3Xӗ��k0��6t�6�+U?_M�����%CmOO���*�|�7t���|�5Bh�e�ɩP�H� -��eJR}}��L��;@.l��1(����yS��e\��<�c7���A`j��E���!lPF�ԩr��;<������,�dI�r�4�٣�N�=)�7�[x�.p�o���x3��'�^���{zэʭ���PU��\����2�s�� �35�;c
����FF×��̼B�]vs/�O���o�81��a�x�w,8��D�w����gc0�����'~/�
�!�]��r��P��j,'<���X>��=vs������+���(^˝ �^��|KY`"j�I轰�C��w�Q�=�^�@��U/�lSR7�+�t{+���5]S���&p��Y[����I"�s���/�?ye�<��[��ӽ�$��FM�6�	�\��)���`7(R���D-���8Xrm��X�A�2�&�u�ז��&�Ğ���\���%�������g���"ed��v�P����^.}��Ʀ�.�
���_��gƟ�Ov7���ޮn=�a+\��%� mm�9A�0��0�U��c㒂�6v�h('�����)/���E)N�_ڱ�"���.�� ��"l�9�wb������ JQw�����2���o�R��,/y�T-+�Nd�'��R��;�Hwi�����>�2Ƥ��7�dA?R�9Y�(ħ� �n���-~��}
���nz�|b�!��B�~�4	�r8g.��Z �*��!�����/�I�N��#��.���hۀ�s��x�C� �mԇ�y{�	7�M'c�˂���7%�%E�a�N�	c�zΞhx}:�B����\�SY(��k2��{|߀7(L�7�d�,�r���W������y$��˂��`���o\|x��]f#���d�zٓ|O.Ѡ�p�_�˨~A)��]t){���c>�d� M'��X坂���#�C��V�oL��b8���8�"��g�I���b�!�'�;=۶]�	S����w�&h��Β+���U�X�����Qǔ�g:s_H�|��<���i�1����p�g��#��<��Af�$"��5/%�=k.� 3�2z?Jj�X���M	-�R&�r��LԺ)]
E>_��_A?DiOtM��nSR��u�q��@���Ss�4�&���x/�y���|I4���W��1S�GB@�W�`%�����M�H!��wY�|fQE[���ͅ!7�'�w��򋣋�[|�xNy8U�3�K���;m�����A�A��\^�T��N�e�>T-'m=h���MG�$U�@���Oƒ&���._��P$5}WC"�t���#�������J`��FlX��Ө�`���}	��(��� 8��;�.���1^�o��ʡ���ts��u[^���׉Gx�*b�ЎƩj&gq�\d����DBaz��#w��u�/��׭01Gտޮ�4�m��}���AG�g-)Bǲ6�HY�nh�He��r��+�~���Q�9��DQ�z0�O�s���2%����cY��P��_iZ9��5��䉮��[Z��3xQ� �dٍ��}D��5!�M6�P-'�/~&����N;�2��� v&>wk�-�~��b\|'M�������&MVYQN��(�)r�3�>:B�5�,O�M��o�pX�xOZ C�4�x(�Y�$�o�7Vh�[�G,tw�c���t��5[�s�B��7�h ���<I?4/uٕ�-���Ŧ�ك8�%�M,J��זJ/��B�T>��@��R��:-yI�E�<�x\#�!5ܚ$|/ �)�����6S��>w� ~w��}�SǠ<��R`�^�Z!�=�y_��:�z���ǔO:P�Y�F{�-ֆr��7Y�a��<�]bQ�KĖ�_�� 3k��\��
r[+}�����Q����{Ze	���#��)�e�?�2�/Q���k���F�%2�L����GU�m�e���`�q��R�e,��.^��&���4���t�������}������ (?f�V�g|o��d�{�2�Lvr�mp%�^���O{E_.>�)@a��ј���w���0�߂���Ͳu!� yf%���%�8&�G�?���~{2ͽ@�"��D��UC�0e9T�$��nf�V�u�~ �$&a� Ι����;}���')i�?��~B�ʹYT� ���L��v�\4��'0�!7��8љy�f{�aN���>����5{Nk�Q���1�P��Z%��FM|��;�F��p)մ^=����=5]Lkg�NY��r���P���<�]��P�q]����h�%Dh�:#�5�P���"0���A�/t�DMp٬|$E��\$��k-�jx���2dh�ΰr
�ȶM�*�iwR`���#TךX�����u�욙M@���j��vұ�W�&XNT�Kݵ����. � �0i��R^�2���d�?Ѫ3Y��-b.�B��F7tI��v/fMC�ݹ��������Y�A9���u�v�-�?�W�J�P�����l1:�$�75
e�o�~a��O�V�ϓd����Ͻ;+�&�;Ikԩ�:�%$k5R�L�I��b��;0+�bحd��~|�4��`��� �zԲ�g]"D�!�`��yp��4i�E��y�$'�Ir�;p:���=��$h���M�D�5D�گ�(JL*�I��SԚό&T�pP�v��WbNvPP�B͇|u::rƁ+����X0c^�d��W"�'��F�	���?�d6�P��"�u4���d���E�,@���j���%�&N�tp��oP��}���u��:�5��!2��"�+m>��2\����~�X�	l&w�{��m�1@�u����Bg�+�cLҸKT�x�;	���sDo�����r&�lP��Q����3�>�sR���3"�J��)���;f�=�B;LXD���^����)p!���g�Rj_��֝L
�e���g�,�%VzS7,A���z5�k�`|�����/Q\����I���%��HX�Q�BV����;v����{��]�)��?���0��*��~��x�7Іm�u����{3��G82J��C�_,�ֱ-�AZ'=�KR�U#�B_g��gJ0����E�ꚇ��aU(�^���o�]*I�@E��9�&p��1Θ�ꉫ��1�I�o����ќ	" ��0���ߙ$�-}' ��:��>dF�����<p�� \�N�U4���N����;��u���V2p�Q�u� }�n=�5��)-��ƺ���sN��� l�����E�T0w��^s�Q���l����%9Z�ݎ����%u؅�1�'\&q��8���|���Wf;�F�$���fG֬�i��߬����������:@Q��{�&}��~�w���b��X�8j������'��4M��,s^�FB�tg.וZ��r�;'e���H��,}��4�w�x��L��*�a�Ŗ��ܛo�M�]�JxC���
�k�����+�H>�@�b~t��#h%�yL��A�ʒ��	��_����Y�<�j��N��_� ���^!Q:�6���z��E�h�af�]��B*1!�{�n�xZo3�m_X����O��d��=^;���+e0��K[c-<���E���F�=P�Z<o߭�~C��1j�`<�
����b�&�nb��w�Ø����J��Z]�C7j�����Njhd�����7N7����$y���.;��ۮ��Vō��A��.�Q�=��G��	��[5���~���e)�-�\�g:=�k0�{c�v|o��wj�r��(J���
L߸�N���GK� �����R5($Ug�� �(��f�c����3��X�L5��mm�6]k~�6q؋`��rT���?�٣Ǘ��k���NCONni�D��/�rK���lKa�*M�l
2О�bi.�k�d�b�{{�#�Ծ�B��
��4��P�O(!�$�z���_B�5g���ϲ���N�%���F�üA_Yu�ct�tD�s�_=�:9�2:�`��￡�4�{hFL���$s	C|{�^Lgm�����N�G�]�U-�~:�5��u||���)��_�\"�w��faW���C����7�4�:'�_pf��%�AK�B��	��;y��cc��e����GU�%���Z��[�W�l}�Ė%��#�.���y/6ӈ��
��4��t�v��X�_���nc6Eӽp#���Ip��֞\��lƷ����Mw�H�
�@�F�w���M�s �T���O�5q�GS����Mf�MB���|GГ]�;,��W������$]���Lz$�@��JG�H����
�o��?
F8~!�s9E��D���#�R�%�a6�\	�$�.��U^�S�����(���% ܈�4*�<�pj�=/؃HD��_�r?>��Y2�1��7���o8���X�;�/f	z������ëx�gr�����!��ݯ�N΃8���5]�?s�ł��=����F���B�9h�g��I��Į,�"�ʐ���*6ª(��r߿��!�6�y��D� j��G���C�Q�q�56ݦ2��;����~����m!�?받��t'R]���Eq�G_�[�6�b�'3;��wv��ʎg�h�Yc�N��q��&3ݮ�V��{B���-D�W W<���Ig3�y�����H|Ww��wW� c�T��5Q��M`4��b���G�e�������$�1�z�PN_�*�s|CEVsL3wP��ϳq�3���u�`����
q�z̭��qx�Çm�@$ �i�t=�-�����r��BW��wQ��"B��	�xZ���|v]tL�~��=�rҳ��u����ݬ26@�Z���A��w'�cB��f&k8Ͽ_n��J�0�Zh9�9#�c:2��_��gOlN��~X�!o;ᇸ�OCv͓���3p�Gi���R�/f���`��,�d2�=��k�[���/v����x�)P�Mx��AB�b��p�9��j�����ş��Q�*�q5�(��]�_'��gF���c��<�v�>l�w߀.Q� ��B�Aw�/�״���?��~N:�w�|�;��à_*}�z���}��T$J���J�L*�\}�z-~��o�:��	�!�Q��.��$�~�	���K��*�ՇG{K�B&�j	@R�5��o��~�-��q|�q��C����k���}PL]̆<�d��̂@)!��Z�Q5F�/qQ!D�5�+C =�X�n�����o��;����Q��9�I��� iī�
!J�̢ts�M ɕ<�J�giR�㎒��S��(��f���h����>�.$��|�:��\Lr�MA��;Ŵd<�]�R�]v:��xjC�`
&���5k�4��.�y
�r��-nYզ��+$f��$"^8^��#�i^�b\ w D�Ùsrn�#uU�n�Exc���P���D��xpyy9 K�Ӭts��ApS{�+�NW,,gj3���*���m`�BXl#��CTZ��ް\z`�Y����`�4�#�A1����+|ñ��Y�����-�?�H״34���|��������8x&8�	���_�aXz�kg��҂b����P6N\fC`y��m��7�c�We?P����C��CU:�MêW��f��g4\Јfy�[d��̍G�E^��&�_e^n��x�`���2g�o4�̫�)������1jS�sQ��p��K��.��a��F��>�̤��o0��r*��C:�=M��p�	��b��O��V��W{��\������N�mJ�-#�.[�zF�8��Kl!���?����Z�f>�]���v�3gv��{#�Uh�+����c�?�ň�1*o:M��.H����Y��uF(�V��-%��W�K�%˛����{�y�<���6mU-��8
�5|��R�����c6y�N ���LƎ�Fn�p������]��L2��,��6��	�upcEjk�����G��n�`�i]�(�^��~w���W��E�;k9+�h�+IT�b��G�zLȗx���� �&�.=���
�+�c�5�;�pEJ���T+N�����r�����E)orL:��ر����.c���H�7�/��5��\�%c�)���&�d���L޿�B@��A���#�^��u���r*<0H�iW�l�������6#2��(S>�j[���0�Fyn�ە���S�],>���ZN�,A*��0y���Lk`��+r���*���h�&���Y��b��j64��_��.�C�@L���$�r6ueD����-J<��m�a��-[�EJc��b�bo�+R9g;~�ͤp�k�q4�R�[��um�>�ǡ���AX��������y��N�V[�i��$���1�+�����u�S$J<���~!$�J�̋�E��<A��K�4`(�p��8��;������v�[�#Sӂ���Y�"Y���݊�q�~K{��_��]]��G�b�5K�lvS��{{����'����N�i�r;.PZ�<�n��M�#����-�v�W�a� ���Q��3Y@6��D���`�r�ۻQ�E�m�h��U2��9w�c��n��f�l�'�d��y,#m�B��t��NN���
�F���vf���b4dx�k~�?+�*ޣ[�#�XW�@�Ĉ�qDG�y��o��ģ�_���7���!e�8I>���]$,��kU�<K�遶��-��Q�2JA% 6�\��ZE/��e��������"�AG�<�+j��O���M�.���rב���$�����Fڝ�*'�d|��+���p���)O���z���ڒUɅ1v����'U�ve$=��<e���,��
b�;%e�Q ��$f;:Y����x�6�Ut�nn��q��P�1X����[^O��)��PIVi��G5*̽7��s��q)�h���HTI��]_7�q!��_�i�v�<I���d�0�{�b9Fi&�<�=���C'�nU�ޔ
�#�S�j�?;o����@FT'�#泞���1%��߸8��s�6�<�֨X��s��a�&�Ʀ?ߴ!�x��J���Xe����=�Z�����x������ k��Z��Ԑ�s�z��&�a	R(���:�~� �WY5�)�Eʇ�����rm�ȓ��L_u�Ǟ�G?3�,��$���~�n�Mt1ϫO��:5��*
�5�o��2|��y�P@B�����q�|8����tK�櫫m(-I�m��
����\fJ�1|�3O��7)��坅���1�@F���8*XͯןĩL3�œ��uǷ�a��G|9�*9�ENaկ�3��ڨ����-?�sI�NV[�c��t_.�_$��.?0�i��H�]�+�qE�5�c�a��e�a!Ä�EX��5I�����mZ�f#6ժ��q�/NET�xs��Xw����?l�8+����yK����D�h]�MM-�/N��QM��&��SI��-�v�낼�����ë��[n���>wԎ���/.�3~vD�5a��&�/i8RnCЈ�Gu�����xHj�6��=c�o:x��qw}}��4q��k@fڕv��k�(�\��E�?{L�nh�eo0�3�R>���jY��hDL����J;�zK_��H�(KY3�L��zcS�PU{ �Àvy��t�i�����<������`V���� L�/�J�9Yn\^(_N% Q���E�1�הKM��dM�H�5�Y��ɋ7p��x�b�b�4��0\��67�І׈D��U��^\���.^������ݱ��������o������oh��@{�.��9���/aA
�ƶ�I��:%�Il�ge���4A�|)���G�_>:zA1�A��N/%����Kz�N$P&�|�SQJ�ix�X�K2��_'�Y��j�!]�����L�c�T�)�(tߞ20ՋBk��P��ܩI��l����HڔLʃ���ZZ���b������[��4ԘU�� O�t�Py���s��K�'y���X���T�x"x�Δ��ّ	��&��B���Ć_[���FY�`��a�#������ڕiJ	�/�v���aO[#�v�qM�����ѵ1�UKH��d��А���tө9\���{�d��T��N�O�Xq���{#�įp��r�������/�>q�w�Q�\��j6v�ܨ��]UF�H�=�'��T��!�Soe�E��H�pW .�z\���,�2�xKh��-��~�nK>'���c3B-�τ�ީ�@�M����ݡ���Z{l%�� ���<?���SO*��銰]E�%�򋲠��Ѓ�:��O��E�vđ�Y�E��,I��>f�|�#���=���`1����$@�)`�F��E����߅>k����b���)���z�%�ĥ[�ZX�CF3���ȗ$�g"/ܗn�Q�R,�����E�\�Q��i������b���vKn5�(��2������ĴP��ծЫn�C�2Yڋ]�b�^��,�L�#	(̞+���8V�b6�ᯉ����!��'��	�͂�zb۟8-jJa0�\��50�H�N]�]D����������4_���N�e}���~`�6Cv��^,ƙ��ͤqa�f�$�eʺ)���W���.ؗ�7�W�o�����j���SO3��6���-LDr���Y{(�2�`ήi��TK,7꾴�s���2�9o�p�V�~V;lF�A�A0�yR,�"7tn�y��⊅6`�Cx�76-�R�Ȏ��}ĭ�j \�l���]�3]���Ķٯ�����q7�.�m�O����W��!\mޢ���v��Ժ&l�lM��?��7�m��?)C�;>��6�,"�&�1{�m�/�{���ԙ������h���/�#h�a��7Z�s��~U�aK�7꼢����H�C������y ��Ṹ��M���m�$ +�-��j��j����q�X2�z���_*������}a=��
_b4��ۨE�6��>���G�����G�se���9U~�FҴ���m_�5��H^�3��J����$�0�q�~Ghm}'V�cH�~gk٬@�g��x���X�����I��r�%ӷ-��'H��O]ґ��g�y��g���~5�e��Z�L�ms�b�H��:tԃktA����7v�+��G�[�n��m�x[[ÿmS����!��|��/�*^G�Wy�=�f�T[�4u����1e�d���:Ovw?��j�� ����;u����Mœ��\ʋx�����h�kݺne��G|���3w�;Bғb�4��7)�[���ݡ;�ڹ֋���wp��]HƁ�t�M��54�-^�/���_��:l�8�b�G���O?S����.4�c��h}�w#�.�|��ᐶў��_��v|���ޗx�G�DK�_�rgd����T�	��A��2���#g^��H���+�Qw�d� ?�Y��S��uЗXAG�-�����R���$�/�M�w�� gm�+=���q�^.d���f��waC޸�U=�:��3��Y�|Ķ�_�qb�G I#@�vsN=�#k�b��lB���ur���&���1� ^ʣ���k8��4��~�<p�u��߱��k��O�R�HB��>�}��ZP��^ߙ�J������,N#��?����.�g��yx�&�$�с���.?�(+}G_jDq7�~��'���$�z��ğa\�l�:������n�o�I?�S�d~�)�+؄ܽ�8U����C%��F����8jsM��7�✌hݯ�|�в{����i�o�ה�ɨMw8�+��Gy��~P�Ju�����̂�nȷ�v��)�^�ڢ4pT�{�GH_��ߢw�/w�5�)"԰�Oym�)���yX�u���̵�es��H���/@��h̅�˻�̻LƟ��uu�aV����M�L��'7v�[z�ͺ����!Q�9��Z<<�(�M�T�^�~��8dR�q���!˃5֨�;Ճ�i�&���}4�`�_��N�ђ2�*%F/�'%���K�i�~_�=�ͩ�]��-K4�Xْc�v�wB$�7&H��?�N}�?�Ues�(�w&~0�� �� ��O��tj�)��ac��&,��;�b;�YE��8���uC���G;Ҟ2���
���'�dF��Ծ����O?���B�A����0����ŽÜ��$ĩ��g[�xL��[wl����s�ӽӳ_c[�)��oo��3���HU^�k46=WY뮧'V�Iy�c�[�����yq�OZ|��m3�3�ZM�9��@*|C����=�V���p����/��~���#�=mŜ��+��Ͻ�s���QI���kRh�i�&��#���^~�f&���Ab�o��V2�GUh�H��'U����?��������[b����z�J��$D�����1�{��������(2�v����oD������AO�χ�������V��	V�y_��[Ƅn��#��^�	��s���u]��n�ڸ/x�/�q���?�(���4�f�uѲ�a�����03�����U珖:�!�;[�۲-���������?U!*IYSꮆ��S�c��/��C"�q�m�_L�2��JT�=�p6�c}����O��Z=k�4)-[0B0����>	�fa�8�3���l`v��jOZ/����l7PX<z<���_��?y7>����>ε]�)�ïI؈6x��p����N�w�>����q���ġ�GƭY�����E�V��O2��4�T��'�'��9���z����t2����m\�y�{�r�0�u���4m|�yo�X֤����9�����?+/���?�iON�ՖS�ȯ�`�w�÷*K#*���4g۝�o%�*���ڂ�:�~=O2�܏������T��8��Ժ��WQ��򀈨7�]^]!M������M�ؕ 8�yh/ J��/I���i]�zlb�-`�+�O���`����[��\�?T��bү�0u�sۆ��$כ��f|�RJ����6��^��r��937���h�^���rY3@�^x����w������xX=l��tó�n�2��p�O{&i!�X�O���쉆)���cB�i���,��&�(X'��F]�ᚨ���Y��B5}1b��7$��n�{g�.�DKհR��?xc9U��
x7�ڧ���*ȩf�����X�D՟ti�g���>/��1Ոt���y@v�0-t
{�i�(��Ћm��CSy��F��| ���ρe�Y�#֙��v�aO�R����%��zP��Hj����P������/@����П:���)�����+Zo�*�M�(-^�L�e(��7�S��-�_oұ,��55S��3��0��ܼ���M8j����N��*�5�Q����H���ǿ=l��%��v��g���"��ǣ o���Z}���GAf��'�\K�`����8�W�q=�욕E,�3�_�T=���NfZ$3j���i��z0���T�Y�pb�%8�%����2Ꮁ�it�f��<�&$t�m��U�Q@�3!�E,of>i=7��h֊ih�S�RxМ��Y�����Z��n��BD����Hi]Iǒ������c�1��QA��!�П�� M���7������R��2�/��_�l�$s6M&�O�1u,�|����|�暥��Q�D���남Qa�޹�0��11w0G�+R�Y�f���6���ᗞ���[r7�J%IN�7��gaǣ0�!��
��K�O���:gbk����P-b��H�x���c�,��q����mBA]�^D�׎�t��w��"�v���d�ϳ��Rz�F����s�o��״	��?�����مJn��5���<�/��.L� )�Ҳ^%�P+f
�^���G{]
�2\�d��<��^x�:>t���M��кD1iMB���:��UC�Sr��oS�:*���U�If�p(0CLy;ܪn��|J#�vԘ[Zv���E[���PT���/�G8x��!5�E7�q�(���\�:�Mgp������ᷟ�s4��;�
�����^��;6t8�؏���w�j_8��`���๐!�>���q�V��x��Q>��u�0��L/.ӊ�%��&����o��Ga��Ay_F�����!��Jn�5܈e�=���/J�cy"���,,����R��q>�B��e���bg�v�An��x���W�mS�DZ�}�0�^I?9
y��hX�O�Niz[7�57$��1�z/���`N�b�[������K�J���6ZN�]\1��!��@��?n���[6.�����"cn�ς�KE�v6V�G��E
l1�7t<�*��=Ng>�W- ���}0�(�oe��I\F�,3�дN�G�"���+*�ɥ>� Be~$��sf,۹@�����;����GS+{���+l��$�<�Q�I���ա���9��/;�i���q]!;���U-��%lZoJ�`M��E��灴^�����6Ϯ#�������v�$Q�4��ZS��j���H����)�Ȱ�s
��i������@�؊i|[�Ѷ�I���������H=薺����w����g�����Uێ�!W����w4R(�x���01��1�S���7P�q���Z�	�i�H�m�-x�o��"Q�
��Z�6���C�/�k��շ^��O�ຘa(�Bri��.}����BD 'w�M�m�_V�;��w�0���������W�I�-b�1#v��<Rz\ִ��J��eUβ����9n�����v2Y�7�-�1�keҾUC���wK��^��~Q�Тe��'?
��˃?//�u��Vha̒�!�q[��Jz��6�]��Pr$_X�����48l|�(����
�E$�>��0��k
��1��ֵA�\���g��Q�S�5pS�����͎�������NA�C7�SG�]v���TH֒�`�|�%�,���4�\���O�A,��4�}�M�q_W�o�w�k��#�
w�����Ts�tXͮa�߆�X)�n��r�xXٞ<����jg�<��{�Qۯ�U셾��������<D��B�B�jYU��`�k��w?��;�U�{�b��vǤhג�
��0����_H�3�SA�[@��JH�)����e�>U�:��)f\���/�"�mF�46`8�T>���^Wt��\�H��N6CV<Xf�j��x��a����5D!��|���*�)Ks��	yC]C�Zr|�P#��n:�x�6��q���*�UEZYϽ��-������j͊BD�-<�2�!�p�ꦞ�m'��1Z�q�L��W�㯉Cow���-�^��au��M��xeR]�;�{��N�r7�u��#����_�>�V�p�^�X>`D��,\�\4g+5�cmg��*K�$�}@*��W��R��q	}}M��u`gi��&&#��~s�r�+{��G���(�T�������y�u'��?�a-M�Q����TT�.��.e;�cx���Y���ՅEX�`�H�}���� /�U�\SP��3�sV�n-���X�ɢ�UU����P�����|��:������}����죷r��_s��7~8a�>��K�+~��	�X����z3�zRQ�QSeu�V�X�k�#V�U)������j�|�����o	�S4N�~�Ί�#aO��(I������9�;yZ��6���$�t��d΋�_�N-fA�T���=���X-Z�&�[�2�H�ot�Sa� 8Փ9 �>�����_��_ ~Y�Ƹ>�Jդ�JO�Y&��>�����QOM������f��;�L>�h�w�iS-��&N�Ḭ�JK�U��x�Μl:�y�D�:Y��e[G!f�	���ǈ�):""b����d g��עy�b����s�MxS����}󈗉�	-�<b�]�SO��c��3j�-�P�z�;��������c-�Sp�&�j�c�������
H�5X���>A�.zfq4!qA����7<AEY
������<f([���J{I�o�;�����r�9Z0*U��a}�� O"�"j\���ĉ��4n͛M�'��F^� �����}�$ø��K����:��"�~�U��}��������|�0*�wW\�.��/�']��c�׷@t�M�~���[�,��a��T�TB�,K��q�Q5�)�ox6����mJ�v��2#&�_�����1��PuJ\���*�"�SE�&���塡[�����,��9�s�
ʙ_�mz�����M�h��Z���֗l��M��@���k�s�&��xT�u��@Wo�9�9�#����6+f��K�G/cZ��ew��լf�e���.Bl+���f��d;�C�g��
����_��$"|r�Z�h&͙�n��0�t?�i�8r�]��
ࢿ�,�x͉�'�ZkuA�ΐ�6����W^�`�0���)��G���f��W���p�gi_HWg,t�"�?���8��\90h��Z�����2j�k��/�r7N�"D���a	��̡�3�S����3�_8;�$$����%2��2�yݫOvh���#ص�U�)�Ò�L�cRd��ʼ!�ūy������Q�*�KI�1Es%}@b�X�C>0'؎���a�-��
��a$�=��	����,@pܝ�%x����`�%@`������>����TM�:gw��^{��G�����,Rk�0C��狍!��aXi���V/k���EA� ������g�1j�L�fB����&s4?l��ٱ.G�D����l#XE�[��Wy��y4�Ž� �&Žc���ٰ��TW@�*K2$�s�������!N�=�����ӪhnԵ)�O�~�w�����T�Wr|��ښ���3a�ǾV���yPE�Â����ݱ�:�,�d�� �I�m,�W�xК�֢�"�6	�Jr�K"����"�Ȣcla�m5�%��`^�,�>��ۧ�@�w:A���MY���<��2�PXAJ���.�_�э}�_ӌz�G���Cr'� ��64�ɓ��9�7��������2D��D��y;��Z�_��኿��i@Oh�5,���"����mh��WJ�(�x�|;�������#����@f{k���_	�]�wd>ԇ���,�Cd������C�k������ ��~7K�?Af ���������T61P#������b5���	���P�5#��g,S�OQ�]���%"Up�/� RB"��װ�{�Km�
����W���4E���+
d�-��~r_�;��!P���%��,�`i��@��_��������&�A��+��e6HiO����w,^2c�Rs[F�F�f�tF��u�E��P���R�*��EqY��V�ց�'�O�Y��6&?�bO���z;�CV2����`����&�4P�0XR�"}�	�`�3�Ǿ2?��7���������TA��if��'�O�(a�����K���������EnY݅;��~�C���F��#�2j��F�R*���N�~�@v]��/ٯdL����h�׽������ֹl���9�!�-6H����߄O3�t�?:�y��pLg��")]�V�mL�@"����{(�h"�7i�2�����I^=0e*�w��W��j�Ɨ�v�/6i�t����N��d�	��`�?5=���D�<���)_�xS��k�sy��m��ϐ�($"I=�L����m��aW8`(�q�o�l�N	��${�,Y[D�������qW�L���0oRJCUx�	�E��N/6��:�E�{�Fq�0��ۍ^�^����˟ȇ�7�Ƿ3^�|Ħ�/��8�ɍ1�z��#�g�k ��`'�܉��؆-�	8|�RE��],�nr�QLW�;t�?�͕
�䛼���`!�|��J�bH��0��%�~܊ �L
��1-�TTЀmH ��*�q� �d�}l}�}��v3�?���������\g�]�����$��c��S��> 	?���V����Rt�骴^��X����'(��pg��Ȟoi[4���d��$���b�A�<��JN�/m2��m��n�]<I��/��}P1"����\���P�RVl�͸~�iP8Y���Q���R���U���Dw���{�%!u�`�a�P���!&`9�( ��0+˂���]�n�{#�Kk��X(%�q:��1�HVY�8ex�qe�G[ʩ���8
�]�j�:𐑋��T*��B��h��#�1�,4�l� �ӿ~�߼�ȳf=k�)�h�q��OR����;�`+q�H+|""N3�����̾1{ikU������5���oj�����\|_�a�T�\����6��պ-!mA�q,�Bf#׊�:3~���� [TT>U/D?��Ǒ�G��q�R�*��o%wǨ��J�%�yP#ʂ�ݵ�w96Ocd�J�� ��тU�׷ˣXT(k�ZH�
>	e���hEvZƏs��2qjw����ɠ�1h���V;�F��g����e����K��,�+����<I�,���C�Yf�+������^ӕ� �����rY��f%�ZCJ�@])�vҀ��	GǚQW'%ƥ!�*�a�.v��է��ۏ�nJ������h��_��Hw�~�0���;PE�7�T�0e�VB�z�1L�=��Ԡ������J�*5��z:WK86>�+��`vp��> ����+L!�V��5#�.�=��la�/<�2WǳFnx�p،��*��;��G��t��gS�T9�X��]�!�E:K�u��Z�_.ɹ��=z]ft�����%�0�R�}U1q�"r�����Y�`�Yf�jmr�=݄���%UGp2�'u����{>��e�Z��&1�,�Lt�&�� &-��x�_��h�3��KW=���)�)'����s�+��>�<bL�3�ڭ�s����6d���-������Iu'Msr�+�]:Ն6�N�vk�s�w�f>����p^g���c��l��e7ѧ?��aG�yJ�<.%Úx�VDVϻ�n�g9��(e�냈=�9��e�l�$C�okĬ�d��ogtE"!d�����nI�N��������i�PJ��L�tu����l��]���>dպ��zHL#�,�a�W�.�L�͇�kD@�_R���!�(`��U���O�K�"!;�u���0�f�#�>�G:����$�3�A �q�����xC,�s����O硸�;�ś4ÆcU���`@:�c�B���	��|�=ͱ�!w�*�A��?��.��{Ǣ��8�;��u"��w9N�IV\��~�[3�����a�?��}5b���`� �`6�lm���w��z�H�Y�O�t,�U!Xy���y�]�Knaqt�d�-����|�"z���A��&cwՅv``���`:�>s�&�6�h��>�Js�1�����#��0syꉂ��9w~%����a��M�")+�
�Gr�o''@�Hp�&��T��A�溡��N�#K�if���MBK���T6�����^�Xl!�6ق6�+4'Q_��6}j�ܡ�Dԙ�/a����ԫ�{�M���)�ĥeo��ܤ���;���B�\��O���<˦�.�G+�rjBԬ�g�����|��U�*ԭ� ��a�ح��f��Є�0�3��C�&�eK��Gh.��]`%�̕�)>�]�ܤoDC0TT��;�I�22�>�L3ph��G�v]4��'�c;ڪ��4{��Xq���+n�Bx�pk�9�*�f{����`���	~x��	��Eį�}ȂF��
Wĥ�R��WS�88��8�m��ëiNzK��"�%#>���K��d���Ξ������wQ���64�M�jn����˕N���+�cX�rI����"�f�D�� ƛs�3��Ȑ���_+n3����?������� �k���.φg�>���g�l �g�P���_��O�X^E�ɠ(.?��)1�����/�苂b��S��g<��s�wy�x�%�~���c������;a|U�}R����x�*��u�H<��U�"G���k�2nMĿD\ɻ�Q��:?���2BQ�?�VT���UBAO�%�m�x����V���||��v���<���jg���r7� �&7!��_7�sN_�<�|Ω�����"j��6�PR�`,ذ��������{���"\PT �:�%�C��F"E�M��������FG��W��w�.�c;�U%��yA7"�F��"��t%tv�)���eޫ]1��4���~�5|��g9�M����ٳ��gU��,�k����)��h�J�gMy���xi^��-��c|7o��bxG%�G���P�_�S�b������ k�[��H��w��p^H��G[�7$��L+R��S�0>rs2�� �\� �\f���]�T�u!eW�0�H�UN8�+l�染rq�~�I����g����ʼ�JrO�	35=
�1bO���j�7�^EF~�[��ҋ����Sh�|m�S�xܒ����FA���^7�d��:��=#�����,tC�wxJYH\g��:<�e�0�ĝ����IO��AH[嶧Kz���ߙ�KQ́~랞�C|�DM�v{0��D�w������e@O�q���F�)�0�iY�����#�	�O��-|�8��#�Ͻ֞��}�c�����;'Hn��^.�x*�T�}�b΢�8���ʈ,��5��J?�����[2���ו��DS�t����gJ	QI��6덞��+<�<�[��N0͞�ڵܤ�q_ ��H���̇Ƈ����^��]uw�m����HwЄ�6T���s�� oQhNѕ�e�?�b$��AQۏ2E�MI���e�u�\p�$D��X:�Ɍ�z�T�h��vk�����{c��'�B�#s��_E�/������w")�XW���G0���w3�2k���m��a�`�Us}~���t�dj-ʭv��˄�R���ܾ�+�N�jb�@��k�]YK�&,�XO,�.�R�Ŵ��ڀ�励-E�u�_�<TH�t��8_��#�,��Q�v"^Ge�=�OWM�ɧb�/�H��������
z�����5S��%'���`�,+`nz�6��2�0��vd��p��͋{�7<L�����c�H']�s<5\��sakb�?a�:h�§�xF�om��]ǭ�0��sн�'ς���0讝Ey�����> g���6�4@i;�!�������X�6!rf:h��UnZK����,M����LO�q�ٓ�х����0�Y�g'5m��ϒ��T�,Pjp���	������'�hg/��1&�SB�Y&��X�] �����(��}mc����_�0�O�����
"�T�Q��dG�cs*X2*��~��[_��o-I��5�G���ďB��.�!H��SklB� U���"��z����~��q���U��JyE>���`H0�ۭ��j�f��컳.�:�Q�<<3=�}�H���I���PS]�\�]!�mp��3�%)·�`�~��e�-���(��w�=�kBY7���mw���U�zSE-�{kL�'62 ���G��Ӻ�sV����Ƽ>���{�n4��O���BF�t'#vsfgq��Gg�,m��������.��E��j�t�Xr������>����{�:9t��^�ϙ�����VQXx_�.��"�N��n
p�3⻸U&�x�\GC���vxT�%��م��ȱ����rSY0 c�?^�~�󮔍^Z�r�;(�a��ij��HI!˥�R��(PRL[��{�2h�&���4�����,��:rC����`3Kl��1���3y]���(A�]����\I�'�-z��7��g��/����@�`V�@�aT.��!ܕ�`��ǖ�c�����R9]��BrC��u�n�ک�=��|�����s�t ���;V��ր�j~~�� ����,0+�, �1��R��H�����Awk�Ly��YKzg0���ן*���i�.%�n:a"]�zT�V$2EW5��虿G�l��qל����>��U��r�Ò��v��cU�Zi�%��Wx�҇R{|��'pҚ3�y:9�L��zm��nU���綶���)�[�n��	@�-�ܾ���/� DhЂ�}	�r&�Q�PW&_ހ���k�Qbg���G����ٔ�n����aʪ�;HQP�!�o��J@e�0�設���S��\�&^�e�������6���{�l�jAJ-���G�t����U�eaw����2B���'��~O����S��oB+?�:��<�Q�IHuzd�H��V��
Sl1I]9ؤy��@���p�H��y�����;th�sR�5S��_[0�ص�fJ>�Z%jG�Vm��5`k�z��8�_P��7����B-�d��C%���L�����伧¿�s��~���~	���Lt�;�tC�������qe�[�m@��&�nlH�e5)�cr�����)qu����w+���'Z�v�Zd_)�%��a�M�2��N{M\oA�?�ODf��Ф�b��屎^�d�nٓuر��X���'�����"0�z�U'��"���ذ�us�8
	�+T.���9����Ѫ@��F]�o%vo3����˳��$3��ut�e���철g5ڴhl�$�9���m�|$l���MA݉ѣ�h�H{���N[;J����&G���ܞ�A�i}��C3��[�>d��VX G�Um�_lI�,
��&����������<h� ��,q���#\��&U�Jrҕ���0�����8y���*��WT�*
�DEw�2gr+��x��H-�yYGP'_�J.ǕJ��Ҙ�Wp=ѻ�ܲGbk>�ۼ�ͭ|?
��hQ'C��k�?�C?ʂs$��H]���Z��Uu��;v �0��{��.�Jz``ʏ����4��i���J[���s&�:g����� �4�}��Z�t%��0o>AMC�d̻�٫����zL��v/�1�5 �C���;r�F� �/��k]��=n�e�����X��?�>J���P�N���amH�9'�ʆ�y�!�Z�KX̶�HGy�4��Ӯ[�9E�ʯA��	��)�{Z��������VnBe ��	��*ˑ�灶�n�r��d7��`�aV�gt�3XW�⿍6s��3R�ʁ{'¤��9��!z��&�ß� ui�����p,1�Y�F�T����.��IG�4N2Uv�4A�ƈ���h �jOk��=���T�T��
��kfgQf��l�O�/�(�.�˷5(��Ĉ�����[e��Z����NR(�bd�=�K+�f��O�G
����7y��� 
�xL��w�܌�I$G�g{����
��+��8~0H��{�x�Lr�drW�Q���,`Bl���(�h���ު��	ךM)s�>��D�ul�om-L�$��D��^D��tߡ�Lubzφ�V��~?�*��_+	f\=KtR>ʼ�QI���x��+�rJ�dR�֐�yF����I��Ym�<莢�����rɾ��ʻ����4���x��`��l�٫���~)�r��r@%�>�ծ��'К"cw��Wm�	���8��]�&Wp";VC�9V~�} E��2�yK�:�����_�����������^jv�P��o�i3����d��k���݄�ٴ�{��rE�I>�[��O��@���]�J�;�+�)�NKz��5�?qL	��ʟ�lȑ���>���2T5�FZ��?��R4z���R򖸑Z��5ˑ�>��2�� q.}}�f�����C���(u��Q��9�ޝ5�^.Uk_o�L�s�h���7)����ƈ��$���I��w
9,�ٕ�YD!$੔-2��]�nz�Ю��;+v�ڐ�o�s|��PNT�m>$�U�'�/���U,V��͢�'r&鎉��L�RU�U_ݔ��ռ�vB�HY:��9H�\�Z��4"~��f1�Ġ���b��J��Bp{���rلU�|N\�lC�g?���K���+�V������
e�9fX�l���S�l]r��k���R��(��B��]n|8PH ��;�E��}�s�v��a�Y%�|aE��I�X��Χ���{MO��C"����y����|�����ͥ'V�ŷ��(��y��ѣM���KYl��k%��S��$��B��c�kI�x�@���8;��l���������ʡcl`4ˢ��4c�ͼY��h%34����[d�i%s��t-Df�)D�u���f��'�52)����\<E��U���󻎅�(�G���+//�@�k�H�9rgX��S�N�4�|R�lٞ��������˴�H*5q��mrͬ�	�lk����0>��w(i�/����p�ӱ��� �F�T����wN½7˛�;OM��z;���d���a�����~w�|��n2����M�_�����������6Bu+�k�����d�Nku��ό��e�n�������������O�� ��SB���MFk�J��v�G5χ���́�>_��5k/�y �0C	G���Y;QߚJ=W���q+X%ƨ�lQ����.�HA��w̡�3��% �^k%�W�F:���Q����A�E֤��p��D=�?ך����O��'f}��v:�����)'��í��92ӊX�]L�z7�����5�X�W�`�W������인J/^r/�Nu[O�[��L�  }�W�Ch��e�F@��\�GԠ��P�O���B�0쌢p��tY�0�u�usZ�d6grxc��1$����{��B���?o� Qg����A{�ڼ��r:%p*�>���B���+תؾ~���^o����0w(Svk���1�1��ӑ����W�L��7�� X!�/3X����X��Jt=,���@���e�Gbbv��I�J��E)�ɽ? UH�*,��T^*i��������̉����(�)2����C�����$ )!�|z�1�7���P^9��OT��X�T�v��:Q�)��Z2������W�S�������@F��,i���?��"?9�}�9��h�B�-����f(Ú�Z�W?�����M�����f���:�3���*�H��e��	���[P�ߑ�b�Hy��uL����
��>��b�~~�G7i'�S!,ʄ(^����9e�'��G^Q"S������H8�BS���GL�C���Ɯʽ:��s4�9�Q�ƨ�Mg����~�,�q����)�.�fX��bz�GN������*]���+�jE)�WT|�;�h��=�\CO�s;yƗ�γ�)W&:�e �x�$��vm��T��B����ki-ߪ-~���$*�Ѱtc�C�L�I�#���a�w`�e��M»fr���6^>
?���g����MF4,��_�!���:YM&����4�`Iu�a�KȢ{�0D�skC����̀�ӯ�=���lߋ�]"C����<���o��n��`c����xұ#A�0]���h�|��*��r��3A�A�S�uA(;�3�o׵�]_Jw<3(U���!�_###�6���4�0�����E��D|���Rz�	m������* ��
�-��y�wI����4���~���6)�x�]T�zW�c��O�����ߟt����!|�z�zzD�&Zc��D<:�)�H�� �or��ޏZ�t?/'#��K��5������w�r���Xֈ?O�
,��+���h���C��?�W67#T�3�`���i5��z3����L�a��U �n8g����eQ�[��e<���I���m�š�>��J�	 ^w�ʯ�S��S��Q ��x�Hi}��}�EB���l9�;LS�:K��o &�צ}����b����H��I���o?~*C>z��yH�0�G��qyYpdɟĜ���s��Ov�;�E��_�ܽ�)'���N��*5ۜ}ӦkD�������.�J�7|.7t�^���3���V{t�������eT�{ڄк�v*�q@nW���?t\y��a.��U�����d+��|B�ɞCj�<�n���M� ���Ȏ��A�.��"2��*tjҸld==[��ly�ܬ����v9���]�F��y���Y~�>�x'tHX�i���+��ט:4���
��nm�������S��Ke��i �~:�&���{���'yl�U�O�<N��[��������}Ijr(Ijc��Z��/��O 6���fX^����}�g���t� `h�C��s��$Q���Dr���N�Ľ߃=R���%Z�~�f�1�jj�r��Z�iT�'f+�ު�2R���Κ
 }4^/	�ls�w���^�������c�>gC�e��k�wa�װ��;C�4�v�a'��W+y��VK�X�|�we�T�x� =�P����&f���X��6�F���!*���6�l�~�S�j�-nZ`�`ç��fe�I�.|�8���sս�b�r���|�b��۽Hf�r9�N���;�9�)W�Yn#$G������dk+h��Z}�����c�2Y�z?+��"�}�)�̈T;�s�~QQ$BYvۙFq؉�P}�CA��3�l�����%fpƨ�jIZb#��6C�-�a���R`.y��%ڃ���]��F�_W��X ���u�9ci��c&�J�[d�$�\�PF$AD�Cٟ�T��k�il!Wvg�J1=[�����М�5�a7n���i�W�+�Q1�Nh>�������G��9��l��0��Z��!�H�@�C�/�ߡ7���V����Z>�؋�aK.L\��$���d�<���*P�c7/@o��9�AI��ZÛ��Q\�G)Jy��Ht�p��I�*O����[��H�d��M���1D�P3�����208�S��k5rJ\��x���G��#YU�٘��1��m7�<���{�l��|��Z�m�j�.�{t���	0,�R�M����_�Mb�9�;��\����;��	a��>��Red?i��7�E�^�'+��M�2j@{B� �
��A���Q��C��K�>����3%Y���4��c0�6����]<����VZW
��9#];�[<��ݪ��%�	s*q͚l�G,�c�����y>�{X�����c���_+�]�ðE���$�����@�>�[���`D	����
��YB��4�c���o��1��u��q-=)����.v�,���3��G. �wg�1�4���~�'��W���9#D�r-`���6�2Ry�r�J#�o@��{Ţrg���5�O���3��z�b2��X}[�p�yBy>xͨjiֈ���gr��b*�fN����q�}�-�)ǺR*4�!�ll�)E	ɼ<18�� M0waa����$_�y�@��z7R�����`��"h��|N�a�^�C\N�G쀀ʄ��̔������u�3�fVY���L�W�a�&��<iRϪw��!D�ֹ�m)L/�]��b��קf��lY��4s�~]x,�H:��)w���9˦-e'�?T���Gs��q�?��gq�gL��ܵ	PQ&�n�#��~�B�Ó�b�2J�r����e��f��#�6b��~2@���9���|< AH�q�P��+4�.7�������Ƅ�s��R�?h#��<}z��g ��&���<4��I�R0�㭷�s�.x�,�1:�;5ϧ����}	�K��;n�.l_G�/��S�b�l��!��~͇��B=3��(ˁ��C�Zc��wV��j�nD��Z�2^���ͳ�tqW��d��E_%`��^��E�����_�Ϛs���sh)yW�]�"	ޟm�w�cL�kM~�`�σE�;
kfh_zѩ.��-^`"l=���}K0��n���,����\ܴ��f+�����2�XF���W�`}&�N(�#�Kѐ�-W{�}����M���	��2<��c��*��kU��}ǻ|,�<�3Iy�ohͱdJyT�LA;@����|�O�E3!p���:�0�#p�;��,ј��O�N��HS?Q��RWO4.�*�/��^p7NJ"$��-��$�t?��:�k���z��]���an'��(�`H�0���ϼrK���s�z)[�����~�vb���5��ݥ��o6#D'�#'j�G�y�}��~�u[H'	���9�c�ӊQ(�����L �V�Pa-#�����jU5=����������[l��Ք~����V8!9�/+�B���,鎅SE��]�xz���S�<H��E=�S3�c�-�9�"H:h��>G�1x�+�-��Z���*�2��������+�W
�pL���,Mo����T��9����1����\ؑ$ZG���oO��.�yVJ�7C��$����z���WD�jC汛��)F������:���u,��QX����IOb3�L��]����8lB�d2��K���d��>�
�[������c���9��d�J���-t�Rb.Q1L8��~��(��{{E>7ӌe��a"Ղ����9�\!��3���~{�y�.�l��m���,'�"��M����?,Z��<4�d�.��#�� @��N1��b������nB�J�m�)��Y��ڊ����hѤ�km���2���� ������56��-f���;q�\鼋�E�]2f����b>����Z�/��$�6~���?��|���ui;"vy�ɥiێח[��D~����x&�%��T)�. I�D	�*�<.�ET��?r6|L�&������C5.���x�o���7�d0��'����k/�q�p���N���w���`��5�0�h��;��z�!	�_ArרOʼb��߼��,*�K;�|l�(1�2nAAV��q���\&��~8���>�v�91�k͈փ�Fz�r�}��¼�wr�tTi.�$���X`�Fj�O�v�r��S5x���1�������Ԥ����\v�*����QUѪ��EJ�mI"ç�����~E[NE��Q�&�>�y��023�&�jt���*H�#�~�3X��ru��"brU絟�"_8�-J��&�����{;��{۫��1�X�|�]��=�X~Q�K�g�V��,�8����_u_m��eX]]������������
߲�u�0%��GK'�O|Y��V�)�RC�Ї�Hc�&��{�O5HW��2i�
'@?�Ϋ��ّ�o,�@F�Øl&��o�҆�vq�����s�!�I��k��aO���c����ϼ�*s��/v+WY�� }c\c�W:Z��,�هW/�[�mO�K�a�{��
PAn��%W�����>���sOK�Ig0�Ӂ�W��Ο������0�C���K=F�"t�=�%4^��'+��5�;!y|:B�]�Ȉ���~�ɇ5=�ݏ����bb�V�Q�Mf����T����Y�	�V�I)F��4z(-��<&~���#Y��b�q��I*��p��ٯ՛w�:ێEb�T��f����͵'"9����þ���]��Ӝ�,�n#��H��$ȗن�vv���`���"����&1�~��.o%�(9�Z9��uv%��ҩ3F���=�}��`�(>�������8-i�V�9E��.�>�3�ȿ*���>u���]��d�}�c�.|��wL@���������`i�IӢ�7o6݆�����0d%≸�!>�-]Oww������ހ���/���/�#�-�V,����t��AZ�/��RqC�t|�7?|��0`@�d�hD��?���d���|H�!䃈!.���a��<�~1�k"��A:f�N����J�4|���&�X��.K׶���JQ��ABe����%���+F��ێ��:��C09�T\�s��m��VV���̶��CB\?�2���ϥw�go���(��.=�$�".>�%�ؽ�f ){��N�s�.WM"2K���Ez��&R��s�8W�nB`8�8�i��VG�v�.�)��K��w���Ǯ��.�<}���ƣ?.s�]�/���U�R���I&��dJ�eL�����F%�50���We�y,�L��`j�S���#%��\�f	?����N^J�u���t�g����˳�@aC�M~�W����tJ	����jw�~�8�r�����]!	2B�)Y���N��M��	&��%�j��o=�u��ִ�So������]�;�ʙ�	��=��6�q�a<+[ۅ�Dl���W��
**�(((G(�˨loIz{N�&Ұ3�:�P�{��g��,Z��/��hKJ翓�8G�:��d�Գܮ�1���Cvke����F,��:�+�T��m2ۚ��3ٚ~��$2�)��(T'���:}�v��ٺ�S�]h����������)�P?�'���g�Ek�N��XTT���)�Vakx����J��ی �# +��n7�Vg���I��ñ ��e2)��B١g�<jAq-��ĸ�x���h�m�]m��B��}l�HF`4�<�D�0η$�=��I�`+�#�L��@4�t4���f<S7�|�,x�{1���K�"�s��GOL�,^���O���|�A��1`YǸ��s_��668
�<��������-P�W@M��e/G�H#�W+�K
H�<Lّr|�
�z�8�X���Ԕw~�!�H�	�^= (E�C��H�d�����q���<$�Ή�D�ƈ~��ȓ,�[�³r����	�-�r#���dt�q?I�?��\+�I''8gd�-< +�!��7��r�垆ag�H��x.+����6^�x1se'AҸ�}���pӸ�i��̭�/�믫������q�X��4,��j7V�Ν��KR�;#�U!�|q�O����Σ�LLR����q�x'�x�&�����58����%Kd]P�]��Hkg� M�K�S*u��S����^Q=[=���v?�G0}�Z���:mu�"Z��e�}I���P�.Ǳ�]�G�kM�a�Q�ٲ=%���=����@"�eA�r�Z���B��Mr�����xd��J{th׳���I3c���!������)�f���m�#\��7��=���W<��R�8aL`hӨ0��Z�lw�쭒�S]�p��p���gK]D5���f�%�����ڑz����;+����[�MB��܏������0Yw	�
��"���`�ٶ궙���S�oY�[�HU�Ӌ�N��W�
�Ŕ�P�y5q&�[���̭��k1
�9`�����Dqi�>��#~إX�i��K�@�J�E�~z1B��QF�>"<Q�}�B��f���^b�y�#�3��S�o~����浊+'�G�N�-P�J>�
�iǹh3@�m]Co����ˎ�;'Q���2~�� �q��y�J�����NTk7��[��~�0��d�)I�6<��_�'�@o��K�Gə�P�hM�eG��JϰgՅ��"s�rj�wo��孶N��L�B���h׊}ފ��cRY�۷����Z���t�sڥS�u���*�/����rv����o2m�S�m�r5�4t	nu�	G�|`�[��������?��:# �:�C���l%]#�*��_nƙO��Q�(�h��ԖŽΈ`Z{�Q����G�Qݭ�R���卍�I'[��4�'�\ؽ��f�"�w���А0�l�on~݂)�^�J&�n��N�/ޢ��in��*s�9>ɶ�H��s���C,�3�q����1�e�g�$�Ӂ�"3��C�MU�&L�u�4�2�����������S���/1v�Ki�U��+�QKlj�%$ĀMe\aBնR���+���b�^��ڞ.�v�q�N����B��e������m� �  ������w��<�����R/���'K�Yx,őY(\��&�����שm|��q���R%8��X[a���X2K���˧��!����6�d,��¡^��i�i��d�$h���U�w��-��AWiL���u]�[�kMC������Ű�3����iO-�Yk^���Dܲ]��Ŝ��S?���S۳��*��;m"Ͽ^�(�G`�ө���v��ϥ�YXc�=�#pG̉.,Ҽ�fT�QX�mƑ�H���Jx��Ug�:�)8a��U��v.��&n	e�uI�u^و
�!1q2�@8�;�Q�Ol��l�e���j]�a$) m�R����PɌ�K���J{�q��Dk��1�ulz���C@�&�}
�����%I-ޥ����,]�a�� ,��VH��+�s���d��+i�����M�ȶ:P�`�	�T#���6«�R�r-�,8��j#�S�I� ���q���]����+�����98��?�*���"	�im�p�r|��v�B��~���I1�B��ӿe�l�F��A�\q.�M�s�M��z�JSÐ;bʠ��}%��Y<͎5b�Sv�W����j�<�&��22v~�vj�aVj���fټ�(�����ʐys4��?�Z�Yki�%gK:�(��3�|���׫����A3R�_oV4ޠ�.^M��gC��oMvK�E�a�ɀ\}GW;��v�}��jhp4z矽�pm�&�-� �������TWN�9i�MÓ=j+��]�m���	q���|0���I��M6��O E�N�C� �1�yD4�g��X���?��Hr2O�[$�*����A��'����7I.��.�#E&��	�k,���n�G�?<=�a�3�s�����y�		�낱����J����$zm���U]���eɕ�,T�Ay��VI���T���}���Hx���R�͂G�w�0r� �����O�ı-�T3�H�t�9�<,�]�Go8��	W����2�i�RE1�3A(! ��ͣ�]�0�����@t{���h���8�BJ�j�
H����#�i������#���ߖ0�j�@)k�r�)�L���V;q���3��h~9VƄ�L�������'1���\�͎�( F�L�Z�s
�`�{��u���I^�_v��\��_�r�hD����Y��d���n?ՙ	M�����i�/��F�5�a@�Δ���N�����oX%���'�/3���s������Z����iA�8�Z��ݪ�?bsF?C�\z?v�V��R��U�z�CIzVp�Ҷ?7��x7����4�?�h����T����.:�h�E���:ˇ��*L��k����u�qQv[��A�kHA�KB�nɡ�;��nQBB��[@�BJ�������?�3��g�}�:�WbF���H�;�U�6j|,j$��K3�j�G�/�����U?M��`F,O3[xz������X�T�5H_s;<Yϱ����<���^�^:�X�[���qt]��GK�@ʞ�D���5�&ʱm���a����z�����k����I��d���!���0;��R�A?�1�ȖG"_�w�Wa���jyu[���n�J��E���1@��v��m=a�k��E5����R����gA��wBV[�3�����rth����v��I#eqS��2�-T:���@��F�@��<؀ȞXHz �M���wg�G�	����m��#j���_W����'�s4�$1|a�M��ɿy4o�/O,�6�uN���V��?o�!�Y������k�l���G��dJ
�ŧJ^x �59�����*&�L�K�9����7	?��{��>DE�����R{%H�}��	���u�-�!�Ⲩ߻m9��=�%v�Z6�O�e���%���u�\z���<��"�����\$ں��j�'��-o����D,�(��k�iG�E�si�+V~ �F<�n��iX0;��A��y,bX�%�ڏ�#�
fD9A\�
�D{����O"n|�� #�Ec�+J�FO(�_�B[�բ��w�SP~c�9g���sJ�ܪ��?AD�W��<MWi�)!��	בή� Y�]n�u��֪ʕ=?����9�ߴN}8w��H����Q�^�U�?���?%��?2j�#Q�Y��o������$��-�ymR�iǇ�$�sL�Zhg=n�8k=E���aQ��C��d�x��0��ꄊ��r1P\���o}f�_��i�	:I��9����憀��Dy����#������\�37�}�.�B>��&�.�aK$��@�߼V.�$v�T2��!jk����I���\M��JIGN���#��g)�m�si�d��/�n{�#6��)%� T�s	E��[�LգX:�UG�ˮ�73-GT�6�c�c�g塀���힠�M;�W}�.�H�áT�7��m��#0}y��t�5��/���s���d��2����5vƨ#����S�6ǚ'*��W���T�$�uՔ}�s������>���1��s�o��Wl?뤅1��9i��������ve��=`�"��� ����p��Uƛ�	qD�8 ��N���l�5�l��뿺,�g�(�`��;6ʡ��C3�_gv�[�v�����3���n�C��!=�y�H,D�����7'`m��rSJ��A����|*�}�M�,Z���������n8^1k�m31Y�iET�|�R��G��T�11�n�5���ܪI�{ =U�XNl{��#w�v���f��L9�+�v�g��)ˎd��&��B����u�A��d���fR'<02^�wG�}\�$@m�u��Df���yS�����X�Ĳl�ڵX����}#p?�X�q8[M���N�{�U����?���nߨ@�El��c$ڈ�r�#��8*~��P5��*.�&�a����Uφ�a��Fb�\5���
�f{�ߡ[ٔ�Q2W��?����y���x��l�<�ir�m�.Y���2u�>r�͓[@۶�8��7�-���u����m������iM�<y�\��/vNJ8�?�Ƴ��z,���$�0����U�Ԫ�>��d�{<m�����Ã��]b�+L҅ԡ����s���x������:��:��pBA�RR	v\/�4���6����To����Vq�if^��=y�ϑ{ͯ��N��{���5�%�;�A��u`amB#�߮�T8�|�u�rX�U8�*^���i����'e#vH���@�b���O�Ǥd�����^�u�Si
��?�7��W�xi/��9e^��1��#�x�- ��鼰`���
.�	_t�$����7�>��w�����P���(�O ���{�VӁ|�(��UA���x��:v��K���P��-0aʬn�lɫJ�2�8�y����k^��YH�\�:I+c�O��7�ث���\��Y֊�ݨ�἖��Uȕ^!Bg�|]����x	@O2��Kg��J(�|'���˃����.V|W�(���T�f4��a�!�i���W���Ϸb5�n������,�!
�yhN:���w�x9G�'e���61�*��S��9����o�RK@�{�s�&��0%�]�6��"����=]@.����mV��w���q�y�2;^�v�K���ʋN7��� �A��k	^f����`�#� a��b8P�EE
[�E�r�.m3PDXy.�2���R=���8�.a;ӧ_��Ew�'ߺ�.���6�Wy����矼��(g�TN�����Ez�М���u�����s����uc�;C0��G�6��X�x��� ϴ����g�B��)��]'���5��/]��d���MQ�*� -���3������j-.�(��`e�9�~T���~�غ:Q5��%0�ؚ(8�ٜ�Rw��y_��c�m����tb�kR3>�yC�Z�ݣLa�>��T�2�5D�Vk,��D�u���W>
���R8�ʙwt �aY�U��@&
�,[Q�1j[��o\�|�J�]o�=���p�"Q=.K��G�#�%��m��oW4��2�v��JP�۫�Bz���'㛢����H�,��嶳�?I�����\f?�2i�����s��Ȣt�ૼT�u�E��9�[=����~L�+S���m�-�_�}Λ�̠��a�ٍ�C޲�٩�fMj�x��}���*�GP5��i�.�3Ҟ3�W{)������<=�^�98)��8����ݶ�*�O�c��v	˻Q�y v��[�4V�w<��	Nrl �fN�rՔ�n��R�]������q���\��r�*�i}�}	��%�4�|'2v� �O\�_}l���R���7�Oڳ!v��w�&O����=M4�E��̣�rW�g,��+��F{lӅ�+3n�<ko�/�Da�V=�O3���@���	#V����7v-�:���*ŏx�R�c�Y|��6A�}D�HKR �ON�+��L�'IG9�?{(x�J7|pYퟷ�|e>g�O�|��d�;8����[4}ْ#�[�c5�ĹɈ�q�|��^�V_���,A���8�+�gKXz����9F��Q���[�Y���X_=��'���f ������s��������jt�S��Ti�Z�*t�L�k�glo��t�+�ӌ~1��ĺs,�3�;G�rD^˗�QS�!��'��k>��P������?&])��[̚�F���s��
Ь��n���Y%�sk��f|��!��r��	�����)��@��]�W��^'�a�Q�,u�ћ�j�C��n�0C��B%��H�"�܆u˲�b[�B ���m��jyǪ9�ܝ�k����3t��*�ڻ���:M��~�cd��y�f�K���*-;c���_)�@�)��9`�~�X
I6bWe��^�>K���Y�ʛ��T����)̘��|QD�����S�S�.���(�:�X2U��Y�c�uKzh'�MVրۇ��K�vs9�{�����N,MϜ;���}q�bw�r��L�����j��b�udsР���;���
�ƾ��+��	����AߏYn�`����p�𾨄V� ]����G�E��65���Vc�,c����o�����T���G7��O�B5B/l-�����֛}��%�EEr��AQ'�x����ߔ���Y\\�`����饵�?}-u���t�Y�E�	���9��Dn��2�x����J�0�4��^�e��������S��
�^̗�`Oz�����Zѻ �,������C�9��s����L���R���1��1��g��t����(㔦�;�3�$�������)6�q���Y3��*��N2%�`̐hu'�l��&��Bu0���\��F;�Tc�3�ʠ������CM�+o���B��x��4D�!���	%u�O2�cY�\;f�a�Ҽ�����_���i�;���9�����w�2�,�(��{zÞ�W�~����C�[�R"�SJ6�^Y��1���{%��w���F�:���)b:��k�2��\����dV\�G��y<��_�fsu�?�k*���	��'�c��Br�v��Ƈ����A@��~�I%�C �@*SG�����x��f?�-<*���u�S����ס�Ɔ�r�1�ei���BXi�5#H�'hx	���)�&2��QP��GK��?�y�:��n�fFN�&5�Њ��x���h�wm��o�Ve�eY(py�ڱچ}�+_���P��F�eK�	����A�/����ʂ��'K
c�� �&�S�OR�`��M�+q[�F��������f���.E�� ^�i@�$j�c��)h���CT�-������d������yL��ͲqD���2���#����ﺾ�v��N���P]w�Y�*&	�H%���@),A_a���k0r.i��v~#>���?�t�@2���wYG�4�&�7:X:���a|C�&c��q��4��\�rg�GK����ejJUa ��S�~�l�m�"�&)	�򗹮�9�?�%Z�٫�ݸ]�����]@z�g�z��`�b�wgq�G��9Jof���O�Ҿo���o*cch�D���4h� ^�'�<�`	$p��y��Ү�?��/qO�кW샇Mo�7�D�b昹�}��Y[W��	I�9G�Z�M�'f�ӭ$��Ǔ3����v��j�"?-�|D����M�6�m�e� q��)��ъ�Gs�#-�]�R���sa_.��_z���z[����YD��e��L/ի�r�11�f����!�;�T)]QG']��#��z�o���kbVгT6��`dLeoܾ����]TT�	�4�	>�Ln��1j���#N���%i�[��ldI���3ޖ?Ν������6j.�����ޮ,Zv���q�2�s���@\���4�i�X��'�-��t�҂O�Y��!A��x�B�`��FZi�>���Rվ���C�T��
��V�L��ږ�+���C�����	-�VV�#B��_�I�,���OA�eoK~;�,:Ru���9�����}3�d��\�8� ��V�{�yA;N�Ԫ;o?�j��?Gˬ���8ϜJY�8q{Ѧ�ྛ��~������>CE��l�B�Jtn�n���Ư���ޑa��б�w�ܢ�Gn�ۂ��Ai��lݱ�m	v|p�e��=R��AY��}���i̺�vop��� Q��J>;Gj�R��nU�,n�b�����v�� ��q*�um�w����BN�-��)c�vl;o��A���܋ �Q���ϵ�
�u+D]Zib�Sn�pd��v����#�T��;{��MYU��]��]q�
׋<�������>C�UF��j�T�{_L<L	���Ů�K���ڗ/e)W^���u�-EM��?�Z_y&&���W�럆�>�z��5�~�s���u1#�}:�7u$uٶv�y3��93�yh�Ԋ/Y������Wl��w���?8�O�Dq��_����9xJ�z{�ځ�_�F'��`�=>�|�LJ0��Y)�"W!-m(�������ͪ����$���cX[�//�Ok)�{+>�{M�����b(�	޺8Wc�ױ�Sa�$��r ��r5�e���k�/����m�G����aSpD�X�\lNN�����-�'-{T���;���-(	�+5��b�(�iCf����'���Ǻ�+ 9u� %�V��e��*���dB����VC���p�cl;�}B�"�`���3�/��f�l�-&�\��G�y[�گ����v/��+��%!&����<5K>��� <�_;�|��л�O���x؇��Ii��-�T��ee��$#hظ?�%;�"��	���q
�K����?jU�����yWP;���V@}�z=�_^a{��z��X4�"�GO���c-��7.7�կ�O�[O����z�{	�=��Mi�`rʢMoF����my�a��_B�a��D�x��o�rA������%yp������@*؏������K�������Mea݈����N�$9�S:��d���Q��i�ZSUX�����߸Ww�z24��(Sz _.鋻t��y�ތ�=�tݦ���:݈r�[j�){�+\����0� z��wp�� Gyj�S�%���a���L�h��ƈ�j�3p.(o�z�����5��ß��~Ǒ!��S*~U�?�+ZIB�\��ĺ8�+�,P����y�VLf�#R�Z�"�L��ȷ�]A>O']l���+}x�ǎl�鈆�blJ�p3�2��� �5g�V4+dXt�{kȷ�VEҨY�4^d�8�U"^K�J�\�p-���ͨ�'ʇ���VsW�f�n���7��ם�Nb��o�Pq�Vܩ2�H1�~@�aa��C�@��zW=��J�n���礯�(��['c՚f�4n�#VZ�EC�Y��h(4�iH4�hl�O;�����9�:^4aW��X]�"�"��zugh�	��OI��mB�����8"�4  +�O�L�d���=o\���@О���>��H_���Sh֒�Z�񌏝�7)�W����*B��1k����;����[���������	=�ԍHT��)���l�+��X>bU.�����Xj��q;����A�Ա����7Ib�YI���^���.�
h(�*AV�Y��S��qO��4u~ff8�^8=�ܫ�RS����F���G��~c��Y?��ƍ��?t�$�HJ���lɽ�UϮ�w�`o<�χ �N�LCc���T��w�3�͇�D����� �'f%b
� c^mޜ��p�ZM z@���\���c��Wk�f�x�H+WwIzWJ�D��3U9(�=RݝȖ��t]��$�'����߮Q\m���ԠF���	����˵�MZ�#���@&���C�LN^�6��spay��hw[�ĥ����\~�-�u\¢N�?|��L�QSŸ��c�f�����캨��ۏK=Mع*���x�����\��+�T����/w|���oU9��>7l�g'����3���&�� �Gσ߶*�Atz�����!���<�5�ߕD�O w�4���Yn�:�D�[���:YA��Z<������6��V�g�a�\�$|�Rl��B+�o�Z�1���W]
�ӹ�U���vclN8�5:�އ�r���ʦ�.�+�:x=�:rq��� �>��A���s�~u�������;'܁ط7r�Y��=s0�F�	� !��{w_:�d=�!Th�AYvZ#�3�)<����$�g�E�UQ�|^�F�	���X��P��J�����(k��}���������Q6�<�=Օ��Q�s�S�^�����&�Ou������q�g��$<�~G^��S�5�)����0���}W�~���C�&	���
w�N�k,��j����I� ���!r���S2�5�9"�
�����!�¦�Z�61���� (�B�F��,`[���%�$ ݙD���������؟��1���v�g㈓[��F�BG�lQ�m9�*O��������z���f��{pwG�O��Dx/��R���"�n��~\;D��1�7ܙ���^�۳Op:˾:��b̥�20�9��TU����aI�?�,Œ���<����o��� ���PA/���vċ߯���e�5�
�C����ߓ��r���8��B�}�f׉+�V��V�<�ۺk�8��.ͫ+�e��%����I�G��Alw
�_�]���<�K�3C	[��e��{������;�j�^��q�4������q-�VN:��j��1��k6�q#�%�|T�li���J;:>�� �]�/;��t��(:y#�����`QO�ǲ�oi��R�9r�x Ҳc����g��g{�\R(0�Kr�~Z�'����/mE/�`���pWc��4�t�\Ow�O�V2�!��6�Z8~ A��֕/�5�	$�h�7'f��x�^,!鳼厞!��A���l�����<^<͡���9�<�C �v��6�
��ņ�0������R$e���,���{��t�v�#����Yn�)!�qW��j6Z�{��k�$g�)d�����=�3�c�Q7*,0z	|���OU�tli������ێ�bH1G������F�����$;Q�?b«?Ѷܝ�)���kP�kn<xE�1d��'��,����Q��>��� ���/{7�0\�;�Z�8��M�6τ�fm/���\�"�W$�����lRq�-�9�̐�$�tqU`��y�聺�W^Z�|�����R;>���U}���%c��/E.}l)�O��,�T�}�q
-iJ�z�(�U9}\䷩V� �a�����tW�W}�����P<I]̺"٠��߇�)�9���7�G��7R(���>Z0��xM==��{IN�a�H�i4��.���E�Z#�|]���!�dDSC��o8?���y֡k�25�.F>����H���+̔�f�Ub�9^�r�aoԧ�t��;���~������y��V��"���~l8^�N�.�(�@������X}�)�v�42�����,B�wp�h1*3�>m�?e��LXx��ʂV��ZՅɴ�\^���|b9��Id%| ㌣"s���&a��`�@��+�#�b�dc�����T�I��E{�:��$�a�]��E�$j���4_�iaI�m`�JI���b:0'�b`}^�_x	��{hzaU�!rk�;�b���T)Qu���z�:��x�t^�p��K}���;��g1Ƒ�á�X�n�i��a�F�ޠ�8�ٓ�S�N%�7�S�!�S�u��)�|�` ���P�_���N{G��P1h=����O��h�r>����O�6�G���fS�O�����m=�a4�j��(%}���<�1D�O��������<�*xߏu�X�a+���q�nY3���Np'����-_�*��:�����"��޲U��Ӛ��]�L�%\O�ɼ��ܔ�Djj��n�g���V	A���čh��W�$.�������t7~�f<�NC[s�N����t������ղc�vPeB���z�ӛ����NN�gCM��y�F���"CU\X���2��CSR��|�!Cdi����o,���ݹe�G��cҌ�(CW6@������S&�N�l3�(�,[n�v�E���)'u�Oln���
G��K=%�e���d���Ǻ��T�&-��@�}�< ���A�l��f6��elzb��m�fq=��Z�����\�ܥ��n�=�~T�>��^��]�����}c����4�!H-��S��Y�]�����鬓�����ӄ�b$�l'{�Z���_��]�҉�L�~{P�9�m�
��tƄc8p���E4��LT��;�-Z7:�T���x�wc��B}n�a`�V�h`��ʰ�p���K�D���c�ѳ)�,+�����(�}풃	c�$��2@�Ggg�j�4@�	�8�ā�L>��=�����_cc������`*�e������aE��
��R���e�n�[c^�R�H���G1�b{�%�k���8:�Ōff���m:
` ���K��iz����N�b�2���m���^��N�����E���.�UMw�R	��T����+��j�N��FD~��2��\�c�'�߿.��f߇�D��!�ך�ٗ�[bMﺵ�S�����A8�!7}�I�	w6�׊���v��ay!�&#�H�����G���V��ϚF�e��p��z��zm��fu6F�ɽ��k�	�%�f���<�P ��#���'�;[[X(�{b�@�ъn�,�kf�
 ��
� ��3&v���ц
��\�gU������c��ڥ�,�I�[�'^�����q�sL�-�Y�녎�'�$�*q�D�< ��J��7*��3�R�I�X�o�b�V��]�JO�n<��h���~a��0A|�kb�:��ג��5��i�x'�<��f�ȝ��G������ ������e�^�&���3���?�B�����5 �x�<Y���WA+c�'��/)���"C�w�\	6�dʣ�j�c�U�MgJ/�J��[�K�4(�����T�f��tżR q9�����N�_ruT&�o\Ԟ8����g�q�9�+k���2L״jF&��2Jt�[��o���%���Smj��l,pAm�~I��8�h�ܖdW.�j	K�	F�!� V��nT�4;�������o��1{�Y�I�f����;JP��سR��"�ȓv���hff��$��l�m��NnL38}2�7�4t1�Vn�ww�N��P-�����hܦ�(�]8�V���b/����O�y�F{��NՅ	���KP�|�t��eM@�@u���n�o��qk`q���P�i��t�޾��Lf��2tyvC�~���o"�酅�������0�,���N	�U�V/H������㥠��.�b�k���[����ȡ_���.4=���_�qd\�[��CG��5(0r#G�#�X�b��$�x8#4�tSӹ`�l�y�ө-"[)`j�r�p�C��:����vϮd10>v�O��Z�'!V�>�aj�-�llv"}7��
��hj�:�hG-������Px��8ޟdl�۔��dcEo��[�d�UM���RJ�$��n9I9���}����l���yS{l�7�����7���^�'j��>"W��P �e!���2���:s2cp�UT')��2�B�j�-������'�d�rhQFfW��$��W+l%���Ol>7zM�n�/ϛ!Q��LFh��7�"b��"��m��@l�H���
rA;���kw��4��}x�Ҙ��.S�L�:"�F&)�^ږl1�Ix��Ϥ�c��T��>5�юt�ȧ���9��S-���m�(��$y��`,>���Iw=���QH_'c0�7��h�e�į[�(Tqhw*s�1�2��~���E9MȹZP['!I�-�`!=Zf�0�?ԡ(�v�q�)�t|���,ȵM$�HR}��n��%��S��"L�uc�6�y��%Ͱ5��rHam��w?�"ĺ&�]2����u�AH��ɦ*�}[�p�<�������W��]��A�:��.y0lk�0�t�Xtm�_*e*,E�t��X�%����R6��QBI�7��{ߡ$(�6�P~v�ő�Åx�kEV.�JZ(�[*!B$e�k�X��7�3�����d��;7�)���7�꧈m+�$%��Aۊ�"e~�	����bJV���ָ�5��E��ϕi�����j���2������Q�O��v�C%JV$3kw�VQ�X櫵|����6	q[�@|�My���e�qzp3{���7�9U;�
����::�=W^����L�9tbN��H��Xu[�(�Lo�oч��j��E�w�
�
�0�cqkǱ�6�x�	�L>$~��.ŏe����j$C}�	Am��S�'V�*��N̡7��?M�n)�����>_�(��ﻡ&Z��&�Q��@+�9Z��I���^�y�顭���sf��>���dd��s��6�pd
�o�*��9��±]ݷ�_���4U2o��������{Sm�����{Y-����^7k/4�ǥ����#�p�����n���x���b"ymbV��������f~6im�;i�j�8�/iSR�3��g^���\b��)	t�b��G9�Ծ$�E�c9����[��hv�w�;�N5�5.�v0�l��ȹ�I�T�hf�-�R0�D:�诎J��
Rɠ��۞^�Ψ�~=���^89��s+++�-�܎o,��N!�4}�b�G�!"ѿ�T��`WZ�X�:����)�>(up�v��^��Wj�c�]]]��5.���6�؛4�遇Y%."ps�s��k1<��W��b4�/��n�'��Ԇ��C��H�'��V�mUF�J �ĦS�;_����U6�Z}�Va��ܳY-�P	E��7ה��/���~�c�٬�8�~!�~��DP�g8�:My��\o����	ƪ�3�ӻ��cb-c'v���0��%��o�<+�U���C�=fI��c_:�o��W,숛�W�Q��-.��9���o4A������w�ED�=<�E���|p�!�RoJ��-˶5�q���r�S���}��������h�<Yi)U{�v��4��Ŝ�Os�J��:�^�(x�tb^׼�2r#&:���$�&����֐U醮-QV2�S��Ȁ�y�N�ܙVh�n���6tc�!ĔMhK�w5��T1��F�u��%Ħ\��a� ;��z4
�͢IƬ���I�P�)(���d$B|ˈش�9�V�$�X1�q�@{�#�'uК Xs�sPO�����v#��R)g"�Tv�*Qjw�e �g�;|y�k��yԴ�Ք`l��4�1�@���^��_��4�)}�j�qe�t�o��r�8�N.wy,���:��
�K�~�b��*߯�sa� �F��̌�����+!��P�R�N}�����&8n������+k�2_�&����ӥ�xw���дy����KL��2�EK����WLtD�F	�܅E���l�b�Nt[d,mpy������,�]E�Vt4�T�	Vwdr�;��EdY���ߔY��nJ�;k�`EK� �W�:�#�ve:��b����-x��C�6�;�)l�N3Z1SN�~�n�(��iٌ[�0�^\�>)E3�HSfi���za^	g�K���ߌg��KRђ-���'P;����� F`wp��(�X��T��H`��=](���ʔ��΁.YPW�Gfu��Ύ4������:���C~Y�-��Q��b<^��m�z8Vk���P���4�-u�V�m0�*�_��д�;��5�<�-�p�Q8�X��ru:N��p�k�KiP���&��X&�9ƣ�,�Yo����nb]!Ŷ�I�wR�a9(���7�
r�]d���u�r�Խs�F�����AT�!qe�t��2ce}�6�0+����4Ժ�N୺�I0a�%�����;�r7�:��)��]$���6��V�6 ��Q8��>/��}����w��NO�§�~�y�8�#B�L�����c+2����o��m.�g��2OV���tWR-v��p��4�	�,�ל=��s��z��݄>	��ޖv�j)n���0&K�C�
�ʞ�7F��o�������m��O�퍯{I��¢Gw�h96`�2)usv�L���?t%��\��1d&�S�����6CC��}Ϗ�~m2��������D�E_/���|��� ��?Et��샌<7�Ev�׵Cz����VO�YcS)���	-����N�c����/�1���c	bm�/�;e-�*S�b�=r��Zp�"M��!�G�]v- 4G�"�Rס~�I>%J�<��,��=6È�$#i?Woy�vI�NR饫��([���{�q&+^������})h���Y�?��\@m�����I���ޑ4��-s�/:_��dV�B�x	�
�v)`�|o"������~���xYD��~��]"\B!��Q�ͺ�i�l���tM㪻>O%&��q;sl�oh�">��ӥ$LE]�x�����4�E�W���tp?^t���a����U����x��U�����u�5gŅPƄE��c_�����Du��l�zq7lU0���a��h@��6~��˫oY�`��"<�L'Qs��֥��#�h�J��|$��爡b����T�'��Y�����i_�su\$}�f��lr�vS�0,NBũ��Ѥ�U�E����	�v�f��I�>�Z��L����_m�vF����(W���a8�<�sl}��
���)ʱ��'h�	P4�'
���\9��\�3���v<�ܭ��`�����H����!�M]�@���95G\���k�q��0_	.�A��pՀ۟���4��̩�Q (�y�ˀY�"����İ���&�'%[���ʻ���D&y�&I'o={F˞�z�iNeN@7:��Լ6�}�@ry
�G@�f��4~�d><=���U�_p >��z�9�!��f�Ie�d?9���f*��ڗ������_f����W�p�(���X�H�	����XL"v9�i��O���sy��N��	���i�I�F�o
D�[-խXg>��{~�8a��l�A��IO���;��]��W	u�f�t�-<=8�R�o�nQ�S$��^�7���TJ���m�g�K�c᧎%d?�#��j�ĝ���������N�������؍��ҭ���s�+�Wl���^6N�*Y�I��?�����]�(�X�B���9�|�{��Yh���� t>��ĕ���W��wxo\8
�:S���!���o6�����FS�̷3�˂����>�gC��=7�+p��m�1�pt]��c"���a�"�BH�NSK�3={�γ�H����xY3��#�&��hD��Q-W��)�VJ��4bߚ�� DZ��646Fhg���L�aI�<S�P��`��^���<�D���O��j���g7��:z�z?� B.@sN��N	���ѭ�sN���=�����/�4+�!�P��f\'���"[� �������;��iM�?nZm���z��VSg��V�9�-y��M��L��6�_�<�<v�5�ʷ5+�B��d�>	��۞U~n-Q����[@5�.'E���v�$�k+@�FK�#���~2�)2l�.\q��q�SB�"�Ԉ�(�r�˥<�h�?dxJ4hI���s遏P�Ҽ����KaK@oWks��!kK�}||z^}Rκ^�U�~չ=���F_�#j	�k&,K��m[�w��V��|S��������j�܄[��U]M�s*|fy��zz�'s����20la�$��@D�%����jy��Ja�i��%.��2��s�)���W��j %u��Q7U	&(�oZk����oU����;h%��(A$�e���������7�R���-4�z�Vt7�2߲X��,8�X��Q�U�f�a�x܈��$�Ⱥ;ۺ���~N��_d��|�.��ѼȰ]L�RH�u�� ���[���G�iB7�����	�,��M�|N���B��lu�:Z�4N�\5��x02f���#��i�*�D������G/�������:(��6x���L
ۊ�����b�Ր�9��� �ͱ�����H����('U+
�')��!S�k���6����я����Z�C��觛� �n�S�~��I�Q�4/6����#}j+�?Ic�0�I2���%D�qt�I4Y"�mp��P>��Ó5����!0���UI9N�LB/�1׍D�Z��ֲ�U�%G�Y�9�IS�WU�D?9(+�L���~��rA�A>O̜i�Y�g��D��ҍ�"�~Y�s ��b�l׻����/"L��-z��j7T��D�~���œ:�����l2�ZR��?�b�(�}��c�w�ǌ�?���Ɂ�-��Eb�ɷ/���<~j7>��p!�����t4��H��k�E
}�F����B�K5��p�����ʄ��u}�ۼM�5)���b�}�[7.v������^��I0��5T_5F,k	SC1i���$�����8&�a>�ޙ��"t������+�QIⲒwm~~>��nA�z��L�w�bo�ЯoU�7��Vה؏p��%�IN�E�)�����N����%p�}@���`�"�B�K�
蓦�Q��V�z���p�����"���=-��eP���kd�O&ɥU�\-��ڥZ���H��&��M��p֎N���~�$ϩ��1���G�~k[��	K}�����C�jmyw��
�ęqn*v�Q!4x[��y����[����XB����cA���E<c֦~B�.�r����¯C���*!ğ�T�xr�(A����c�t�-�M�E�֋��Ƕ]X ڲ��u�r�3����fuS%�IV���9��x3�Ho��=Bt�`�m�r^u[���t��N)�,��h�ӹ�L~z,�Zg&�	�.��x�t���U���f��"wuE3^�<*hB�F�.�>C�r.�|��Yn���Gf9갳�$-q�H�-��U��Bp�`?g�<�v#�--R ��0����Dl�n51u�k@$�^wKD&bd�|~��ݺ"��A���26���+	��������&�@�հ�������z���Y�l�MH�/��4�m�|��� ��6,���ʓ�7�8Ǡ�DU<l�+���юa��zF�O���.	-'+��X%`D�TD��)9N���6�F��xSH}��۞�>���L:M�9݂�py)깬I#E�x���x7;���Y�3>�|^����a3� �w����?d�*C��^���#��x�(�9
�(7�*}(����Ej�M�?>|o��Ļ���{E�2�|���V�7�����>(W�?��2.�'Z��t��)�)"ҽt�����%�ݵ��.Hw�R�q�������r�s�<g�3�̌N6�"$� �A2�cL9�c�|�^���������=�^�=x�$>������G�ƥ(��[��%Jh$�CLKL..FC啽���zD=r���v�̀�~*�q�sƈ0L����e0�еٴd�{C��d���R���Y�L�I���?ԩ+�ǯ��` %e����O��\��@�֍*%7\]�l-=��-�l.������ V`�J�;�q�v����v,���+4��Ca� &� 	w��J[v]$���Q�����U�w@U����a.=h�	g|	d J��<\����w�tO@��Z�-s.b.�����"E�3�'��g�+��	���jt��C"I5z���}�~Bak���]���T�x�OQ���������2T\���r´�s����t�8Q>�?�H�E�ר^�[mI�����>C��r$e��C">@��2��j2$�k�Kr	��������~��j���|WB)F��:�� ����� @�K�4� �A`�ϴW�b���*u���(�^��������2O�a���+ڬ��Da^O��\Z7��j� 5�ȸ!x4����o���V�7��ͫ^
3A)��DG��>S߭�C�L_�2�v߆x��۷7�(Y}u��ٌXwe�7n�zڞR����s9m$�ǈ��-"�O�D�b�"T��y�	Q�2#�X�Z �Ԟ}@]�08gjsD0��)�S6�,��x+��X�~�5K��*P��c	�/�|+���=B�M������#��*����ź��*�=�{�k��U���j�8��z J���+2��v;�����#�ø
n	b4	��eN?�U3$�Na�H�i���q�Ő�_7/�k�,�G��ǵ��"�*V�k��p���窆ՃH\��bCw�FO͊���i�R���En�	��K4I��h�o@��;�U�1����G�q��OH�t������1P1�
�Ǖ"Q���Uv���Iփ�C
��]Q��v3"�@���X�x�+����Z���n�� �.$����8 #��m�t��k3rq�"� grƹ�kcJ/�X�i��os	oG�Wj�-(:���̂��
�{<�\��,�e�����o�������%<�����A��'�����q��g�u��Sh��nuLk��G��X#���!k?�@[%̙��1����4�K�A�ן����B�� �'fec	!WE���H-�8	H0U²UI�uL�����/�$
4"6+M�a��0�'ądc�~�0hO� Fx��H53�G�G���Y ��R��u��r�̻e��h�x@�N�3��K�K��S+Ga)9,(<��ݟ��ANMt�H\]?�$����*����C�A���Uj���
��v\�5K7���6�2��Iy�.�+��!�Rnz?���"z,K��\�+�WbwJ$�#g'�����)��AV/b�� ���v���+�I��'̕s�g�3Dƶ�D%vM��MO��r�N�W�(�z%���\�I����F˘=�:T�aZ��}}~�θ�'���ݚ��KJ%e���}��I��}��a�a�=�"j���ɵ���oｩ��6�ҹ̗2�c蹓d�.eH��(���u��9g�g#|l�D~�gl�D ��8��;Vg>�h��4���"����E��zM��}[|�F�����*c��:8��5�0������?�R�{�&v�L��yU9��89hǝ�g?O�<7�SÃ&�!ق1t��	��x?,g����R�DT��1�+�}X�����nbJ|���7�?.��<��{�\U�r�������+�e����@����I�<v�x�/|1}0Ƿ 2�e����i��G�+lT�I$Z r47�����HEC�s��C�y�»"� *雈<�' IcW�'���ލ���9C����Їo���-��#�gk�S������Q�4&�>ϫbw��ƽ�:�
�V�
jZ�]���I��K���;xG��62y4���m�[���o[T4䥠�RF�$:�]L�1�w4l~�p�J1�*K���t�*����G1�/����P���V.Ed��T�J��!Ϧ��z�i��$E���$ߣWc�ԝ�eD�91��0^�b��u�{.6D'f,.>��
�2cLX~X�&���*��~,�d��Z!��Qű�D��l���(T�ߟ�[Wug��ԛ��"����*G����n�`�A��.�N�C\|l(&+���_Ŕ���q:����t���k��a=��u»��㜩���9@��I%��LH��D=���%���4��Ո2�o�6y.����� |9S���9��a�&��z�)��v5#�f�I^z? w�=�>�)ƹ����<?������R�F���I�:z{&y]�ƚ�(oު������A}�_���e�����F����ܯ�.���]}?�o� <~'	���E��x�bjq�H�Ϊ���}�`��&*-��+hI��]`�,�WKX�>���?�qB�\��v�=D9ﻼ@�����0���{	�Ǌ���$r�}�)�b!��8���8�~�O���9�o�-����q.^[�"�������o���U�e�bio	"����&����NP!�9����f��V`,3�Ou%{��� ����
*�(�=��8)I�=��Z�a>U�E	����i�ud�Dl��0�
"��pJ�#��Ļx�Z����;���[?�)`{� )�����	&�|*��2˦|�p3e=i�1��4ȘʼU�����	�
>UZ"s_v�g�y����i��k��>\v�c��ت��ݧ��R��#v��H;�G	��q �Bg�߸��U�=r'���$]��U�m*D���~7�\��oF-�����n7����z]���PP'Ñ�*ۊ>#��d�|`p��7!7(���/ݼ��x��-�>�۽(����˫����6cQ��$fV&�&bY8D��b��P��։����O	;�F�s�tF�.�*�'����U�u�.�I-g���B��.�3��������*5s&jD��JI/S�qC'���]��'uTD>8�T�Ay��k�9�=WՊ@֯B���V_�|���VFB;��=����\�l�Я�z�M�S���[���Џ#Y�2��-�Bs�ߏ%ֵ�F�wֳ�}�]sc�5k�*�x\/XDN����+���9<���W~�_q_;��3����UDYV����
5X..�Hd��F��H�R��3�>l9z�v�~���[�ao.B]:/�L~4�"�DPP�b[�VGs3w?���O7U���ȉ�ؔ{`b��������&h�1��I�DJ�v��99��ܓr���2��������=Nb���Gڙ�NϜ��i1w;9�ܷ�}ec��|C�d��mךf�_�e&���;%�y�\������SS.s�#g���Ό�,I�����=�t`��~��2ظ�~�]j�	}L�����ź�^��Fh����n��_xD���\֎.	��|�^uRN�<,-hc1��B�s�?(�^nuYZ��O�shՏ���<�,�K�)�����C��'	��&"8N��e��X��>�L��[��@��L����쩴��M:������$�Sp�LgU�I!�젅&~nմl���V�i�J��!J������g��R��=U�%��˹��{��O��R��zڮ�റ���~�"H9��/,�7��"pF�kr>T~qI�ehfTL��J6/���W8�2<�d(�9ţ�kV�CA��t��a�pc��_�2-���d�`tſ�d�-R�?����U���D�p�Ĩp���b�j�xU��Q���4/�ެ�G�.��9�9*��;�[�2ͪ_&��#���>�����$M8N��@�ꥱ�����\�t��_������ � q'�ۘT9����@܍����Ϛj�ښ��O�/}�ԐG��hpi�-�E)r�i�4';qT,����.����x2"V��ycV���Q����Q�mS��9<	@Zi�/ѕ�V���mo/��GK�
0WL��S�}g\3}�3)D���A��!f!o�qq�����P�
��c��~Y!4�.��b(QH1�+LB���$���'�� "��x��j�W߳s��zO��̌���o.���Jc'���5}����KϔD[�;�Y����\����|��)$kN���N�����Ї����C��v�ԗ���^W�V��pĞ1UwАa<V��Đ1��%Z����V	�����R��	头{y.� ߄�"����J���z�,�{{�UO��6yR��s�܎��TSrf�	��Q�t����B���п[���8���/����p��1<(�!I�G3��濠p�5W���ϰkb�=2��\�M��a-L�<CG]����(��?-�) +l���Yr'�+k�,�
?��I��_M�L)k��6>��<]$M*e�vX��Ͽ8��؀�F}):�6�3 ,�%G�Z���=0U��2��F	��4���AţS�S�����_v-b��tpVD��O�]w�,��7+sM�H���Z2='��3`*��m�h�kQ��%��6��}@��
/i�.�V@����Ѐk��7���`eW�� �S��=�}Ic�8�8o-_'>S��_��J^K(,*����oC���	����$�j����u�XvO/ uxxP���g�a�;�M��';�ܠP�Pe꠫e�Mb
_�rt��񳹷̽f��}t<o�ϥy�/u�U��z4���~>�lj=�ͨK����C�]\�����<��z�O�h-�4806I_�����}ʹ��*a�ztɩ�V�̦k�1�76�0<'���g�|�~��xJ�XA�y������.��ڞ�[��� �l]����MN�Ͱ�����Num�Xƹs��X��7k�>0z���W�rml�Sw_����5��^Y�c���Ԓ�(8� ,5|�b� B:�������>�B2*
�:��-]���'�LwZo����:+,��=�Ń��tL;WAL���M�g*���2�c0ϱ�����:e�E�>n/^�>&�%p��T�<��Y'!BM��UK��Fԭekۧ��~�{���,I�/@h�C[!-����O�fX̋wE��|�����t6���F_���c��X@�NU�-@�p@J	��$�v=<POV`�Ɩ�6k7@`�7 ""���s����~���6S�z�
o!�ɋ���L�19�T+�(�Ԕ���`����:(u\�zɘz��eg<�=�S��qJ�2��Yc�o#���Bkd�`��'vP�3'(x9���	
�Y�<�Q[ו�O�ā�ż���g�����`�R���4��������hX1���[�l�����.�`�Q8��֡���E�݁���P��Ub�g�<bw	���~�� �E�sA��g���*�=�$����s]������#�g=<���\0d)R]~�ZnJrH��f	h�nr����8��U����FH�B�󅆊p�	���J�s�0xo@������g��[+VR�|L���'����rg}�S�&�\�Rr-�Ug�T��k{EçZ^*bz{�>��xZ~�x��i�����k��>�`R���q3<ptP��ٯg��Xs�sP�d��K{*^�Rz�^u���
r��(Õ����呚�Go�'$��r�|�������p�d#G���5ù�^*�{,�Έ�o��Z�B���flHQ+wj/p�����70��Djf��8)E��qE���s��W��UMU�?x���B"�D��A��x��P��<���a����-���4�6���>'�s?�(����-u��di���/����`@��왷����s+�3|b��� �����d��a��{,~]�@g<�f.�H�b(���+v���
��?7L2wx�:�T��4���`��� h�è%�|��sE��Vޓ����������L:�N�Pl��5�����!|s��=֯���E#�a�IQ��]�f�Ԃ�mld|ʙ�����1X+�؁S�4�?���o���B�TX�޶�E�3�،�x�A���oh��_��=�?g#���!_,��L�E��:�s �
�'a�R#���3��8*���l���r��=س߉\�`K,KU��j�i� �Z
��]n���tGycRn�G`ڦ�W���$�S<D.���F��o�#����W6�p�=~�l;���B�����2�d_n�!!����b"(C^���\�]�l;7�CN�ZNk��\��Ww�@�Na���`,��ϖ՟��=�k��911�Պ�/ψah� P�K_�CM�&���7�%�wݲZE��p���]���Y���w�18���rw���KSۀS+�qY0���He��l�HB���x�}���qzgnU�򧞎�G���p��D�%���\.v ���,�u^��!�X�}V�D���ǮWc,�,�t�*D����O"��_���?��M ����8~�/����]5j)��m�*go���U�CW�a,moiU	�N��HoBx���P��?���ŃQ���zT��ɠG�����Ԕq�`n�����%a������#�N9b:���'�O)�_�f�sQa�g:hn�D�
h*ʍ�bq|��O�H�m��������t�ϩ��r}��{&6k�.,9���	�fF9��fhɌ�*��t=���
�n+�i_�������fy����/�E�*�KW�Qq�.{�J���"�7~Zۥ?�-���O����R1�w��+չX�EV%2��3s���E�Q��P���!��zq{i���_Q�s��{��O��j��.'�k@f����v�3��,�����]*$ED����Ԍ_�4��%׆�@D�"�K������=��6(2��ӍB�ka<�;喪�>�a��[��eZÆ�>�󹞓Qw���kf�鎵�&<��V�%����Y	�O�|�����w�)���g���#����"�~2�q�E�/�~�+��K��d�C��Se�#�Ћ�}yx��ng��Jɨ��J��HX����<b���4�O�ճ����0��}�]ny�ݬF�UՑ6}u���5�r6���_��_�jwqv�|��pj������'�X�
��EJ�ԈYJ��	���'8�l|C�[�:0`}}�@/����^;d�=O���,�u3���OqO���
�i3�;zÛ�:��\�o;�f��G��3���%]�2��P��=�����=��|�{n�i�!���HԈ#+�n�vA�bv���'�vp�����ys�����r$��Y����wWˡR��\G�hae�E�d�	�I'p��M�]��1��_�;�m�qE^��74�}O8���.ώGd�d��@;t�1��T5�k���t!"\m�WhO�>j&ĳ�;�\���l֤�T��[6��\f����a��z�C�,)VY����	|q����im��o��i����n���x����hK����J��8jf����y�U{Ã�E����<���#���	�eoT~Ԯ]gg������te0�iU` ��XK>K����p�s��+������5��(���lIfg=?��vkqw��7�����b�1V%���
?�m���u��D�x��q��'9�Wi�5��!�����W�KlTYSŴ$��0X�� ���"0�tߏi������5���14!_�-������A�^[11^�i�W$���x��%��ь�sj����k��� �M��GU�g���_T�5���ص����1Bfs?������"�=�n9{f�NX>�� ��n&��b��1��<0�/ȏ����వ�1|��\�t竡Ԩ����	өl]b�Y���2�p��Be�LYy�D�3j+����A��\<�2~�����mk�l+\l�[�Y�|G#��3��i�Z��� ��w�Ȧ�F�',(xa���~����_͉"{=��r�D��!性r�*B�}�\��,,����^=C��ڏ��	*�du��a��2���8oI#�f~�	��
��y+�$�\��hR�J�f�ϯ��a&[�u��l��%��JL���t7{h0<$�r�8.hV�U�Ɏ^�O0���;�&���#�(}ht겉b��U�&�����?�"�ۑ�Q�nm��O�	�<pU��t�A��ѭ�tv>����i�E����n��\�z����}��xG�b�����ӌ(=�^�Q<hU��MD\�cr���2a�)���QMD�;�
e�����e��K�o����1�H�(z�4�nYo����)>��-��d�Dك��r</4�����,�V6	ZS�꨹}��Nq{�_%t�ݬ��ͷf�܇fnJ��(����}�o���qL�\�g%�|��f�o�����Q(i���-�j�U�Qq{߆��Y�n03��P��ViɎ+*��pP��z�fL
k�W����%v����1���92�Y{��-�%����G��Y�H����0R-Gck뻩�T�4M见m�D����$�9��������`�S��Ђћ�%y��)�`Ȗ�\`�jJD�).r<������q�o��[�I�(�@��<����Z��(�,=ȕ��M�r�P����
V�X�}|o��m��C4����?�J��W�$o�d�]!v~�6^މ.]��Tt�������=��ܫ��[6E�cխ?��_r�g�D����0͊K���H��3m��͜7%i��ȕ�480��w^����Pdu�mƩ�(��	�Ud箸R�j��s�g��Y	���փ8F#��3�t���x��_0�CBӻ�%6@ �	�l��x��� �@^bM��̆����I���jd*<��>��d#���r��[�w�<��T1�j�Roߋ��G/�U�$t E�ط��(?��"sbߪ+�=����ӌ���k��;�r�ow&(������!�g8('#���bmE	{Z?���e���t��o�S3� ���H,CLp� W���˩�*9�O$����?�p�˟fx}`���,&W}o�h��*��W?t�
���hi�*���/��7#3Z�J�+��b�?8��G�h�v��k�[F�s��m=�o���b�һ�/���e���R�Lm���7d�hM�z������-�/�P��Ld�w}��S9ˀ����8��x\:ԹMU����Y�w������z~���򬕙?C��)٬��>�$3���N���#ژ��9�O����֫�A��Z.��"(IQ���6$g�f�7�o�ait2a��ǉ%꼞ٲ��M��u֋�w~:�Wi��UΤӞ^�ݮ�d�z��)�au�'VA3�4��
�m<`���Q��v��{�8F����V8��5�+'0]�7�a�}�B9�O�5&u<d3�5�̷{[�]a�;H]z��mԃ>�,3�~�q���#3ʬݖt�L���֦z�x�����?s?�0g��c9����s$��Q��+���7KC�� ?�_�Y�j"w	8Y�w�B�J:ٿ��V��r�c�0������ܪ����ڼ�FWщ�K;�R���1e���'�Q����˻�x
@h��5�,Y�`������BR���E1���4�S=3���� BC�#���C.k(Ξ���"Es�/ј�5��)Ή�/���W���,xK��_�g%'�]���l�$(�����/`�Ë��f�����D�A�h���Jd�E�6�\�τq%g�h,kz?ΞM';��ƾ������:_��9O��G�ٛ���co)��#7��fC�����,��J` ��JI"�_���O6ʔ���zО_�'�\b1i �o�����&h�ZWaM[��Qç}���Q�l��X��0�Q.u���0��aGT(�C�b��`��%Y���+kvDm^O�9�YD�:�ֆKe`6�a����ӐuB�Xʓ���Y���(}/�W�����e�&Y���X�>�SE)I&��Ɉ+���Q�L+��HN��ף�rY�(���`[1��&i)�V�5���'��h�^��(c(�������+����8(.0����K?��X�)n�!��*¸/��T�����K`l+O��H�|n*.�u�U9�O+0���PB�	��Я�Px�Q�@U_�	Zű���t�h>\��y�T��En</����"�2�?�[2��=�4�}믯�}�G^pD�ゴ��	���^H�ы%�h%���\�p�d4�Gq�����0s*x�eIc�p�*/���1��|~6����=�pԾcҳH�*d��f@��H���C8��s�CU���F|��,�+N'�?$�9��^b�xK;�H��1���	wǧ5������w]-JvX�Օ������Ww�xf��)�Q#��O�!����!�b �q�闙��"��9��l��̑ue]~����L	���ncc��A���I���N>	�yM��:����~����;<-��Yfᒐ ��ھA(.ĳ3��GS2,��s�{4��K�F<�ZB��������AqL����F��;~c�V�����(@����g���V�*w�ϫ����Ֆ�p�[����n�C�s*�Uc<�H�o�_��9���9�&�iC��O��g$�8��_��v@L�L"5x��� ?��5���W.��A���<O��;-5�}��D�U@��������<0���q�	�nJ�c�l��y �]v��_��Xˮ�<F��A�WLv^��2TtD�Q�_H��h�韫�q�����D�5j[@ܴ��Gt�Aq�
Ì���4.�<�ڨ�j]t��X08��~�t:>��{�I����ߨ�y`��u��n��9������mF��QH�R]0��N��T|�⿪SG�ۓ���jΒo+��#���َLM\,XR̦G���V�`�]�l������~���.��< :�}8;��MC�*�t����%_�����o���dM$���׿TBC$8�_H{�4�d����N��p�ucX��D�.P��$��8����<��]z�$h+dS��RJ�p%�.��/���=/��F��d4k��6p[%+�aC�q��o%ݷ����K�$x�i\̵$�%IF&�c�s����(�.#�+fp���	�ߢq��D_�i���Cyy���o��i:�$	�7�.��ݼZ��1 �˙���n���&�$'�C'Pr/ۍ
�2���iU�b���{J��
�%�|��y%l��j�/��pX��z�8b�<D�	�S�"{���x0��r	C�^��U���ܖ��I�^.�憤e4Vg���]�h�M�$RL���H"�sX۷�;>� �µ�})� ���Y�����m�'�"s�����T�N�D��k�P�罫"E*l��I1�R���N(hC�^�k�ɾ��S���7slB^��G��z3Q��iB#���a*51L���Q�cR��?�c�$I� Q��""���o�f&a�KQ$b�F�S�	�f��vƇ,s�K���wr���bgc&���[�-;��E�^�f������ލ�5F;̡7���Qx�³;��!u��?�ѣ�\�k��?Ɇi���s�����%ȳ���ܹ�Ey��߁H�a:��#�Ş���PI�f�r�Iy�'�|ad@܌D������ʳ#W�`W�l6��R��j�kӲ�v����D��tJݘr� $�m� �V�z �kp\��8� .�l�O�o���;4�"�-�U���E3��y��jeL���n}�΍ap^�}�Q� �T*S��v�`�<�#baZK�8?��w�y��j� �$�ڠX%,�L�[,_mMO0��p�[W$����x%��������Wd=@$�v{��0��խ�AX1��j�H7���. C���K*y�RyW�P1��e����� UGPqj2�C�' �=��aÚ֮1�h^�1�H�2z�߬���5��d^���2N����FX~2�&`Օ��c-��ʒ�O�AV�K����#�W��}%��ܓ����p[�D�s��Ա���AN2����׉���]J٢��V8��2�	'��G�w��ߋʹywV��+�l�B�~���m�Ň���}�p��p�bۢ�*ÿI|��qTr�R9I�1������(�ʢ�H�� '��L��{-��!F	��xxx�;�%���ϭ"�����,E C�wƋ�w!�.a�m�����M��p���Q�c��?��F�9Ă�5���	��*4��!����ˢ�C��~��IF65��Ѯ����R��F�zÚl�xE����+��O�xҭf�?�l�ߕf����� ���^ο��m6�3�]Y��Y0!&0p���
��m�	.Q�RW�O��o_�������Ɣ*V���\@���@�`�o���c�r�V,���HL���&�m�1�����,�|G6CF�h|7'�5J��~2�dN�	q�!���f!����|~��j��Q��.�[%�����˜����;j� 9ڪ^m �U�d:(s�0��'�A�o�N�?3�qjZ+��V,2Yػ�^�W5J�I%�����b8�=�R�X��A���sd�6)���cI�$��[
i�c�(�.�=-p�����\�gi����<�W��<�S���TN���|� ��<��M�]�m�~��s:�ֱ��ȘБMyf���x*R�(�Q�Y����K{N+>AY-^8*`�+�8�HC�&۾�7u:�ERK�*��>�t�XS`K'M"��V�8�5�U�"�A�c"=�Ѡ�4�I�k�c�Vsi��NZ��y��R�ᇛ��B)l?��ę����r��}�T��c���g��IT��q�FRR����8��?���n�y֓���)��v*"ֱ�]!O�����T�c�j�މ��&�xԉ�>�]��>9���bC<�� ��H��~ȇ���(�_�~�F���,��ԩis� �,|�Ł"��8�۫��Y�!?Xq��dY9�{K��7U�Ʀ�s��w]��P'���C��?����"\к.LA����d�>��ڲ�eI+�>"C)�'���욬@��l:Fu�ph�\�oT�C�ǘ�F����%��ԡ���MX�=��L�n�d���m~&f�t��L�8�-'�C��I)��|��KB/���Ҷ1���)C�f�)Ig�Ka�����H�e���VF�R����^k�mG�.��WF{��q#��F0�x(9���9վ㩻�����<�aR(s՝�����G��8Bd͜��z��j*۲~EV�����+/~�a9�^X���jr�BI<�$��^�&"�P%���g�v���f�E�J�Q�5��!�&{#l�,J�]w���{���b���������I���LQ~7�R��������A��8�cvcֻ�it�5�r aDՁx���l�>+X�Y�d՘�Ϫ����fp�	���Z-z/�� 	�7���{�AJ��]r��h�<?s�9[/ӧ-�rᏉ����P�A��� 
.�PK�k��-"pWj4�rm�qz
�|���L*_�N؛��YA��K��F6k:�:N˃Q!�_v"��lx�(��O��F%��Z3}�~=1Z�H�#����b��6��n�	�X]�-�n����d�i�P1[�qv�����n����ͬ���w��k<�8�n-�@��g�Hē��٫N ����w\���r.>�K�	o4nsA W��$$��ye��NtUS���ؿ�߱��������d�^�I��a��!z:"M 	(4틬ͻ�Y��@���|W�;T�4��jV�^J�pcd���%�H伤�z�Հ�@�g|�(�Գ��z5�ɦh����y�����GLIiNI�Y3�j�1��{S%h�3��ޛy4��U`�N�U�C��B+k��c��	��p�qP���_���h����=���>�]�$^x�o�ɒ�Gn�dk0 m��a�yд��$2\�U�����;0�p����/��`4��Mz4������.V�� ��f���	α����i���C�G��ǹ��5p:]`;:�#��aw�����/S�r7�h1����}o�%����v1�a�~�-���K��G^�޲J�=��ެ^���Č��i�Jy�	�#).J����|UD|d.����]j�Rl2�FŊ�4��- �}pM7���~��xu�h5�D��#���ۮ}���s?���W��j����A��^bN�X��b�����S�H��2Ѳ����`W7
 ��r��w!�6���o����� #���x^�n^�}9��!#RzD�fڕ�b��xB���J-R�)ي%Q��2$~Q��]�A�37?�A�ل@�3s�3�Qu��5����
0=wy�j�'(�&H\�'rwH{mE2~.�֎���!q��+Pܫ�wq���b?�:G-�^�d�����|ڂѓ{��a�W�h'�U��$������ue`���k;���L�-f�e��'Cc�B������G#Q	X�>����~�Z����b�нiDd�}���*߯H���;BB�� o�;B=�IBs��%��+k��Z���w���>�\ʑ��M�&�b��:M���}��h-B�,h�Լ����-k+O㢷�O5;j1��#���tJY�d~���,Y�,�c��A��Ha ������>2��pa�ȬԾ��C�&5�}��ZF�UG���-�7���ju��<*�^�v��u��7�Zm�r&H=�Pb�=K�X�I܊Ն�z�@������ջ��� r��-\���@��]��
\��3$���dl����j,Y�o�P�_�%JaX�l~�����-:B���O"Ξ<=Oj��;Տz$��� ��V	�I6��TS�݌)���K�G�%_K^I�!�������y<�1�p��-�$��Ά�Tw�Zx�����#0b*Ce!�0AX�0g�j"i�!�W]m�h��O�C/�����LUWe�`��&P��$l9�!�ٞ����f��+�G�P���ٞ%�K�&�:2����ئ�O"O�����}�8��>lҥQ���G('{isLi���/A
ƾ�Jy�ϧ������m)�8j��W�ڻں)��\L���߅P�-�h��\x��f�f��eZ 2��Ki��,�]����&]3���?4�D?�6���[���%�Z4�-"�ʾ�[�*f�k �RY�{�����i�5��:ہ��'D�䅲3Bf���,�.��aўs�G��YU[��� ^|gO�p�re��yl��"P���
��Ȧ�px���~G�1w�4N��BW1!���^tZ�����7%���D>Q�����逘���5B��U/�E��¿�۶m�4f����!_��@�<�ؘ�b6^��wd��ב��|�@m�c���~�œq� �﹎�糠����*���P��xeCx|s+��ڄƽZ����LYDD�~���*��߃�����'T�g�݂��K$ �ebk�7r��#a��s������_)���C�ԋ�jH������/���Ь"�DG����1}l�~=	�'tY�sj5ҟ�q���6-1�B�sF�<��њ1�b.M�!T��2cm(Mu(�E�8�����hD$��S�ٺ���B�2:��-�t�2V���J�p���Em�Gݟ�ך�7�w/��s��1���o6*�~9�ѡ��S=|��{�6Q�!%D(��v��a�3œ�-���}z?��J�����%�h1.P���q�C��Ԃ#ٲQ���d��eH)YZ�|PL�D��oV� ����Z��Yp|9��_u��.��'c���Оغ��Y�������kyS�E��k�V���A����T?U��ԟ��On�J*1�)�
~?T��$~O�	��Y�tY���,��VG�.��d�����~��/�[L�+�_���9��ɼ��m��Jɽ���αܐ��$�L��`of�5�k7őA��p��H#r�f�1�����s�v�<jj�M���4^t}�y2'��^�
$�uw�7<Đ�պ���:'~���X���*t����iғ%d�r�,�(�c{!��������x^��.=��)�o �M ��V��	$����-��%ů�	R�U���l7!m,���1�%{�29�n��� 
1��n.��Px��P�%�W���k�L�NS�l��ZJ�;U�b}�]V�ׅ�Ѱw88�6R����}n����N������DN���B1Y4s���+<eT�VuTngS!��8��S���+���n�4�����ƈ��\���l-�����A�g�	6�9{浄�D{Z�����EH��K�J��A�ޕ[�>�p;<��w["���J)$7O-'��~2#W���\1���g卓ړ���h�[���-�;�l�aM����!m�:�^�A,�����Jp � H@��n�B�uX�D�z�5_�у�0�S`$sy�:;���b,v&�@>*�Xw`�#�a���)���ղ���U���ŋ�h�\h��F��`9-Z�Ⱥ�R�̂E+i��Vv�1SE*�(roP�w��bA�s1����3���g���dĔ/z����=�����l�N�~�KO��xF��;@�q�ӯ�F�6r�`��23[�GV�r��9�3���f;=��,߬N��m8˿��E�(�45��BO沾��e�JZ\*_f-o�Vv��,Y�L�l�C�E1]od�M�Ȯ�̂���@�0�{q4.���|Tx�4f��m�]蹗��������������#*ꤣw*P8�Ut4{hLc�n8�Rk���ޚ���gblx�8L�VTQ�9�=�o7��L�z@dpΫ�4P�0ҹ<�)�BtH�BD�L���f6�o�z��s&E�����q.m<�d�<��eG��	�-�l�;����	��l�# C��w]���B��9�=o-\��&��!�8qN��4;�y�B��N�m��0=r8;I3�IiT�,q�@F��u��H#��r,[)aT�UȎ���t�5��|)%c��#�p�ۯ���2:5���Z���)E�!*�0�[g�\g�EW���v-� �<�ˣ��м�W�듦�ĩEm��R�U�9��m$��������MYE��pL�5�����z!�{�u��t��k�.�-eZٹIY�eLZ�4�/�s�K�R(:��ZO�\~&��`km�L������f9EeT�X��LZL�
�0NC���,;C."�h͜����ʛSi�%Ʌ�&�e:�I	��}���4j� �t���\�\���k��	�w�������g1����a�1���rG����UE��Ƿ�ׁ�*zT���vt�9R\)�v��@Xl�Dj�xW���I�O��0{�J}��o���s��ہ��Ut�-�9t�����ΧDzf�R���$��(�,.h�"P�m�s�d9)�8sԪ�ә���Z�RE�r�u������P�e[�rrl�  �y^�{�ǰ��h��<�\z�RX�[����YD���ף�b%a8�؝h����6�L86~1�w-㘲	-&&Jcz~⌳�� V�aR&j���Gut�u�М����G�) ���{�r�<e�Vj��)밑�F<d��K��U�|�L�l�Þ�B�FWu���[DL�C���m>e�-h}�,�5T�}���i�1#h��F������n���z���8�1aƦ��Q:�P�Yt	���]���֭�**uQt8H#6H���t�7��!.�=��f4��l�2$DE�/�,!���@ey�4��U�+�e�������� ��k"	mI��=s_�r�Mi���Dy��m�0~l���k���C>�h)���{|_6?Q��˖���)����.ޗ�3����Υ���E��GM˰�X,��~�J��M�������ت9w�������w����Q�����b��P�#n��{�n�^v�[N�·��9.`�Iϣ�hU��%R\87�KiUk�.��=*5{�w\s:���;
���06�41l��D���`N}OtC�c����轅����h��{��!CGw�~~ٗh��ǐ׺�l�=�t*򝙼fs����k#��ƆEa����^~)9vH�`0}�����<�Z���o/�:+G���-v*b��91� ;�X�h�cC]C�3;�A�f���&}0s1��gh��֒��$��d0]p�i�-,*zp�1�~�̀�8C��e��N��J�Z!Q�G���-�-t����Z���&���?~w!�8z0�q2�d�ݙTZt7���덞"nW�dJ?������g7�.�<[����&t���6N�_ v8�qo&;��O��r���K�#q�s)��pyL_��n�?��������ѐ�)2uΔ1|@w؁���pH��St���j+����o�_x�����qޭ��J�F;*�����_�y�n�ڇ�6�r�5Z�	������E���I/������T1� s����Ш�3��_v��]� �f��Tt�E��YZؘ�?�3��N_Ы���_qm=j��&vvء�7h�@�+v�b?	^�v�"}i��&v�1���~�f%c����ΣA�,t_eǶX�p�+��E%-KUTj}�\���,������`�K���=,��������x՗i�����7��G��&p����4�#؛�|`�J�.��v�/���_~})5��V��G�*�+�<�p�!g�di�DaH;�vְ֢���l������w+M�3��y��4�Τ.7t��Q&���{�B���C`P�r^��1�y@�bӡ��
�]�s�/=�o�q(���l����6�N&Y&���9���(EgAcG�+lW�Q0���o��K�GxWKr�b]$�����9O־{�4��!��̌���O�<�h��}����Fa�9�4�@�m�@�?^J�����*zM��8�~�a"
m�[T,!�=�Xb�6L1���W�ZB)g8iz��<���l�����H������+�Т�Ki�]wA�,����0����;b,_���	���)6���H�]��ؓ�xn�2����Ɵ�E�ޜ�:��'��Aƌ�p��X=�0v�fg#`=�7�cOO�_��	��ޗ8\�q�H�6ۄo��%C����}t=����$�a�T�xp'���;mI/����2�P�T��z�Y4x@J8�,i�G#Z�E����d��b��}���Z��q��t�?^Nxo���@�{~2m��@�x����,����Mg3�����"�u��2N��y ����P}}D[�E��5�O��V@EϞ;���O8�����䋼9�YG�<�*㑹):M�Ɍ�b/�������K�<͛�${�rĻN�qS�c?���:+<3�m�������b�LStLW�E>e�����3;�Cj~��1��@��+��#�3o8����b!�&�e��aҲ�t�ew�kSf�������~j<��4`�`jm]Ei�9�n�!6�"v�,]�5#���Ɣ�!�?o1f8�2A�3��z8��}i��G�ج@ib�/�� 7*�S�9��i��<
X;L{ -X�J�^~����>�\{�E�����������(6����u�<$,��| F�e�40��:���	���yG�[a��ْG�Q��W!Z�0FL����-�̱�&����.��4s�*�۷%��wfӿ�;�?pwr��l�9�B�l�#1*�}�lQ�b�2x\+
hĈaԚ+����@r�n������=�wa�,S,G�RHC�=Χc.���/�B�L;f?�9e���e�c\�$^�b�b�@Ť�k��e���?x6"g��X2\�IS�9G�f�.Q��Q��'�L����ל'j7����~���I��a����G7A�%��8�خ�&����g��?�C�*��9����M/��lA���ˎK��H��1}?J�����_��&�����HUL+:d��):��Ȍ|����{.�[�i*�+Iˤ�xVC��(�(�F�e��S��7v����8B���ͫ��f�%�1)�-��	]Gk�t�ee\��dk>�x�>������w���[�C�eG��|ˊ���3�B &����X��}i:}����X�В��]\��Y�(�θ�d�ev�M���A>5R$�Q.U��6 �-Щ_�G����;��9��Y�'s���= �}��H35��)���Y!���g_��<���r�C�ި��!�8uΊ���u�L�Fn*`w�s�ؙ)9.��ak�j�N!�uV�3֐6�h ���ӝ�f��\D�g�S|��1i��cH'�a'C�zu�4��w�Z[y��&N�M-M���v[Q�i��ʻE��4���^���@2u�}w����-�g����'TuŚAg'��Т��E��r֋z��:j��8�8�B��<96@�b`ѓ/�M��i�D3����h��,��x0i�AQ�9��{�`m�z~3;�E:��}�'�''R(ځ���+�$+�Q�j���c�>v����w�t��#a�D�2w�}��ߞx�e��rb����G�7HÇ����Ʀf.[�b��ޥ�@��s�G�O�E�?pWz��I"_Pt��o�s$m��P�C�<�"CGWtγ cl��+>�Qi�iXnc/L����S���c7sR"J�
���(�{`o���6�}����M72cG��B�m�(:I���Q���kh�I���tӍhΜE�`Ys�@EW9��=h�v��9�ie(Լ��"J�#qi��a�y]_y{:�����CgƼ崪��v�=;L-�E.:��Mg��f��_d�,_)�X�"����mz��wJgR(��~�(�f��"�3�D:+��锸h�֧(�z���;�� ��n��<������<�����Q*eЖ�7�g��(�*��`���b.eL?��4���M��k�Ԭ5�O��I���`�Ie2�c�.;�p����KL;��H�-9��ޗ�7�RX�^{k&��lc��1�	�Ե =�5�B�lv���#/d;�)��͘.gޟ��tEW�{���c���gyA%;������+��(���*~ؐD���S����|����sw���M�d�bCP]ӻe�;i�¥��f���9�fcK�e�Ub=M��(��Y�C�Q$/�Ȉm����JG)�
���#	2C�D�W�`��bm�
|���`�x�ٲ�rϿ9����sdg��)�`Z�(��a�ǠPϐ�5���ToL#G�aU�[�'����.���{��[YƲ�Jk,S��C�yj1�~臢r��ޠ���56�+�gp��<2�^zu"577�����-��K:j�x���8�00>�k�=v޼t�b5C��i���YsL3K��@���+�b�d*1� �&��syz�����ޯx'�o���ֻb�G�O��P&�l�r��L����g���d��{�!��&�'���D/��Q�X���DZ@!/A��6�)�<Z���y��E�W5�o�7L�^��Z�����{����'��vdl�E]s؀/ո�%�FL	lW��9��.�:'%��0J���b������o��� $��?�m4]
��或qҲ�92��֬mQ!�чs�@%h��Q��̜���5��c6�ZA����W -m	cJBJǎO�9��s�a��C�{;9�B�s���F�F����Gb.}4�{�)� ���)�S4���{�2�_���om��(�tp��-�\�Xw-�ذu����2L��4eR}�����g�$'Q�<(_�r����d:���&=�)d'��¨@^�S�j �,Г/Ϥ��;����kg�.;lIC�fXU�d7��<u.W�"نN���A�uj�=�nCϼ�~rE��M��?\�i��2�n�i~�FP���o�T�ä�}���N"���hw#'%��@5ۉz1��I����G���y�#���?��.0�֛/�4g|`�.�-���+v��FK"��Ȯ��{������^��Ea��H��#G���d�&o`'�I�:6п.M�F�L�4Z\�����7>ȿ�?N�����34m�v��b|}}��bAt���i¸ET�����m���h���qW(X[L�;�aa&�6�^bu���ԐBDl���ј9k9��ǅ������描д��d;u<v,2d8Y�ِ�K}�1ϸia�6���X+`�m6�tڡ������3��4,L�D�fyʘ��4�����ϲ~�NЏ�6����b�s���"�(K�)��b�?г$
<�N4��g�P p�~�et� =�ȶ2b���h�T��%#�:˺��Cn1�Z��7f�·�Ƌ��#��̹��/�[��'��4'�-�2Ѝ��U\�y��K[�B��Ci�bC�D�p�\��dia0�乁�2��9r�:\?L�q��]�{*~�kG�x��7RS��g�`Zl:�.S��Qar�x����o}QU�(�����ɶv$8���"ݦ���zcPʱ����)���������k�N-���(v�c�r�=š/ʶ8֨>3���|t56��Ƌ�+j�?����.�[��3�G�A�7��y�I��S�7]u�?��[�ϗ��.�쬨��/��1�?�a��o�(��c�
�?=��J��
��ȃ��1���)�,����ٴ�����QO�MKѹ�L�lh1�lXX�L��o�^�Cf'G*:����'R�귮��^��XdŘ'38�hyK�(Ӿ��a�y��z���ň��������M��ݱ!�ٴ-�pHm�d�ܥB�@~�ӋoL��zfK��ӿ�n�`6�"N�V?鵂
�'�:��16Gc�|)��e�����Z�B�j��`��$zA�6�t�������
}�I�ׇ_��@kwL)��@7E[8T;�a�ΰ��L&Rc�4j�:�-��b2����pvBo�N�S�yk]�5��|����	�˳����Yyt�3��i��Ȫ�䴀�S�.ՐS�.�o�@�r8��.Y���qb�΃�@�@]%&������6a�}�(��h�7~r�,�o�!��HEgQ�x���S4u���K�!?�.YC'�r̸������=J��W�F�fi�b}�晟#=v)�M��%2*zq���(��y�[�{�t�K��EV�^BϽ�6���~b:�ePT�������#���g?8M8�ZE�?������,;�I��q,--M�?!e�u��B�\LϾ2�*��K��s�����(��ʪ�l9N2����i�V��>��KE-���?8�b��`��L8��TZ4D�%<��:��I���)�飏��s��?��^��"v�1?�9!��P1v�9LK�BS��8/��׎�4S���Ґ1�7W~�S�'/�r^l�� �T�0
(�j(��,Q\ L'��|}U�R�3v���%oE}Ȼ���]Ay�=�5��亇no
��,�."��"[��.[�]�7�X3�3`;��Ͽ:O�J�	�i�ݷ�e��!�a�^�b*�y�u�,�b'<"�a OU�S!��]ϑ�� /�ŋ�1}p��ec��0C)+�,Z5	�"n2�f�)�u���R%+�~�";�1MQ.�Q��誛���V��\y�?��4�[�U��[�S��-�
GåA���A)�f���e�m�����|s9��\V�S
�O�wq�F��鉪��0u���2$C��"y��	[淮�͒�֓��1v3�E���=���ʟ��6�Y�8����l1�*p�)Nz�)�F�z�l[��䤴ª��+���kv��]B9�=GK�;<��c\�,c�;����Z�$R�x��8�-�C��;�Di.Я��	��Tt�f��S]&�BK@N�XG�.�iK�n��ӈ�02h�si����_Vh����j�L�V�'�m"�ڄ�]�X��|�ޥ_*j���ޒ��NZ��Y'�v���x�:}�����wX_�V�Xx}�,
�,9�b��e����Cn;�Cv�]:x��K�T�(�t�~�X:�[�����)��D	�2)���,=��GU�-��_D�O�G��)?]ጛ�A;��!*'��"�D�xt�Wt�_^v2�Q#����655�by��Dtz?E�� v ��wE_��p��Bs`�E{���ٷ��*@[7��eJӓ/~�Ȓe+&��*�
.��� ¢��Q�3`����	(�b�f������*}�Z��y�I\h�P}�jjA��H���S
����豧�#�NUr�=O�Ӷ���ٱJz��+N��kN=�>�=h;�N�_*j]3��S�B���Ɖ����%��S��Z�XWL����z��������B��]~v����G1�3����e��<���ШA�Cu���TW� ���U��ф��Æ�e����z.�a��"�ѧ^e=	(���Nf�0ty�|1E\	˰y�C߼���U�t��'H[�ٔ�&��#x�N��y!'��8KŢON�J�^$����Ql;�ٳ�������p�U�v�|�Y0w�ۗ���S���eEF����&Mus�2;����4|6��ˤc�؏�1�HT|L!3fS�b-�FR39��Q�D��ޥs��S:k�b�����/�t!|��T�1O&���
��2�u.9>��Jv�Ҵ� ��KE���cJg-J�DE�'���7Ywع�#WT\i��OH�ߛK.��JKΥwߟAk���%�u�"��D���n�ȏ,��9�Ը�Zc�!)2�f��u�M!����>�G0?� �<;��'L���k׏��1�Y���H#������)��<�R��C#4h����Cŧ8`�h��g�'#^E�Q=&�x{�,qJtS'��4ݣ�W���8�F��s��k:�D�"�I��sY>]�I��w�����'�yQs�w#J�{��7�xf�#3d��Ǳ_�)�I���`#F�5н_L�����b�ۤK��"m?f0g.��mPǶQ�_"{i -�g��y�\�ڪ<�3���D�ż�\�I��!GE1�� UL�ا����a � 1P|0R��C���":��j�W�DϽ�i0qʇb�k2�7J������ȡW;^[�A�����s�mX����1��Q>'eND:ˉf����N~T�Lyo��zJ����(�8dW< J�M�;h7< ]��B�"D�n>��y��"� Ei1ݨ�kz(z>��Չ�"�G��P��'KO��(�Fv髯�;����Fэ()����ϗ�3k~�0�
6g�n䑙aC��bt��i*u�ӄ��Z��)�N�O�u"˥�m�����~��B:�HGi`�,��_����Vb�2m�XU`'�f�Ӡ`�8j���;]�M1;\���^��E�q�{�+��%gوʋ�
��A
Q�|j�$*x1=��V7O��>��I�*��©��\B�!Сc>�Gi���y�n��>h�3&놔Y�� +[\z�E�s5s�#��@End�e�Xȶ�aO�|�	�/�i�gܹ�+�6���;�,�H"[�KX���zX6��/�i:����3s9�u��eނƗo��'��Yɯ݉r�{�ez��|�y�0�S���{e�G�eD�k��<"��@����B���)��5�(ǩ���9O��xn�̘���;�������6����8F�x���B�%i��S*���w�a�!x��7�rN.Z�В�<(���ĩ3Xz�9|�B�#��OZ>�	�m�f��S�o�`:m2| �uC�%b����ʊ���ή��%���p�|�/�*�+��v~�`�v	�bR�1r�N\F+�� %n��<v[��q[g�Hl�)���7zF�C�׭�f6�|4��
���f������e�T>\��� ʒ�=��Z�j³���b!�Z9�8�ـ�0rEW@���e��]$Sj��\4��������&{�C�d(B��58� F4����[�<�;�N�{E��Yj0f*q00Z��ȣ�Tt�Z�!��
[�0X0�{�L$�/X�A��"5�ձ��4}΢�����y"�@�+����k8��i!�4T�#�fؑLz�ű�& kT����CSޯ�F6���^�z����F�k�X��d &��q�Ѡꦬ�T��n��؎���5��
T?���W~aW�X�0��e�����2ؖ�]jjY:��Ƨ�������蒾,����Q�x�>43o����.k���hjV�hYQt�p�0~�s�gDa����L�qD��,��$E��ug쪀k�bL=b�t�H �t�aH�����q,^�8�l'M��T�p�A�
3LI�4��46�xߐA���D��'�;$#�L����c^ә:jmm�l��^����M��<�շ>"�qD^��CV��;�|����E֗�ا�~�n�w�	9�~@6PA��匈�����h��o���F� �r^���M��c�q8m8O����u��$,��O?��=�b�A�M=�yJDE����(�Fly,�\��T�u������xiӔ���i>
�����!�#޻4����}�A��,%?l�+���4
y��{�OE�3��mv��u���X�)���}v�ߵ���e��z6|6�V�0��H`0�\�1yviK��)vV�j�S2q!�b�e;z�2��"8������~��v6�h��Ft�H��Kc�\gg�B���0������ȗ~U�,Z�B�BA|.w�d>��O��aL��F�6E�3f�p�'�a
p�Q}���)��І��V�����xs
*��oؔʤ�.�-.g��|[�ܱ0���Z��B��/|vg:�]��b2l�Z�f�����H�XW�l�J�m�i]E��\c+�gƳ�����ǋ�������A�#��,�����ʄ7L'lT��.c��h��dw�4i�e����Gi��.g�*�髧H��UM��2x �\���d���j0ʇ�g�h�膎9��#�$( �F^D��V�����x���C|a!���w �2�#v�cӢ�K��K�.�)����8>�;��Ð��Z`�ȡ�-��pO��	�
�eƥ9s$�k�|�Y�-�_$;��N�Yw��v�9]�ko���/j�f�9�����������"?l,	�K��)�D�6z>��.SO��`ի����������NE����%ђ�w��k���[�01`�D��"Mq��!V�A��%��a$���$�ۢ^�^�bˤPT����<]|�Q���!5�o5r0ivș �Ӆ+��N�f�4mn���KW��8q�#3Nq:D�!���	�5,�7���Q��jg�k���D�"Y�T�~����fX�<�b�f/hI~PC�����l=a�YL�d�aܡ<C8���)t5�q����v�1:y�Kċ��aǢTbӠo6��-\U{�͇���u����;G~n ;��N;�z�і#��~Q[�&�z�`���/P���B�TbF���)r8Oɲ�� �,_z-���a8MN�X�sZ�� ��5���=O����fYUw�0��j��<���83ּ KgS�z"�����������u�n��ʴ�ɲb��7N)�ܔ�!�]��N��� *4 ֨�onɉ﵄��m����u6����
R_�HF��3Q�q�УB���o���)�^dz }�.��4��ꧾ.�����u�ŉm�b�9⭭9�/@�� k�|��$>V{1H &?�.>�|��e�g�4�ö[&�e�t]ڬ��{aK�[�Z"���,[T�"�対�������A,3u���Yr,[���ȬE�]%e9�	Oَ誎B��Zx{@�]{nMf3�F��爐��+�V�\����X��\^��4��4��'T��5#c\A�,Hy���j/�����"��l����IÌ1�9j�x�������zH�#�I���+_Pq%^8Q�������eN��k�k:'��>����d�:z��C�S�E�O�1%ܲ���`����z�w�;�JE��>��{�0��xq춴4���Fj���|?�t�I�VtB
Ծ�� ׏�)�i@Ʀ��~�5��+��c�l������p40��p=O��J2�4D�Q��LbB�HG���X˖�Z"
�8�NP�Nb\=�/٬�AR+H]H�M�.U���c)����%���y	Ht'�L���PH�M?9�FOQX��r:$� =�nX�J;������z�ߞ�7��K"��G9�}K+�0������k�u4'��u6�rE��4�R*K�*:�ibz]�+��؁��O[�"�6a�Ͽw�(j����4�ړ����#+ց^V�6��E]I���g�(kۯ�>��-?�	U�|������^<�/�sm�q=^��laHf\{5�N�P��ǎ��7���Y�I��M�NEo��g���+�{���b�jF��Y�D�DZ�x�*����@���F��T9�z��J��햃��Y3
��q���2+@�<��-�'��h��/%� �Kт՞Y��x��N��	 ?�FUc M�k��.�Xjq�K-�^U�c���H���϶]{�Oey��Od� �ì���x�o�}��p����:
���(����'���|+�R�����7i��'y��d���P�x߃�Ss�y��ǃ8�v��R����gR*#�2�j(dC1�ȱu*�����Ԕo&3͎h�������نN9z�ҏ����V.�a(!�N�`#)N>G����84]h˝,PnHJ��m*E�������=)2���f��1L~�����!I�0]���6��N$"�G���1򡡢7��x�8N���C�XCti�s�i�2�ځ(�~��t�>;Q1(��D:[�	�,��R:R�sr�9�|�?�e6/ʰ�e�#^�y��_��O�JO+��i�h��C�w�0J��9�I!HW���NT��?&�Rz��V���Ӂ{oQ�e���1ǆPҒ'Z�8+�Kߥ!�tB��Z�4厸4�������Jcs�߹|��~�3�+�ˇ�Ԟ#�gƼ�x~� �+Х0��Q9�5Ck.��<T��I����mȈ�m��$�/l�`��T�3��Ƕ�����8i 7�X.�11h�!_/��₝����5�����ڛ&�P�x��2ki�ѻ|y�cfeB=�#6�D�M��J?�.Gi�A���Z'F���υ[$�:���1�Nf�9���i�O�;�X�j���;g�
�4�l~� r�\�h�C�Y�E�Q��;j�!�X���D+��KLy�ڌ(��FӬ��J�PT;�/�6&yo���i��x��l,�-��^��5�0#�9�y�VyaqO��0Q��r�;c��wR+L_\d-�)D+8��d'+OzO��x����,t���e��6�^����Ov�<�"���N��� �,���3g�VW/[n6�.��!�&v��l�����\���(k]B����z�7"�lm�m�]�����ၩ��Y���q�k���r�+�E���yf�»�8j�� Na|���34I$ktd�1`��Xlk�Qt�ʻ^����O������7m�-ofg�3i=�w���C�R�4����gϲޱ�&-�a)� �&��xۜy�K�PT;��3$yB�l.Zl4C=B�'�;�6[n.��#7ۘ��4;XIF���%�p̡?����Ϭ9�E���MT����#���ź4z�&|tm0Æ!/`�ӄ���k-FZy��$�G�})��ՋN7��D1,P���y�
^۔M�)d������RnIM}�������ʋ�0�������H���l������cR]s����C�i�^׮�Ƌ\Nw�:;�1�Z@}z���Vm]��U#�N�Ci�SJ#I^�5zӁ�s-���j���|J���GA����>���a�Ѭ�K�)��y؉�Q	�	��[i�1�8����P���R;�|���z.�8ʜ�DO�n����.R�x�0�����5���=�do>Ȅ�y*�����a�&�Jg8���CLJQ�^�6��!�I�O"F��U�9�=����s��Ŕ�U ǞJ�MT�T̻Tg����Q!������y���J�*��W��b��U7��hX�	���+�F�	K������=�͊��m�s,̋��)�����_�Y����HI��O:Im|bT���}wߦ*�`Ml��P2u�yeW��\��sX�!�B��1`#��[,�,_�B�eS%N���	�,I+�@#?vy:h��J��n�L�ǖI^d˧,���@gR�C�W�1�²M�N@W������DL! }�Sm;f��^���"[��y�P0
��Ӌ���-�V5W_8������Xij�=rk�Ҳ��<EA�RY�u�b��(ې���_��7� *��Wș�7c���,9ҭ\��E�$�Q�a�'im���p��gL���BާL&K��S�ʥdi>����NQ
,O�"g vP�@А/�͘Mź����5vS�l�!E��i�i�k,�F0,��'�,-^��ZaE���A��?�D�˲�^4��v��y�����4��"߀��|�;8`h��c�V4������-d�ia�`�l	��H���r^[�}vے�%��f��c6F)'CͭMT�͒$�Z`�G�9�4�8O	B�
ޚ�� o�禯� ���"�Q�إ���´9�M�
�b�e�|8s���X�*�^��j��c�#^��ya�7���Vʌ�Ri5Y�B
���I~��<�fS�'���r��b6 B6t(9�E���7]�fx5���wf�c����A��"�(YG;l5��H|�n��w�v�DB�+����%Ƌ�W
�%�壩U���J�pq����BA`\'zG �#6%Ψe��P-��q��c���(���H��:�X|<9q)j��VO8�1睉(�.W��|�����[n"*u�$�;�!�����t�k������YwB�'S�ή�$�)qߍgQ�t�]��D���ʹ��9��9��ȋ�\�0'^~��1.|/�1Y}��ܸ�e�{o|���=�Z\������:�d�n��eR���G>��O���je
.�}�օt�/�;�'��$"A���8��s6�ӡ�n-��f���֛�q�g�s�%�S�%5�g�^�NUJ����~��I��ís�Z�4h�J��(f�a�:�=6,M[mV��m�5�5Xmy�h�.���i�+fG����.�JQ@_^}��G�E��C&�~�L����Y���{mCi��Y1s�A���#�����qC�<���RJ�`3����ɰҔ�0M�E��<Kg��WW�F%�S�߁OZx~lϿ��[��%�k�kEr���Q�x�|x����'^~m�Ė��U��ǲ��0zT��.�N�p�,5�\(rـP�	E���^SH������U�O���L��D+�t��Y~�
-�׮�������:�Pr.�Ƈ��i��y�!i�%Zƣ��7��;E�0a�4�XWX-��S�%b#:q85<	���5��<x/���V:�=�-���D�ȏ����6dߞ��jq-��S/NNfrY�y�t��L�gȇ����=�0�S����^��﵈a-���e���g�����"2m�>�U=�@��l~�:���F:��!9N@Ma#9l�ǉ+#֍�_�2i�
��
S�C����}_������;К,b�)�ȱ2�V��浢K���,�<�B��`TFl^�!�@Y2R6�~HC�0����U��xaD��il(!b��(�:� Z��NE�B&�h�cXު�PB;��{oAN�����ɆQ�����M�Q [˰�h��E�rSQK,k�(2��:r�p���
�
M*�y2��h�2<��wK���u<ѭ���'����΄��m9�pQ�q�x1�)��9	榨�,̳}�"�e�u}�L��h@`��0�"{��h߽�;�셽ǎ�⸅
1�����q���ee���kE�9?)�����q�To��|�!^ �6:qv`"L�/t��ԫ ^��.�9_�0:�Ҝ�Q*lZT��������%oAQ!(G����I�~��:M�b�`�ir�f�`谣��Y"v����5��@7��\�r�_�n��~�y2ف��ّ��;�]��Zz1"��OYdF&}���K��.` �����.��a�	��h��S)N�";�l(-\����*�k���a�[sY.r��ى@ �Xgyis2�u�]pvJ���AU�\���;� 
<���#*�Pq��#�K]��c*�^z�-N�ꭔP����a��,�/�0��l�S�y�?�m�q5��/~n��uƿy��l��b��rDe�i���F)�Z��BJ�������ۮ�it�5���L�D��+L�sO��������l��\!��p��n�GW>U�Qa(G���������Þ����!1x��S�,~�B�4rE��&2Ȥ�~rV�W��^�J.�^���R�I�E*eS���CkF��#���!{�����3z������
.�*-�b��U1el�Bͣ?ލ8'�Z�����2��d�l�����b�;���:���kU�*��wk�عn����c!Z�9=4V"���E�Cw���)�a5����t����:�Xg���ꜿ�����<t��՗��މ��g'<%z��ވE����r4*�E2ɦ���~����7��ڨnۧ�����"���5;�[lv��l��/�)k�_���8VGDIWs�V ��?|��3ǽ$�[\ׅ%$�����R�AJ����b�!�����f�n�n���>����9k�u־�#�9�y϶����*�o��i��]i����&�e����g��DJ����냧%�۟w���Wv;#��,f��|���=�ȁ� �s~��jR��t^Zь(�o�1]��̰nK�=S���o�iLؿ�~,��Up��#z��`rd3�[ǚ�����X���y'�ųx$�-���soq��Ƞ(�C���z|-�n5�Pv#��6}��Y���M�縖������ϵ?���˄H��d���݅�z!�|�$[��^>d����~�*��ZĴU������=��gUۗhce�ǁ^�G�w]Z��@��5�_JEؑ���s<�,F�7Ԍ���Z��ĳ���ٽ��gZ���bq>���5M���T���j,��8��Mz.(�P�#��.�C=��`���*�Oy�.%�'y��/b@c\X�0����&I��ƔC�c|�]��\�����P_ϝGGa_@�.x����Hz�lQ�����)�,�s�hHC�y�����^�rX�ލa҇�S�B�|"�"����d�8��%���E�������	U�Wz���ty��ٵJ�����`��������o�e��5CX���1SG,ѻ;��-Y�O���.b��Gc*ZPk#�|� ��n��@:��ƫ�;����$_ �)Ƒ�¢�E%�b�4���֥9�ڗH$�(3�k#�wf�W6����W�����cJ����"�%����7/(����B1���+�܅9dc��݃�\-�f�$:w���I߬X��ԤU�j�E�;LK}�3vf@3/�:%P,��/#�� ���8��|Wn��p�+b�,��Wt�l�f�B%�Bg����3�P�K�n9NFag��q#�|��ir�z�@�]0��'�s�Ώ�I߭��9�?)��EQd�O�@G�y�Z��9O�U�ڤY�үşBq��hUzЧ7A~�a��}$��&�J�<��Bo���	Xg{�V��
��QX�`�y��*G*^���v��B�,_>W��>B�s^�}���+���Ol&��G~����G��_o0�fW!!C���7�������{9��8��=�
�Q���Q]=m�n<���Zಎ��.�c�N�Z	�O���\�'e�������󼁏�_�<����v&�]��꭮����8�Y���#E�5qOU�w޶�1g���j�k�#' �����Q������	2gf}��� PW�ڣ������&���O����]�7\�r#�W�Iĥ%@U�r�6�(v:I&���&V�Q ~�����y����X쫴=�E�����#����S{e:�:=X��4ܤ]rj{�X#�D�O6^yP9
���.��y�{
��LIŘ׷��U�,���W3���T�ͯ6�d��Y�bH��|����ä�SR�� ��[6&�C^(E�"�����ˬ6���&ry��<�+�Y2�T|�D|pd�<���t��Zb�;�ͅ�ׅ�r*�"R�I��'��yآ������NT�~~l0��9�h~�&V�\����5g�����)U�]m��X�|���Z)C��3��|UU�tN��������Nw�¾/��_�\J������)ibB�@�S����}�\���c��R^�Z����l��|�	ZF�hsUU?�G�R>n��Z��ba�,;�;%�����pbK��u�,AA�����!H@��zI�ɀi�4�ϖ��{"��A;�ڲ��!X�R�k-?�4�x?���0���k#�x���s;�����%Q'��r�S𷷤ʝ�{T�y���?�b��͉��N�A�ͱJ�ǌ(g�=����~Gh{x�2�kئC(&]mA=U��QO��vB�6���1b��J���|�"�l���c�o��w��Kc޽<wT\����3�.����pe炯8�Vl#}�&wW9�fX���!�Q���u����7�}�Ij�SǢV�α�G3[̧׮'* N��<�5iS����Tg]��~�������}h�\5��ͣ��ug����M�)T��Q��ly�S�ib��I��%�ՎF�E��-n�<���˙�Ԣ=���i�S��/W�M\0.n�I��
�n�7){)�$�_$��e�N6�GHt��K,g+lk�f�$�z�V��	���m��+����1}��L?��r������rj^ʣ��BPn�XX�v�B�OX�1^��A)�j�%��	5��ͻ%mU.8п�H>��xzO��0��)���3)h�D���nR_�QE�!�]�+$|�q|+�.�b�x29��m�^�~g���
�������}�����Ow#��@?N~�a��%H���&G�@�=�)����Uʩ�g h�8��kO�2���ʉє]��K~p/�![��F��?�&'��������\�jK0��j�b*t��������Z��ZAǕ޼�+��¢��Ґ��	������#3��?8����fAl��XN��B�s>Ҩ+/�����L�S�ݢ��*Bc��s4jk"�h#tZ���~��eF�	ZJ�=m/b�L���
AR�=�񡿱Vm���;�♁��󋱹����g
JcB�@p�/������gTI:I����gTY��>�V��1��#x�N�8�����:+X:������I��q7'Ϲ���.�RƇ��5d�0	U1*�<�.��3R�ܪRG�{�N�B;�٭tۑj�0^�'��5�F��^oIr��O>�:����Z�����9[�N�h���l�*jZ����QB�i(����vE��r��ws��@�%A�&?�F�� ns㗁�.�ސֺ�¾���j��C+R���Z��
r��l�ƬC�P�v�������i�������C�'���Y��L<��W���퇋�԰���'z���	�m�;��7�הF娟�&��z~�r-z�wt[�J�
�̉���r���g�(�9����<����2�)<���&�/��Ο���'�F�n��g����F�J�&��9e�*[�_*�" 
i�nu<������ޮ�Gֲ�D�G
���$�]I�"v5��r�k�t�
�ЛO �n�$2gݜ�9U��2�:�c�'���}NWt̂�%Ue�&H
U4�U�}[Z�[Ϋ%�pq��/C�y����1�g&q���qK��݂ ܤ�+/��ŋe��"*����n���nO�I�f�Ac#�W�� �/��H�KnW5Y�uf�}aJw�ſ��.�Z�Pekl]�mF�c����u������&MCU�D�B}�^��~��b�F�S ѽr�F��Ʌ	Mקs=��������H���o�8s�~*r��r�r�-�HՍ�>�"���z�6�A���6��r�����ˊ�:5���y"�d�-z�#ErB�'�q���'K-����? 9O�sѶ�NY��za�O���֣44�Ǧ<������ʩ����Z����{�ޚ�2��[�f�L��(nTti�렷�}��]<����f��"ޒ�i�������0Id¬w`ύ���ԞR�[�4�#���p~������MO�{t}u��� �Ҙoп��n����L��:��͇�J��~�!�	z�'S��F?��j��$,2��:gj@�Gb�X���cs�[L�� ��vn�2�Y(��L�/�Z{��20�T��x6U@�;�GP��[�����ZX�[��#A�&t�f^2�f��>h�.����5�5p�y�	�J(��k	o��m<���jy�ٮc�e�°[�+�n��0p���1��/A��ē|W���s-	��Um��I�L�j����(�g���S翼�Q���D���gb{-�)��x%���l_�l�Xl0�{I����׉V�'t֡o�����.����z:��$�%w�����E=6$c���ζ�G^��3*b�协&�Sy�J��*1C1�h�C������N�5{0�I4�I��:��+$��'����=C\_�r��$ČY����3�xr��t�����mW��Z�:H�#'�R��s+M��L�ú��S�Qy$�b�8��i-:L���^�鱇��Q��NfW�3RC�V��|���ޞ`�,߅*�7��'�2� ��6�F� 7w��_�ſ<�P���yhޱ��BK> V���9�\�����aT���w�ڮ�^(X����������4��MA��n�	�i�8����� ���L�g�������솙�s��8+7B'h���r���;=�����x��Z���W��
mk�7����Z��5�2#@ū}�ʴq�F�G�m�T��z�/�YF͸,FϺ�ч����m	F����(>�HQQwʜ��(,��E�֬�8>k��h�=O�n��z5YMΫ�[���-K�nU?����P~��ﺍ���	�w}*��x�Yf�0�|Ғ&�H�>`"Ŗ�D�5��b0q��i�㶿b�U��4�F�������^)m�km��/��m���z�"{e�4�b�nf�w��eR�O��?�*��x�p"��&h?���q%63%$���@�%)��#e��k�8��r2�����Ҡ�!�"�ŵ���G�%��?|���^��o[���ezZt6����_nD�_�5���+r���e�mZ����2���p�Y�3-_T�I���w�L���1��W����O\�O�F��kْ� )�{=��#�.e�����^����^�;�n�!���K�9.�`����gc
��}&a�\\�TI��e2��۳���i���m4� �;C�Ė�FEа��[*�?�V ���ۡa�K.�wE֘�|H�a�X3�m�b��9߻��s��`iIy�J�?c�9"ض��(x��醹�;��"��8�=DsM
ˍ;ʆ��� �T���#5*�%�hxVT*.3[����f�]�yM�b*ڣ<�(%%�Wa����"�C��M�����;�������D�y^iW�-��GAHV��X.ᴒ8CH�������p^?�I��d�=N'��p�2��྇�$�/�1N�.g�Q�4Dy�����Kjzf�I3��@�,c�"���S#K �W����J-���$0���i/ǃ��I�Z! r���<�ʆ�[�#�ÚL5��jF���𵥛��'Ѧ&�46�ŭ��u�[<�e����d?�tr)3
+f`�O3с��x�20n�i��l*�x�q�4%�_�紧��߄��]ݾ�9�4�'ؔGw	���hzߡ*�b8D������t�g�Z,�2��R��	���A���3�To�s)�-��-�|+	G�p}F��_}����:�����R�F'ť<	w������c�A�(�v�s��BS��mlQE�^��}�wi�Hh��~���<�WF)�v3�i�tL���R��IV9)Y���U�h�CO?�:EtQ^Su�����1� l��b�����W*�L*�PMڠ9��]��0<U���lR�b5_�w"�0,}��q~�׎|y�ކ!6P�@��JQiȋ��x+?_S�nf�<AC�bhC9s-��ȚA�ny��#j�nPZ����@U�w�e��
�}�1�'+C@��*� :JY�B�A/R�;���Zm�nx���1��%#�A��#A����A*uQ#/9���_�D�|c~ش#|7��g�m�.�-B4�Nٚ�E
ǃ@�FA����U�>\��� q��eBR��]|�5�1]��G�����eN��.������ż��@���f�bj9�D�E!��_���xO3��_��^?�aW���J�HP/�6C��:��_�qP�c6��_L��k��i��S�3/�9� ����3
C�i[N�g�����4+p��Y�+���i�v ���d�k%������aN��7S���Ѧ��#  �W�oH���Oi"�w���h҈�K���BJk�������ua=�)�0^ɍz�DBT�46:,��	���H{+����/�T��$���8��X
�JrC)rW:�/�� WrI� �l�o�m��{~��&)i��8-����(ulÊoK�|i�$=8�p�^3�]f/���.n��^�;vaW��%~?R	��$�~}��C�M�����U���'��E�(�^�!�"?��1��Y��	Bl7��f�rqg����ͤ��n�ʍ��;1鸘o��b�����E��͒�=�m ��bמC���h�[��w.U�s��QZz���}~�U���qmvFى��ᣭ�r�Y�E���R�Pī�!ɺ��Ě���(Lty#X��C�0�Z�µ�o����Sn�޳|т�|y����'[����*��L&=�j5��˪�ϔk�G��"XO(ge�Lv�3�uɚ�6�w�2=K�Rmc��p��G�Rت�8�l2����iuw52{���a\�=W �Il������\f��w |_܊��TX�i)��* �r%l�q���4�9�j��:+�hz���;(�0�sS����%�M�ʔ��'.q<�I��b����1ۧ�q2��i�2$����;����{��+��Zq�&�S����qUv��������ˏ�����S�5��S��0a�?j�w_��tۢƳ�����D�2z����@��Y�6<37H��p
�q��y҆���F��ߎ�q��o��f6�N���� �ً��k�۬;�͐儝�E�]"�܎a����<�6l�#��q����F'g|燳9�N1��P[
P�7�|J�w�]�Del� �]R�_���3j�*1��f��/���+f�;��M�#�_��n����i�+ϖ��&�_O�O�?TPpnK���@��'��B�HJ?�O2KA����e+������y�U�Gy8��W�p��t���5�K�"�>}�:��U#[���x��~*n�>�0�Xk׿��nA�a��ID���/�<���/$�2ڗ#��EyZ�.��lq͛�J9sI?�\���S �l�xW�w	^��c�b�q�L���X�Cr��C%��%m�~�M1!&��Z�u%�Y�����F��Wu���,����jw����Ʊ�'!��g�6Y9���-Ix��)�Gj��u�V����ۻ�XB��%yT�F�J�HI�j�j���S���bQ�B0�:����U��$�[��l.�8k@J�(��ӾN���	
�4
^壓�<�{��������db�L�XOY���9��k�L^��RX �W	"�RW�b��{i�\�k�Mǐ�0(*)�~�Au�O��碝�q�j Y\�v3Uݵ?�g����e�o�����F�%���<w���J����J%[��F�����.~�KEf?�w�^�7,B?���3e�~\��_r������=�1 4I'����������tx�e�����@�ɬ�x����� ��9�����,�I��p�g���`KR�~W�L�U�S�7��,Ɣe��#
�8�Z�tX�+V��(��Ү����U�V�M�~��/jw�L8�5G%�����"�:W�G�T�@-;`5�W��T_�c!�����$���?��[i���8
��.o$�6�������u&�KrЃ�d��:,BH��	P���Qo$��*!�����BHc�5��IvC������D@�y>��)�0
_j��^p��l�ddBO������#kk�K^� m�c���I�*W�[*�%5��pLv���U=U�\w�|��&2�on|�F�x��fy�N����%$����Թ��H%����9W��C���xꖶ�I�@x��-+�ռ��V�3`Q�LL;���=�� ����+a��A�s���}�Mq2�����xt�4�kD0q Մ�m��*yC�%}R������_Q�at�_�.3Hߌ�0��܇!n�=ɭ�Rb��E�0���.�Qʺs!b�	k��3zݕ���in�H?3�lg�E_��"���M����}��=��sx��k��k��7C]�M�d�
�OZ3�a�
0K�#�=�Ʌ��(�[�; ��_LCު<��"<��afgoPB�����p/�ԅSM���^Z��=�1�g!�7��1�T�5��>'�_9�EӃ��L�����o�7�S	��Wd�O9z�����?Bq:7���t�R�\%����`���ƕ#�-F�����k��!\�Pi_f�q/*��w�@�f��>�?#֒�e�.�f��a�#FR�����&�l��h��:�p)��_�6�O�^�r) ��B�Pb����Z*c�Q�K� ~�&��Vv�Di���)�@�����dm��7^3u��qPQ�"��-SxI����/J4konޛ�ز�B޿	�nΨ�KGO���hЅ({wB���z`��b�b��1�2a�ZU���%7?X�Ö0��5{{w&+�)њ�Ǭ9BX�2�
�l��#̡�](R��]#���[0B�q�&W�N1wy*~�
�Q��rR� �3�۝���RVbq�Q.բ�����b|F$L��ؘ2V���S�^g6�Z�K�h��M��)	g��!B�QL%G4���~[Zx�N���A����Q�YX�IȜ��;�J�R��:��:6��3�,��b�qd�Q��̇�~��z�q�Ȍ���[r1B��
���&S�[�&S�'F��>@��M:.�B��B����*"�6���S̿t81KB�JP�}i�6`W;��.���F�����"QHxxoD|����59��7'��q��� �u�Fk)�c~vq!�m�M�M'y���z�-�B:�%�ӽ�|�+&�%�z΅��--<m���I+���Y�nwg��&��7	���~���Ɏ��Mq����.����{a<Y�ԚWO�!�3Dڌ;�<H_Og��F�E-���r���2��%w�Ԥ�^�+z=d�M~'<`�B�Jʥ��1�P�j]���
<�@e?��U�1H(j���:G�ݪ$'�	�z��~_���m�EI,Rr �h�^V�U�7������SwK:z��=iwI��=�*��*K���ݿ���O�g]=��6�`ZVs�5t�����9��"�>����ò�[
޵֏^̨q�?��[d��I�y�|�愗|Ng0PP.�|��@�|����w����m;�@1r%�Eo�p��;��@r��}V>pf��ك;r��b���֡2���!�<C�)��q�Y����l7Qi��A~>���c��`B�C缄��.��u��u7�ծ�(N�"r���D�g�}���qr^
n1���W��"�r{����=�<ڏ�d������$��T������Z�Ԍ�{����� �@���t���$l)������cЫN�f�¥f�U�[��E{�<sh�&��!��1r����"|�d������������k�+���U���X�YH��s����+�Q��{��38�hȲe$���mg�_�C�
W�L]_��!J,���s��/f�d���{������/UE���U��V��nԄ(E������Pl����y�o�����aKw�[���������F���+���52lZ��o��u�tn���T�b֦�e�T��oI±<����Yn�I�P�}l��-	bZud!���H���b��$t�o���ۋ��(&s��'����q�W����c�Is��t S�d+\�!iJg��`:���w&E���*S$�AM�B%пѩJN��m��}��"hZQ�jH'T�7�P5�5�ܷ*�6 ����/��� Gb;���j�� qI8m���(s9ܯ\�j@��[{y�+�(�ܱF����"l�܊�+2qݹ���i�g�_��},��3�pQyU#o &~e;�I���9�ѭ�- A�W:>��>�K���8���7��XC"I�m��d�\]Ć0c��Jt��J�u�;pJ�W����V���pm���L����V������`�9}׵Yv����� ӦOJ��mUш�Dao/�^�AJϵ}0��p�	�H_����)�mvk�fI �ȑ���|B��H��C�l��O������%�֬U����VX�b��[]�t�����$���D�_�L֋�H/�0��:�5��YΆv�p3�K��Vn��d�{�_�Xv��d>�7�"�\��f7��4�����#�s�İ{�%�h�鶂���d����]����|"s���=�#�P����+�<&�f���-��Ķ���\����T8�}��k�M4L-[%��B�L5�~̽0����<�+,��:�!����"5����YS��f�%�ulf�f��]{`6��i1�_=߰�C��6!�<��W*����Ib��~���<�7���0G���3w���H����Fj�q�9C�OF�J�G���S��E6#鈞����Dnc�D��M�rݜPh���o/�-gY�F�c�p��ۖ'\>d{�;���`
U�m�4x�0lea
2�J��5aYg��]�^ןۮ���|�o�4t��@�t.?3��\$k���9G�W�\[��<�d����k�����\ � {��&8I�L��9�·?��5�YO{��S�!�a��=]�o^�)������?��(Ro�8���d��0��O�.cT1��C��(�p�������[h�V��R�ɇ2��z&�v;W��ޓ-�/��C�z?�"7(1eV
��c�/9��*I�,���=��&0/�!b���*^�e����~�-�/P�Zܑ���f����"t;�*� �^K����] `H�T.-sK��vFHb:��>C�;���ިL�>�[�*۰Q*D�����#�6B��v����Ǥ�3��jnKb�����+�p��R �L��uѓӓtf�>*�#k��y���k��!����e,�2ȸ2+i�g)�@�(��"1\�y5�ֈ��/���	ރ쁈���\";hOV�(+��K��+�Aw�l�����:/�J:j�䇚�.��g���+"���=�H���D��>�H�t<J�z�l2��qr�q������K���5����fW���N]�cke�'�]L�9�6Jߍ��]�z-�r�1�c��u�3���N���I���H��vXӆ��A�*[4Ro��s�(�{*�ӂK>�~�6�E� �<>ȊJl�R�?�\7_��O7ϴe� ��\�n�u��ɾ6"LTKH�&�n�=�2���6��+`����r��)��;x�s@���^�\�f�%H�)��>}�gV����j���3�.�$��m��"��FsT�m���8��Q,?qt)�&��f����	hc���Wv��
P�:p�p�6f�|Pe3����X��b�Z���p`��l�)g�����&L�MZx�����h�/л&�k}E@T��|��M�o���Z���H��n�vJ,���3�0q'j-	����O]k0��~�Cݦ;ݹS���Hȟ(��>ͺ�ʄL*hU4��� �Y�r`�79�A�ӝNA����S^������<?�O-� z:Vn���o��Ã������d��p|U�a�rw�8�Zԟ)�DA�(���55֦��/6��n��ة��O��Ut�����������έ��{���8ɿ�98�FZ[V[��²��(Զ��pn~��;'C]'�R��Vހ|Nq{�(r�k�5 ��wY?�Z�o�.	�	��U<k�I�F3��u��I��@~$ʒ�
��pk����`�r���4��'�ƎMX�^o={���P�R��L�ն�/;����5��dko,�>gE �m����UC�ן�u+��ZI)�T�6�~I\�o�s����"���ZYĹB+���܉挧�ƭ�����\K��Xޔ��!�?��MV���G�|���u��ٱ}E�äc�s�P����Q�.��Г�
��������E�hO�{Lpl��"z�j 7��	 ������N$�~�$p�_��ƒu���ȡ���
\[W.X�xq؄W�Z��%�����Yi�Z)�D=k8	�z'"l_�i�u��U�$&	>nǼ�|ϟ�q���z��� �T�rפ8�W�5���>��x	�>�E�4����N��`͟[U|�
i�χ꜐$��5
 S��bk�!��J	��I�譸2R�߇�r>q����'7`��q�F<�}�1g�_x�q	��X|!��[��&FC=�{��� �+�UE��.�>_e]́��;����^z��ۜռ��·^����9E���3Fz��A��x�s�n6�=�w#�5F�e��I;7S7� ��e	U�Y^{��7���`��>��箆Y?�5�e��'��D��(��y����1x/�%��J|�=\V�"�^J��m�.���I
��х*�{8��J5�R���0���W/E+���#�H��̸��e&-�ڶT�ǣ���ѤS�q�Ns!G��)r+efW�1�:aS�CÀQ�n~��,�%x_^9�ui�~�ItNG��*~����'����ؓ���.\+��'��s���!��w����(�^h.�ʽ/�3#���f�?�P��f�qU����|�pX#<o+�gc����3�:�u���}�b��O+��w&p_���DG��*�g�n�
�l��
䚶���~���vl:A����GI�R��J_��l)[3�m�2A�i�S���/$�,����Ez�Ys���D��G�p���b��1���=����U�[?Y Tm��Kޞ_��R�����N{�U =T�Z)�Ɛu+&��K�l	@�������*Y���+E�x��5���ǚ����"�����L�����	k�}��p�΅}�����2%�0z ޖ��(�^�l<�ߏ��ї/禣�	Mk�O�ؗ>CS�_6D}����5o�`*�bb���z�^��}��=޿X(��S8��*T��e[��n�d�/خ���3�)����0S��NcID������F�a��a�E���w�|� B�bZ1J�\eDh��u��-�kD������$�W+/�\ͮ)�S��yZ>�`��<jZmr����+0��1�s���5(b���o��������^y_F�uʑ�US��I.��Jl�/��hI�}Fg��8Π���6:H��v`�PƝ�$	�j��b� %XI{���$��T9ʪ��W1� �RFT�
êu�yt��6�I��2���Oq�qM���tJ��.5�F	}���J/F6�`o���tgԋ^.�˽C=$��g���.����~��F��Mo�ꇶZ��/a��3�䈢ЂoN��=<5cĆ?�GR��o��11�+&��Ky%Z�S�`��X��̌�麚�M4��!���[�.Ϛ��rGT���e�	�Z�:�L�/���;�>z'�۲X<�(V����w�D���'��:�A׍h��J���}:^g�Hj����	ɍ�Q���Ҵ����������P8�x��6����z� ���� �GT��5�tޠ3�`m�n����؞
1X��49ˁ��I?3��m�M�mq�S�nİdI� ͚��?��GM���=r)���Iw�V��?�@��?݈A)����i���1�����Q�?���vb��������d-i��}��&JcK�}��"�,u���}yZ�O֟q�/�V��E���z�/8�sv|8},���VL��J��m�W� [��	u���J��$���ݤ��\/U.�ߦ�☗O��/Y&��n��~
��.S������Գ$Tl`�>)1;�m��1_�H2ه����1/V�i�xd�щ/��J�[i�N]��<~?��9�n��GM�������������p_�?/�m�����T�3-(��ڻ�����}wOI���v�~�F��tYVd�jf3�� .37�.״�I�����9�n�b���	������EW��X��}�d�O��@sSM�+�SD�2���<���t>f�K�}_`M�Z*��\��/27�(��4X��@-A�;��Chu�ק��h� G������K��e$��'sXAa�b�oĥ�����W�GY�!)�h^�ڻ^+m�N��0�����
���Y� �e�L5�u�~�p�&PZF����g�;b1΂ADo?��(u�!�4�(b�uǛ��,�P6=C�-ns�W=	a��6���atr�w]���'���Y���*��zh��B�2�7�Y aF�N��tC��Y�mZ��2�I������x7X�"���8��׺�S���U���-��:��su����.���JDf� )d>�Vk(�Y�W���zb������U�V��!�~�-x.��y��� @&�5��Z���kc��1�ïr¼A�h��m=lg�*������ 7�a~�~�.F�͞�N'��ˋp�ܹ
�ft��d�}W�;l�^/�����9:G�q�ܟ|�����`z��O�����_�Ӵ��a��S�8��~�i����g��F����'ܢ�F�������5ﰙ���TC#~��-B9�i�C�g�n2HI��ڐ�yK��w3JKuLA:�yMY#�Lſ3z�T��{�>��-T�0߉c�P�G���X��$CA���~������\[ɫ�����8ʓz���,�|.Q�f�k�*��39jM��X�yR
�[e�6�����5ґ���:ù�D4��5�Q7���%ue7���IB����j#H<^��B�sd��t�u�D�/��"�Ro�E;Q�Nfl%�քn�wQI��19���j�D��[6S�=F�at��2EQy�O��4���M�Ǉ�M���BW9EHM�gm[�/T~�i��N�jI� A�p-T��X�Zk�1�6�p��/U#�^8�#�����ڛ���O8�S!_��b���(x�Y�a\��&����k�e=�1*��Nq�!����'��Lǘ�,���曲#+�^*~��F+��f0��/�sm�2G��{e��(�\j4���[�pFĐo��S�Y~S�w[��KFG��7��j���˹\��e����:!=�a?��I�u�:� ����������rh���)>���&�n8s=B��.֊BP��mi����)n^�ds��7Qq��g�]@�� �P��-=I	���=����4i��@�����X�_�4�5���sR�}�i����K��)H�n�T+�?��O_'DֱS�lZ���BY�
��ɫ@�[X���Ljܳ������v����J�IU�D4x8( <��s�'����ԍ]k���c�,��b�[ݳ$��g������f����#a'1�����hC���渵�������	ܕ�F-5Yb�Q�-���q�t�����'�Y�C?C�nlDq�:��ņ;�PDӊ��}��9�c�O�v�� s��d;�� ?s�?_j�";��O�|S\�Y+���9\"K"=����:�&��Jsv�`����Tr�uY� Ϥ<��ڛ{�$��Uk�Hx�㊮������#��	 �^`)Mx$�������"rE����nmo="6��L=��gy�Ϳ=U����������Yk(���c��ִ��X�c�kʆ��
�)��Q��x��W��6,�,���5/��P�Tҏ.��i�L�5��C�i�.]�Z%�<;`0�\���׈9+�n{���|�zhs�,m�ҮZ�O{�1k��ȇ59�G\�uEBa|����N��j%�u/���l7p��2�: ��x�j����;˫�j��	���:z�qVY(����azL��ʑ�ocOMS��צK`w�{Q�i��O�m<��C�s��R���"�Ǚa�*2L6ETU�Q7������b�T4 !����*o�����e�֛1�̩�/���f�����/^��6���_&��_P���5�r4b+5i���ԫ����K��R��� ��ZT_>Y�q�}���2#���a����������h>�������m�|,���c����Wd����9�~X�c!��&�Η������CmW�������H��J�@Tf����q��va��Z��;�9\���p��A�y|V�#(+􂸪&.�Q�� �5��2�y�;%z�gԗ7�������?.C�_��Į˾��*H�ጟD̽�	J(�y>�92�L��-]C�6�Cn|
��|wt	�/�0k��z�ɞG�=R���!�G�x�]LT~�$�(V�Kv/��kD�k1H���}���(�ڏ�O,�/���Ґc�Bh~�Z�Od�9n�_��xB���n<������;�	��c��|�~��.�;��Q�'}1C�3�I�����AT�k@�*0ƶ�6����5�Z!�y¢�{��n���P�b��~��F �88Y��n�7�'�7D=�䠸���B����6v�3L�g�u��J�Y�M���xzˀ���i�-��]����V�Hq���ݭX��N�Bp����n��~�����Z3kfN�I"h��rc}̣z��B�1?�����AF�6��
����W��Si``�ġ&�-��v̢8�$����M�?�w�p�����\�M��dZ0�/.�nc��g�j���a好���o���N��)��j�e֯�].�w8L�7)>cx�,��������<~���tn�ʮ�Mun��e��Yl��q,U�/��'���I�]ׅϿ\3�
H}��X�L����_�$�E�]po�̐1��8���x�S��i�5<O��R��WWz�@9�C���7ߚ۾A�#�+�f�t?A�X�H�i�'h�X��Y��`@2p�?#�0W5���������XS�z;<��ᾑ7(!�t��^`�˒vD��̝vh��Cıi�ln�=O !Yēr)/U��)�������aҜ����@�Ô.���&1	��o
��j���d�Ͼ��A�'��1&
�I��9Hx�l�>���n-8��l���VD��P�f�h�� ��%���*���{��szLi�X'NO���� h`	F���NB/�Y�Q�ZCXXА�.T���w7��Z���5���P�|k�b��>$2�-�+uf�β ��N)��H���1V��D�#mq֚��O���1�jKٻC}t�� �{�K�D]L��	���>��,X���E>��'f�~f5�u��M�5��LV�%:�&htnl���JBxiND�m�\Q>������k��@�,H��h��v#*M���{��-o��2�o�2	���m��l25����s���*Ĳ鱄�9��/zg���G���-b�]]c�Y>x��V����g6�ð�&�iDx������I���x��"���EQ0{�q_��=<�2A����,�K�{��=�/4��b�;�dMh,~��n���Su	��A�X1μ�$|�dW(��w�I`WOY�ɗ�{0���n��fa���p�y��@���װ� !x��;��$�^���AW��w2��۳�Z�W�Y�S-gspE�4)$�k���Z��O���P/K䮡]P"A��_�J��/����[�:�W����S,�g�U���9��b�����#� � ���$wG����'2Fy#�d77�s���v���כg���x1V%�"���v��1�푒��0 <��d�Y��oH�~T����g$᯻㭑O_	c&��[l'*DڎAC2A,��o%}b�w����k77�Ҧ9��(�i3�*]'A���y�~���9jȗj�X�ԕ�?a�Q�,�9޳?���}zN�2I�v�Z{��<�\g���l5��*��)�	�Q��;�z=ј���9&�޾V��_������`�=�q��G�+�=��:[�i��å�&�w�k��p�SP���`�jQ��`���#�w���:־d�,o��?hζ°�1+fNWx�t!����̒f�n͗%�[�Q?�@7&nh�@��C�w���ݝ��o����:��-i����+
�ф�_����ҊLVP�Z�i��)
�awݩvs���V��뚹[uZ�F�M��dN찁���Y�����){�tn�� VF$i�M&5�mM\���Y�!���8��0�U�M�\�3�bF��5_Ur���������T�(��4�^�}ޟ3�e+��Ҕr��Ɨ"�4����@"�1[C����$�I�{��,ɷ�୻�(U.��-Ŵ����zH��H��R��B2b4)K旅�䔤�ڣ��ߣ�]3'0�5���7�}J|w0^����+��5?���O�h]��4��_J8K����GI �YE���u����f8"s��s�E�h�c���j�u�Y�Iw�u�.�%�e�sR�2�������ݸ�1��y�"�)QE
!��剧�~����f^�&�w��H���ix�_��ON�I�mg�_#�8.G�I'�$��Ő��K3N���n��y��Lɷ�K~~[j�4x4X�`p'��"�H%�Ys��U���G�C�x��ůhלV���Qބ(V]�����,L� ���V��?7kt�/ﷂ��fS<]��	����'��8"�ai[�S��~�W��؄�ݕS�J`.}6�r���{�K��$��@��ܲg ��C�u~�ǡ������]��T��6��p+'i�[ׂȝ)�;��:#�N�6�_���ʆ�����jb7*|��f��ǍGD�}}��������g�ZH�h5�Kæ*����M���!�u��\T�=
v?�Lr����T��@_5p���n�@Rnح� ��� �����������9�޻6��P�&��+Sm�Q\+%$��b#������ �IBys�X���?�0)~��3��i])2���]/ �F[�],��'�D�ĕ���`�"�T2fd�����r�Ԗ��� ʋon�V��IS�k;�Z%�!_ώ���V���r�Д#T��O��nă���<��4��0�I�%7+6�9p og�3!��XyD!2���5�	���3s_y��|��	�� kiu�e'�V�ם�i�.`v�h�8盅~�e��u\��o��P݅��e��>�r�/�'������ �����������EŞ�Vm�G8A�fL����Z��Ut�c:O��1*ӪN\�qa'ܙ\�"

�� �UH��EH�.�h��y�:�����^������g!+J�Lh~��Ũ!afO0��Z[ꍰY�1�Hx�+�/)(�b�[k�!]w��}Ꭹ�H}_9�����IJ��E�{r�.�uW J�?)��e)�%�R��V�A�J^����o��u��`ib�ïFyauv��;�`�gOp[OHG�1^ocjY=La>.D�g��
����7��'�(U&t	�y��S�D�.��:�e��Fq�`�
��d?�ׂ3����S:�A���g�檖��1*�l���g�.�к�Rܢ%X�_����W����(� C�����������m��1�x\O�U�Mqe��ˎ��k8�.T�kQ��F
y�*9	�v��; 3p�h68%����E>&4�(?jL9�!Ұ]���皱�5����Ŋ�q��&�r�ӱv�N��>%�d��Y�����Y{�m�LC��4���i��8Z5%����?��TMՉ�eC�z�BO��v�z�b+��6կ���"!O��~S��C^q�������,���(��W��I|���Oc�G�0�F��t%�d��W����V���4鶟���7�)�G�!Br��UJ�}`l��V�RV���A����<.�[f��Ӂ�Zjx��"��Y���	�ifA}I�6z���,ۭ��N�Б�hw�?G�@�}�:m���u0F��kȑ���qx1[9��(����3qUʂ�:8۟C�,���Fl��r���n�W��=�P'�1n�߁����w?ٚ(��K)���)�1ZjeG�aT���bd�Baa}P�B��c-�1�N��b@�)������Ȧ��;��7x�8&e�a�5�2�#�{�2�+y�}�xv�g��9�Z��QxMiM
/TԵ�X	���M�o�B��u�Q���#{�.ط�=M_�t��Һ}���k�3""��h��a?��o�����Z7����L�f
V6\�ӝ��Y�J���!vA1nsЃ�e1vkЍ�?
��|�@���f���@@�1I_!�a���{э3�'��1rV��k����3�N��&����c9%��@�z���_�P;���:��bG�ԜյZ�rCm7y��������u�� �~tr�:~"%�Ѻ�"ߓ�*����F_h��eE{~�c��L��8���	����	��3!LD,��E�]o���+�z���u	"I�K��Xo��9��P"o��B�g$mȴ�.5��X
��2�wS�o���:�ѲX��Z�V���ӌ���4X�M�������߆�I�1���!�<���	Nc:qi�*�e>|'��/�;{�]��W�����6�[��{�3@���[�dFp���^
��+a�)\sPY�vS;�퍱�X
%�(X:);��k�1l(�i�<8Jׂ;z�xr.�|���=^��bQG7��5\�C���J2p���z\�|Z��Ռ��(�m�G�����}���[t��S����D��|��y��C��e�3�PX�jq�ɨA�c�-9���p,e*�-����,5��,�ۚ{�,r�9?��$j�&�(_9f�~�R��3�g�t"�;���q8�"�B�\wBH�%��%���+�U�v���ϥs�1�kx���{g��a��$�U�}P:|�j޺�=��(�h���O�1���b��	�����f�{O$��7ir.���Rݏ.a��O��C��L���͂�OPK��kd�]��;Ě�|�/�/p�m1�%�;-���w��{cl�R��;��N�(�S)��Ӌf��o�A廼�Ftx0�Ɯt4�Nh%RǼ�U���2�U���=�To4�1��N�5��jI#Ҋ���I^rBq�s*�{4����&Uh�`�1�2-�&����/�gm��"RR�V��5o�&����{��| � '�ú*��J�e{Ƕr�cK�9.��5RD.+���$�۸�J��\O�w���,/1q��59+1��z�bsV:��>B�v`i~�rv�����y���XZ���z�UR�P M��oIZ1a�Q��1G�Gkը8���JWL$6A�����wm����z���=0>)�J��C�W��1<���>.��i �!Z����y��m)�}1��O�2�e�vX2Ɍ.u(,�_!�ŝo/���$���u������>�dHh�)/�ȑsw�b��H�����5u~~�X+e�)a����+tp�r���bl>.����hC��\�7�=�~n(��O������¯�'m���������y��]A�jX���+,mj0�xڲBN�S��,@�	J��
X(٨.�T
G/�K�6��Q�ţ�"�S�p#����������#
�0a�vdI�UԻ��M�DZ�����:o��\�Vy��G�Xf�K���lu}nD�V��t�����w����F��v!���Dr�sz:����a3�w���d,.��P�g���R����ש����M��5�r���-@j@ϱ��8��j�g�m�6����dq�)X����b�f��M9/X�|zv$9�a�n�%���ҧG��iIu���ޔA���k�g���×��q�ޠ�Z�j����6N�§��;�O�rF����!b���1|�(n��T��K�������s&%󙮃��X�G֎�-�����{ 9�iB6�j��T����u�W�O<��� �B�=��Z�C��T=��%1������`���0Įh���ж��QЬʩ�)PYL�b��?G��������@Q^ġh
#�H�������[C�~#!��[���V���a�'�%i&��r������k-�*��M%N���tv���Ho�Y�ժN�c�ߗ~b:��#�8��A3�`s��tb5}S>$�R�۴���D����,[[p�ƀu��[|:	^F�69�
;J��d��U��jt$��5�x?�Q�U�����|��d�� a���\����Ƥ\���]�2�`8Fo;�g?*��9����="�]��_P���TP ~/�r��:0�{SJ�S<U����Eg��#0X�"�����ˈ{��.�Ǣ�应#r�jɯ�:D�7,��h[��Xl�K�K��l��:Y��Z{��~�g��S|/�	�hK����qQ8�*�U�N���rw���g>J�Tjvxu��"���.|�~M �6���f0j9�Z����|efklS�����]�ˊO��S=S�Gxd}\~�r�i�gF`�N� ?��U���Љ���<��߭@d&����ق�1�4h|Q�q?v��ˤ�
s@�$9����ކ7B����|t��4��A�K�#��SL�ϋ� �H))�w�N)DՒɸI���m�8'}��)�jP�ϱ�T��Y�7�є������H�^r���gdu��
&��p�o��h�QϜEה������`�f	)��i>�����BN��B��/��㻡D#���'�ÇI�zq\s�X���j��R}���3/�]� �.u�K�1S-��E8ґdx�g3����~����Q�s���ss���q�޺(��v�*�V/`<��ռ}{���mǵ(WZ`��^"F�9�2��+������2t�|#�CQ����/�$�v�a�|��3���j�/&������yC?,� v��|���j�	�K�
����gOK ҕ�4��,�r�Q|t���Q:A�������v�@U`gAIX~�C��C�GwUD�7�K�^���-j�������R{�UDƙס&K����[K)��$P�5K�r����B�D��z��YԵ�m"�0�`��ET�!���G���w����/c���jn_�ۜ4��xc2�d�-�о��j��k��GJ_��ee��o��EF��H���TB�䩕�T��L�8Y�I�6m������E��UJש��A��Fi�>�=��7�U޸6`=F�!��aR�O+��=k��XC��O	��J�Ru�A����vXƂ�(C����_�����<�ٞ�c̵*�h���f(Q�F�� P�y�����X:��\����k=��LM�3_�)F(��meʋi��G��㖠+g��#�n��vn�*�����Gf�:�'ް�TKz��޿n�mX�E�l�f
��z�k�����Ѡ��Q�Omh��MB�\�;��8Ȇ�U�����%^%���w�2_����;I����"��%�sY/�P;����X3���F�u�yc�"��~`�m=�c����~&������\,V�#�TV��2!�� 嗣���&�fB�d�σ����ќ����cdȰ ���oJn���H�HV|�DyP6Ӝ�lPg�d���8��������a�R5}!�6߁����nϛ�tg�Ҭ�W�����wh�P�7*ħ�e���������q�o���Ÿ����N}J��금�eK��M�,�V��S�\q���U�#&	&C��@�����
���m㊜7���^i,X�YR�	*v��z�87A�Ix�}6�כ�'Id�L�Ě�h�O�&io����Ԇ��3{~���-�&���)�@���'��xN��|ߢ*dT�5d*GRAU�J���	�$��M ��u�:�'���4H
��z'�xvY*���M��m������~���ԋj����o+��o��d�s��:�c?B5	k�	b�k��W�a�$J��|�<�F���c�|��)����}���`�?���q�_��w�j�M��� _CL@�~ ����}�Xt^�.ɰ0P�Ϛ��$���_T`��|E朅|���q6�u��s��-a�nƋ]�**t湤S{��@)�{�G�5?�B1��mPC�E��t 
�QU$��i�-?*t�o�Y', �O�_;�Q��3�M�+ X��i�26rI�q�v-Yp���`S��2���WC�s�����Z0�����N����v(aD�G�b��Z~��y��}�懱���� �b�*��D-~������H��G��Ǵ�"��{�3ls� Dӑ��� ��2��$�]UQ����v�w�Z"�%@��7�'�"z�t^<���䲙*�ܤ&��T%��n����9L��O	���+VL-LR>5o[���Jm�16������JJ�i�� 0�nh����|��n�R�(V�/��=���]Ů:���n�Ry��q��I�ǜe��A�B��F�a���P��$�di���S���4�߳�̶'�?�ީt�!��)b�?dt�5y�P�m�)
K[�QE��(��@��a��Z:����z�ww3ZE�Xܥ�Q^���՛��V#�c��w{�3q���	�<�v�UBB�+�]c��M�ɷ�Bĵ����S%�t��m\�H������XQ��bt�`�k�" =�%j��
]�2g�}ß�`�'���]U=��S�40�#��
�*j5$\�m�6�R�
�o�K(pN����K�W�-��ۉ�N���w���eAQ�G�Yp6m��:�c?/�LGr�a6`~�Ӗ�吸����<=�A���"�;+o82
�	�2�C��j�UJ�g�g6���K�H�JJ��҄��U\b�f���j���p-�����_K����
yܹ���5���VY;��"���O�>[jEQ�"Τ-��ㅡ�e�&�*,uj!y^�M2Z=��?���\vL�i���-��3���������_b����M1�o�x�<��kQ����pl�͔H�k���h܌o��-\nȯ}$4�w�r��Z�7��>9��#'glr@o����H�Ʒ�aǿ`��yl�� q�?�p=����_���li�Ϩ��bN��m���1�Oc/?[{I��vOoiԄ�-��OԜ3'�p�Xb��P0T��(���}��&">�C�D�R���U�/GY�n�	�V
�N-喝����K�ˑ��e�ȳ���i��X<ce��� ���]�Or��l<�� �o����!�M�Tb��4������,�����TY�����B"p�⚄$�1<d��[S�x�;�c�SJ�G���Q�z���8�r\�����Xf�0�2�x�H�zC_�.3�T�d/��o
i�u��e��a2g�IY�oت��	��c%#�;�t�Cuq�hCA�&ZH4�h�x
<QW^��P��,T$
G]̈�=�$8�
���O��r�P���H �wN��uU�X�-l/���������EC�Z��R �lc�r���?��|?pFU�B(���ް�����Uo�	x�^��~M/p��݄yV�%������(�+}�9�8zk�W~���-B�d���M.�"�4��:^.#<Z��/}2�	@a�o��E����ȳ
͎'�x}p�P���(��C=	�'ƾL�������L�^rBs�]��3����܏_Ӑ�t���z���@ۖ�=w%'�(�.�����sR7p+��%�0�l�&En�Q/����R��q��M3C�޲�z/�ًXd��0&�LD{*�T�E$�Z���EdNn��u���-�"�G/�� ��B��$?�؟��aI�p��	�tko�MK�4���bi�k�a�&uY�u��8\hv��a�`��@ȝ�ס̾�.����|l6���Ǌ5�9�3��B���G�Ƴ�����|�j�cg��g]��MI�>f�s���(��8�P���h&��#{����'��6i�ӏ�v j Q�ר��@7�*L�����ӝ���Nr����pD��L=�B7�3q�ԨǠ�	��NY���"���īIu���D�&��l"~)EAi�ݦ��ɨ@a����;�&c�X�6�����ϭ={o�Ǐ����.+ �.#J��{��lob�C�IB���ZIfvEĞ��f�={�L�{��;�ʠ�n�ˊ	}̺�=.��ߨ��Q��m����)�j�Vn��띖H���g�o�j�!�Ao��7�fH$��OK�b��Pi_pb�D�ȢIO�MT>�\.�Se�W~���^d��-Q�fua�����'��{m&'d��ը�%`�pk�F��#��/.&�t(i�&��⧔yDȗN�R�������*����\ƛ;�qA�W���+�ۇ�3����c�����)��p�癏�H̀�M��^�Nl8e�o�ڏ�=���k�Z��3NY��v[2�Q%,�<�0I] �[ ���.����v�e���6�"�xp��>!�T@����+n(�jɐl��`ȴ㏯����u<("@�:�_T��K1Lѕ�֕Q�π��n{�u[D&�Y��!�`�J�2wY<���fx�h�mGkl�qV��R�g"Ԧ��K.���`�D�ɭ@��PC�_é �mԜ�Ν-]pV5J��b�g��<���Ӯ�/d>����?�x3�-W��7�M�T���g�o��:˯��ڍgmOE"��u�;�~qFX&�������w6'�y���v����U���2b�"�& k�?��GT�� |�\�2,�oaT̎�y(�̂��xߗ'�F�9�{��0��Ȼ���F&�{�"u?ŧ%vp�f��S�M3D�Ǩf���� ��k��6j�,�˯��m*��lN�(���2�*��n��7<�Hq���Â�i��5l��d��Zٶ=V�!QD���g��[�>��u�w'��T"z��w��W�a3��b@� ��OBR.Wb:�X� �|��Ԃ�1�5q��}5H����RV��4�T�&_��km����װ�Ŀ��/���^��ގ�F^+>��]��H�g��`>PС�;@�F2%�1 i&.V����~�!����@�-���� �X#�Ӹ!���o1?���6�$t�e���
�Y����˝�d5_���Z��ƾ;��5AY"�#m$-T<*����(y��h8m�WO������:x��Y�$���7�w4�QY��F���Qk]�4�a�-���X���}gi�H3/�mO��~qvu_�Iy2B�E�[������{�r�" �S���cQel�\5}�
�C�������#���=�����D$�Av��H�ZE��/	h��dڅ-[0P�a�u�r�gٯ��:y�}#=�vۈy��@vg�Ti�����p��D8ZV�qs����23V7��c	���\+x4K�:�A�����P[�t�+�-��^��=�# 8�ơw׈�lI_Mv��i�߃pl��4��5�L�O$�U���#���5�F0{$*2,DC����!u?f���zu�͠��)�D]j��K՛�C��m.ػ����p��mo�d�G�n&��@Q}��Hu���.K8�Q1:Q3���Je'�c��X��g����S�:���J��߄�aJ�h�2�**b��~a��#���M�K]�M�����i��?�é)�y�����א/�뻝dP�F�X�Lpe�^��2����9�z���avD'���o�����L�(k*x�,,���uC14ؠB4���I��&���:t��}7��"���X��7�6��7r�Qt�9tL�p����n�?��ԩ^��+���}�� @]�gNI[ɷ�?�3^v�1O�9�-c�i��Ѓ��_,Ce,�6lWp�E0A��	��'��*�b�E�<�� �ێ��(��(��-$d?�{}}m4Pc�8h}��q�M�$��n� z���=����J�V�݅*k:�$X�����Ǡ�Ǡ��Z�X6�R���{0��� Dg�+X��㹛q����
2�a��1�!��kb�������9(9���+[nwzay4)��Q�:=(���4��=�nXzt9d`A`�wX��y�xXػ}�����Ml�����խ6���P��s0�y�����da���4u�&��3{"d	��<ZE�S\��\��oJ�V�S���x�Pۭ�f�r�O���x�دj.�O��x�`�l2Ըx��2��
.���XmUjT�f����
��'��i,�{����R�X�&G�߬(t�!��~Ӝ���x�Mj~�ߒ���!M�◓k��M�.9�(��A��ιf�eMq�g*���lmejJ��0����>�<�J���S0'Ts�o���<=�d»��yl0�*����5��^KE�B�z�>��z<����&7cW��a����Y�ٰ�a�ben*����G��D矫��d%D����z`kп���>��}�͊@���l�R^�+����o�P�˸���c��r�3F�MX|3�͈�SZ�u��G��"���N�*�C!����9i�QI����2Z4�r쩝\��fU�`�\�-A�]��]���������K���o\��%)6���:93 �F�AȚǽ��y�&��Z!K�Գ~�t^���a��w>ƝO_љ���ت�m�/6�a��2�|��C��15t��ݜ����=��[$�at馇�tw��m�#�j):�s��{�:f��nd��ĥ��#�$C��_�B�˛���<.�t���N���\�h�\�,�y��?J�w���'PI�21������C��9W #���1��k�t��ܧQ�͑?�4t����*�hM���zkN�OR����y\7���"�����Ё.N����4�@ �f�8�9�vw�н�尾�ǵ^�8��=)�KpܟK���&ik��9��� ��2{[�����Q�N)��>?�xU{kS|6*���X�mW��$XIC�n�H�t��an7��=��TR�(� Cb��G�BꚂ����L+�klF��nA;5�D4\Z�V���P���Ȑ4�qRV�;[6���p�:���J4�2�A���k�fZ��P�Q�����ZZf��z���9:/*i�	c��tP5g�ܮ�SV�����q]'�!1��s��Z�;��!s�OC�M1d��{��â�&4֍zm$[�<	cT��l�"X<�׿n�2p���w��Ե.	��$�O���\vl���{L9���k�^U0�nY͡�����P;�;��ӟ�|��O*�c�Ũ��0��$�$��ǱY����E칀��j�]"1��O:� �{��T:�R0�ªޠ�8i�����k�$>���O�g�B���(���iL�i��g���]M� �����g��vA ӽ��^�v���↊�z�X�����&EZ�0�$;���%�<%��dutL��ca�h��qh{��ob�C�z���@G���.���~�{���k�b���I�m
�#���iX3I�� \��j�iKf%0N؎�>_ ��aC`�W�4�Wj6�uI��-�����&��J2�=ƈ1��T!5�t����Ϙ��Ӹ0tp�7���7ŎL��chʋ�T�J/x7���A:�a��FbK(��<�� /�J�˖a�nH��}s��#C�<���;S���mi\F�b+u{n���G��M���y��lm�����#1̠�G��红�뽟i��R�;�^��XK1.^�L��g��k\�M8AN�㸲{��|��{�nRf��>F��n���V�w����D����Y�k:P� P��u�q�\^�;�L�ͤ�n��%vD!�~�6���6���z��їؙi��Y�A�����C�v������[R���D�e����7�	�c��P��y��m��\hO��E�L-(�{}5���-"��Qt�!����}�u����(H8�,��� �N����1%G0�d�,q�C��lϢ�h���2@�@�cF�!�������A^���"�����L1�����2"duL(g�����ɝ�\��g�!�Z~g�����b�	�����<��)
]��+.4r�`R/��?5��q=�{ZS&�1L������������ud6p�L-_���2%��4�L�N
R���HC'���?ރ"���#����Z���B�]鶷�⦮yA��7�!�χ �v�)(�+�ں�}nV�k)O�|N;�oƹN���;})7@
�����)�:5e�TK��L3��K�b�Ci�υ	�m(g����U���D�Q����H{��ė$��4L� ���}��K�|3��|<Y�^*6�"��P�1P�3���t;[�r����x�+���]�2��,ı�����"�D�J%B�l��V��f��;D�|����D$��ޏ���I
�%�@��b�|qp��O���G�y�s���c��l��<s�~�A��v".�سY4�/KzA���
��ߚ�ڲ!�Q��}m��}F4"�M�����ia?��T�Tt�c�Q-	��H��6�'���Jf$A�z�L�{����d�ft:�Kev�`c�~��N����2&�<z�u�K]�6�(��2
 8���R�{�&���BU��t�{((ȴB�;T`��]f'v��EHK�����H���]�8;ϙ�v-5�RJ��,9����7j��WM^�W�Ӊ�',ǔ-��e��] m5����m�?;�t�A��,㙴�#��>�5�pH�ߢ;�P��yL{�$QĿ���0&\X�fs�{�SH�a�'T�E�-����i��ݶ�WKsz+�;)��� =q��[� ?/�V��K��Y�Htb�z"�ZQ_��FJ��lB�9$.32ʀ�+����u�w^��Me����U��2���4�[���Z�j�[/�y��>B�'$"BX��,D�@�����{��NQR�����c.W�YZ�ߑ%/�&s/��ϊ8oy?aj��v�������D5q�ۖ)R�g����Jf��j��Ly�g�EɉI�Ӊ���ހs��4~GSܚ�*�MTZ�U>4O����#�ї��OLm|����Yz|�\�m�mmE"��|�x�e��3�lR���]1 ��p.�юpc$~��k�W�e�������f��~'���uyq��m�*ΘHı��_l�-���q.�w�򿺍���B�����o��'�N:J�5-b������f����^�82������R?H���#=�}0�Cm�����sfC�����ѫ�=˂*����J������,�=*Y�FpLH��̽��U�Z�r���nNC}E�6��BK��1/���e����zwj���wa�9JƳ"����h� i4�r�j2 K��A,�㻄�;�m.�C����&�YG�_��T�_�������D��l����PRS�ĝC�O�?�+v&�����>�:ųQ)z�k����-�b
=d����z���iU����n�8o''y��K���e��ϭh_��+�A���-`^�8*�_��ezs�E>�ښ��L|��.������ٜ���G]3�s�\x�e���f֕Mv�[����q�Oy��Q`���Z.b��v��8�1����(ؾ�f?z4��F��w�I����钹��������}*�6a?T�Еo�h�9`�o�\���/:k��Z3qYd`PE���x�H�P���W��G��l�YY��A�:����2,�Cc�ur"� Y����#�S�ɖ��z�[���v��۷k���R�~SP��|��8i5��Q���5��˥6-�ǸJ��bh��G��BO8�?�����Ds�!qw��m�S����u�Se�bo��R�9�K�w ٳ�;(sE6�C�N$��y��-SJ�׀��&��d�2�f����Ta����.�B��WPJ�������p)�Ս��#�_ yL>���xچz��K��\�ˉ+"w�@��u�#��~�l�;��`��>i���A���1�ע=���<�o� �у���ęx�֮��p�O������Lg^�tޭ��Arݎ������<�;�qk�#�i:�
���|toO��̤��av`?�t���RϝH�m���}�6�e�zX|Cf�f���+��@lh#%���F٧֓ߘ���%p�χ�}M�W�!��ɷ���φ� ,4-D@�(���NL���uQ�l���Qo��͒tL�q`��D�g��:bm�&�U��U��p+�$��
��	��$�7.��uv�&�܁B�|\1\y�`	\�?�Aŀ݇{��9V/�q�����R���WZQ��I����܁�����]�,�l)����_",E�S�T~���Dl��̍(��F��$�WHz�ݩ�/�t�"�β��f+d�cSU�S���i̝U���Y�S�]�4�ekOK(���.YA=
:w�?��v�0�?����a�_$��0>�D�s����u׮�KF�E�:�D����\��l��w����Bt�w�ҥ#?6e���@77(�*���$� ��'u��B��)u��l7amg�5�*�C�3��࣎��������c����oq�y�7?[i�o{�@������+�4f�7��'I6����:��HJ�[Y���\C[�F����[��UQ5���u�:)�+��6���Q�~������)�H��D���Y�: ��E���Ȑ��]!�SD��m���Y��e�uū\������d#gd�y?���9k�R9ʡ��W�%�G\>}��DY�o]��մ[Ũz87gn���{�򰈦~�y���[E��^�Ew������5��LsB
6k����WT����@x/�!I͡�]��9l��m�%X�Y4� ��������3���H�s�F%�J�/�B
� 2 T̻���8*)��ok(�y��:��l�d	F�0�6
�����R��OȔ8	=D=�RN��^�'C��L|p֨ ��om�y/Y�r4O�����@Q����(>�-	�-喎�p��^��0��W��S��"�6�^(�עAj��ݚR�)��2��b|JT�c�U�MD؞�M��ղ�^u�����ì����a��mD��4oA���R۵���.2{х��"Ru�K`�7�be&=	��<��2^v��G&4x��
+��lKq�d��Y$�u1��ЫC2�ȳRȮ��ܟ�����Լ��-� �8�����lh��(( H�"� 5*A:>�H	R�J｣����ނ��!t�#%��;!� ��$�z��}���|;�ff�5k�5g�f�@h|�����|��[�2�d��K�d�#o�7ת���̹
΀?;��3��/O��n6\����xI��p˶���������J���z���j�?�}��Gj��Ճ赋˟��I�"��_�'Tm+����m֥|7K�<��S	����wS��nx�[��x4�}�m��܂�2<_�
��u��ffE�H��!W%��k/I�z�k��J%.�m�%ʟq[��H>p��E���g��G2ۿ^����o~��a�ῐ���?�M �<D�e:���<���5L-���Du�{:���u��w��+s~���Z�.'L�K��0d�j�� ��7�l��� �Kfs�NN4hu=�t�^[ݜ%�f�.|ё�/X ��I;�9�r�+���U�9�,�N���S�ߠ&N���B��hV䨾$^�&�K����V��j�\�
G��}�Qj�[����Ȋ?)��wKd}�S\~��Y3:��5��a�;;77�C���p9�D�-�o�4gTBr�\�Xj��NГ�%f!V{��i��r��s����Σ"�*VjE�J�f�iK�N����޹�uY Dw�Q{$�|�x�gӠ�5jmPx��4�H��M�-+��
%C,xk���l���=��޾V
���Tr�2�H�G�6/�9^�rF��jJF8����ֳ���O^���ޑjK�@��LƵ�~y���S�[�t|Uk�"����ֽߧ��n���3L,�Y ���B�0�0�-|(���Fd)��	 �?˩Q�!u�IB.�`�?���)�ov��A����=�����]�[_QW廭����BN�YF������h����D檉�l���l�:�~���ו�d����\ZE�~�"��kYd���RA3e�DU���d�ef�J��6�L����������ZL����x���\�D�o�`�4��s>�6�4Y=d��1�D�c���sg�Ds�`Jo���=:� P�H-OZ#̺&]2`TүZ�^��H�X$y����@aED�������-�@�5Zb�d"Z"����3�%о �HcM�R�z=݁�\i���
�)�4WM�Pm�,�]#E�</�x6�����R�g�������x�lL����U�5Ʋ�l{M�W��E�iS��ʄl�T�@t
Q�d�F��ի���)
���~�.͘$���e� �)��,)B����X�^�R�O���g��r8��r����%W
�̺-I��E�I� ��=ΎF�^Sw���f
�_"I�C��GҲ�t-Y"�I{�i˔K#��y���n����<�e�q�U�8y�(Y����7�SJW�5��y�;�$����+\��$�T<k!k�7�v�j����c{�<�ͱi�?�������v�-yMaG8_Z�a���I%�vX�1�m��5��UwL�h[���G0��,�@F_�;���@�RN����5̶l�6���z��H5�6��͈�D�ה�W��E
�8]�w�b;��-���(�Q�ՇX�E��Q+�U�WFް#��A|��z�[������S#JZ�����b	s��A�������6'���,Rz'< %�G�H�p�;�8j����{�P�{At
D��*Η�T��d0k�=�
ˋ"	̀&E��8���}�<{�q��h���L1���p_�0�ܙ�.a�@�s����5蹋J/��,���`^% �A�j�>�I�!���a�:3��LحN����)�{X���7:�i`�Z�<e�g���$�<T2���.=p�>������q���B%hG̐����
�&\Mb�O9o�Ȯz���y�"�WxƙP��������gk��(�cE�Y�&��C�˃�Z0��DA�1x��_�D�k@�ǎ+'�D��AG$�u�(�p�W~>��U_tX�����yw$�S!�M6ؔN����A¡�(��F���	��I=h���am��؈Қ��X�g��9����a���X�&��f���+�8E0���K?�G���; �Wc��Ri�@��j���c�ϩ�_N������")��dBf���!k-�ٍud;;��)��[���ǵ�7]���J��m����=1�C��������Ҩ1�wr!���-��W������Ȏ�/��n�T�%�\pᅦK������'JsۿW66�*0�~[.�i��"���ދiG��4X�)��]�c���̧Zl��d���@5��&��w���e�.O���/�j�7�9�Mdh�?��<BP�#><����Y����ܵa�mʔ�6*&l�"�J/�St�v�B��� �t�T��n�ݑ�����IL�����S7�4���U��)���F��m�#��֬��=ʖ��8�箤�����T�c[�2�!Ԣ�sL�9!�gA5��@���GA���r2,b���}랰ST'S������@*��iu�^1W�!�8'��%�+j�
�x�a���"�ݕb2U/�IX>{>�{I�p�Zݖ3Y�Rի*���-��6 �Τ>��o�5Z�^�x����t��L�Q誄j�$O�x�"�-�2e��!��1Vi:��Sn�̤Vz��oF�bc�ئX�8��x.; ���N�(����6��~5^>MI}�NZX٫A`Έ�ң�D�Ÿ?k����7�܇3�B��z8w��-1�T���E�c�;NO7�{���#�u��,Q&&�_��7�	K�E<�%��b��}�z�{	ߎ���л�aC��k9�?��<�?��Od�7S�v&L�X:��+[ܬv�4��c@�3�>����5�����K�+���*eJ��I_̔~�AZ�W��
�XJJ�!���X�e'�''�K��Z�C�ŉ��^�p='��ջ������M~H�ŭ�,n��^���'Y��}�Ӝ׵a����M�]1&|!9ƞ@����o�q��~XY�N��Z�u刍�Ό	�Ẅ�$7A�sZ�J��@T[�[w��A]õ��.m��5���'��nc�-��-����<�ƍBם�L���rc/Gq�̧Z�M���쮝a�!�_#���fk�oE�~m��ǎ�M؅����8�U�$���B�Y�l|ME�8�`�H;�y�)ܑ�\]Z����o1+���1���EQ�m����0\ɪ�L��$�������\�$�[X@���K�a��m{nF��AEk��z��˄����{|MM�bm�0������_�P�����Mm:��Պl�.�p�&@�O���hE������ݣGDף���7S�_��G7���sx�Y�_k��с��! :~_�9k̥�N&��cT~��A�T/"GtY���1c���Q&��u��.Q,�	��rD�ڻ�T�����^�������4t?��R)7!�@��$�I!Y�{X�6&ݵH��ݓ�}^��d����JSCMQ�<��"���Z�e�wSM�C�V�j1�4���ҩ�fa ��0hD��԰����/R�*�><5�h�S�ƺ-��Ox{��o�ڂڋ�͢�Y��P�gA��`��q��R��vʷ����m9 ��؉���	j�2n�)��s����:���T�i����.��i}��3�D]0!z�Oi�=𖧰�l�1���k0|Y����؃� ���֋�ߨ>	&��dR˭&��}�~st��w%F[�9����l����u�-v���9�����O��oYCKj��YՏ|^�����z���ޓ�͛��`;�����&�_�cM�(Qh��c�����|5�_�e@@�4�)Z�6��Ƕ��/NhR� �O^��'��܋��+ڶWj������so�ZQ�k+*>�.~V)%k��	](�X�i#��<	��-��ɱˣ�A��:q9��6�-)�����<��v*�y�J>��~sk����&_V�(�5�D�0>�i�S/[!��o��k�*��1D��BZ\�U���k��J.v9�����L
�h �j�*����M�Юնfa��H
W]O��=�P�[؀g�)ָ5I)��=�:���H�*���*%��Ū|�㱱�ݬ�7�|�F]'����ՆO�ls/�˩��Cr@d�̸���Sp�%���๚@C��a����yy"V���K15 �on�X�F!�Ǥ�Sg�h�R��.�l�ø�W^�ksAz�E��+�aJ�qmAL��Υ���G�Z��R�PW���W`mN��Vmo�pã}��%�3kh0
��m؁�r�ӄ���L>ǵ��6&����ݠ[���x�xn�Δ C�y�U2�)%V�񁆌���%��E�2yVQ���I�i�d�^m�l�	� ߉fOd�<��@�j �o����{���"2&����	�t�*�P�ܻR�m��6C���8��DK��l�]1ͭշ�$��fV�l�R��ψY��7����p����F �����_B C� %�ֱH&�8X�+�SJ=7~��FLe߆���y��Xc�Q�hp2�A�|@�SH n��q�g��f�.�~�����'���I.i��gx�^�o�j��5��R=N*��}�Gf��G*�KV��Ѹ��a�D����E�o�!Cd������ý 3q�2��}n��6n`Z��B�W6i�񡛨s��l�M����b�?�`
:�/�;X�C"�^9]W��̈�)^:����/�Np��;�s��N�5����
)�������Y��xy�x�)��5PwK���+��Պ5�%��{���-��z��#�7���߀X��|�c^�Ģ0�C;��K<�R��ڝ����r�p{�"X�|SP�'�ug�Ŀ'A�u��IUI?��}��H�E�u��xfoK�O��E	�H�MҀdG�xu���*���ԣ��Aqc_��
E�?�j?j�����@� `K�c
��*p��W�μĲ�z�>�$8�d���y�r5��`=����Z�5XA�zZ]�F�y�͊����P��ђ)h'�y�i0k��I'&�U�F䄾�� �/�(%">��V#&��W���c�o�����_�]+5rc,+��F��+�Wu�kn���t�K*S\#�7x���3V�`Q�O����-USj.)�AO�t q�͗S����.g�G�i�c��y޹�M�y'4�HZC�{�i�˒T_4��Y��~g3�r�a\i@��u3l��*���s�%/�?a?>�$M	�uLq��"�[ IDs��W�x�Q+�����<d���E7����{�����;X�'|G�c<gN��./Z2v��As�qcᾞ�c�R�<:^��/%���Y��]=[��<g���ѕ�U�����M��= ��(�F�E� �p��[G�����}��IukW�K�$��W�e�������7Ҏe�pĤ���Ճ�������?��+=�*�]+g�)!$�xv^
����
�������n�H��Tmr�K�]~�%��{2�� s:r�+&.�
a�ɣ�F�
}}P�����J���+�Z�pN��n�c��*�~8�xj�O)�{��ǟ �Ub~LFHWB�2���i����6�:S{e�!Co��t��\��^�X��+Xb$lk�>8���k��m��FM�(T@ڡ ��E�ɍL"s�~T���e����m�ig��������-�=dÁ��XL�<4W5=z��ZO�Ƙ��!��%Ţ1U��r�N��qz��6��������t�`����{go{����IGWM���`�t����p�%T_B�����t��3:���xx�w_�v+�G�
����8�_���e��$py��~��=Dx*��/Y��k�mң]x�AC�;�$�꘧���2|�톨#���;i���!�ߡ졒oǭK��El0�� l�<�ȴ�}����������O{H�x��*A:_��b��?���A��S�����:�8.!&��ƽZb�d1
����E�Y�>Ŵ�&��6��l�{�e���W�U� ���,��ל��AM�_Ѻ��o�8oi�&�6H2�V��$���f�Y��o��9���m�u�u�hl��$��Kq5�����	m~�{y��5��cr�Z菖���oB�3�a�xJ�}�����L3L�Ę[������\�H|���G����|���[_)�v�fw����f��!h�A�n)X�9������&Y�B�x�@����
e����3\ɮA�g���	�����J�=
(�I��C������w%y�We/��PK   vOX�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   vOXu}6x  
&     jsons/user_defined.json�Z�n�H�A��ũ}��Jg����n``�1&F&�Z:���)Z����r�1���I"���Z�9U��:^}����x��ΗU���`��_,��7`�,צm�����s}�>{�t�XW�����J&�B{�W�S���?5�< M�8���-���
_ǥt�!�Q'��
���E����]���j��$��~Y��[!��e�X2�5U���*e�"Z��Sxn^�'uٌ������Z�g��q3����jw����Ő x`3(��c�O�t��B�0zm�fY�y�U�p�SU��s�6_dhR-�j{�,�����b�d��o�ߜ����GG��l]D�o��1���I4<>	�?�|<����B��B��%F�v��m|���:����?���ϻ<0��U*���0��b��AX�)F����D����Q �����>��z�U��E�o�Ң��Ūڪ�Vʖ�@ڍ<���V��l��"���]m���|Q7��'�V�n�eef������~�}�g����ץ����/�p�D�v�����ƥ�M�Q=�)e�+��-��2��
o<f~�z6�4��W7�B�B�{�ɟ6A�7�:_g��w�a��W���K�GD�.A���_C�G��}�w�J��iB�(�5`�K͡�AVz3��Lc��Y>��J
��
P�PY@XYR.���lGd7��j_+\)(���a�Vذr�%F,m-��#����C��K�ҕ�+ R�|[2���2�������w P�= �	����sp4~�������)��1����@|���_�Ƨf/�ʞa>�a� �FQ�D@��E����.�H�!�R��ZсPq��Z�\�H�GQR/P�`�"��b�\ɸ�=ы$�Q.��SIZ�l^��$�Q6�1�C$�����ZQ]rc>T��M�A�����e��Y��%� ߢ㓀����2n:�/$�%� ۢQ�=g@>�BS��.�w �\C�!��y�o�q��]2� �M�M���p�� NQ9�DqܧI���J�K��؜o�$��H���J���s��~ ��JR����i��CR��v��e E�l�|��A����InK�Kh1�l�U׹�.��;�^���Y�ᤞ��Uf)�G��@
� &$����R�K��ͭ2S�)�%�!TM��Z���Uf\P�do����&bX�cT@��	I;+�*v�.���]�^�}@�yCy6�-}�G�^�L���8J�L��/x�v����)�lz� ��ӟ�E���o����po^���k�شeJ�8P�	ꡆ\hޮLy�~r8��܌��z�i�}��8�7�J#<A� ˘���Ry JF<u�x�<�UBz��Ǳt�R`=��v�	(Y�JM�$�ve�EX��bu���&\HѮh���}�"m ����E���k�O�DO.( )�B2�F�l��P����	+�\�
+- �l+�[��7�v����:=��A�W0��E�]`�[sU:�0�p/4�FX�U�9� v��R�7�����%�h���������x��^�il�E I:����Zm\,�׾W��Q��׾i�� 6e��F��{A��4��𒆇L�=(xP)Kv%��~��
���o��n�L �
>"��h��"/H��?��l"$~)�3��6�y a*�����xA�煵zL�f�?��z�6B3���=>M.�8+�C-�����M�^��A��.�h��?qX���@!��@��QωIt��Up�������P��H���+�l��A�a*N9߮@�aWDY�d!�D�?�XA1c*�ʮQ<�gK"��=8�U�?4� J��	﹐

+\�x��kd�r`����<�)�B?�^��h����0܊o��PK   vOX���l  %�             ��    cirkitFile.jsonPK   vOX��g  n  /           ���  images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.pngPK   vOX�j�� 7q /           ��M(  images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngPK   vOXhT���� ċ /           ��� images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.pngPK   vOXS��lG  bG  /           ���� images/52445b69-20cf-48af-a05a-7b7247ebe25e.pngPK   vOXإl˨6 �= /           ��@	 images/734bc482-36f4-48b6-9076-7f88fee16b3e.pngPK   vOX	�\  \  /           ��59 images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.pngPK   vOX�R�{� �� /           ���U images/8b783ee3-b9bb-4285-aa49-cf7c99b593a7.pngPK   vOX�1.:�  )  /           ���� images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK   vOXǐ]zd� K� /           ���� images/972a987d-5ae9-491b-9c1c-35ff468aee03.pngPK   vOX@��)  /           ��v~ images/b4aefdef-6992-46c6-bd27-cdaf728c7c35.pngPK   vOX��n�% �, /           ��� images/c1d4a215-2c3d-48ac-b15d-f6239b4c4b94.pngPK   vOX�GDU7� �� /           ��W� images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK   vOXu}6x  
&             ��۝ jsons/user_defined.jsonPK      �  ��   